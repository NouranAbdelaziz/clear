magic
tech sky130A
magscale 1 2
timestamp 1650894151
<< viali >>
rect 2605 20553 2639 20587
rect 3157 20553 3191 20587
rect 4721 20553 4755 20587
rect 1501 20485 1535 20519
rect 2237 20417 2271 20451
rect 2789 20417 2823 20451
rect 3341 20417 3375 20451
rect 3985 20417 4019 20451
rect 4261 20417 4295 20451
rect 1685 20281 1719 20315
rect 2053 20281 2087 20315
rect 3801 20281 3835 20315
rect 4445 20213 4479 20247
rect 2605 20009 2639 20043
rect 3249 20009 3283 20043
rect 4261 20009 4295 20043
rect 3801 19941 3835 19975
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2789 19805 2823 19839
rect 3065 19805 3099 19839
rect 3985 19805 4019 19839
rect 4445 19805 4479 19839
rect 4905 19805 4939 19839
rect 1501 19669 1535 19703
rect 2053 19669 2087 19703
rect 4721 19669 4755 19703
rect 2053 19465 2087 19499
rect 2789 19465 2823 19499
rect 3617 19465 3651 19499
rect 3893 19465 3927 19499
rect 4537 19465 4571 19499
rect 1685 19329 1719 19363
rect 2237 19329 2271 19363
rect 2605 19329 2639 19363
rect 3433 19329 3467 19363
rect 4077 19329 4111 19363
rect 4353 19329 4387 19363
rect 1501 19125 1535 19159
rect 4261 18921 4295 18955
rect 10517 18921 10551 18955
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2421 18717 2455 18751
rect 2881 18717 2915 18751
rect 3985 18717 4019 18751
rect 4445 18717 4479 18751
rect 4905 18717 4939 18751
rect 10701 18717 10735 18751
rect 1501 18581 1535 18615
rect 1961 18581 1995 18615
rect 2605 18581 2639 18615
rect 3065 18581 3099 18615
rect 3801 18581 3835 18615
rect 4721 18581 4755 18615
rect 5825 18581 5859 18615
rect 6929 18581 6963 18615
rect 2513 18377 2547 18411
rect 9689 18377 9723 18411
rect 11529 18377 11563 18411
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 2697 18241 2731 18275
rect 2973 18241 3007 18275
rect 3617 18241 3651 18275
rect 3893 18241 3927 18275
rect 4813 18241 4847 18275
rect 6009 18241 6043 18275
rect 6745 18241 6779 18275
rect 7389 18241 7423 18275
rect 10057 18241 10091 18275
rect 10977 18241 11011 18275
rect 11713 18241 11747 18275
rect 6837 18173 6871 18207
rect 6929 18173 6963 18207
rect 8401 18173 8435 18207
rect 10149 18173 10183 18207
rect 10333 18173 10367 18207
rect 6377 18105 6411 18139
rect 1501 18037 1535 18071
rect 2237 18037 2271 18071
rect 3157 18037 3191 18071
rect 3433 18037 3467 18071
rect 4537 18037 4571 18071
rect 5365 18037 5399 18071
rect 8033 18037 8067 18071
rect 9413 18037 9447 18071
rect 6745 17833 6779 17867
rect 9965 17833 9999 17867
rect 2605 17765 2639 17799
rect 6101 17697 6135 17731
rect 6285 17697 6319 17731
rect 10517 17697 10551 17731
rect 1685 17629 1719 17663
rect 2145 17629 2179 17663
rect 2421 17629 2455 17663
rect 3065 17629 3099 17663
rect 3341 17629 3375 17663
rect 5181 17629 5215 17663
rect 7021 17629 7055 17663
rect 7941 17629 7975 17663
rect 9045 17629 9079 17663
rect 11069 17629 11103 17663
rect 12909 17629 12943 17663
rect 21097 17629 21131 17663
rect 4914 17561 4948 17595
rect 5733 17561 5767 17595
rect 10333 17561 10367 17595
rect 10425 17561 10459 17595
rect 12541 17561 12575 17595
rect 1501 17493 1535 17527
rect 1961 17493 1995 17527
rect 2881 17493 2915 17527
rect 3801 17493 3835 17527
rect 6377 17493 6411 17527
rect 7665 17493 7699 17527
rect 8585 17493 8619 17527
rect 9689 17493 9723 17527
rect 11713 17493 11747 17527
rect 11989 17493 12023 17527
rect 13553 17493 13587 17527
rect 21281 17493 21315 17527
rect 3433 17289 3467 17323
rect 5733 17289 5767 17323
rect 9413 17289 9447 17323
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2605 17153 2639 17187
rect 4077 17153 4111 17187
rect 4353 17153 4387 17187
rect 4620 17153 4654 17187
rect 6377 17153 6411 17187
rect 6644 17153 6678 17187
rect 8033 17153 8067 17187
rect 8300 17153 8334 17187
rect 9689 17153 9723 17187
rect 9945 17153 9979 17187
rect 11529 17153 11563 17187
rect 11796 17153 11830 17187
rect 3157 17085 3191 17119
rect 1501 17017 1535 17051
rect 2421 17017 2455 17051
rect 11069 17017 11103 17051
rect 1961 16949 1995 16983
rect 7757 16949 7791 16983
rect 12909 16949 12943 16983
rect 2697 16745 2731 16779
rect 2973 16745 3007 16779
rect 13277 16745 13311 16779
rect 6653 16677 6687 16711
rect 4353 16609 4387 16643
rect 5273 16609 5307 16643
rect 8401 16609 8435 16643
rect 9505 16609 9539 16643
rect 10057 16609 10091 16643
rect 10977 16609 11011 16643
rect 11897 16609 11931 16643
rect 1685 16541 1719 16575
rect 2237 16541 2271 16575
rect 2513 16541 2547 16575
rect 3157 16541 3191 16575
rect 4169 16541 4203 16575
rect 5529 16541 5563 16575
rect 7573 16541 7607 16575
rect 8217 16541 8251 16575
rect 11253 16541 11287 16575
rect 12164 16541 12198 16575
rect 6929 16473 6963 16507
rect 9413 16473 9447 16507
rect 1501 16405 1535 16439
rect 2053 16405 2087 16439
rect 3801 16405 3835 16439
rect 4261 16405 4295 16439
rect 4997 16405 5031 16439
rect 7849 16405 7883 16439
rect 8309 16405 8343 16439
rect 8953 16405 8987 16439
rect 9321 16405 9355 16439
rect 10333 16405 10367 16439
rect 11161 16405 11195 16439
rect 11621 16405 11655 16439
rect 2145 16201 2179 16235
rect 2605 16201 2639 16235
rect 4629 16201 4663 16235
rect 6745 16201 6779 16235
rect 7849 16201 7883 16235
rect 11529 16201 11563 16235
rect 4997 16133 5031 16167
rect 8984 16133 9018 16167
rect 10149 16133 10183 16167
rect 1685 16065 1719 16099
rect 1961 16065 1995 16099
rect 2421 16065 2455 16099
rect 3229 16065 3263 16099
rect 6009 16065 6043 16099
rect 7113 16065 7147 16099
rect 9505 16065 9539 16099
rect 11897 16065 11931 16099
rect 2973 15997 3007 16031
rect 5089 15997 5123 16031
rect 5181 15997 5215 16031
rect 7205 15997 7239 16031
rect 7297 15997 7331 16031
rect 9229 15997 9263 16031
rect 10425 15997 10459 16031
rect 11989 15997 12023 16031
rect 12173 15997 12207 16031
rect 4353 15929 4387 15963
rect 1501 15861 1535 15895
rect 6469 15861 6503 15895
rect 11161 15861 11195 15895
rect 2697 15657 2731 15691
rect 4261 15657 4295 15691
rect 6561 15657 6595 15691
rect 8953 15657 8987 15691
rect 5365 15589 5399 15623
rect 8309 15589 8343 15623
rect 3157 15521 3191 15555
rect 3341 15521 3375 15555
rect 4905 15521 4939 15555
rect 5917 15521 5951 15555
rect 7941 15521 7975 15555
rect 1685 15453 1719 15487
rect 2145 15453 2179 15487
rect 7685 15453 7719 15487
rect 10333 15453 10367 15487
rect 11253 15453 11287 15487
rect 3065 15385 3099 15419
rect 3801 15385 3835 15419
rect 10088 15385 10122 15419
rect 10609 15385 10643 15419
rect 1501 15317 1535 15351
rect 1961 15317 1995 15351
rect 4629 15317 4663 15351
rect 4721 15317 4755 15351
rect 5733 15317 5767 15351
rect 5825 15317 5859 15351
rect 2329 15113 2363 15147
rect 2789 15113 2823 15147
rect 4629 15113 4663 15147
rect 7205 15113 7239 15147
rect 8217 15113 8251 15147
rect 8769 15113 8803 15147
rect 9137 15113 9171 15147
rect 3709 15045 3743 15079
rect 5742 15045 5776 15079
rect 1685 14977 1719 15011
rect 2513 14977 2547 15011
rect 3433 14977 3467 15011
rect 4353 14977 4387 15011
rect 6009 14977 6043 15011
rect 6377 14977 6411 15011
rect 7573 14977 7607 15011
rect 10894 14977 10928 15011
rect 11161 14977 11195 15011
rect 7665 14909 7699 14943
rect 7757 14909 7791 14943
rect 9229 14909 9263 14943
rect 9413 14909 9447 14943
rect 6561 14841 6595 14875
rect 1501 14773 1535 14807
rect 2053 14773 2087 14807
rect 6929 14773 6963 14807
rect 9781 14773 9815 14807
rect 5733 14569 5767 14603
rect 11805 14569 11839 14603
rect 4077 14433 4111 14467
rect 6929 14433 6963 14467
rect 1685 14365 1719 14399
rect 2237 14365 2271 14399
rect 3433 14365 3467 14399
rect 4353 14365 4387 14399
rect 6653 14365 6687 14399
rect 7196 14365 7230 14399
rect 10885 14365 10919 14399
rect 11161 14365 11195 14399
rect 2789 14297 2823 14331
rect 4598 14297 4632 14331
rect 9137 14297 9171 14331
rect 10640 14297 10674 14331
rect 1501 14229 1535 14263
rect 2053 14229 2087 14263
rect 6009 14229 6043 14263
rect 8309 14229 8343 14263
rect 9505 14229 9539 14263
rect 2421 14025 2455 14059
rect 5273 14025 5307 14059
rect 5733 14025 5767 14059
rect 8769 14025 8803 14059
rect 9781 14025 9815 14059
rect 9137 13957 9171 13991
rect 10793 13957 10827 13991
rect 2145 13889 2179 13923
rect 2605 13889 2639 13923
rect 2973 13889 3007 13923
rect 3893 13889 3927 13923
rect 4160 13889 4194 13923
rect 5549 13889 5583 13923
rect 6377 13889 6411 13923
rect 8042 13889 8076 13923
rect 9229 13889 9263 13923
rect 10149 13889 10183 13923
rect 10241 13889 10275 13923
rect 1501 13821 1535 13855
rect 8309 13821 8343 13855
rect 9413 13821 9447 13855
rect 10333 13821 10367 13855
rect 6561 13753 6595 13787
rect 3617 13685 3651 13719
rect 6929 13685 6963 13719
rect 2789 13481 2823 13515
rect 5549 13481 5583 13515
rect 9965 13481 9999 13515
rect 12265 13481 12299 13515
rect 3893 13413 3927 13447
rect 4813 13345 4847 13379
rect 8309 13345 8343 13379
rect 1593 13277 1627 13311
rect 3433 13277 3467 13311
rect 7297 13277 7331 13311
rect 8125 13277 8159 13311
rect 9045 13277 9079 13311
rect 11345 13277 11379 13311
rect 11621 13277 11655 13311
rect 7021 13209 7055 13243
rect 11100 13209 11134 13243
rect 2237 13141 2271 13175
rect 4169 13141 4203 13175
rect 4537 13141 4571 13175
rect 4629 13141 4663 13175
rect 7481 13141 7515 13175
rect 7757 13141 7791 13175
rect 8217 13141 8251 13175
rect 9689 13141 9723 13175
rect 1501 12937 1535 12971
rect 2237 12937 2271 12971
rect 5733 12937 5767 12971
rect 9873 12937 9907 12971
rect 6377 12869 6411 12903
rect 7849 12869 7883 12903
rect 10241 12869 10275 12903
rect 10333 12869 10367 12903
rect 1685 12801 1719 12835
rect 2881 12801 2915 12835
rect 3801 12801 3835 12835
rect 4077 12801 4111 12835
rect 4333 12801 4367 12835
rect 7113 12801 7147 12835
rect 11897 12801 11931 12835
rect 6929 12733 6963 12767
rect 7021 12733 7055 12767
rect 10425 12733 10459 12767
rect 10885 12733 10919 12767
rect 5457 12665 5491 12699
rect 3157 12597 3191 12631
rect 7481 12597 7515 12631
rect 9321 12597 9355 12631
rect 11529 12597 11563 12631
rect 1869 12393 1903 12427
rect 2145 12393 2179 12427
rect 3157 12393 3191 12427
rect 3893 12393 3927 12427
rect 4813 12393 4847 12427
rect 8953 12393 8987 12427
rect 9781 12393 9815 12427
rect 12081 12393 12115 12427
rect 2789 12257 2823 12291
rect 1685 12189 1719 12223
rect 3341 12189 3375 12223
rect 4537 12189 4571 12223
rect 6193 12189 6227 12223
rect 6653 12189 6687 12223
rect 6920 12189 6954 12223
rect 11161 12189 11195 12223
rect 11437 12189 11471 12223
rect 19717 12189 19751 12223
rect 5926 12121 5960 12155
rect 8401 12121 8435 12155
rect 10916 12121 10950 12155
rect 12725 12121 12759 12155
rect 2513 12053 2547 12087
rect 2605 12053 2639 12087
rect 8033 12053 8067 12087
rect 9505 12053 9539 12087
rect 12449 12053 12483 12087
rect 13185 12053 13219 12087
rect 19901 12053 19935 12087
rect 1685 11849 1719 11883
rect 2697 11849 2731 11883
rect 4353 11849 4387 11883
rect 4813 11849 4847 11883
rect 6745 11849 6779 11883
rect 7113 11849 7147 11883
rect 12173 11849 12207 11883
rect 12449 11849 12483 11883
rect 2237 11781 2271 11815
rect 6377 11781 6411 11815
rect 9680 11781 9714 11815
rect 13645 11781 13679 11815
rect 1501 11713 1535 11747
rect 2329 11713 2363 11747
rect 2973 11713 3007 11747
rect 3240 11713 3274 11747
rect 4629 11713 4663 11747
rect 5457 11713 5491 11747
rect 7205 11713 7239 11747
rect 7757 11713 7791 11747
rect 8024 11713 8058 11747
rect 9413 11713 9447 11747
rect 11529 11713 11563 11747
rect 12633 11713 12667 11747
rect 12909 11713 12943 11747
rect 19257 11713 19291 11747
rect 19717 11713 19751 11747
rect 2053 11645 2087 11679
rect 5549 11645 5583 11679
rect 5641 11645 5675 11679
rect 7389 11645 7423 11679
rect 5089 11577 5123 11611
rect 9137 11509 9171 11543
rect 10793 11509 10827 11543
rect 11069 11509 11103 11543
rect 13277 11509 13311 11543
rect 14105 11509 14139 11543
rect 19441 11509 19475 11543
rect 1593 11305 1627 11339
rect 3249 11305 3283 11339
rect 9321 11305 9355 11339
rect 11897 11305 11931 11339
rect 8953 11237 8987 11271
rect 10977 11237 11011 11271
rect 13277 11237 13311 11271
rect 19441 11237 19475 11271
rect 3801 11169 3835 11203
rect 9965 11169 9999 11203
rect 14841 11169 14875 11203
rect 1409 11101 1443 11135
rect 1869 11101 1903 11135
rect 2125 11101 2159 11135
rect 4261 11101 4295 11135
rect 4629 11101 4663 11135
rect 6745 11101 6779 11135
rect 7021 11101 7055 11135
rect 7288 11101 7322 11135
rect 9689 11101 9723 11135
rect 10333 11101 10367 11135
rect 11253 11101 11287 11135
rect 12173 11101 12207 11135
rect 13093 11101 13127 11135
rect 13553 11101 13587 11135
rect 19257 11101 19291 11135
rect 4874 11033 4908 11067
rect 9781 11033 9815 11067
rect 12817 11033 12851 11067
rect 14105 11033 14139 11067
rect 14473 11033 14507 11067
rect 6009 10965 6043 10999
rect 6561 10965 6595 10999
rect 8401 10965 8435 10999
rect 3065 10761 3099 10795
rect 3341 10761 3375 10795
rect 5457 10761 5491 10795
rect 6745 10761 6779 10795
rect 7113 10761 7147 10795
rect 8217 10761 8251 10795
rect 9413 10761 9447 10795
rect 15025 10761 15059 10795
rect 6469 10693 6503 10727
rect 8585 10693 8619 10727
rect 9873 10693 9907 10727
rect 13461 10693 13495 10727
rect 1685 10625 1719 10659
rect 1952 10625 1986 10659
rect 3525 10625 3559 10659
rect 4077 10625 4111 10659
rect 4344 10625 4378 10659
rect 7757 10625 7791 10659
rect 9781 10625 9815 10659
rect 10425 10625 10459 10659
rect 13737 10625 13771 10659
rect 14381 10625 14415 10659
rect 14657 10625 14691 10659
rect 18337 10625 18371 10659
rect 5733 10557 5767 10591
rect 7205 10557 7239 10591
rect 7389 10557 7423 10591
rect 8677 10557 8711 10591
rect 8769 10557 8803 10591
rect 9965 10557 9999 10591
rect 11713 10557 11747 10591
rect 13921 10489 13955 10523
rect 15761 10489 15795 10523
rect 7941 10421 7975 10455
rect 11069 10421 11103 10455
rect 14197 10421 14231 10455
rect 15393 10421 15427 10455
rect 18521 10421 18555 10455
rect 2605 10217 2639 10251
rect 5181 10217 5215 10251
rect 14105 10217 14139 10251
rect 15761 10217 15795 10251
rect 2329 10149 2363 10183
rect 9781 10149 9815 10183
rect 11897 10149 11931 10183
rect 1777 10081 1811 10115
rect 3157 10081 3191 10115
rect 4261 10081 4295 10115
rect 5825 10081 5859 10115
rect 6837 10081 6871 10115
rect 4445 10013 4479 10047
rect 6193 10013 6227 10047
rect 7104 10013 7138 10047
rect 8585 10013 8619 10047
rect 11161 10013 11195 10047
rect 11621 10009 11655 10043
rect 13277 10013 13311 10047
rect 14289 10013 14323 10047
rect 15025 10013 15059 10047
rect 1869 9945 1903 9979
rect 5641 9945 5675 9979
rect 10916 9945 10950 9979
rect 13032 9945 13066 9979
rect 14565 9945 14599 9979
rect 16129 9945 16163 9979
rect 1961 9877 1995 9911
rect 2973 9877 3007 9911
rect 3065 9877 3099 9911
rect 3801 9877 3835 9911
rect 4537 9877 4571 9911
rect 4905 9877 4939 9911
rect 5549 9877 5583 9911
rect 6377 9877 6411 9911
rect 8217 9877 8251 9911
rect 8953 9877 8987 9911
rect 9413 9877 9447 9911
rect 11437 9877 11471 9911
rect 13553 9877 13587 9911
rect 15393 9877 15427 9911
rect 3617 9673 3651 9707
rect 4721 9673 4755 9707
rect 8401 9673 8435 9707
rect 6009 9605 6043 9639
rect 7573 9605 7607 9639
rect 9873 9605 9907 9639
rect 10793 9605 10827 9639
rect 11796 9605 11830 9639
rect 13829 9605 13863 9639
rect 2625 9537 2659 9571
rect 2881 9537 2915 9571
rect 3525 9537 3559 9571
rect 4629 9537 4663 9571
rect 5365 9537 5399 9571
rect 8769 9537 8803 9571
rect 9781 9537 9815 9571
rect 11529 9537 11563 9571
rect 13185 9537 13219 9571
rect 14197 9537 14231 9571
rect 15117 9537 15151 9571
rect 15761 9537 15795 9571
rect 16037 9537 16071 9571
rect 3709 9469 3743 9503
rect 4813 9469 4847 9503
rect 6929 9469 6963 9503
rect 7665 9469 7699 9503
rect 7849 9469 7883 9503
rect 8861 9469 8895 9503
rect 8953 9469 8987 9503
rect 10057 9469 10091 9503
rect 10609 9469 10643 9503
rect 10701 9469 10735 9503
rect 14841 9469 14875 9503
rect 16681 9469 16715 9503
rect 1501 9401 1535 9435
rect 4261 9401 4295 9435
rect 9413 9401 9447 9435
rect 15301 9401 15335 9435
rect 3157 9333 3191 9367
rect 6377 9333 6411 9367
rect 7205 9333 7239 9367
rect 11161 9333 11195 9367
rect 12909 9333 12943 9367
rect 15577 9333 15611 9367
rect 1593 9129 1627 9163
rect 1961 9129 1995 9163
rect 9689 9129 9723 9163
rect 12909 9129 12943 9163
rect 6837 9061 6871 9095
rect 14105 9061 14139 9095
rect 17233 9061 17267 9095
rect 2513 8993 2547 9027
rect 4721 8993 4755 9027
rect 5641 8993 5675 9027
rect 6285 8993 6319 9027
rect 10241 8993 10275 9027
rect 12357 8993 12391 9027
rect 15485 8993 15519 9027
rect 1409 8925 1443 8959
rect 2329 8925 2363 8959
rect 3249 8925 3283 8959
rect 6469 8925 6503 8959
rect 8493 8925 8527 8959
rect 10701 8925 10735 8959
rect 11805 8925 11839 8959
rect 13645 8925 13679 8959
rect 15761 8925 15795 8959
rect 17049 8925 17083 8959
rect 5549 8857 5583 8891
rect 6377 8857 6411 8891
rect 8226 8857 8260 8891
rect 10149 8857 10183 8891
rect 11345 8857 11379 8891
rect 12541 8857 12575 8891
rect 13185 8857 13219 8891
rect 15240 8857 15274 8891
rect 16405 8857 16439 8891
rect 17509 8857 17543 8891
rect 2421 8789 2455 8823
rect 3433 8789 3467 8823
rect 4077 8789 4111 8823
rect 4445 8789 4479 8823
rect 4537 8789 4571 8823
rect 5089 8789 5123 8823
rect 5457 8789 5491 8823
rect 7113 8789 7147 8823
rect 9137 8789 9171 8823
rect 10057 8789 10091 8823
rect 11621 8789 11655 8823
rect 12449 8789 12483 8823
rect 16681 8789 16715 8823
rect 17969 8789 18003 8823
rect 2329 8585 2363 8619
rect 6377 8585 6411 8619
rect 8125 8585 8159 8619
rect 9045 8585 9079 8619
rect 9413 8585 9447 8619
rect 13001 8585 13035 8619
rect 15025 8585 15059 8619
rect 15945 8585 15979 8619
rect 1409 8517 1443 8551
rect 13912 8517 13946 8551
rect 2053 8449 2087 8483
rect 3453 8449 3487 8483
rect 4445 8449 4479 8483
rect 4701 8449 4735 8483
rect 7490 8449 7524 8483
rect 8769 8449 8803 8483
rect 10333 8449 10367 8483
rect 11897 8449 11931 8483
rect 15761 8449 15795 8483
rect 16681 8449 16715 8483
rect 17325 8449 17359 8483
rect 17601 8449 17635 8483
rect 3709 8381 3743 8415
rect 4169 8381 4203 8415
rect 7757 8381 7791 8415
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 11621 8381 11655 8415
rect 11805 8381 11839 8415
rect 12817 8381 12851 8415
rect 12909 8381 12943 8415
rect 13645 8381 13679 8415
rect 15301 8381 15335 8415
rect 16221 8381 16255 8415
rect 5825 8313 5859 8347
rect 10977 8313 11011 8347
rect 17141 8313 17175 8347
rect 17969 8313 18003 8347
rect 18337 8313 18371 8347
rect 18797 8313 18831 8347
rect 12265 8245 12299 8279
rect 13369 8245 13403 8279
rect 2421 8041 2455 8075
rect 3801 8041 3835 8075
rect 4997 8041 5031 8075
rect 5733 8041 5767 8075
rect 8033 8041 8067 8075
rect 8493 8041 8527 8075
rect 16405 8041 16439 8075
rect 1869 7905 1903 7939
rect 3249 7905 3283 7939
rect 4445 7905 4479 7939
rect 7481 7905 7515 7939
rect 10977 7905 11011 7939
rect 14473 7905 14507 7939
rect 15301 7905 15335 7939
rect 3985 7837 4019 7871
rect 7021 7837 7055 7871
rect 8309 7837 8343 7871
rect 8953 7837 8987 7871
rect 9220 7837 9254 7871
rect 12633 7837 12667 7871
rect 12909 7837 12943 7871
rect 14565 7837 14599 7871
rect 14657 7837 14691 7871
rect 15945 7837 15979 7871
rect 17785 7837 17819 7871
rect 18245 7837 18279 7871
rect 18521 7837 18555 7871
rect 1961 7769 1995 7803
rect 3065 7769 3099 7803
rect 4537 7769 4571 7803
rect 12388 7769 12422 7803
rect 17540 7769 17574 7803
rect 21005 7769 21039 7803
rect 2053 7701 2087 7735
rect 2697 7701 2731 7735
rect 3157 7701 3191 7735
rect 4629 7701 4663 7735
rect 7573 7701 7607 7735
rect 7665 7701 7699 7735
rect 10333 7701 10367 7735
rect 11253 7701 11287 7735
rect 13553 7701 13587 7735
rect 15025 7701 15059 7735
rect 18061 7701 18095 7735
rect 19257 7701 19291 7735
rect 21373 7701 21407 7735
rect 4261 7497 4295 7531
rect 5549 7497 5583 7531
rect 6377 7497 6411 7531
rect 6745 7497 6779 7531
rect 9873 7497 9907 7531
rect 10241 7497 10275 7531
rect 11529 7497 11563 7531
rect 16681 7497 16715 7531
rect 17785 7497 17819 7531
rect 18981 7497 19015 7531
rect 2022 7429 2056 7463
rect 4629 7429 4663 7463
rect 5641 7429 5675 7463
rect 12664 7429 12698 7463
rect 15402 7429 15436 7463
rect 4721 7361 4755 7395
rect 7573 7361 7607 7395
rect 8116 7361 8150 7395
rect 10517 7361 10551 7395
rect 13369 7361 13403 7395
rect 15945 7361 15979 7395
rect 17325 7361 17359 7395
rect 17601 7361 17635 7395
rect 18705 7361 18739 7395
rect 19165 7361 19199 7395
rect 19901 7361 19935 7395
rect 1777 7293 1811 7327
rect 3985 7293 4019 7327
rect 4813 7293 4847 7327
rect 5457 7293 5491 7327
rect 6837 7293 6871 7327
rect 6929 7293 6963 7327
rect 7849 7293 7883 7327
rect 9597 7293 9631 7327
rect 9781 7293 9815 7327
rect 12909 7293 12943 7327
rect 15669 7293 15703 7327
rect 18061 7293 18095 7327
rect 9229 7225 9263 7259
rect 14013 7225 14047 7259
rect 16129 7225 16163 7259
rect 18521 7225 18555 7259
rect 20177 7225 20211 7259
rect 1501 7157 1535 7191
rect 3157 7157 3191 7191
rect 3525 7157 3559 7191
rect 6009 7157 6043 7191
rect 7389 7157 7423 7191
rect 11161 7157 11195 7191
rect 14289 7157 14323 7191
rect 19717 7157 19751 7191
rect 20545 7157 20579 7191
rect 21005 7157 21039 7191
rect 21373 7157 21407 7191
rect 3801 6953 3835 6987
rect 5549 6953 5583 6987
rect 8953 6953 8987 6987
rect 18797 6953 18831 6987
rect 4813 6885 4847 6919
rect 8493 6885 8527 6919
rect 4353 6817 4387 6851
rect 7665 6817 7699 6851
rect 9505 6817 9539 6851
rect 10609 6817 10643 6851
rect 11069 6817 11103 6851
rect 12633 6817 12667 6851
rect 13093 6817 13127 6851
rect 18521 6817 18555 6851
rect 20637 6817 20671 6851
rect 1409 6749 1443 6783
rect 3249 6749 3283 6783
rect 4261 6749 4295 6783
rect 4997 6749 5031 6783
rect 7021 6749 7055 6783
rect 9965 6749 9999 6783
rect 11345 6749 11379 6783
rect 11989 6749 12023 6783
rect 13369 6749 13403 6783
rect 14105 6749 14139 6783
rect 14372 6749 14406 6783
rect 16221 6749 16255 6783
rect 17877 6749 17911 6783
rect 19441 6749 19475 6783
rect 19901 6749 19935 6783
rect 20177 6749 20211 6783
rect 1676 6681 1710 6715
rect 7757 6681 7791 6715
rect 16488 6681 16522 6715
rect 2789 6613 2823 6647
rect 3433 6613 3467 6647
rect 4169 6613 4203 6647
rect 7849 6613 7883 6647
rect 8217 6613 8251 6647
rect 9321 6613 9355 6647
rect 9413 6613 9447 6647
rect 11253 6613 11287 6647
rect 11713 6613 11747 6647
rect 13277 6613 13311 6647
rect 13737 6613 13771 6647
rect 15485 6613 15519 6647
rect 15761 6613 15795 6647
rect 17601 6613 17635 6647
rect 19257 6613 19291 6647
rect 19717 6613 19751 6647
rect 20361 6613 20395 6647
rect 21005 6613 21039 6647
rect 1685 6409 1719 6443
rect 2329 6409 2363 6443
rect 9781 6409 9815 6443
rect 11069 6409 11103 6443
rect 12265 6409 12299 6443
rect 14473 6409 14507 6443
rect 14565 6409 14599 6443
rect 15945 6409 15979 6443
rect 16681 6409 16715 6443
rect 17049 6409 17083 6443
rect 17141 6409 17175 6443
rect 17877 6409 17911 6443
rect 18153 6409 18187 6443
rect 19073 6409 19107 6443
rect 19993 6409 20027 6443
rect 2237 6341 2271 6375
rect 1501 6273 1535 6307
rect 4086 6273 4120 6307
rect 4353 6273 4387 6307
rect 5753 6273 5787 6307
rect 7001 6273 7035 6307
rect 8657 6273 8691 6307
rect 10701 6273 10735 6307
rect 13389 6273 13423 6307
rect 17693 6273 17727 6307
rect 18337 6273 18371 6307
rect 18613 6273 18647 6307
rect 19257 6273 19291 6307
rect 19717 6273 19751 6307
rect 20177 6273 20211 6307
rect 20913 6273 20947 6307
rect 21373 6273 21407 6307
rect 2145 6205 2179 6239
rect 6009 6205 6043 6239
rect 6745 6205 6779 6239
rect 8401 6205 8435 6239
rect 10425 6205 10459 6239
rect 10609 6205 10643 6239
rect 11989 6205 12023 6239
rect 13645 6205 13679 6239
rect 14381 6205 14415 6239
rect 15761 6205 15795 6239
rect 15853 6205 15887 6239
rect 17233 6205 17267 6239
rect 2973 6137 3007 6171
rect 4629 6137 4663 6171
rect 15209 6137 15243 6171
rect 2697 6069 2731 6103
rect 6377 6069 6411 6103
rect 8125 6069 8159 6103
rect 14933 6069 14967 6103
rect 16313 6069 16347 6103
rect 18797 6069 18831 6103
rect 19533 6069 19567 6103
rect 20729 6069 20763 6103
rect 21189 6069 21223 6103
rect 2421 5865 2455 5899
rect 3801 5865 3835 5899
rect 5733 5865 5767 5899
rect 9137 5865 9171 5899
rect 13369 5865 13403 5899
rect 14749 5865 14783 5899
rect 15209 5865 15243 5899
rect 16129 5865 16163 5899
rect 16681 5865 16715 5899
rect 20177 5865 20211 5899
rect 21097 5865 21131 5899
rect 19257 5797 19291 5831
rect 1869 5729 1903 5763
rect 2789 5729 2823 5763
rect 2973 5729 3007 5763
rect 4353 5729 4387 5763
rect 7849 5729 7883 5763
rect 8033 5729 8067 5763
rect 9597 5729 9631 5763
rect 18061 5729 18095 5763
rect 2053 5661 2087 5695
rect 4813 5661 4847 5695
rect 7021 5661 7055 5695
rect 7481 5661 7515 5695
rect 8953 5661 8987 5695
rect 12449 5661 12483 5695
rect 13553 5661 13587 5695
rect 14105 5661 14139 5695
rect 15025 5661 15059 5695
rect 15485 5661 15519 5695
rect 18521 5661 18555 5695
rect 19441 5661 19475 5695
rect 19717 5661 19751 5695
rect 20361 5661 20395 5695
rect 20821 5661 20855 5695
rect 21281 5661 21315 5695
rect 1961 5593 1995 5627
rect 4261 5593 4295 5627
rect 10425 5593 10459 5627
rect 12173 5593 12207 5627
rect 17816 5593 17850 5627
rect 3065 5525 3099 5559
rect 3433 5525 3467 5559
rect 4169 5525 4203 5559
rect 4997 5525 5031 5559
rect 7297 5525 7331 5559
rect 8125 5525 8159 5559
rect 8493 5525 8527 5559
rect 9689 5525 9723 5559
rect 9781 5525 9815 5559
rect 10149 5525 10183 5559
rect 13093 5525 13127 5559
rect 18337 5525 18371 5559
rect 18797 5525 18831 5559
rect 19901 5525 19935 5559
rect 20637 5525 20671 5559
rect 2881 5321 2915 5355
rect 3893 5321 3927 5355
rect 4261 5321 4295 5355
rect 5365 5321 5399 5355
rect 8033 5321 8067 5355
rect 8401 5321 8435 5355
rect 9229 5321 9263 5355
rect 9505 5321 9539 5355
rect 16681 5321 16715 5355
rect 17693 5321 17727 5355
rect 18613 5321 18647 5355
rect 20453 5321 20487 5355
rect 3249 5253 3283 5287
rect 7512 5253 7546 5287
rect 10640 5253 10674 5287
rect 13001 5253 13035 5287
rect 14749 5253 14783 5287
rect 1961 5185 1995 5219
rect 4353 5185 4387 5219
rect 5457 5185 5491 5219
rect 7757 5185 7791 5219
rect 8493 5185 8527 5219
rect 9045 5185 9079 5219
rect 10885 5185 10919 5219
rect 11529 5185 11563 5219
rect 12357 5185 12391 5219
rect 15025 5185 15059 5219
rect 15853 5185 15887 5219
rect 17049 5185 17083 5219
rect 17877 5185 17911 5219
rect 18153 5185 18187 5219
rect 18797 5185 18831 5219
rect 19257 5185 19291 5219
rect 20177 5185 20211 5219
rect 20637 5185 20671 5219
rect 21097 5185 21131 5219
rect 2237 5117 2271 5151
rect 3341 5117 3375 5151
rect 3433 5117 3467 5151
rect 4445 5117 4479 5151
rect 5273 5117 5307 5151
rect 8585 5117 8619 5151
rect 12173 5117 12207 5151
rect 12265 5117 12299 5151
rect 15577 5117 15611 5151
rect 15761 5117 15795 5151
rect 17141 5117 17175 5151
rect 17233 5117 17267 5151
rect 19533 5117 19567 5151
rect 5825 5049 5859 5083
rect 6377 5049 6411 5083
rect 12725 5049 12759 5083
rect 16221 5049 16255 5083
rect 18337 5049 18371 5083
rect 19993 5049 20027 5083
rect 2513 4981 2547 5015
rect 11713 4981 11747 5015
rect 15209 4981 15243 5015
rect 19073 4981 19107 5015
rect 20913 4981 20947 5015
rect 3341 4777 3375 4811
rect 7757 4777 7791 4811
rect 10149 4777 10183 4811
rect 11897 4777 11931 4811
rect 1685 4709 1719 4743
rect 7481 4709 7515 4743
rect 13645 4709 13679 4743
rect 1961 4641 1995 4675
rect 5181 4641 5215 4675
rect 6101 4641 6135 4675
rect 8401 4641 8435 4675
rect 9137 4641 9171 4675
rect 9597 4641 9631 4675
rect 18061 4641 18095 4675
rect 19257 4641 19291 4675
rect 8125 4573 8159 4607
rect 9781 4573 9815 4607
rect 10517 4573 10551 4607
rect 12265 4573 12299 4607
rect 12532 4573 12566 4607
rect 14105 4573 14139 4607
rect 16405 4573 16439 4607
rect 18521 4573 18555 4607
rect 21106 4573 21140 4607
rect 21373 4573 21407 4607
rect 1501 4505 1535 4539
rect 2206 4505 2240 4539
rect 4936 4505 4970 4539
rect 6368 4505 6402 4539
rect 9689 4505 9723 4539
rect 10784 4505 10818 4539
rect 16160 4505 16194 4539
rect 17794 4505 17828 4539
rect 18797 4505 18831 4539
rect 3801 4437 3835 4471
rect 5825 4437 5859 4471
rect 8217 4437 8251 4471
rect 14749 4437 14783 4471
rect 15025 4437 15059 4471
rect 16681 4437 16715 4471
rect 18337 4437 18371 4471
rect 19993 4437 20027 4471
rect 4629 4233 4663 4267
rect 5641 4233 5675 4267
rect 6009 4233 6043 4267
rect 7021 4233 7055 4267
rect 7941 4233 7975 4267
rect 9137 4233 9171 4267
rect 10517 4233 10551 4267
rect 11805 4233 11839 4267
rect 14105 4233 14139 4267
rect 17049 4233 17083 4267
rect 10149 4165 10183 4199
rect 11897 4165 11931 4199
rect 14648 4165 14682 4199
rect 17785 4165 17819 4199
rect 3341 4097 3375 4131
rect 3801 4097 3835 4131
rect 4721 4097 4755 4131
rect 6929 4097 6963 4131
rect 8033 4097 8067 4131
rect 11161 4097 11195 4131
rect 12725 4097 12759 4131
rect 12992 4097 13026 4131
rect 14381 4097 14415 4131
rect 16221 4097 16255 4131
rect 18061 4097 18095 4131
rect 18705 4097 18739 4131
rect 19165 4097 19199 4131
rect 19625 4097 19659 4131
rect 20085 4097 20119 4131
rect 20729 4097 20763 4131
rect 21005 4097 21039 4131
rect 1961 4029 1995 4063
rect 2237 4029 2271 4063
rect 3065 4029 3099 4063
rect 4813 4029 4847 4063
rect 5365 4029 5399 4063
rect 5549 4029 5583 4063
rect 6745 4029 6779 4063
rect 7757 4029 7791 4063
rect 9229 4029 9263 4063
rect 9413 4029 9447 4063
rect 9873 4029 9907 4063
rect 10057 4029 10091 4063
rect 11713 4029 11747 4063
rect 16865 4029 16899 4063
rect 16957 4029 16991 4063
rect 3985 3961 4019 3995
rect 4261 3961 4295 3995
rect 7389 3961 7423 3995
rect 10977 3961 11011 3995
rect 19441 3961 19475 3995
rect 19901 3961 19935 3995
rect 20545 3961 20579 3995
rect 8401 3893 8435 3927
rect 8769 3893 8803 3927
rect 12265 3893 12299 3927
rect 15761 3893 15795 3927
rect 16037 3893 16071 3927
rect 17417 3893 17451 3927
rect 18981 3893 19015 3927
rect 21189 3893 21223 3927
rect 4399 3689 4433 3723
rect 6837 3689 6871 3723
rect 10885 3689 10919 3723
rect 16773 3689 16807 3723
rect 3341 3621 3375 3655
rect 6561 3621 6595 3655
rect 8953 3621 8987 3655
rect 10149 3621 10183 3655
rect 19809 3621 19843 3655
rect 2789 3553 2823 3587
rect 5181 3553 5215 3587
rect 7389 3553 7423 3587
rect 8033 3553 8067 3587
rect 8125 3553 8159 3587
rect 9505 3553 9539 3587
rect 12817 3553 12851 3587
rect 14289 3553 14323 3587
rect 15301 3553 15335 3587
rect 4629 3485 4663 3519
rect 8217 3485 8251 3519
rect 9321 3485 9355 3519
rect 9965 3485 9999 3519
rect 12173 3485 12207 3519
rect 12909 3485 12943 3519
rect 13001 3485 13035 3519
rect 16129 3485 16163 3519
rect 17049 3485 17083 3519
rect 17693 3485 17727 3519
rect 18613 3485 18647 3519
rect 19625 3485 19659 3519
rect 20177 3485 20211 3519
rect 20729 3485 20763 3519
rect 2544 3417 2578 3451
rect 3157 3417 3191 3451
rect 5426 3417 5460 3451
rect 7297 3417 7331 3451
rect 9413 3417 9447 3451
rect 13645 3417 13679 3451
rect 14473 3417 14507 3451
rect 17969 3417 18003 3451
rect 21281 3417 21315 3451
rect 1409 3349 1443 3383
rect 7205 3349 7239 3383
rect 8585 3349 8619 3383
rect 13369 3349 13403 3383
rect 14381 3349 14415 3383
rect 14841 3349 14875 3383
rect 15393 3349 15427 3383
rect 15485 3349 15519 3383
rect 15853 3349 15887 3383
rect 18429 3349 18463 3383
rect 19257 3349 19291 3383
rect 20361 3349 20395 3383
rect 20913 3349 20947 3383
rect 2697 3145 2731 3179
rect 2973 3145 3007 3179
rect 4629 3145 4663 3179
rect 6377 3145 6411 3179
rect 8953 3145 8987 3179
rect 13645 3145 13679 3179
rect 14565 3145 14599 3179
rect 15485 3145 15519 3179
rect 17325 3145 17359 3179
rect 18429 3145 18463 3179
rect 8432 3077 8466 3111
rect 10609 3077 10643 3111
rect 1961 3009 1995 3043
rect 2513 3009 2547 3043
rect 4097 3009 4131 3043
rect 4353 3009 4387 3043
rect 5742 3009 5776 3043
rect 6009 3009 6043 3043
rect 7021 3009 7055 3043
rect 8677 3009 8711 3043
rect 10066 3009 10100 3043
rect 10333 3009 10367 3043
rect 10977 3009 11011 3043
rect 11989 3009 12023 3043
rect 12532 3009 12566 3043
rect 13921 3009 13955 3043
rect 14841 3009 14875 3043
rect 16037 3009 16071 3043
rect 16957 3009 16991 3043
rect 17509 3009 17543 3043
rect 18061 3009 18095 3043
rect 18613 3009 18647 3043
rect 19165 3009 19199 3043
rect 19717 3009 19751 3043
rect 21373 3009 21407 3043
rect 2237 2941 2271 2975
rect 12265 2941 12299 2975
rect 20729 2941 20763 2975
rect 15853 2873 15887 2907
rect 17877 2873 17911 2907
rect 7297 2805 7331 2839
rect 11161 2805 11195 2839
rect 11805 2805 11839 2839
rect 16773 2805 16807 2839
rect 18981 2805 19015 2839
rect 19901 2805 19935 2839
rect 7389 2601 7423 2635
rect 7849 2601 7883 2635
rect 10149 2601 10183 2635
rect 10425 2601 10459 2635
rect 11529 2601 11563 2635
rect 15761 2601 15795 2635
rect 19349 2601 19383 2635
rect 13553 2533 13587 2567
rect 16865 2533 16899 2567
rect 17325 2533 17359 2567
rect 17877 2533 17911 2567
rect 19901 2533 19935 2567
rect 1961 2465 1995 2499
rect 2237 2465 2271 2499
rect 3341 2465 3375 2499
rect 4353 2465 4387 2499
rect 5457 2465 5491 2499
rect 6837 2465 6871 2499
rect 8493 2465 8527 2499
rect 9597 2465 9631 2499
rect 10977 2465 11011 2499
rect 12081 2465 12115 2499
rect 21097 2465 21131 2499
rect 21373 2465 21407 2499
rect 3065 2397 3099 2431
rect 4629 2397 4663 2431
rect 5733 2397 5767 2431
rect 6929 2397 6963 2431
rect 8217 2397 8251 2431
rect 8953 2397 8987 2431
rect 9689 2397 9723 2431
rect 11989 2397 12023 2431
rect 12541 2397 12575 2431
rect 13737 2397 13771 2431
rect 14105 2397 14139 2431
rect 15301 2397 15335 2431
rect 15577 2397 15611 2431
rect 16129 2397 16163 2431
rect 16681 2397 16715 2431
rect 17509 2397 17543 2431
rect 18061 2397 18095 2431
rect 18613 2397 18647 2431
rect 19533 2397 19567 2431
rect 20085 2397 20119 2431
rect 7021 2261 7055 2295
rect 8309 2261 8343 2295
rect 9137 2261 9171 2295
rect 9781 2261 9815 2295
rect 10793 2261 10827 2295
rect 10885 2261 10919 2295
rect 11897 2261 11931 2295
rect 13185 2261 13219 2295
rect 14749 2261 14783 2295
rect 15117 2261 15151 2295
rect 16313 2261 16347 2295
rect 18429 2261 18463 2295
<< metal1 >>
rect 1486 20748 1492 20800
rect 1544 20788 1550 20800
rect 4706 20788 4712 20800
rect 1544 20760 4712 20788
rect 1544 20748 1550 20760
rect 4706 20748 4712 20760
rect 4764 20748 4770 20800
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 2593 20587 2651 20593
rect 2593 20553 2605 20587
rect 2639 20584 2651 20587
rect 2774 20584 2780 20596
rect 2639 20556 2780 20584
rect 2639 20553 2651 20556
rect 2593 20547 2651 20553
rect 2774 20544 2780 20556
rect 2832 20544 2838 20596
rect 3142 20584 3148 20596
rect 3103 20556 3148 20584
rect 3142 20544 3148 20556
rect 3200 20544 3206 20596
rect 4706 20584 4712 20596
rect 4667 20556 4712 20584
rect 4706 20544 4712 20556
rect 4764 20544 4770 20596
rect 1486 20516 1492 20528
rect 1447 20488 1492 20516
rect 1486 20476 1492 20488
rect 1544 20476 1550 20528
rect 8202 20516 8208 20528
rect 3344 20488 8208 20516
rect 2222 20448 2228 20460
rect 2183 20420 2228 20448
rect 2222 20408 2228 20420
rect 2280 20408 2286 20460
rect 3344 20457 3372 20488
rect 8202 20476 8208 20488
rect 8260 20476 8266 20528
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20417 2835 20451
rect 2777 20411 2835 20417
rect 3329 20451 3387 20457
rect 3329 20417 3341 20451
rect 3375 20417 3387 20451
rect 3970 20448 3976 20460
rect 3931 20420 3976 20448
rect 3329 20411 3387 20417
rect 2792 20380 2820 20411
rect 3970 20408 3976 20420
rect 4028 20408 4034 20460
rect 4249 20451 4307 20457
rect 4249 20417 4261 20451
rect 4295 20448 4307 20451
rect 8662 20448 8668 20460
rect 4295 20420 8668 20448
rect 4295 20417 4307 20420
rect 4249 20411 4307 20417
rect 8662 20408 8668 20420
rect 8720 20408 8726 20460
rect 4154 20380 4160 20392
rect 2792 20352 4160 20380
rect 4154 20340 4160 20352
rect 4212 20340 4218 20392
rect 1673 20315 1731 20321
rect 1673 20281 1685 20315
rect 1719 20312 1731 20315
rect 1854 20312 1860 20324
rect 1719 20284 1860 20312
rect 1719 20281 1731 20284
rect 1673 20275 1731 20281
rect 1854 20272 1860 20284
rect 1912 20272 1918 20324
rect 2038 20312 2044 20324
rect 1999 20284 2044 20312
rect 2038 20272 2044 20284
rect 2096 20272 2102 20324
rect 2314 20272 2320 20324
rect 2372 20312 2378 20324
rect 3789 20315 3847 20321
rect 3789 20312 3801 20315
rect 2372 20284 3801 20312
rect 2372 20272 2378 20284
rect 3789 20281 3801 20284
rect 3835 20281 3847 20315
rect 3789 20275 3847 20281
rect 4430 20244 4436 20256
rect 4391 20216 4436 20244
rect 4430 20204 4436 20216
rect 4488 20204 4494 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2590 20040 2596 20052
rect 2551 20012 2596 20040
rect 2590 20000 2596 20012
rect 2648 20000 2654 20052
rect 3237 20043 3295 20049
rect 3237 20009 3249 20043
rect 3283 20040 3295 20043
rect 3970 20040 3976 20052
rect 3283 20012 3976 20040
rect 3283 20009 3295 20012
rect 3237 20003 3295 20009
rect 3970 20000 3976 20012
rect 4028 20000 4034 20052
rect 4154 20000 4160 20052
rect 4212 20040 4218 20052
rect 4249 20043 4307 20049
rect 4249 20040 4261 20043
rect 4212 20012 4261 20040
rect 4212 20000 4218 20012
rect 4249 20009 4261 20012
rect 4295 20009 4307 20043
rect 4249 20003 4307 20009
rect 2222 19932 2228 19984
rect 2280 19972 2286 19984
rect 3789 19975 3847 19981
rect 3789 19972 3801 19975
rect 2280 19944 3801 19972
rect 2280 19932 2286 19944
rect 3789 19941 3801 19944
rect 3835 19941 3847 19975
rect 3789 19935 3847 19941
rect 2958 19904 2964 19916
rect 1688 19876 2964 19904
rect 1688 19845 1716 19876
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 6546 19904 6552 19916
rect 3068 19876 6552 19904
rect 3068 19845 3096 19876
rect 6546 19864 6552 19876
rect 6604 19864 6610 19916
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 1673 19799 1731 19805
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19805 2283 19839
rect 2225 19799 2283 19805
rect 2777 19839 2835 19845
rect 2777 19805 2789 19839
rect 2823 19805 2835 19839
rect 2777 19799 2835 19805
rect 3053 19839 3111 19845
rect 3053 19805 3065 19839
rect 3099 19805 3111 19839
rect 3053 19799 3111 19805
rect 2240 19768 2268 19799
rect 2792 19768 2820 19799
rect 3602 19796 3608 19848
rect 3660 19836 3666 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3660 19808 3985 19836
rect 3660 19796 3666 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 4430 19836 4436 19848
rect 4391 19808 4436 19836
rect 3973 19799 4031 19805
rect 4430 19796 4436 19808
rect 4488 19796 4494 19848
rect 4522 19796 4528 19848
rect 4580 19836 4586 19848
rect 4893 19839 4951 19845
rect 4893 19836 4905 19839
rect 4580 19808 4905 19836
rect 4580 19796 4586 19808
rect 4893 19805 4905 19808
rect 4939 19805 4951 19839
rect 4893 19799 4951 19805
rect 2240 19740 2728 19768
rect 2792 19740 4752 19768
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 2038 19700 2044 19712
rect 1999 19672 2044 19700
rect 2038 19660 2044 19672
rect 2096 19660 2102 19712
rect 2700 19700 2728 19740
rect 3878 19700 3884 19712
rect 2700 19672 3884 19700
rect 3878 19660 3884 19672
rect 3936 19660 3942 19712
rect 4724 19709 4752 19740
rect 4709 19703 4767 19709
rect 4709 19669 4721 19703
rect 4755 19669 4767 19703
rect 4709 19663 4767 19669
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19456 1952 19508
rect 2004 19496 2010 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 2004 19468 2053 19496
rect 2004 19456 2010 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2041 19459 2099 19465
rect 2777 19499 2835 19505
rect 2777 19465 2789 19499
rect 2823 19465 2835 19499
rect 3602 19496 3608 19508
rect 3563 19468 3608 19496
rect 2777 19459 2835 19465
rect 2792 19428 2820 19459
rect 3602 19456 3608 19468
rect 3660 19456 3666 19508
rect 3878 19496 3884 19508
rect 3839 19468 3884 19496
rect 3878 19456 3884 19468
rect 3936 19456 3942 19508
rect 4522 19496 4528 19508
rect 4483 19468 4528 19496
rect 4522 19456 4528 19468
rect 4580 19456 4586 19508
rect 5902 19428 5908 19440
rect 2792 19400 4108 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19329 1731 19363
rect 1673 19323 1731 19329
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19360 2283 19363
rect 2314 19360 2320 19372
rect 2271 19332 2320 19360
rect 2271 19329 2283 19332
rect 2225 19323 2283 19329
rect 1688 19292 1716 19323
rect 2314 19320 2320 19332
rect 2372 19320 2378 19372
rect 2593 19363 2651 19369
rect 2593 19329 2605 19363
rect 2639 19360 2651 19363
rect 2682 19360 2688 19372
rect 2639 19332 2688 19360
rect 2639 19329 2651 19332
rect 2593 19323 2651 19329
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 4080 19369 4108 19400
rect 4172 19400 5908 19428
rect 3421 19363 3479 19369
rect 3421 19329 3433 19363
rect 3467 19360 3479 19363
rect 4065 19363 4123 19369
rect 3467 19332 4016 19360
rect 3467 19329 3479 19332
rect 3421 19323 3479 19329
rect 3326 19292 3332 19304
rect 1688 19264 3332 19292
rect 3326 19252 3332 19264
rect 3384 19252 3390 19304
rect 3988 19292 4016 19332
rect 4065 19329 4077 19363
rect 4111 19329 4123 19363
rect 4065 19323 4123 19329
rect 4172 19292 4200 19400
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 4341 19363 4399 19369
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 9674 19360 9680 19372
rect 4387 19332 9680 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 9674 19320 9680 19332
rect 9732 19320 9738 19372
rect 3988 19264 4200 19292
rect 2682 19184 2688 19236
rect 2740 19224 2746 19236
rect 8478 19224 8484 19236
rect 2740 19196 8484 19224
rect 2740 19184 2746 19196
rect 8478 19184 8484 19196
rect 8536 19184 8542 19236
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 2038 19116 2044 19168
rect 2096 19156 2102 19168
rect 5994 19156 6000 19168
rect 2096 19128 6000 19156
rect 2096 19116 2102 19128
rect 5994 19116 6000 19128
rect 6052 19116 6058 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 4249 18955 4307 18961
rect 4249 18952 4261 18955
rect 2746 18924 4261 18952
rect 2746 18816 2774 18924
rect 4249 18921 4261 18924
rect 4295 18921 4307 18955
rect 4249 18915 4307 18921
rect 8202 18912 8208 18964
rect 8260 18952 8266 18964
rect 10505 18955 10563 18961
rect 10505 18952 10517 18955
rect 8260 18924 10517 18952
rect 8260 18912 8266 18924
rect 10505 18921 10517 18924
rect 10551 18921 10563 18955
rect 10505 18915 10563 18921
rect 5626 18884 5632 18896
rect 1688 18788 2774 18816
rect 2884 18856 5632 18884
rect 1688 18757 1716 18788
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18717 1731 18751
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 1673 18711 1731 18717
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2884 18757 2912 18856
rect 5626 18844 5632 18856
rect 5684 18844 5690 18896
rect 3142 18776 3148 18828
rect 3200 18816 3206 18828
rect 3200 18788 4476 18816
rect 3200 18776 3206 18788
rect 4448 18757 4476 18788
rect 2409 18751 2467 18757
rect 2409 18748 2421 18751
rect 2280 18720 2421 18748
rect 2280 18708 2286 18720
rect 2409 18717 2421 18720
rect 2455 18717 2467 18751
rect 2409 18711 2467 18717
rect 2869 18751 2927 18757
rect 2869 18717 2881 18751
rect 2915 18717 2927 18751
rect 3973 18751 4031 18757
rect 3973 18748 3985 18751
rect 2869 18711 2927 18717
rect 3068 18720 3985 18748
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1670 18572 1676 18624
rect 1728 18612 1734 18624
rect 1949 18615 2007 18621
rect 1949 18612 1961 18615
rect 1728 18584 1961 18612
rect 1728 18572 1734 18584
rect 1949 18581 1961 18584
rect 1995 18581 2007 18615
rect 2590 18612 2596 18624
rect 2551 18584 2596 18612
rect 1949 18575 2007 18581
rect 2590 18572 2596 18584
rect 2648 18572 2654 18624
rect 3068 18621 3096 18720
rect 3973 18717 3985 18720
rect 4019 18717 4031 18751
rect 3973 18711 4031 18717
rect 4433 18751 4491 18757
rect 4433 18717 4445 18751
rect 4479 18717 4491 18751
rect 4433 18711 4491 18717
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18717 4951 18751
rect 10686 18748 10692 18760
rect 10647 18720 10692 18748
rect 4893 18711 4951 18717
rect 3142 18640 3148 18692
rect 3200 18680 3206 18692
rect 4908 18680 4936 18711
rect 10686 18708 10692 18720
rect 10744 18708 10750 18760
rect 3200 18652 4936 18680
rect 3200 18640 3206 18652
rect 3053 18615 3111 18621
rect 3053 18581 3065 18615
rect 3099 18581 3111 18615
rect 3053 18575 3111 18581
rect 3234 18572 3240 18624
rect 3292 18612 3298 18624
rect 3789 18615 3847 18621
rect 3789 18612 3801 18615
rect 3292 18584 3801 18612
rect 3292 18572 3298 18584
rect 3789 18581 3801 18584
rect 3835 18581 3847 18615
rect 4706 18612 4712 18624
rect 4667 18584 4712 18612
rect 3789 18575 3847 18581
rect 4706 18572 4712 18584
rect 4764 18572 4770 18624
rect 5810 18612 5816 18624
rect 5771 18584 5816 18612
rect 5810 18572 5816 18584
rect 5868 18572 5874 18624
rect 6914 18612 6920 18624
rect 6875 18584 6920 18612
rect 6914 18572 6920 18584
rect 6972 18572 6978 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 2130 18368 2136 18420
rect 2188 18408 2194 18420
rect 2501 18411 2559 18417
rect 2501 18408 2513 18411
rect 2188 18380 2513 18408
rect 2188 18368 2194 18380
rect 2501 18377 2513 18380
rect 2547 18377 2559 18411
rect 2501 18371 2559 18377
rect 2590 18368 2596 18420
rect 2648 18408 2654 18420
rect 9674 18408 9680 18420
rect 2648 18380 3648 18408
rect 9635 18380 9680 18408
rect 2648 18368 2654 18380
rect 3234 18340 3240 18352
rect 2884 18312 3240 18340
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 1673 18235 1731 18241
rect 1688 18136 1716 18235
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2685 18275 2743 18281
rect 2685 18241 2697 18275
rect 2731 18272 2743 18275
rect 2884 18272 2912 18312
rect 3234 18300 3240 18312
rect 3292 18300 3298 18352
rect 3620 18281 3648 18380
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 10686 18368 10692 18420
rect 10744 18408 10750 18420
rect 11517 18411 11575 18417
rect 11517 18408 11529 18411
rect 10744 18380 11529 18408
rect 10744 18368 10750 18380
rect 11517 18377 11529 18380
rect 11563 18377 11575 18411
rect 11517 18371 11575 18377
rect 2731 18244 2912 18272
rect 2961 18275 3019 18281
rect 2731 18241 2743 18244
rect 2685 18235 2743 18241
rect 2961 18241 2973 18275
rect 3007 18241 3019 18275
rect 2961 18235 3019 18241
rect 3605 18275 3663 18281
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3878 18272 3884 18284
rect 3839 18244 3884 18272
rect 3605 18235 3663 18241
rect 2976 18204 3004 18235
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 4522 18232 4528 18284
rect 4580 18272 4586 18284
rect 4801 18275 4859 18281
rect 4801 18272 4813 18275
rect 4580 18244 4813 18272
rect 4580 18232 4586 18244
rect 4801 18241 4813 18244
rect 4847 18241 4859 18275
rect 4801 18235 4859 18241
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 5997 18275 6055 18281
rect 5997 18272 6009 18275
rect 5776 18244 6009 18272
rect 5776 18232 5782 18244
rect 5997 18241 6009 18244
rect 6043 18241 6055 18275
rect 6730 18272 6736 18284
rect 6691 18244 6736 18272
rect 5997 18235 6055 18241
rect 6730 18232 6736 18244
rect 6788 18232 6794 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 6932 18244 7389 18272
rect 6822 18204 6828 18216
rect 2976 18176 6408 18204
rect 6783 18176 6828 18204
rect 4706 18136 4712 18148
rect 1688 18108 4712 18136
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 6380 18145 6408 18176
rect 6822 18164 6828 18176
rect 6880 18164 6886 18216
rect 6932 18213 6960 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 10045 18275 10103 18281
rect 10045 18241 10057 18275
rect 10091 18272 10103 18275
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10091 18244 10977 18272
rect 10091 18241 10103 18244
rect 10045 18235 10103 18241
rect 10965 18241 10977 18244
rect 11011 18241 11023 18275
rect 11698 18272 11704 18284
rect 11659 18244 11704 18272
rect 10965 18235 11023 18241
rect 11698 18232 11704 18244
rect 11756 18232 11762 18284
rect 6917 18207 6975 18213
rect 6917 18173 6929 18207
rect 6963 18173 6975 18207
rect 6917 18167 6975 18173
rect 6365 18139 6423 18145
rect 6365 18105 6377 18139
rect 6411 18105 6423 18139
rect 6365 18099 6423 18105
rect 6638 18096 6644 18148
rect 6696 18136 6702 18148
rect 6932 18136 6960 18167
rect 8202 18164 8208 18216
rect 8260 18204 8266 18216
rect 8389 18207 8447 18213
rect 8389 18204 8401 18207
rect 8260 18176 8401 18204
rect 8260 18164 8266 18176
rect 8389 18173 8401 18176
rect 8435 18173 8447 18207
rect 10134 18204 10140 18216
rect 10095 18176 10140 18204
rect 8389 18167 8447 18173
rect 10134 18164 10140 18176
rect 10192 18164 10198 18216
rect 10321 18207 10379 18213
rect 10321 18173 10333 18207
rect 10367 18204 10379 18207
rect 11054 18204 11060 18216
rect 10367 18176 11060 18204
rect 10367 18173 10379 18176
rect 10321 18167 10379 18173
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 6696 18108 6960 18136
rect 6696 18096 6702 18108
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2225 18071 2283 18077
rect 2225 18037 2237 18071
rect 2271 18068 2283 18071
rect 2958 18068 2964 18080
rect 2271 18040 2964 18068
rect 2271 18037 2283 18040
rect 2225 18031 2283 18037
rect 2958 18028 2964 18040
rect 3016 18028 3022 18080
rect 3142 18068 3148 18080
rect 3103 18040 3148 18068
rect 3142 18028 3148 18040
rect 3200 18028 3206 18080
rect 3326 18028 3332 18080
rect 3384 18068 3390 18080
rect 3421 18071 3479 18077
rect 3421 18068 3433 18071
rect 3384 18040 3433 18068
rect 3384 18028 3390 18040
rect 3421 18037 3433 18040
rect 3467 18037 3479 18071
rect 3421 18031 3479 18037
rect 4525 18071 4583 18077
rect 4525 18037 4537 18071
rect 4571 18068 4583 18071
rect 4614 18068 4620 18080
rect 4571 18040 4620 18068
rect 4571 18037 4583 18040
rect 4525 18031 4583 18037
rect 4614 18028 4620 18040
rect 4672 18028 4678 18080
rect 5350 18068 5356 18080
rect 5311 18040 5356 18068
rect 5350 18028 5356 18040
rect 5408 18028 5414 18080
rect 7006 18028 7012 18080
rect 7064 18068 7070 18080
rect 8021 18071 8079 18077
rect 8021 18068 8033 18071
rect 7064 18040 8033 18068
rect 7064 18028 7070 18040
rect 8021 18037 8033 18040
rect 8067 18037 8079 18071
rect 8021 18031 8079 18037
rect 9401 18071 9459 18077
rect 9401 18037 9413 18071
rect 9447 18068 9459 18071
rect 9490 18068 9496 18080
rect 9447 18040 9496 18068
rect 9447 18037 9459 18040
rect 9401 18031 9459 18037
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 6733 17867 6791 17873
rect 6733 17833 6745 17867
rect 6779 17864 6791 17867
rect 6822 17864 6828 17876
rect 6779 17836 6828 17864
rect 6779 17833 6791 17836
rect 6733 17827 6791 17833
rect 6822 17824 6828 17836
rect 6880 17824 6886 17876
rect 9953 17867 10011 17873
rect 9953 17833 9965 17867
rect 9999 17864 10011 17867
rect 10134 17864 10140 17876
rect 9999 17836 10140 17864
rect 9999 17833 10011 17836
rect 9953 17827 10011 17833
rect 10134 17824 10140 17836
rect 10192 17824 10198 17876
rect 2593 17799 2651 17805
rect 2593 17765 2605 17799
rect 2639 17796 2651 17799
rect 3142 17796 3148 17808
rect 2639 17768 3148 17796
rect 2639 17765 2651 17768
rect 2593 17759 2651 17765
rect 3142 17756 3148 17768
rect 3200 17756 3206 17808
rect 6914 17756 6920 17808
rect 6972 17756 6978 17808
rect 15746 17796 15752 17808
rect 7576 17768 15752 17796
rect 5718 17688 5724 17740
rect 5776 17728 5782 17740
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 5776 17700 6101 17728
rect 5776 17688 5782 17700
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 6273 17731 6331 17737
rect 6273 17697 6285 17731
rect 6319 17728 6331 17731
rect 6932 17728 6960 17756
rect 7576 17728 7604 17768
rect 15746 17756 15752 17768
rect 15804 17756 15810 17808
rect 9398 17728 9404 17740
rect 6319 17700 7604 17728
rect 9048 17700 9404 17728
rect 6319 17697 6331 17700
rect 6273 17691 6331 17697
rect 1670 17660 1676 17672
rect 1631 17632 1676 17660
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 2133 17663 2191 17669
rect 2133 17629 2145 17663
rect 2179 17629 2191 17663
rect 2406 17660 2412 17672
rect 2367 17632 2412 17660
rect 2133 17623 2191 17629
rect 2148 17592 2176 17623
rect 2406 17620 2412 17632
rect 2464 17620 2470 17672
rect 2774 17620 2780 17672
rect 2832 17660 2838 17672
rect 3053 17663 3111 17669
rect 3053 17660 3065 17663
rect 2832 17632 3065 17660
rect 2832 17620 2838 17632
rect 3053 17629 3065 17632
rect 3099 17629 3111 17663
rect 3053 17623 3111 17629
rect 3329 17663 3387 17669
rect 3329 17629 3341 17663
rect 3375 17660 3387 17663
rect 4522 17660 4528 17672
rect 3375 17632 4528 17660
rect 3375 17629 3387 17632
rect 3329 17623 3387 17629
rect 4522 17620 4528 17632
rect 4580 17620 4586 17672
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17660 5227 17663
rect 6914 17660 6920 17672
rect 5215 17632 6920 17660
rect 5215 17629 5227 17632
rect 5169 17623 5227 17629
rect 6914 17620 6920 17632
rect 6972 17620 6978 17672
rect 7009 17663 7067 17669
rect 7009 17629 7021 17663
rect 7055 17660 7067 17663
rect 7282 17660 7288 17672
rect 7055 17632 7288 17660
rect 7055 17629 7067 17632
rect 7009 17623 7067 17629
rect 7282 17620 7288 17632
rect 7340 17620 7346 17672
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 9048 17669 9076 17700
rect 9398 17688 9404 17700
rect 9456 17728 9462 17740
rect 10505 17731 10563 17737
rect 10505 17728 10517 17731
rect 9456 17700 10517 17728
rect 9456 17688 9462 17700
rect 10505 17697 10517 17700
rect 10551 17697 10563 17731
rect 10505 17691 10563 17697
rect 7929 17663 7987 17669
rect 7929 17660 7941 17663
rect 7800 17632 7941 17660
rect 7800 17620 7806 17632
rect 7929 17629 7941 17632
rect 7975 17629 7987 17663
rect 7929 17623 7987 17629
rect 9033 17663 9091 17669
rect 9033 17629 9045 17663
rect 9079 17629 9091 17663
rect 11054 17660 11060 17672
rect 11015 17632 11060 17660
rect 9033 17623 9091 17629
rect 11054 17620 11060 17632
rect 11112 17620 11118 17672
rect 12894 17660 12900 17672
rect 12855 17632 12900 17660
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 21085 17663 21143 17669
rect 21085 17660 21097 17663
rect 13320 17632 21097 17660
rect 13320 17620 13326 17632
rect 21085 17629 21097 17632
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 2314 17592 2320 17604
rect 2148 17564 2320 17592
rect 2314 17552 2320 17564
rect 2372 17552 2378 17604
rect 3418 17552 3424 17604
rect 3476 17592 3482 17604
rect 4902 17595 4960 17601
rect 4902 17592 4914 17595
rect 3476 17564 4914 17592
rect 3476 17552 3482 17564
rect 4902 17561 4914 17564
rect 4948 17561 4960 17595
rect 4902 17555 4960 17561
rect 5721 17595 5779 17601
rect 5721 17561 5733 17595
rect 5767 17592 5779 17595
rect 6730 17592 6736 17604
rect 5767 17564 6736 17592
rect 5767 17561 5779 17564
rect 5721 17555 5779 17561
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 9490 17592 9496 17604
rect 6840 17564 9496 17592
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 1670 17484 1676 17536
rect 1728 17524 1734 17536
rect 1949 17527 2007 17533
rect 1949 17524 1961 17527
rect 1728 17496 1961 17524
rect 1728 17484 1734 17496
rect 1949 17493 1961 17496
rect 1995 17493 2007 17527
rect 2866 17524 2872 17536
rect 2827 17496 2872 17524
rect 1949 17487 2007 17493
rect 2866 17484 2872 17496
rect 2924 17484 2930 17536
rect 3789 17527 3847 17533
rect 3789 17493 3801 17527
rect 3835 17524 3847 17527
rect 3878 17524 3884 17536
rect 3835 17496 3884 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 3878 17484 3884 17496
rect 3936 17484 3942 17536
rect 5810 17484 5816 17536
rect 5868 17524 5874 17536
rect 6365 17527 6423 17533
rect 6365 17524 6377 17527
rect 5868 17496 6377 17524
rect 5868 17484 5874 17496
rect 6365 17493 6377 17496
rect 6411 17524 6423 17527
rect 6840 17524 6868 17564
rect 9490 17552 9496 17564
rect 9548 17592 9554 17604
rect 10321 17595 10379 17601
rect 10321 17592 10333 17595
rect 9548 17564 10333 17592
rect 9548 17552 9554 17564
rect 10321 17561 10333 17564
rect 10367 17561 10379 17595
rect 10321 17555 10379 17561
rect 10413 17595 10471 17601
rect 10413 17561 10425 17595
rect 10459 17592 10471 17595
rect 12526 17592 12532 17604
rect 10459 17564 12532 17592
rect 10459 17561 10471 17564
rect 10413 17555 10471 17561
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 6411 17496 6868 17524
rect 6411 17493 6423 17496
rect 6365 17487 6423 17493
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 7653 17527 7711 17533
rect 7653 17524 7665 17527
rect 7524 17496 7665 17524
rect 7524 17484 7530 17496
rect 7653 17493 7665 17496
rect 7699 17493 7711 17527
rect 8570 17524 8576 17536
rect 8531 17496 8576 17524
rect 7653 17487 7711 17493
rect 8570 17484 8576 17496
rect 8628 17484 8634 17536
rect 9677 17527 9735 17533
rect 9677 17493 9689 17527
rect 9723 17524 9735 17527
rect 9766 17524 9772 17536
rect 9723 17496 9772 17524
rect 9723 17493 9735 17496
rect 9677 17487 9735 17493
rect 9766 17484 9772 17496
rect 9824 17484 9830 17536
rect 11701 17527 11759 17533
rect 11701 17493 11713 17527
rect 11747 17524 11759 17527
rect 11790 17524 11796 17536
rect 11747 17496 11796 17524
rect 11747 17493 11759 17496
rect 11701 17487 11759 17493
rect 11790 17484 11796 17496
rect 11848 17484 11854 17536
rect 11974 17524 11980 17536
rect 11935 17496 11980 17524
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 13538 17524 13544 17536
rect 13499 17496 13544 17524
rect 13538 17484 13544 17496
rect 13596 17484 13602 17536
rect 21266 17524 21272 17536
rect 21227 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 3418 17320 3424 17332
rect 3379 17292 3424 17320
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 5718 17320 5724 17332
rect 5679 17292 5724 17320
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 6914 17252 6920 17264
rect 4356 17224 6920 17252
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 1673 17147 1731 17153
rect 1688 17116 1716 17147
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2590 17184 2596 17196
rect 2551 17156 2596 17184
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 4065 17187 4123 17193
rect 4065 17153 4077 17187
rect 4111 17184 4123 17187
rect 4246 17184 4252 17196
rect 4111 17156 4252 17184
rect 4111 17153 4123 17156
rect 4065 17147 4123 17153
rect 4246 17144 4252 17156
rect 4304 17144 4310 17196
rect 4356 17193 4384 17224
rect 4614 17193 4620 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17153 4399 17187
rect 4608 17184 4620 17193
rect 4575 17156 4620 17184
rect 4341 17147 4399 17153
rect 4608 17147 4620 17156
rect 4614 17144 4620 17147
rect 4672 17144 4678 17196
rect 6380 17193 6408 17224
rect 6914 17212 6920 17224
rect 6972 17252 6978 17264
rect 7926 17252 7932 17264
rect 6972 17224 7932 17252
rect 6972 17212 6978 17224
rect 7926 17212 7932 17224
rect 7984 17252 7990 17264
rect 11054 17252 11060 17264
rect 7984 17224 8064 17252
rect 7984 17212 7990 17224
rect 6365 17187 6423 17193
rect 6365 17153 6377 17187
rect 6411 17153 6423 17187
rect 6365 17147 6423 17153
rect 6632 17187 6690 17193
rect 6632 17153 6644 17187
rect 6678 17184 6690 17187
rect 7006 17184 7012 17196
rect 6678 17156 7012 17184
rect 6678 17153 6690 17156
rect 6632 17147 6690 17153
rect 7006 17144 7012 17156
rect 7064 17144 7070 17196
rect 8036 17193 8064 17224
rect 9692 17224 11060 17252
rect 8294 17193 8300 17196
rect 8021 17187 8079 17193
rect 8021 17153 8033 17187
rect 8067 17153 8079 17187
rect 8021 17147 8079 17153
rect 8288 17147 8300 17193
rect 8352 17184 8358 17196
rect 9692 17193 9720 17224
rect 11054 17212 11060 17224
rect 11112 17252 11118 17264
rect 11112 17224 11560 17252
rect 11112 17212 11118 17224
rect 9677 17187 9735 17193
rect 8352 17156 8388 17184
rect 8294 17144 8300 17147
rect 8352 17144 8358 17156
rect 9677 17153 9689 17187
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 11532 17193 11560 17224
rect 11790 17193 11796 17196
rect 9933 17187 9991 17193
rect 9933 17184 9945 17187
rect 9824 17156 9945 17184
rect 9824 17144 9830 17156
rect 9933 17153 9945 17156
rect 9979 17153 9991 17187
rect 9933 17147 9991 17153
rect 11517 17187 11575 17193
rect 11517 17153 11529 17187
rect 11563 17153 11575 17187
rect 11784 17184 11796 17193
rect 11751 17156 11796 17184
rect 11517 17147 11575 17153
rect 11784 17147 11796 17156
rect 11790 17144 11796 17147
rect 11848 17144 11854 17196
rect 2958 17116 2964 17128
rect 1688 17088 2964 17116
rect 2958 17076 2964 17088
rect 3016 17076 3022 17128
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17116 3203 17119
rect 4154 17116 4160 17128
rect 3191 17088 4160 17116
rect 3191 17085 3203 17088
rect 3145 17079 3203 17085
rect 4154 17076 4160 17088
rect 4212 17076 4218 17128
rect 1486 17048 1492 17060
rect 1447 17020 1492 17048
rect 1486 17008 1492 17020
rect 1544 17008 1550 17060
rect 1762 17008 1768 17060
rect 1820 17048 1826 17060
rect 2409 17051 2467 17057
rect 2409 17048 2421 17051
rect 1820 17020 2421 17048
rect 1820 17008 1826 17020
rect 2409 17017 2421 17020
rect 2455 17017 2467 17051
rect 2409 17011 2467 17017
rect 11057 17051 11115 17057
rect 11057 17017 11069 17051
rect 11103 17048 11115 17051
rect 11146 17048 11152 17060
rect 11103 17020 11152 17048
rect 11103 17017 11115 17020
rect 11057 17011 11115 17017
rect 11146 17008 11152 17020
rect 11204 17008 11210 17060
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 7742 16980 7748 16992
rect 7703 16952 7748 16980
rect 7742 16940 7748 16952
rect 7800 16940 7806 16992
rect 12894 16980 12900 16992
rect 12855 16952 12900 16980
rect 12894 16940 12900 16952
rect 12952 16940 12958 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 2685 16779 2743 16785
rect 2685 16745 2697 16779
rect 2731 16776 2743 16779
rect 2774 16776 2780 16788
rect 2731 16748 2780 16776
rect 2731 16745 2743 16748
rect 2685 16739 2743 16745
rect 2774 16736 2780 16748
rect 2832 16736 2838 16788
rect 2958 16776 2964 16788
rect 2919 16748 2964 16776
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 6914 16776 6920 16788
rect 5276 16748 6920 16776
rect 3878 16600 3884 16652
rect 3936 16640 3942 16652
rect 5276 16649 5304 16748
rect 6914 16736 6920 16748
rect 6972 16736 6978 16788
rect 13262 16776 13268 16788
rect 11072 16748 13268 16776
rect 6638 16708 6644 16720
rect 6599 16680 6644 16708
rect 6638 16668 6644 16680
rect 6696 16668 6702 16720
rect 11072 16708 11100 16748
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 10980 16680 11100 16708
rect 4341 16643 4399 16649
rect 4341 16640 4353 16643
rect 3936 16612 4353 16640
rect 3936 16600 3942 16612
rect 4341 16609 4353 16612
rect 4387 16609 4399 16643
rect 4341 16603 4399 16609
rect 5261 16643 5319 16649
rect 5261 16609 5273 16643
rect 5307 16609 5319 16643
rect 7834 16640 7840 16652
rect 5261 16603 5319 16609
rect 7576 16612 7840 16640
rect 1670 16572 1676 16584
rect 1631 16544 1676 16572
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2501 16575 2559 16581
rect 2501 16541 2513 16575
rect 2547 16572 2559 16575
rect 2682 16572 2688 16584
rect 2547 16544 2688 16572
rect 2547 16541 2559 16544
rect 2501 16535 2559 16541
rect 2240 16504 2268 16535
rect 2682 16532 2688 16544
rect 2740 16532 2746 16584
rect 3142 16572 3148 16584
rect 3103 16544 3148 16572
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 4154 16572 4160 16584
rect 4115 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 5350 16532 5356 16584
rect 5408 16572 5414 16584
rect 7576 16581 7604 16612
rect 7834 16600 7840 16612
rect 7892 16640 7898 16652
rect 8389 16643 8447 16649
rect 8389 16640 8401 16643
rect 7892 16612 8401 16640
rect 7892 16600 7898 16612
rect 8389 16609 8401 16612
rect 8435 16609 8447 16643
rect 8389 16603 8447 16609
rect 9398 16600 9404 16652
rect 9456 16640 9462 16652
rect 10980 16649 11008 16680
rect 9493 16643 9551 16649
rect 9493 16640 9505 16643
rect 9456 16612 9505 16640
rect 9456 16600 9462 16612
rect 9493 16609 9505 16612
rect 9539 16609 9551 16643
rect 10045 16643 10103 16649
rect 10045 16640 10057 16643
rect 9493 16603 9551 16609
rect 9600 16612 10057 16640
rect 5517 16575 5575 16581
rect 5517 16572 5529 16575
rect 5408 16544 5529 16572
rect 5408 16532 5414 16544
rect 5517 16541 5529 16544
rect 5563 16541 5575 16575
rect 5517 16535 5575 16541
rect 7561 16575 7619 16581
rect 7561 16541 7573 16575
rect 7607 16541 7619 16575
rect 8202 16572 8208 16584
rect 8163 16544 8208 16572
rect 7561 16535 7619 16541
rect 8202 16532 8208 16544
rect 8260 16532 8266 16584
rect 8294 16532 8300 16584
rect 8352 16532 8358 16584
rect 2866 16504 2872 16516
rect 2240 16476 2872 16504
rect 2866 16464 2872 16476
rect 2924 16464 2930 16516
rect 6917 16507 6975 16513
rect 6917 16473 6929 16507
rect 6963 16504 6975 16507
rect 8312 16504 8340 16532
rect 6963 16476 8340 16504
rect 9401 16507 9459 16513
rect 6963 16473 6975 16476
rect 6917 16467 6975 16473
rect 9401 16473 9413 16507
rect 9447 16504 9459 16507
rect 9600 16504 9628 16612
rect 10045 16609 10057 16612
rect 10091 16640 10103 16643
rect 10965 16643 11023 16649
rect 10091 16612 10916 16640
rect 10091 16609 10103 16612
rect 10045 16603 10103 16609
rect 10888 16572 10916 16612
rect 10965 16609 10977 16643
rect 11011 16609 11023 16643
rect 10965 16603 11023 16609
rect 11054 16600 11060 16652
rect 11112 16640 11118 16652
rect 11885 16643 11943 16649
rect 11885 16640 11897 16643
rect 11112 16612 11897 16640
rect 11112 16600 11118 16612
rect 11885 16609 11897 16612
rect 11931 16609 11943 16643
rect 11885 16603 11943 16609
rect 11146 16572 11152 16584
rect 10888 16544 11152 16572
rect 11146 16532 11152 16544
rect 11204 16532 11210 16584
rect 11241 16575 11299 16581
rect 11241 16541 11253 16575
rect 11287 16572 11299 16575
rect 11974 16572 11980 16584
rect 11287 16544 11980 16572
rect 11287 16541 11299 16544
rect 11241 16535 11299 16541
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 12152 16575 12210 16581
rect 12152 16541 12164 16575
rect 12198 16572 12210 16575
rect 13538 16572 13544 16584
rect 12198 16544 13544 16572
rect 12198 16541 12210 16544
rect 12152 16535 12210 16541
rect 13538 16532 13544 16544
rect 13596 16532 13602 16584
rect 9447 16476 9628 16504
rect 9447 16473 9459 16476
rect 9401 16467 9459 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2038 16436 2044 16448
rect 1999 16408 2044 16436
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 3234 16396 3240 16448
rect 3292 16436 3298 16448
rect 3789 16439 3847 16445
rect 3789 16436 3801 16439
rect 3292 16408 3801 16436
rect 3292 16396 3298 16408
rect 3789 16405 3801 16408
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 4985 16439 5043 16445
rect 4304 16408 4349 16436
rect 4304 16396 4310 16408
rect 4985 16405 4997 16439
rect 5031 16436 5043 16439
rect 5718 16436 5724 16448
rect 5031 16408 5724 16436
rect 5031 16405 5043 16408
rect 4985 16399 5043 16405
rect 5718 16396 5724 16408
rect 5776 16396 5782 16448
rect 6546 16396 6552 16448
rect 6604 16436 6610 16448
rect 7837 16439 7895 16445
rect 7837 16436 7849 16439
rect 6604 16408 7849 16436
rect 6604 16396 6610 16408
rect 7837 16405 7849 16408
rect 7883 16405 7895 16439
rect 7837 16399 7895 16405
rect 8297 16439 8355 16445
rect 8297 16405 8309 16439
rect 8343 16436 8355 16439
rect 8941 16439 8999 16445
rect 8941 16436 8953 16439
rect 8343 16408 8953 16436
rect 8343 16405 8355 16408
rect 8297 16399 8355 16405
rect 8941 16405 8953 16408
rect 8987 16405 8999 16439
rect 9306 16436 9312 16448
rect 9267 16408 9312 16436
rect 8941 16399 8999 16405
rect 9306 16396 9312 16408
rect 9364 16436 9370 16448
rect 10321 16439 10379 16445
rect 10321 16436 10333 16439
rect 9364 16408 10333 16436
rect 9364 16396 9370 16408
rect 10321 16405 10333 16408
rect 10367 16405 10379 16439
rect 11146 16436 11152 16448
rect 11107 16408 11152 16436
rect 10321 16399 10379 16405
rect 11146 16396 11152 16408
rect 11204 16396 11210 16448
rect 11609 16439 11667 16445
rect 11609 16405 11621 16439
rect 11655 16436 11667 16439
rect 11698 16436 11704 16448
rect 11655 16408 11704 16436
rect 11655 16405 11667 16408
rect 11609 16399 11667 16405
rect 11698 16396 11704 16408
rect 11756 16396 11762 16448
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 2590 16232 2596 16244
rect 2551 16204 2596 16232
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 4246 16192 4252 16244
rect 4304 16232 4310 16244
rect 4617 16235 4675 16241
rect 4617 16232 4629 16235
rect 4304 16204 4629 16232
rect 4304 16192 4310 16204
rect 4617 16201 4629 16204
rect 4663 16201 4675 16235
rect 4617 16195 4675 16201
rect 5994 16192 6000 16244
rect 6052 16232 6058 16244
rect 6733 16235 6791 16241
rect 6733 16232 6745 16235
rect 6052 16204 6745 16232
rect 6052 16192 6058 16204
rect 6733 16201 6745 16204
rect 6779 16201 6791 16235
rect 7834 16232 7840 16244
rect 7795 16204 7840 16232
rect 6733 16195 6791 16201
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9306 16232 9312 16244
rect 8864 16204 9312 16232
rect 4522 16124 4528 16176
rect 4580 16164 4586 16176
rect 4985 16167 5043 16173
rect 4985 16164 4997 16167
rect 4580 16136 4997 16164
rect 4580 16124 4586 16136
rect 4985 16133 4997 16136
rect 5031 16164 5043 16167
rect 6638 16164 6644 16176
rect 5031 16136 6644 16164
rect 5031 16133 5043 16136
rect 4985 16127 5043 16133
rect 6638 16124 6644 16136
rect 6696 16164 6702 16176
rect 8864 16164 8892 16204
rect 9306 16192 9312 16204
rect 9364 16192 9370 16244
rect 11146 16192 11152 16244
rect 11204 16232 11210 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 11204 16204 11529 16232
rect 11204 16192 11210 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 11517 16195 11575 16201
rect 6696 16136 8892 16164
rect 8972 16167 9030 16173
rect 6696 16124 6702 16136
rect 8972 16133 8984 16167
rect 9018 16164 9030 16167
rect 10137 16167 10195 16173
rect 10137 16164 10149 16167
rect 9018 16136 10149 16164
rect 9018 16133 9030 16136
rect 8972 16127 9030 16133
rect 10137 16133 10149 16136
rect 10183 16133 10195 16167
rect 10137 16127 10195 16133
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 1762 16096 1768 16108
rect 1719 16068 1768 16096
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 1762 16056 1768 16068
rect 1820 16056 1826 16108
rect 1949 16099 2007 16105
rect 1949 16065 1961 16099
rect 1995 16096 2007 16099
rect 2130 16096 2136 16108
rect 1995 16068 2136 16096
rect 1995 16065 2007 16068
rect 1949 16059 2007 16065
rect 2130 16056 2136 16068
rect 2188 16056 2194 16108
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2590 16096 2596 16108
rect 2455 16068 2596 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 2866 16056 2872 16108
rect 2924 16096 2930 16108
rect 3217 16099 3275 16105
rect 3217 16096 3229 16099
rect 2924 16068 3229 16096
rect 2924 16056 2930 16068
rect 3217 16065 3229 16068
rect 3263 16065 3275 16099
rect 5997 16099 6055 16105
rect 3217 16059 3275 16065
rect 5092 16068 5957 16096
rect 5092 16037 5120 16068
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 15997 3019 16031
rect 2961 15991 3019 15997
rect 5077 16031 5135 16037
rect 5077 15997 5089 16031
rect 5123 15997 5135 16031
rect 5077 15991 5135 15997
rect 5169 16031 5227 16037
rect 5169 15997 5181 16031
rect 5215 15997 5227 16031
rect 5929 16028 5957 16068
rect 5997 16065 6009 16099
rect 6043 16096 6055 16099
rect 7101 16099 7159 16105
rect 7101 16096 7113 16099
rect 6043 16068 7113 16096
rect 6043 16065 6055 16068
rect 5997 16059 6055 16065
rect 7101 16065 7113 16068
rect 7147 16065 7159 16099
rect 7101 16059 7159 16065
rect 9306 16056 9312 16108
rect 9364 16096 9370 16108
rect 9493 16099 9551 16105
rect 9493 16096 9505 16099
rect 9364 16068 9505 16096
rect 9364 16056 9370 16068
rect 9493 16065 9505 16068
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 11146 16056 11152 16108
rect 11204 16096 11210 16108
rect 11885 16099 11943 16105
rect 11885 16096 11897 16099
rect 11204 16068 11897 16096
rect 11204 16056 11210 16068
rect 11885 16065 11897 16068
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 7190 16028 7196 16040
rect 5929 16000 7052 16028
rect 7151 16000 7196 16028
rect 5169 15991 5227 15997
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2976 15892 3004 15991
rect 4338 15960 4344 15972
rect 4299 15932 4344 15960
rect 4338 15920 4344 15932
rect 4396 15960 4402 15972
rect 5184 15960 5212 15991
rect 4396 15932 5212 15960
rect 7024 15960 7052 16000
rect 7190 15988 7196 16000
rect 7248 15988 7254 16040
rect 7282 15988 7288 16040
rect 7340 16028 7346 16040
rect 9214 16028 9220 16040
rect 7340 16000 7385 16028
rect 9175 16000 9220 16028
rect 7340 15988 7346 16000
rect 9214 15988 9220 16000
rect 9272 15988 9278 16040
rect 10410 16028 10416 16040
rect 10371 16000 10416 16028
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 11974 16028 11980 16040
rect 11935 16000 11980 16028
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12161 16031 12219 16037
rect 12161 15997 12173 16031
rect 12207 16028 12219 16031
rect 12894 16028 12900 16040
rect 12207 16000 12900 16028
rect 12207 15997 12219 16000
rect 12161 15991 12219 15997
rect 12894 15988 12900 16000
rect 12952 15988 12958 16040
rect 8018 15960 8024 15972
rect 7024 15932 8024 15960
rect 4396 15920 4402 15932
rect 8018 15920 8024 15932
rect 8076 15920 8082 15972
rect 3878 15892 3884 15904
rect 2976 15864 3884 15892
rect 3878 15852 3884 15864
rect 3936 15852 3942 15904
rect 6457 15895 6515 15901
rect 6457 15861 6469 15895
rect 6503 15892 6515 15895
rect 6546 15892 6552 15904
rect 6503 15864 6552 15892
rect 6503 15861 6515 15864
rect 6457 15855 6515 15861
rect 6546 15852 6552 15864
rect 6604 15852 6610 15904
rect 11146 15892 11152 15904
rect 11107 15864 11152 15892
rect 11146 15852 11152 15864
rect 11204 15852 11210 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 2406 15648 2412 15700
rect 2464 15688 2470 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2464 15660 2697 15688
rect 2464 15648 2470 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 2685 15651 2743 15657
rect 2774 15648 2780 15700
rect 2832 15688 2838 15700
rect 4249 15691 4307 15697
rect 4249 15688 4261 15691
rect 2832 15660 4261 15688
rect 2832 15648 2838 15660
rect 4249 15657 4261 15660
rect 4295 15657 4307 15691
rect 4249 15651 4307 15657
rect 6549 15691 6607 15697
rect 6549 15657 6561 15691
rect 6595 15688 6607 15691
rect 7282 15688 7288 15700
rect 6595 15660 7288 15688
rect 6595 15657 6607 15660
rect 6549 15651 6607 15657
rect 7282 15648 7288 15660
rect 7340 15648 7346 15700
rect 8941 15691 8999 15697
rect 8941 15657 8953 15691
rect 8987 15688 8999 15691
rect 9306 15688 9312 15700
rect 8987 15660 9312 15688
rect 8987 15657 8999 15660
rect 8941 15651 8999 15657
rect 9306 15648 9312 15660
rect 9364 15648 9370 15700
rect 11698 15688 11704 15700
rect 9416 15660 11704 15688
rect 5353 15623 5411 15629
rect 5353 15620 5365 15623
rect 3160 15592 5365 15620
rect 1946 15552 1952 15564
rect 1688 15524 1952 15552
rect 1688 15493 1716 15524
rect 1946 15512 1952 15524
rect 2004 15512 2010 15564
rect 3160 15561 3188 15592
rect 5353 15589 5365 15592
rect 5399 15589 5411 15623
rect 5353 15583 5411 15589
rect 8018 15580 8024 15632
rect 8076 15620 8082 15632
rect 8297 15623 8355 15629
rect 8297 15620 8309 15623
rect 8076 15592 8309 15620
rect 8076 15580 8082 15592
rect 8297 15589 8309 15592
rect 8343 15620 8355 15623
rect 9416 15620 9444 15660
rect 11698 15648 11704 15660
rect 11756 15648 11762 15700
rect 8343 15592 9444 15620
rect 8343 15589 8355 15592
rect 8297 15583 8355 15589
rect 3145 15555 3203 15561
rect 3145 15521 3157 15555
rect 3191 15521 3203 15555
rect 3326 15552 3332 15564
rect 3287 15524 3332 15552
rect 3145 15515 3203 15521
rect 3326 15512 3332 15524
rect 3384 15512 3390 15564
rect 4890 15552 4896 15564
rect 4851 15524 4896 15552
rect 4890 15512 4896 15524
rect 4948 15512 4954 15564
rect 5902 15552 5908 15564
rect 5863 15524 5908 15552
rect 5902 15512 5908 15524
rect 5960 15512 5966 15564
rect 7926 15552 7932 15564
rect 7887 15524 7932 15552
rect 7926 15512 7932 15524
rect 7984 15512 7990 15564
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1854 15444 1860 15496
rect 1912 15484 1918 15496
rect 2133 15487 2191 15493
rect 2133 15484 2145 15487
rect 1912 15456 2145 15484
rect 1912 15444 1918 15456
rect 2133 15453 2145 15456
rect 2179 15453 2191 15487
rect 2133 15447 2191 15453
rect 7673 15487 7731 15493
rect 7673 15453 7685 15487
rect 7719 15484 7731 15487
rect 8570 15484 8576 15496
rect 7719 15456 8576 15484
rect 7719 15453 7731 15456
rect 7673 15447 7731 15453
rect 8570 15444 8576 15456
rect 8628 15444 8634 15496
rect 9214 15444 9220 15496
rect 9272 15484 9278 15496
rect 10321 15487 10379 15493
rect 10321 15484 10333 15487
rect 9272 15456 10333 15484
rect 9272 15444 9278 15456
rect 10321 15453 10333 15456
rect 10367 15484 10379 15487
rect 10962 15484 10968 15496
rect 10367 15456 10968 15484
rect 10367 15453 10379 15456
rect 10321 15447 10379 15453
rect 10962 15444 10968 15456
rect 11020 15444 11026 15496
rect 11241 15487 11299 15493
rect 11241 15453 11253 15487
rect 11287 15453 11299 15487
rect 11241 15447 11299 15453
rect 3053 15419 3111 15425
rect 3053 15385 3065 15419
rect 3099 15416 3111 15419
rect 3789 15419 3847 15425
rect 3789 15416 3801 15419
rect 3099 15388 3801 15416
rect 3099 15385 3111 15388
rect 3053 15379 3111 15385
rect 3789 15385 3801 15388
rect 3835 15385 3847 15419
rect 10076 15419 10134 15425
rect 3789 15379 3847 15385
rect 8404 15388 9674 15416
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 1670 15308 1676 15360
rect 1728 15348 1734 15360
rect 1949 15351 2007 15357
rect 1949 15348 1961 15351
rect 1728 15320 1961 15348
rect 1728 15308 1734 15320
rect 1949 15317 1961 15320
rect 1995 15317 2007 15351
rect 1949 15311 2007 15317
rect 4154 15308 4160 15360
rect 4212 15348 4218 15360
rect 4617 15351 4675 15357
rect 4617 15348 4629 15351
rect 4212 15320 4629 15348
rect 4212 15308 4218 15320
rect 4617 15317 4629 15320
rect 4663 15317 4675 15351
rect 4617 15311 4675 15317
rect 4706 15308 4712 15360
rect 4764 15348 4770 15360
rect 5718 15348 5724 15360
rect 4764 15320 4809 15348
rect 5679 15320 5724 15348
rect 4764 15308 4770 15320
rect 5718 15308 5724 15320
rect 5776 15308 5782 15360
rect 5813 15351 5871 15357
rect 5813 15317 5825 15351
rect 5859 15348 5871 15351
rect 8404 15348 8432 15388
rect 5859 15320 8432 15348
rect 9646 15348 9674 15388
rect 10076 15385 10088 15419
rect 10122 15416 10134 15419
rect 10597 15419 10655 15425
rect 10597 15416 10609 15419
rect 10122 15388 10609 15416
rect 10122 15385 10134 15388
rect 10076 15379 10134 15385
rect 10597 15385 10609 15388
rect 10643 15385 10655 15419
rect 10597 15379 10655 15385
rect 10778 15376 10784 15428
rect 10836 15416 10842 15428
rect 11256 15416 11284 15447
rect 10836 15388 11284 15416
rect 10836 15376 10842 15388
rect 12434 15348 12440 15360
rect 9646 15320 12440 15348
rect 5859 15317 5871 15320
rect 5813 15311 5871 15317
rect 12434 15308 12440 15320
rect 12492 15308 12498 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 2314 15144 2320 15156
rect 2275 15116 2320 15144
rect 2314 15104 2320 15116
rect 2372 15104 2378 15156
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 2866 15144 2872 15156
rect 2823 15116 2872 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 2866 15104 2872 15116
rect 2924 15104 2930 15156
rect 4617 15147 4675 15153
rect 4617 15144 4629 15147
rect 3620 15116 4629 15144
rect 1670 15008 1676 15020
rect 1631 14980 1676 15008
rect 1670 14968 1676 14980
rect 1728 14968 1734 15020
rect 2501 15011 2559 15017
rect 2501 14977 2513 15011
rect 2547 14977 2559 15011
rect 2501 14971 2559 14977
rect 2516 14940 2544 14971
rect 3326 14968 3332 15020
rect 3384 15008 3390 15020
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 3384 14980 3433 15008
rect 3384 14968 3390 14980
rect 3421 14977 3433 14980
rect 3467 15008 3479 15011
rect 3620 15008 3648 15116
rect 4617 15113 4629 15116
rect 4663 15113 4675 15147
rect 7190 15144 7196 15156
rect 7151 15116 7196 15144
rect 4617 15107 4675 15113
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8205 15147 8263 15153
rect 8205 15113 8217 15147
rect 8251 15144 8263 15147
rect 8251 15116 8285 15144
rect 8251 15113 8263 15116
rect 8205 15107 8263 15113
rect 3697 15079 3755 15085
rect 3697 15045 3709 15079
rect 3743 15076 3755 15079
rect 5730 15079 5788 15085
rect 5730 15076 5742 15079
rect 3743 15048 5742 15076
rect 3743 15045 3755 15048
rect 3697 15039 3755 15045
rect 5730 15045 5742 15048
rect 5776 15045 5788 15079
rect 6914 15076 6920 15088
rect 5730 15039 5788 15045
rect 6012 15048 6920 15076
rect 3467 14980 3648 15008
rect 4341 15011 4399 15017
rect 3467 14977 3479 14980
rect 3421 14971 3479 14977
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 5902 15008 5908 15020
rect 4387 14980 5908 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 5902 14968 5908 14980
rect 5960 14968 5966 15020
rect 6012 15017 6040 15048
rect 6914 15036 6920 15048
rect 6972 15076 6978 15088
rect 7926 15076 7932 15088
rect 6972 15048 7932 15076
rect 6972 15036 6978 15048
rect 7926 15036 7932 15048
rect 7984 15036 7990 15088
rect 8220 15076 8248 15107
rect 8662 15104 8668 15156
rect 8720 15144 8726 15156
rect 8757 15147 8815 15153
rect 8757 15144 8769 15147
rect 8720 15116 8769 15144
rect 8720 15104 8726 15116
rect 8757 15113 8769 15116
rect 8803 15113 8815 15147
rect 8757 15107 8815 15113
rect 9125 15147 9183 15153
rect 9125 15113 9137 15147
rect 9171 15144 9183 15147
rect 10410 15144 10416 15156
rect 9171 15116 10416 15144
rect 9171 15113 9183 15116
rect 9125 15107 9183 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 11146 15104 11152 15156
rect 11204 15104 11210 15156
rect 11164 15076 11192 15104
rect 11790 15076 11796 15088
rect 8027 15048 11796 15076
rect 5997 15011 6055 15017
rect 5997 14977 6009 15011
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 6365 15011 6423 15017
rect 6365 14977 6377 15011
rect 6411 15008 6423 15011
rect 6454 15008 6460 15020
rect 6411 14980 6460 15008
rect 6411 14977 6423 14980
rect 6365 14971 6423 14977
rect 6454 14968 6460 14980
rect 6512 14968 6518 15020
rect 7561 15011 7619 15017
rect 7561 15008 7573 15011
rect 6647 14980 7573 15008
rect 4246 14940 4252 14952
rect 2516 14912 4252 14940
rect 4246 14900 4252 14912
rect 4304 14900 4310 14952
rect 6546 14872 6552 14884
rect 6507 14844 6552 14872
rect 6546 14832 6552 14844
rect 6604 14832 6610 14884
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 1762 14764 1768 14816
rect 1820 14804 1826 14816
rect 2041 14807 2099 14813
rect 2041 14804 2053 14807
rect 1820 14776 2053 14804
rect 1820 14764 1826 14776
rect 2041 14773 2053 14776
rect 2087 14804 2099 14807
rect 2314 14804 2320 14816
rect 2087 14776 2320 14804
rect 2087 14773 2099 14776
rect 2041 14767 2099 14773
rect 2314 14764 2320 14776
rect 2372 14764 2378 14816
rect 5074 14764 5080 14816
rect 5132 14804 5138 14816
rect 6647 14804 6675 14980
rect 7561 14977 7573 14980
rect 7607 15008 7619 15011
rect 8027 15008 8055 15048
rect 11790 15036 11796 15048
rect 11848 15036 11854 15088
rect 10870 15008 10876 15020
rect 10928 15017 10934 15020
rect 7607 14980 8055 15008
rect 10840 14980 10876 15008
rect 7607 14977 7619 14980
rect 7561 14971 7619 14977
rect 10870 14968 10876 14980
rect 10928 14971 10940 15017
rect 10928 14968 10934 14971
rect 11054 14968 11060 15020
rect 11112 15008 11118 15020
rect 11149 15011 11207 15017
rect 11149 15008 11161 15011
rect 11112 14980 11161 15008
rect 11112 14968 11118 14980
rect 11149 14977 11161 14980
rect 11195 14977 11207 15011
rect 11149 14971 11207 14977
rect 7650 14940 7656 14952
rect 7611 14912 7656 14940
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7742 14900 7748 14952
rect 7800 14940 7806 14952
rect 9214 14940 9220 14952
rect 7800 14912 7845 14940
rect 9175 14912 9220 14940
rect 7800 14900 7806 14912
rect 9214 14900 9220 14912
rect 9272 14900 9278 14952
rect 9401 14943 9459 14949
rect 9401 14909 9413 14943
rect 9447 14940 9459 14943
rect 9447 14912 9812 14940
rect 9447 14909 9459 14912
rect 9401 14903 9459 14909
rect 5132 14776 6675 14804
rect 6917 14807 6975 14813
rect 5132 14764 5138 14776
rect 6917 14773 6929 14807
rect 6963 14804 6975 14807
rect 7282 14804 7288 14816
rect 6963 14776 7288 14804
rect 6963 14773 6975 14776
rect 6917 14767 6975 14773
rect 7282 14764 7288 14776
rect 7340 14764 7346 14816
rect 9784 14813 9812 14912
rect 9769 14807 9827 14813
rect 9769 14773 9781 14807
rect 9815 14804 9827 14807
rect 10778 14804 10784 14816
rect 9815 14776 10784 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 10778 14764 10784 14776
rect 10836 14764 10842 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 4982 14600 4988 14612
rect 3804 14572 4988 14600
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2406 14396 2412 14408
rect 2271 14368 2412 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 3421 14399 3479 14405
rect 3421 14365 3433 14399
rect 3467 14396 3479 14399
rect 3804 14396 3832 14572
rect 4982 14560 4988 14572
rect 5040 14560 5046 14612
rect 5721 14603 5779 14609
rect 5721 14569 5733 14603
rect 5767 14600 5779 14603
rect 5902 14600 5908 14612
rect 5767 14572 5908 14600
rect 5767 14569 5779 14572
rect 5721 14563 5779 14569
rect 5902 14560 5908 14572
rect 5960 14560 5966 14612
rect 5994 14560 6000 14612
rect 6052 14600 6058 14612
rect 6052 14572 8800 14600
rect 6052 14560 6058 14572
rect 8772 14544 8800 14572
rect 10870 14560 10876 14612
rect 10928 14600 10934 14612
rect 11793 14603 11851 14609
rect 11793 14600 11805 14603
rect 10928 14572 11805 14600
rect 10928 14560 10934 14572
rect 11793 14569 11805 14572
rect 11839 14569 11851 14603
rect 11793 14563 11851 14569
rect 8754 14492 8760 14544
rect 8812 14492 8818 14544
rect 4065 14467 4123 14473
rect 4065 14433 4077 14467
rect 4111 14464 4123 14467
rect 4154 14464 4160 14476
rect 4111 14436 4160 14464
rect 4111 14433 4123 14436
rect 4065 14427 4123 14433
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 5534 14464 5540 14476
rect 5368 14436 5540 14464
rect 3467 14368 3832 14396
rect 3467 14365 3479 14368
rect 3421 14359 3479 14365
rect 3878 14356 3884 14408
rect 3936 14396 3942 14408
rect 4341 14399 4399 14405
rect 4341 14396 4353 14399
rect 3936 14368 4353 14396
rect 3936 14356 3942 14368
rect 4341 14365 4353 14368
rect 4387 14396 4399 14399
rect 5368 14396 5396 14436
rect 5534 14424 5540 14436
rect 5592 14464 5598 14476
rect 6914 14464 6920 14476
rect 5592 14436 6920 14464
rect 5592 14424 5598 14436
rect 6914 14424 6920 14436
rect 6972 14424 6978 14476
rect 10796 14436 11192 14464
rect 4387 14368 5396 14396
rect 6641 14399 6699 14405
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 7006 14396 7012 14408
rect 6687 14368 7012 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 7006 14356 7012 14368
rect 7064 14356 7070 14408
rect 7184 14399 7242 14405
rect 7184 14365 7196 14399
rect 7230 14396 7242 14399
rect 7466 14396 7472 14408
rect 7230 14368 7472 14396
rect 7230 14365 7242 14368
rect 7184 14359 7242 14365
rect 7466 14356 7472 14368
rect 7524 14356 7530 14408
rect 10796 14396 10824 14436
rect 10336 14368 10824 14396
rect 10873 14399 10931 14405
rect 2777 14331 2835 14337
rect 2777 14297 2789 14331
rect 2823 14328 2835 14331
rect 4586 14331 4644 14337
rect 4586 14328 4598 14331
rect 2823 14300 4598 14328
rect 2823 14297 2835 14300
rect 2777 14291 2835 14297
rect 4586 14297 4598 14300
rect 4632 14297 4644 14331
rect 4586 14291 4644 14297
rect 5718 14288 5724 14340
rect 5776 14328 5782 14340
rect 9125 14331 9183 14337
rect 9125 14328 9137 14331
rect 5776 14300 9137 14328
rect 5776 14288 5782 14300
rect 9125 14297 9137 14300
rect 9171 14328 9183 14331
rect 9306 14328 9312 14340
rect 9171 14300 9312 14328
rect 9171 14297 9183 14300
rect 9125 14291 9183 14297
rect 9306 14288 9312 14300
rect 9364 14328 9370 14340
rect 9582 14328 9588 14340
rect 9364 14300 9588 14328
rect 9364 14288 9370 14300
rect 9582 14288 9588 14300
rect 9640 14288 9646 14340
rect 10336 14272 10364 14368
rect 10873 14365 10885 14399
rect 10919 14396 10931 14399
rect 11054 14396 11060 14408
rect 10919 14368 11060 14396
rect 10919 14365 10931 14368
rect 10873 14359 10931 14365
rect 11054 14356 11060 14368
rect 11112 14356 11118 14408
rect 11164 14405 11192 14436
rect 11698 14424 11704 14476
rect 11756 14464 11762 14476
rect 19978 14464 19984 14476
rect 11756 14436 19984 14464
rect 11756 14424 11762 14436
rect 19978 14424 19984 14436
rect 20036 14424 20042 14476
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 10628 14331 10686 14337
rect 10628 14297 10640 14331
rect 10674 14328 10686 14331
rect 12250 14328 12256 14340
rect 10674 14300 12256 14328
rect 10674 14297 10686 14300
rect 10628 14291 10686 14297
rect 12250 14288 12256 14300
rect 12308 14288 12314 14340
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2038 14260 2044 14272
rect 1999 14232 2044 14260
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 5997 14263 6055 14269
rect 5997 14229 6009 14263
rect 6043 14260 6055 14263
rect 6914 14260 6920 14272
rect 6043 14232 6920 14260
rect 6043 14229 6055 14232
rect 5997 14223 6055 14229
rect 6914 14220 6920 14232
rect 6972 14220 6978 14272
rect 8018 14220 8024 14272
rect 8076 14260 8082 14272
rect 8297 14263 8355 14269
rect 8297 14260 8309 14263
rect 8076 14232 8309 14260
rect 8076 14220 8082 14232
rect 8297 14229 8309 14232
rect 8343 14229 8355 14263
rect 8297 14223 8355 14229
rect 9493 14263 9551 14269
rect 9493 14229 9505 14263
rect 9539 14260 9551 14263
rect 10318 14260 10324 14272
rect 9539 14232 10324 14260
rect 9539 14229 9551 14232
rect 9493 14223 9551 14229
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 18138 14260 18144 14272
rect 11296 14232 18144 14260
rect 11296 14220 11302 14232
rect 18138 14220 18144 14232
rect 18196 14220 18202 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 2406 14056 2412 14068
rect 2367 14028 2412 14056
rect 2406 14016 2412 14028
rect 2464 14016 2470 14068
rect 4890 14016 4896 14068
rect 4948 14056 4954 14068
rect 5261 14059 5319 14065
rect 5261 14056 5273 14059
rect 4948 14028 5273 14056
rect 4948 14016 4954 14028
rect 5261 14025 5273 14028
rect 5307 14025 5319 14059
rect 5261 14019 5319 14025
rect 5721 14059 5779 14065
rect 5721 14025 5733 14059
rect 5767 14056 5779 14059
rect 8662 14056 8668 14068
rect 5767 14028 8668 14056
rect 5767 14025 5779 14028
rect 5721 14019 5779 14025
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 8754 14016 8760 14068
rect 8812 14056 8818 14068
rect 8812 14028 8857 14056
rect 8812 14016 8818 14028
rect 9214 14016 9220 14068
rect 9272 14056 9278 14068
rect 9769 14059 9827 14065
rect 9769 14056 9781 14059
rect 9272 14028 9781 14056
rect 9272 14016 9278 14028
rect 9769 14025 9781 14028
rect 9815 14025 9827 14059
rect 9769 14019 9827 14025
rect 2314 13948 2320 14000
rect 2372 13988 2378 14000
rect 5902 13988 5908 14000
rect 2372 13960 5908 13988
rect 2372 13948 2378 13960
rect 5902 13948 5908 13960
rect 5960 13948 5966 14000
rect 8570 13988 8576 14000
rect 6564 13960 8576 13988
rect 2130 13920 2136 13932
rect 2091 13892 2136 13920
rect 2130 13880 2136 13892
rect 2188 13880 2194 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2958 13920 2964 13932
rect 2639 13892 2774 13920
rect 2919 13892 2964 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 1394 13812 1400 13864
rect 1452 13852 1458 13864
rect 1489 13855 1547 13861
rect 1489 13852 1501 13855
rect 1452 13824 1501 13852
rect 1452 13812 1458 13824
rect 1489 13821 1501 13824
rect 1535 13821 1547 13855
rect 2746 13852 2774 13892
rect 2958 13880 2964 13892
rect 3016 13880 3022 13932
rect 3878 13920 3884 13932
rect 3839 13892 3884 13920
rect 3878 13880 3884 13892
rect 3936 13880 3942 13932
rect 4154 13929 4160 13932
rect 4148 13883 4160 13929
rect 4212 13920 4218 13932
rect 4212 13892 4248 13920
rect 4154 13880 4160 13883
rect 4212 13880 4218 13892
rect 4430 13880 4436 13932
rect 4488 13920 4494 13932
rect 5537 13923 5595 13929
rect 5537 13920 5549 13923
rect 4488 13892 5549 13920
rect 4488 13880 4494 13892
rect 5537 13889 5549 13892
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 5994 13880 6000 13932
rect 6052 13920 6058 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 6052 13892 6377 13920
rect 6052 13880 6058 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 2866 13852 2872 13864
rect 2746 13824 2872 13852
rect 1489 13815 1547 13821
rect 2866 13812 2872 13824
rect 2924 13812 2930 13864
rect 6564 13793 6592 13960
rect 8570 13948 8576 13960
rect 8628 13948 8634 14000
rect 9125 13991 9183 13997
rect 9125 13957 9137 13991
rect 9171 13988 9183 13991
rect 10781 13991 10839 13997
rect 10781 13988 10793 13991
rect 9171 13960 10793 13988
rect 9171 13957 9183 13960
rect 9125 13951 9183 13957
rect 10781 13957 10793 13960
rect 10827 13957 10839 13991
rect 10781 13951 10839 13957
rect 8018 13880 8024 13932
rect 8076 13929 8082 13932
rect 8076 13920 8088 13929
rect 9217 13923 9275 13929
rect 8076 13892 8121 13920
rect 8076 13883 8088 13892
rect 9217 13889 9229 13923
rect 9263 13920 9275 13923
rect 9858 13920 9864 13932
rect 9263 13892 9864 13920
rect 9263 13889 9275 13892
rect 9217 13883 9275 13889
rect 8076 13880 8082 13883
rect 9858 13880 9864 13892
rect 9916 13880 9922 13932
rect 10137 13923 10195 13929
rect 10137 13889 10149 13923
rect 10183 13889 10195 13923
rect 10137 13883 10195 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10686 13920 10692 13932
rect 10275 13892 10692 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 8297 13855 8355 13861
rect 8297 13821 8309 13855
rect 8343 13852 8355 13855
rect 9401 13855 9459 13861
rect 8343 13824 9260 13852
rect 8343 13821 8355 13824
rect 8297 13815 8355 13821
rect 9232 13796 9260 13824
rect 9401 13821 9413 13855
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 6549 13787 6607 13793
rect 6549 13753 6561 13787
rect 6595 13753 6607 13787
rect 6549 13747 6607 13753
rect 9214 13744 9220 13796
rect 9272 13744 9278 13796
rect 9416 13784 9444 13815
rect 9582 13812 9588 13864
rect 9640 13852 9646 13864
rect 10152 13852 10180 13883
rect 10686 13880 10692 13892
rect 10744 13880 10750 13932
rect 10318 13852 10324 13864
rect 9640 13824 10180 13852
rect 10279 13824 10324 13852
rect 9640 13812 9646 13824
rect 10318 13812 10324 13824
rect 10376 13812 10382 13864
rect 11974 13812 11980 13864
rect 12032 13852 12038 13864
rect 19058 13852 19064 13864
rect 12032 13824 19064 13852
rect 12032 13812 12038 13824
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 9950 13784 9956 13796
rect 9416 13756 9956 13784
rect 9950 13744 9956 13756
rect 10008 13744 10014 13796
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3605 13719 3663 13725
rect 3605 13716 3617 13719
rect 3292 13688 3617 13716
rect 3292 13676 3298 13688
rect 3605 13685 3617 13688
rect 3651 13685 3663 13719
rect 3605 13679 3663 13685
rect 6917 13719 6975 13725
rect 6917 13685 6929 13719
rect 6963 13716 6975 13719
rect 7006 13716 7012 13728
rect 6963 13688 7012 13716
rect 6963 13685 6975 13688
rect 6917 13679 6975 13685
rect 7006 13676 7012 13688
rect 7064 13716 7070 13728
rect 7374 13716 7380 13728
rect 7064 13688 7380 13716
rect 7064 13676 7070 13688
rect 7374 13676 7380 13688
rect 7432 13676 7438 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2777 13515 2835 13521
rect 2777 13481 2789 13515
rect 2823 13512 2835 13515
rect 4154 13512 4160 13524
rect 2823 13484 4160 13512
rect 2823 13481 2835 13484
rect 2777 13475 2835 13481
rect 4154 13472 4160 13484
rect 4212 13472 4218 13524
rect 5534 13512 5540 13524
rect 5495 13484 5540 13512
rect 5534 13472 5540 13484
rect 5592 13472 5598 13524
rect 9950 13512 9956 13524
rect 9863 13484 9956 13512
rect 9950 13472 9956 13484
rect 10008 13512 10014 13524
rect 12250 13512 12256 13524
rect 10008 13484 11652 13512
rect 12211 13484 12256 13512
rect 10008 13472 10014 13484
rect 3786 13404 3792 13456
rect 3844 13444 3850 13456
rect 3881 13447 3939 13453
rect 3881 13444 3893 13447
rect 3844 13416 3893 13444
rect 3844 13404 3850 13416
rect 3881 13413 3893 13416
rect 3927 13444 3939 13447
rect 4430 13444 4436 13456
rect 3927 13416 4436 13444
rect 3927 13413 3939 13416
rect 3881 13407 3939 13413
rect 4430 13404 4436 13416
rect 4488 13404 4494 13456
rect 5258 13404 5264 13456
rect 5316 13444 5322 13456
rect 10226 13444 10232 13456
rect 5316 13416 10232 13444
rect 5316 13404 5322 13416
rect 10226 13404 10232 13416
rect 10284 13404 10290 13456
rect 4798 13376 4804 13388
rect 4759 13348 4804 13376
rect 4798 13336 4804 13348
rect 4856 13336 4862 13388
rect 5902 13336 5908 13388
rect 5960 13376 5966 13388
rect 5960 13348 7420 13376
rect 5960 13336 5966 13348
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13308 3479 13311
rect 5442 13308 5448 13320
rect 3467 13280 5448 13308
rect 3467 13277 3479 13280
rect 3421 13271 3479 13277
rect 5442 13268 5448 13280
rect 5500 13268 5506 13320
rect 7282 13308 7288 13320
rect 7243 13280 7288 13308
rect 7282 13268 7288 13280
rect 7340 13268 7346 13320
rect 7392 13308 7420 13348
rect 8018 13336 8024 13388
rect 8076 13376 8082 13388
rect 8297 13379 8355 13385
rect 8297 13376 8309 13379
rect 8076 13348 8309 13376
rect 8076 13336 8082 13348
rect 8297 13345 8309 13348
rect 8343 13345 8355 13379
rect 8297 13339 8355 13345
rect 8570 13336 8576 13388
rect 8628 13376 8634 13388
rect 8628 13348 10364 13376
rect 8628 13336 8634 13348
rect 8113 13311 8171 13317
rect 8113 13308 8125 13311
rect 7392 13280 8125 13308
rect 8113 13277 8125 13280
rect 8159 13308 8171 13311
rect 8754 13308 8760 13320
rect 8159 13280 8760 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 8754 13268 8760 13280
rect 8812 13268 8818 13320
rect 9033 13311 9091 13317
rect 9033 13277 9045 13311
rect 9079 13308 9091 13311
rect 9122 13308 9128 13320
rect 9079 13280 9128 13308
rect 9079 13277 9091 13280
rect 9033 13271 9091 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9674 13308 9680 13320
rect 9646 13268 9680 13308
rect 9732 13268 9738 13320
rect 7006 13240 7012 13252
rect 6967 13212 7012 13240
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 9646 13240 9674 13268
rect 7484 13212 9674 13240
rect 2222 13172 2228 13184
rect 2183 13144 2228 13172
rect 2222 13132 2228 13144
rect 2280 13132 2286 13184
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 4246 13172 4252 13184
rect 4203 13144 4252 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 4522 13172 4528 13184
rect 4483 13144 4528 13172
rect 4522 13132 4528 13144
rect 4580 13132 4586 13184
rect 4617 13175 4675 13181
rect 4617 13141 4629 13175
rect 4663 13172 4675 13175
rect 5166 13172 5172 13184
rect 4663 13144 5172 13172
rect 4663 13141 4675 13144
rect 4617 13135 4675 13141
rect 5166 13132 5172 13144
rect 5224 13132 5230 13184
rect 7484 13181 7512 13212
rect 7469 13175 7527 13181
rect 7469 13141 7481 13175
rect 7515 13141 7527 13175
rect 7469 13135 7527 13141
rect 7558 13132 7564 13184
rect 7616 13172 7622 13184
rect 7745 13175 7803 13181
rect 7745 13172 7757 13175
rect 7616 13144 7757 13172
rect 7616 13132 7622 13144
rect 7745 13141 7757 13144
rect 7791 13141 7803 13175
rect 7745 13135 7803 13141
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 9674 13172 9680 13184
rect 8260 13144 8305 13172
rect 9635 13144 9680 13172
rect 8260 13132 8266 13144
rect 9674 13132 9680 13144
rect 9732 13132 9738 13184
rect 10336 13172 10364 13348
rect 11238 13268 11244 13320
rect 11296 13308 11302 13320
rect 11624 13317 11652 13484
rect 12250 13472 12256 13484
rect 12308 13472 12314 13524
rect 11333 13311 11391 13317
rect 11333 13308 11345 13311
rect 11296 13280 11345 13308
rect 11296 13268 11302 13280
rect 11333 13277 11345 13280
rect 11379 13277 11391 13311
rect 11333 13271 11391 13277
rect 11609 13311 11667 13317
rect 11609 13277 11621 13311
rect 11655 13277 11667 13311
rect 11609 13271 11667 13277
rect 11088 13243 11146 13249
rect 11088 13209 11100 13243
rect 11134 13240 11146 13243
rect 12066 13240 12072 13252
rect 11134 13212 12072 13240
rect 11134 13209 11146 13212
rect 11088 13203 11146 13209
rect 12066 13200 12072 13212
rect 12124 13200 12130 13252
rect 15286 13172 15292 13184
rect 10336 13144 15292 13172
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 1486 12968 1492 12980
rect 1447 12940 1492 12968
rect 1486 12928 1492 12940
rect 1544 12928 1550 12980
rect 2225 12971 2283 12977
rect 2225 12937 2237 12971
rect 2271 12968 2283 12971
rect 4338 12968 4344 12980
rect 2271 12940 4344 12968
rect 2271 12937 2283 12940
rect 2225 12931 2283 12937
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4522 12928 4528 12980
rect 4580 12968 4586 12980
rect 5721 12971 5779 12977
rect 5721 12968 5733 12971
rect 4580 12940 5733 12968
rect 4580 12928 4586 12940
rect 5721 12937 5733 12940
rect 5767 12937 5779 12971
rect 5721 12931 5779 12937
rect 5810 12928 5816 12980
rect 5868 12968 5874 12980
rect 9858 12968 9864 12980
rect 5868 12940 8064 12968
rect 9819 12940 9864 12968
rect 5868 12928 5874 12940
rect 4614 12900 4620 12912
rect 2884 12872 4620 12900
rect 2884 12841 2912 12872
rect 4614 12860 4620 12872
rect 4672 12860 4678 12912
rect 5902 12860 5908 12912
rect 5960 12900 5966 12912
rect 6365 12903 6423 12909
rect 6365 12900 6377 12903
rect 5960 12872 6377 12900
rect 5960 12860 5966 12872
rect 6365 12869 6377 12872
rect 6411 12869 6423 12903
rect 6365 12863 6423 12869
rect 7006 12860 7012 12912
rect 7064 12900 7070 12912
rect 7837 12903 7895 12909
rect 7837 12900 7849 12903
rect 7064 12872 7849 12900
rect 7064 12860 7070 12872
rect 7837 12869 7849 12872
rect 7883 12869 7895 12903
rect 7837 12863 7895 12869
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12801 2927 12835
rect 2869 12795 2927 12801
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12801 3847 12835
rect 3789 12795 3847 12801
rect 1688 12764 1716 12795
rect 3142 12764 3148 12776
rect 1688 12736 3148 12764
rect 3142 12724 3148 12736
rect 3200 12724 3206 12776
rect 3804 12696 3832 12795
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 4065 12835 4123 12841
rect 4065 12832 4077 12835
rect 3936 12804 4077 12832
rect 3936 12792 3942 12804
rect 3988 12776 4016 12804
rect 4065 12801 4077 12804
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 4154 12792 4160 12844
rect 4212 12832 4218 12844
rect 4321 12835 4379 12841
rect 4321 12832 4333 12835
rect 4212 12804 4333 12832
rect 4212 12792 4218 12804
rect 4321 12801 4333 12804
rect 4367 12801 4379 12835
rect 4321 12795 4379 12801
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12832 7159 12835
rect 8036 12832 8064 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10226 12900 10232 12912
rect 10187 12872 10232 12900
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 10321 12903 10379 12909
rect 10321 12869 10333 12903
rect 10367 12900 10379 12903
rect 18874 12900 18880 12912
rect 10367 12872 18880 12900
rect 10367 12869 10379 12872
rect 10321 12863 10379 12869
rect 18874 12860 18880 12872
rect 18932 12860 18938 12912
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 7147 12804 7880 12832
rect 8036 12804 11897 12832
rect 7147 12801 7159 12804
rect 7101 12795 7159 12801
rect 3970 12724 3976 12776
rect 4028 12724 4034 12776
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7742 12764 7748 12776
rect 7055 12736 7748 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 4062 12696 4068 12708
rect 3804 12668 4068 12696
rect 4062 12656 4068 12668
rect 4120 12656 4126 12708
rect 5442 12696 5448 12708
rect 5403 12668 5448 12696
rect 5442 12656 5448 12668
rect 5500 12656 5506 12708
rect 6932 12696 6960 12727
rect 7742 12724 7748 12736
rect 7800 12724 7806 12776
rect 7852 12764 7880 12804
rect 11885 12801 11897 12804
rect 11931 12801 11943 12835
rect 11885 12795 11943 12801
rect 10410 12764 10416 12776
rect 7852 12736 9674 12764
rect 10371 12736 10416 12764
rect 8018 12696 8024 12708
rect 6932 12668 8024 12696
rect 8018 12656 8024 12668
rect 8076 12656 8082 12708
rect 3145 12631 3203 12637
rect 3145 12597 3157 12631
rect 3191 12628 3203 12631
rect 4430 12628 4436 12640
rect 3191 12600 4436 12628
rect 3191 12597 3203 12600
rect 3145 12591 3203 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 7466 12628 7472 12640
rect 7427 12600 7472 12628
rect 7466 12588 7472 12600
rect 7524 12588 7530 12640
rect 9214 12588 9220 12640
rect 9272 12628 9278 12640
rect 9309 12631 9367 12637
rect 9309 12628 9321 12631
rect 9272 12600 9321 12628
rect 9272 12588 9278 12600
rect 9309 12597 9321 12600
rect 9355 12597 9367 12631
rect 9646 12628 9674 12736
rect 10410 12724 10416 12736
rect 10468 12724 10474 12776
rect 10873 12767 10931 12773
rect 10873 12733 10885 12767
rect 10919 12733 10931 12767
rect 10873 12727 10931 12733
rect 10888 12628 10916 12727
rect 11514 12628 11520 12640
rect 9646 12600 10916 12628
rect 11475 12600 11520 12628
rect 9309 12591 9367 12597
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1854 12424 1860 12436
rect 1815 12396 1860 12424
rect 1854 12384 1860 12396
rect 1912 12384 1918 12436
rect 2038 12384 2044 12436
rect 2096 12424 2102 12436
rect 2133 12427 2191 12433
rect 2133 12424 2145 12427
rect 2096 12396 2145 12424
rect 2096 12384 2102 12396
rect 2133 12393 2145 12396
rect 2179 12393 2191 12427
rect 2133 12387 2191 12393
rect 2866 12384 2872 12436
rect 2924 12424 2930 12436
rect 3145 12427 3203 12433
rect 3145 12424 3157 12427
rect 2924 12396 3157 12424
rect 2924 12384 2930 12396
rect 3145 12393 3157 12396
rect 3191 12393 3203 12427
rect 3145 12387 3203 12393
rect 3881 12427 3939 12433
rect 3881 12393 3893 12427
rect 3927 12424 3939 12427
rect 4154 12424 4160 12436
rect 3927 12396 4160 12424
rect 3927 12393 3939 12396
rect 3881 12387 3939 12393
rect 4154 12384 4160 12396
rect 4212 12384 4218 12436
rect 4798 12424 4804 12436
rect 4759 12396 4804 12424
rect 4798 12384 4804 12396
rect 4856 12384 4862 12436
rect 8941 12427 8999 12433
rect 8941 12424 8953 12427
rect 4908 12396 8953 12424
rect 3050 12316 3056 12368
rect 3108 12356 3114 12368
rect 4908 12356 4936 12396
rect 8941 12393 8953 12396
rect 8987 12393 8999 12427
rect 8941 12387 8999 12393
rect 9769 12427 9827 12433
rect 9769 12393 9781 12427
rect 9815 12424 9827 12427
rect 10410 12424 10416 12436
rect 9815 12396 10416 12424
rect 9815 12393 9827 12396
rect 9769 12387 9827 12393
rect 10410 12384 10416 12396
rect 10468 12424 10474 12436
rect 12066 12424 12072 12436
rect 10468 12396 11468 12424
rect 12027 12396 12072 12424
rect 10468 12384 10474 12396
rect 3108 12328 4936 12356
rect 3108 12316 3114 12328
rect 9030 12316 9036 12368
rect 9088 12356 9094 12368
rect 9214 12356 9220 12368
rect 9088 12328 9220 12356
rect 9088 12316 9094 12328
rect 9214 12316 9220 12328
rect 9272 12316 9278 12368
rect 2774 12248 2780 12300
rect 2832 12288 2838 12300
rect 2832 12260 2877 12288
rect 2832 12248 2838 12260
rect 7742 12248 7748 12300
rect 7800 12288 7806 12300
rect 9582 12288 9588 12300
rect 7800 12260 9588 12288
rect 7800 12248 7806 12260
rect 9582 12248 9588 12260
rect 9640 12248 9646 12300
rect 1673 12223 1731 12229
rect 1673 12189 1685 12223
rect 1719 12220 1731 12223
rect 1854 12220 1860 12232
rect 1719 12192 1860 12220
rect 1719 12189 1731 12192
rect 1673 12183 1731 12189
rect 1854 12180 1860 12192
rect 1912 12180 1918 12232
rect 3329 12223 3387 12229
rect 3329 12189 3341 12223
rect 3375 12220 3387 12223
rect 3878 12220 3884 12232
rect 3375 12192 3884 12220
rect 3375 12189 3387 12192
rect 3329 12183 3387 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12220 4583 12223
rect 4798 12220 4804 12232
rect 4571 12192 4804 12220
rect 4571 12189 4583 12192
rect 4525 12183 4583 12189
rect 4798 12180 4804 12192
rect 4856 12180 4862 12232
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 6181 12223 6239 12229
rect 6181 12220 6193 12223
rect 5592 12192 6193 12220
rect 5592 12180 5598 12192
rect 6181 12189 6193 12192
rect 6227 12220 6239 12223
rect 6638 12220 6644 12232
rect 6227 12192 6644 12220
rect 6227 12189 6239 12192
rect 6181 12183 6239 12189
rect 6638 12180 6644 12192
rect 6696 12180 6702 12232
rect 6914 12229 6920 12232
rect 6908 12220 6920 12229
rect 6875 12192 6920 12220
rect 6908 12183 6920 12192
rect 6914 12180 6920 12183
rect 6972 12180 6978 12232
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 10410 12220 10416 12232
rect 7892 12192 10416 12220
rect 7892 12180 7898 12192
rect 10410 12180 10416 12192
rect 10468 12180 10474 12232
rect 11054 12180 11060 12232
rect 11112 12220 11118 12232
rect 11440 12229 11468 12396
rect 12066 12384 12072 12396
rect 12124 12384 12130 12436
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 11112 12192 11161 12220
rect 11112 12180 11118 12192
rect 11149 12189 11161 12192
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 11425 12223 11483 12229
rect 11425 12189 11437 12223
rect 11471 12189 11483 12223
rect 19702 12220 19708 12232
rect 19663 12192 19708 12220
rect 11425 12183 11483 12189
rect 19702 12180 19708 12192
rect 19760 12180 19766 12232
rect 2314 12112 2320 12164
rect 2372 12152 2378 12164
rect 5718 12152 5724 12164
rect 2372 12124 5724 12152
rect 2372 12112 2378 12124
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 5902 12152 5908 12164
rect 5960 12161 5966 12164
rect 5872 12124 5908 12152
rect 5902 12112 5908 12124
rect 5960 12115 5972 12161
rect 5960 12112 5966 12115
rect 7098 12112 7104 12164
rect 7156 12152 7162 12164
rect 8389 12155 8447 12161
rect 8389 12152 8401 12155
rect 7156 12124 8401 12152
rect 7156 12112 7162 12124
rect 8389 12121 8401 12124
rect 8435 12121 8447 12155
rect 8389 12115 8447 12121
rect 8662 12112 8668 12164
rect 8720 12152 8726 12164
rect 10904 12155 10962 12161
rect 8720 12124 9628 12152
rect 8720 12112 8726 12124
rect 2498 12084 2504 12096
rect 2459 12056 2504 12084
rect 2498 12044 2504 12056
rect 2556 12044 2562 12096
rect 2590 12044 2596 12096
rect 2648 12084 2654 12096
rect 2648 12056 2693 12084
rect 2648 12044 2654 12056
rect 4062 12044 4068 12096
rect 4120 12084 4126 12096
rect 5994 12084 6000 12096
rect 4120 12056 6000 12084
rect 4120 12044 4126 12056
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6914 12044 6920 12096
rect 6972 12084 6978 12096
rect 7742 12084 7748 12096
rect 6972 12056 7748 12084
rect 6972 12044 6978 12056
rect 7742 12044 7748 12056
rect 7800 12044 7806 12096
rect 8018 12084 8024 12096
rect 7979 12056 8024 12084
rect 8018 12044 8024 12056
rect 8076 12044 8082 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 9306 12084 9312 12096
rect 8628 12056 9312 12084
rect 8628 12044 8634 12056
rect 9306 12044 9312 12056
rect 9364 12044 9370 12096
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9600 12084 9628 12124
rect 10904 12121 10916 12155
rect 10950 12152 10962 12155
rect 12158 12152 12164 12164
rect 10950 12124 12164 12152
rect 10950 12121 10962 12124
rect 10904 12115 10962 12121
rect 12158 12112 12164 12124
rect 12216 12112 12222 12164
rect 12713 12155 12771 12161
rect 12713 12152 12725 12155
rect 12268 12124 12725 12152
rect 10226 12084 10232 12096
rect 9600 12056 10232 12084
rect 10226 12044 10232 12056
rect 10284 12084 10290 12096
rect 12268 12084 12296 12124
rect 12713 12121 12725 12124
rect 12759 12121 12771 12155
rect 12713 12115 12771 12121
rect 10284 12056 12296 12084
rect 12437 12087 12495 12093
rect 10284 12044 10290 12056
rect 12437 12053 12449 12087
rect 12483 12084 12495 12087
rect 12986 12084 12992 12096
rect 12483 12056 12992 12084
rect 12483 12053 12495 12056
rect 12437 12047 12495 12053
rect 12986 12044 12992 12056
rect 13044 12044 13050 12096
rect 13173 12087 13231 12093
rect 13173 12053 13185 12087
rect 13219 12084 13231 12087
rect 13446 12084 13452 12096
rect 13219 12056 13452 12084
rect 13219 12053 13231 12056
rect 13173 12047 13231 12053
rect 13446 12044 13452 12056
rect 13504 12044 13510 12096
rect 19889 12087 19947 12093
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 20530 12084 20536 12096
rect 19935 12056 20536 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 1670 11880 1676 11892
rect 1631 11852 1676 11880
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 2498 11840 2504 11892
rect 2556 11880 2562 11892
rect 2685 11883 2743 11889
rect 2685 11880 2697 11883
rect 2556 11852 2697 11880
rect 2556 11840 2562 11852
rect 2685 11849 2697 11852
rect 2731 11849 2743 11883
rect 2685 11843 2743 11849
rect 2884 11852 4108 11880
rect 2225 11815 2283 11821
rect 2225 11781 2237 11815
rect 2271 11812 2283 11815
rect 2884 11812 2912 11852
rect 3970 11812 3976 11824
rect 2271 11784 2912 11812
rect 2976 11784 3976 11812
rect 2271 11781 2283 11784
rect 2225 11775 2283 11781
rect 1489 11747 1547 11753
rect 1489 11713 1501 11747
rect 1535 11744 1547 11747
rect 1578 11744 1584 11756
rect 1535 11716 1584 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1578 11704 1584 11716
rect 1636 11704 1642 11756
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11744 2375 11747
rect 2866 11744 2872 11756
rect 2363 11716 2872 11744
rect 2363 11713 2375 11716
rect 2317 11707 2375 11713
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 2976 11753 3004 11784
rect 3970 11772 3976 11784
rect 4028 11772 4034 11824
rect 4080 11812 4108 11852
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 4341 11883 4399 11889
rect 4341 11880 4353 11883
rect 4304 11852 4353 11880
rect 4304 11840 4310 11852
rect 4341 11849 4353 11852
rect 4387 11880 4399 11883
rect 4614 11880 4620 11892
rect 4387 11852 4620 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 4614 11840 4620 11852
rect 4672 11840 4678 11892
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 4856 11852 4901 11880
rect 5184 11852 5580 11880
rect 4856 11840 4862 11852
rect 4522 11812 4528 11824
rect 4080 11784 4528 11812
rect 4522 11772 4528 11784
rect 4580 11812 4586 11824
rect 4580 11784 4752 11812
rect 4580 11772 4586 11784
rect 3234 11753 3240 11756
rect 2961 11747 3019 11753
rect 2961 11713 2973 11747
rect 3007 11713 3019 11747
rect 3228 11744 3240 11753
rect 3195 11716 3240 11744
rect 2961 11707 3019 11713
rect 3228 11707 3240 11716
rect 3234 11704 3240 11707
rect 3292 11704 3298 11756
rect 4062 11704 4068 11756
rect 4120 11744 4126 11756
rect 4617 11747 4675 11753
rect 4617 11744 4629 11747
rect 4120 11716 4629 11744
rect 4120 11704 4126 11716
rect 4617 11713 4629 11716
rect 4663 11713 4675 11747
rect 4724 11744 4752 11784
rect 5184 11744 5212 11852
rect 4724 11716 5212 11744
rect 4617 11707 4675 11713
rect 5258 11704 5264 11756
rect 5316 11744 5322 11756
rect 5445 11747 5503 11753
rect 5445 11744 5457 11747
rect 5316 11716 5457 11744
rect 5316 11704 5322 11716
rect 5445 11713 5457 11716
rect 5491 11713 5503 11747
rect 5552 11744 5580 11852
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6733 11883 6791 11889
rect 6733 11880 6745 11883
rect 5776 11852 6745 11880
rect 5776 11840 5782 11852
rect 6733 11849 6745 11852
rect 6779 11849 6791 11883
rect 6733 11843 6791 11849
rect 7101 11883 7159 11889
rect 7101 11849 7113 11883
rect 7147 11880 7159 11883
rect 7466 11880 7472 11892
rect 7147 11852 7472 11880
rect 7147 11849 7159 11852
rect 7101 11843 7159 11849
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 12158 11880 12164 11892
rect 7852 11852 11744 11880
rect 12119 11852 12164 11880
rect 5994 11772 6000 11824
rect 6052 11812 6058 11824
rect 6365 11815 6423 11821
rect 6365 11812 6377 11815
rect 6052 11784 6377 11812
rect 6052 11772 6058 11784
rect 6365 11781 6377 11784
rect 6411 11781 6423 11815
rect 6365 11775 6423 11781
rect 6638 11772 6644 11824
rect 6696 11812 6702 11824
rect 6696 11784 7788 11812
rect 6696 11772 6702 11784
rect 6914 11744 6920 11756
rect 5552 11716 6920 11744
rect 5445 11707 5503 11713
rect 6914 11704 6920 11716
rect 6972 11704 6978 11756
rect 7193 11747 7251 11753
rect 7193 11713 7205 11747
rect 7239 11744 7251 11747
rect 7558 11744 7564 11756
rect 7239 11716 7564 11744
rect 7239 11713 7251 11716
rect 7193 11707 7251 11713
rect 7558 11704 7564 11716
rect 7616 11704 7622 11756
rect 7760 11753 7788 11784
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 1946 11636 1952 11688
rect 2004 11676 2010 11688
rect 2041 11679 2099 11685
rect 2041 11676 2053 11679
rect 2004 11648 2053 11676
rect 2004 11636 2010 11648
rect 2041 11645 2053 11648
rect 2087 11645 2099 11679
rect 2041 11639 2099 11645
rect 2148 11648 2774 11676
rect 2038 11500 2044 11552
rect 2096 11540 2102 11552
rect 2148 11540 2176 11648
rect 2096 11512 2176 11540
rect 2746 11540 2774 11648
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 5537 11679 5595 11685
rect 5537 11676 5549 11679
rect 5408 11648 5549 11676
rect 5408 11636 5414 11648
rect 5537 11645 5549 11648
rect 5583 11645 5595 11679
rect 5537 11639 5595 11645
rect 5629 11679 5687 11685
rect 5629 11645 5641 11679
rect 5675 11645 5687 11679
rect 7374 11676 7380 11688
rect 7335 11648 7380 11676
rect 5629 11639 5687 11645
rect 4706 11568 4712 11620
rect 4764 11608 4770 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4764 11580 5089 11608
rect 4764 11568 4770 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 5644 11608 5672 11639
rect 7374 11636 7380 11648
rect 7432 11636 7438 11688
rect 7852 11676 7880 11852
rect 9674 11821 9680 11824
rect 9668 11812 9680 11821
rect 9140 11784 9536 11812
rect 9635 11784 9680 11812
rect 8012 11747 8070 11753
rect 8012 11713 8024 11747
rect 8058 11744 8070 11747
rect 9140 11744 9168 11784
rect 8058 11716 9168 11744
rect 9401 11747 9459 11753
rect 8058 11713 8070 11716
rect 8012 11707 8070 11713
rect 9401 11713 9413 11747
rect 9447 11713 9459 11747
rect 9508 11744 9536 11784
rect 9668 11775 9680 11784
rect 9674 11772 9680 11775
rect 9732 11772 9738 11824
rect 11716 11812 11744 11852
rect 12158 11840 12164 11852
rect 12216 11840 12222 11892
rect 12434 11880 12440 11892
rect 12395 11852 12440 11880
rect 12434 11840 12440 11852
rect 12492 11840 12498 11892
rect 13633 11815 13691 11821
rect 13633 11812 13645 11815
rect 11716 11784 13645 11812
rect 13633 11781 13645 11784
rect 13679 11781 13691 11815
rect 13633 11775 13691 11781
rect 10594 11744 10600 11756
rect 9508 11716 10600 11744
rect 9401 11707 9459 11713
rect 9306 11676 9312 11688
rect 7484 11648 7880 11676
rect 8956 11648 9312 11676
rect 7484 11608 7512 11648
rect 5500 11580 5672 11608
rect 5736 11580 7512 11608
rect 5500 11568 5506 11580
rect 5736 11540 5764 11580
rect 2746 11512 5764 11540
rect 2096 11500 2102 11512
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 8956 11540 8984 11648
rect 9306 11636 9312 11648
rect 9364 11636 9370 11688
rect 9030 11568 9036 11620
rect 9088 11608 9094 11620
rect 9416 11608 9444 11707
rect 10594 11704 10600 11716
rect 10652 11704 10658 11756
rect 11517 11747 11575 11753
rect 11517 11744 11529 11747
rect 10796 11716 11529 11744
rect 9088 11580 9444 11608
rect 9088 11568 9094 11580
rect 10796 11552 10824 11716
rect 11517 11713 11529 11716
rect 11563 11713 11575 11747
rect 12618 11744 12624 11756
rect 12579 11716 12624 11744
rect 11517 11707 11575 11713
rect 12618 11704 12624 11716
rect 12676 11744 12682 11756
rect 12897 11747 12955 11753
rect 12897 11744 12909 11747
rect 12676 11716 12909 11744
rect 12676 11704 12682 11716
rect 12897 11713 12909 11716
rect 12943 11713 12955 11747
rect 19242 11744 19248 11756
rect 19203 11716 19248 11744
rect 12897 11707 12955 11713
rect 19242 11704 19248 11716
rect 19300 11744 19306 11756
rect 19705 11747 19763 11753
rect 19705 11744 19717 11747
rect 19300 11716 19717 11744
rect 19300 11704 19306 11716
rect 19705 11713 19717 11716
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 9122 11540 9128 11552
rect 6696 11512 8984 11540
rect 9083 11512 9128 11540
rect 6696 11500 6702 11512
rect 9122 11500 9128 11512
rect 9180 11500 9186 11552
rect 10778 11540 10784 11552
rect 10739 11512 10784 11540
rect 10778 11500 10784 11512
rect 10836 11500 10842 11552
rect 11054 11540 11060 11552
rect 11015 11512 11060 11540
rect 11054 11500 11060 11512
rect 11112 11500 11118 11552
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 14093 11543 14151 11549
rect 14093 11509 14105 11543
rect 14139 11540 14151 11543
rect 14274 11540 14280 11552
rect 14139 11512 14280 11540
rect 14139 11509 14151 11512
rect 14093 11503 14151 11509
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 19429 11543 19487 11549
rect 19429 11509 19441 11543
rect 19475 11540 19487 11543
rect 20162 11540 20168 11552
rect 19475 11512 20168 11540
rect 19475 11509 19487 11512
rect 19429 11503 19487 11509
rect 20162 11500 20168 11512
rect 20220 11500 20226 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1578 11336 1584 11348
rect 1539 11308 1584 11336
rect 1578 11296 1584 11308
rect 1636 11296 1642 11348
rect 2774 11296 2780 11348
rect 2832 11336 2838 11348
rect 3237 11339 3295 11345
rect 3237 11336 3249 11339
rect 2832 11308 3249 11336
rect 2832 11296 2838 11308
rect 3237 11305 3249 11308
rect 3283 11305 3295 11339
rect 3237 11299 3295 11305
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 7190 11336 7196 11348
rect 3476 11308 7196 11336
rect 3476 11296 3482 11308
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 8478 11296 8484 11348
rect 8536 11336 8542 11348
rect 9309 11339 9367 11345
rect 9309 11336 9321 11339
rect 8536 11308 9321 11336
rect 8536 11296 8542 11308
rect 9309 11305 9321 11308
rect 9355 11305 9367 11339
rect 9309 11299 9367 11305
rect 10594 11296 10600 11348
rect 10652 11336 10658 11348
rect 11885 11339 11943 11345
rect 11885 11336 11897 11339
rect 10652 11308 11897 11336
rect 10652 11296 10658 11308
rect 11885 11305 11897 11308
rect 11931 11305 11943 11339
rect 11885 11299 11943 11305
rect 8662 11228 8668 11280
rect 8720 11268 8726 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 8720 11240 8953 11268
rect 8720 11228 8726 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 9030 11228 9036 11280
rect 9088 11268 9094 11280
rect 10965 11271 11023 11277
rect 10965 11268 10977 11271
rect 9088 11240 10977 11268
rect 9088 11228 9094 11240
rect 10965 11237 10977 11240
rect 11011 11237 11023 11271
rect 10965 11231 11023 11237
rect 13265 11271 13323 11277
rect 13265 11237 13277 11271
rect 13311 11268 13323 11271
rect 15838 11268 15844 11280
rect 13311 11240 15844 11268
rect 13311 11237 13323 11240
rect 13265 11231 13323 11237
rect 15838 11228 15844 11240
rect 15896 11228 15902 11280
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 19610 11268 19616 11280
rect 19475 11240 19616 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 19610 11228 19616 11240
rect 19668 11228 19674 11280
rect 2866 11160 2872 11212
rect 2924 11200 2930 11212
rect 3789 11203 3847 11209
rect 3789 11200 3801 11203
rect 2924 11172 3801 11200
rect 2924 11160 2930 11172
rect 3789 11169 3801 11172
rect 3835 11169 3847 11203
rect 3789 11163 3847 11169
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 9953 11203 10011 11209
rect 8076 11172 9015 11200
rect 8076 11160 8082 11172
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 1397 11095 1455 11101
rect 1412 11064 1440 11095
rect 1762 11092 1768 11144
rect 1820 11132 1826 11144
rect 1857 11135 1915 11141
rect 1857 11132 1869 11135
rect 1820 11104 1869 11132
rect 1820 11092 1826 11104
rect 1857 11101 1869 11104
rect 1903 11101 1915 11135
rect 1857 11095 1915 11101
rect 1946 11092 1952 11144
rect 2004 11132 2010 11144
rect 2113 11135 2171 11141
rect 2113 11132 2125 11135
rect 2004 11104 2125 11132
rect 2004 11092 2010 11104
rect 2113 11101 2125 11104
rect 2159 11132 2171 11135
rect 3050 11132 3056 11144
rect 2159 11104 3056 11132
rect 2159 11101 2171 11104
rect 2113 11095 2171 11101
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 3234 11092 3240 11144
rect 3292 11132 3298 11144
rect 4062 11132 4068 11144
rect 3292 11104 4068 11132
rect 3292 11092 3298 11104
rect 4062 11092 4068 11104
rect 4120 11132 4126 11144
rect 4249 11135 4307 11141
rect 4249 11132 4261 11135
rect 4120 11104 4261 11132
rect 4120 11092 4126 11104
rect 4249 11101 4261 11104
rect 4295 11101 4307 11135
rect 4614 11132 4620 11144
rect 4575 11104 4620 11132
rect 4249 11095 4307 11101
rect 4614 11092 4620 11104
rect 4672 11092 4678 11144
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 6638 11132 6644 11144
rect 4764 11104 6644 11132
rect 4764 11092 4770 11104
rect 6638 11092 6644 11104
rect 6696 11092 6702 11144
rect 6733 11135 6791 11141
rect 6733 11101 6745 11135
rect 6779 11101 6791 11135
rect 6733 11095 6791 11101
rect 3970 11064 3976 11076
rect 1412 11036 3976 11064
rect 3970 11024 3976 11036
rect 4028 11024 4034 11076
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 4862 11067 4920 11073
rect 4862 11064 4874 11067
rect 4488 11036 4874 11064
rect 4488 11024 4494 11036
rect 4862 11033 4874 11036
rect 4908 11033 4920 11067
rect 6454 11064 6460 11076
rect 4862 11027 4920 11033
rect 5828 11036 6460 11064
rect 3418 10956 3424 11008
rect 3476 10996 3482 11008
rect 5828 10996 5856 11036
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 6748 11064 6776 11095
rect 6822 11092 6828 11144
rect 6880 11132 6886 11144
rect 7009 11135 7067 11141
rect 7009 11132 7021 11135
rect 6880 11104 7021 11132
rect 6880 11092 6886 11104
rect 7009 11101 7021 11104
rect 7055 11101 7067 11135
rect 7009 11095 7067 11101
rect 7276 11135 7334 11141
rect 7276 11101 7288 11135
rect 7322 11132 7334 11135
rect 8846 11132 8852 11144
rect 7322 11104 8852 11132
rect 7322 11101 7334 11104
rect 7276 11095 7334 11101
rect 8846 11092 8852 11104
rect 8904 11092 8910 11144
rect 8987 11132 9015 11172
rect 9140 11172 9812 11200
rect 9140 11132 9168 11172
rect 8987 11104 9168 11132
rect 9490 11092 9496 11144
rect 9548 11132 9554 11144
rect 9677 11135 9735 11141
rect 9677 11132 9689 11135
rect 9548 11104 9689 11132
rect 9548 11092 9554 11104
rect 9677 11101 9689 11104
rect 9723 11101 9735 11135
rect 9784 11132 9812 11172
rect 9953 11169 9965 11203
rect 9999 11200 10011 11203
rect 10778 11200 10784 11212
rect 9999 11172 10784 11200
rect 9999 11169 10011 11172
rect 9953 11163 10011 11169
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 14826 11200 14832 11212
rect 10888 11172 14136 11200
rect 14787 11172 14832 11200
rect 10321 11135 10379 11141
rect 10321 11132 10333 11135
rect 9784 11104 10333 11132
rect 9677 11095 9735 11101
rect 10321 11101 10333 11104
rect 10367 11101 10379 11135
rect 10321 11095 10379 11101
rect 10410 11092 10416 11144
rect 10468 11132 10474 11144
rect 10888 11132 10916 11172
rect 10468 11104 10916 11132
rect 11241 11135 11299 11141
rect 10468 11092 10474 11104
rect 11241 11101 11253 11135
rect 11287 11101 11299 11135
rect 12158 11132 12164 11144
rect 12119 11104 12164 11132
rect 11241 11095 11299 11101
rect 8202 11064 8208 11076
rect 6748 11036 8208 11064
rect 8202 11024 8208 11036
rect 8260 11024 8266 11076
rect 8404 11036 9076 11064
rect 8404 11008 8432 11036
rect 5994 10996 6000 11008
rect 3476 10968 5856 10996
rect 5955 10968 6000 10996
rect 3476 10956 3482 10968
rect 5994 10956 6000 10968
rect 6052 10956 6058 11008
rect 6546 10996 6552 11008
rect 6507 10968 6552 10996
rect 6546 10956 6552 10968
rect 6604 10956 6610 11008
rect 8386 10996 8392 11008
rect 8299 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 9048 10996 9076 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 9769 11067 9827 11073
rect 9769 11064 9781 11067
rect 9456 11036 9781 11064
rect 9456 11024 9462 11036
rect 9769 11033 9781 11036
rect 9815 11033 9827 11067
rect 11256 11064 11284 11095
rect 12158 11092 12164 11104
rect 12216 11092 12222 11144
rect 12250 11092 12256 11144
rect 12308 11132 12314 11144
rect 13081 11135 13139 11141
rect 13081 11132 13093 11135
rect 12308 11104 13093 11132
rect 12308 11092 12314 11104
rect 13081 11101 13093 11104
rect 13127 11132 13139 11135
rect 13541 11135 13599 11141
rect 13541 11132 13553 11135
rect 13127 11104 13553 11132
rect 13127 11101 13139 11104
rect 13081 11095 13139 11101
rect 13541 11101 13553 11104
rect 13587 11101 13599 11135
rect 14108 11132 14136 11172
rect 14826 11160 14832 11172
rect 14884 11160 14890 11212
rect 15194 11132 15200 11144
rect 14108 11104 15200 11132
rect 13541 11095 13599 11101
rect 15194 11092 15200 11104
rect 15252 11092 15258 11144
rect 15286 11092 15292 11144
rect 15344 11132 15350 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 15344 11104 19257 11132
rect 15344 11092 15350 11104
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 9769 11027 9827 11033
rect 9876 11036 11284 11064
rect 9876 10996 9904 11036
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12805 11067 12863 11073
rect 12805 11064 12817 11067
rect 12124 11036 12817 11064
rect 12124 11024 12130 11036
rect 12805 11033 12817 11036
rect 12851 11033 12863 11067
rect 12805 11027 12863 11033
rect 13722 11024 13728 11076
rect 13780 11064 13786 11076
rect 14093 11067 14151 11073
rect 14093 11064 14105 11067
rect 13780 11036 14105 11064
rect 13780 11024 13786 11036
rect 14093 11033 14105 11036
rect 14139 11033 14151 11067
rect 14458 11064 14464 11076
rect 14419 11036 14464 11064
rect 14093 11027 14151 11033
rect 14458 11024 14464 11036
rect 14516 11024 14522 11076
rect 9048 10968 9904 10996
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 3050 10792 3056 10804
rect 3011 10764 3056 10792
rect 3050 10752 3056 10764
rect 3108 10752 3114 10804
rect 3142 10752 3148 10804
rect 3200 10792 3206 10804
rect 3329 10795 3387 10801
rect 3329 10792 3341 10795
rect 3200 10764 3341 10792
rect 3200 10752 3206 10764
rect 3329 10761 3341 10764
rect 3375 10761 3387 10795
rect 3329 10755 3387 10761
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4706 10792 4712 10804
rect 4212 10764 4712 10792
rect 4212 10752 4218 10764
rect 4706 10752 4712 10764
rect 4764 10792 4770 10804
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 4764 10764 5457 10792
rect 4764 10752 4770 10764
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 6733 10795 6791 10801
rect 6733 10792 6745 10795
rect 5684 10764 6745 10792
rect 5684 10752 5690 10764
rect 6733 10761 6745 10764
rect 6779 10761 6791 10795
rect 7098 10792 7104 10804
rect 7059 10764 7104 10792
rect 6733 10755 6791 10761
rect 7098 10752 7104 10764
rect 7156 10752 7162 10804
rect 8202 10792 8208 10804
rect 8163 10764 8208 10792
rect 8202 10752 8208 10764
rect 8260 10752 8266 10804
rect 9398 10792 9404 10804
rect 9359 10764 9404 10792
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 15013 10795 15071 10801
rect 15013 10792 15025 10795
rect 13872 10764 15025 10792
rect 13872 10752 13878 10764
rect 15013 10761 15025 10764
rect 15059 10761 15071 10795
rect 15013 10755 15071 10761
rect 1762 10724 1768 10736
rect 1675 10696 1768 10724
rect 1688 10665 1716 10696
rect 1762 10684 1768 10696
rect 1820 10724 1826 10736
rect 4614 10724 4620 10736
rect 1820 10696 4620 10724
rect 1820 10684 1826 10696
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10625 1731 10659
rect 1673 10619 1731 10625
rect 1940 10659 1998 10665
rect 1940 10625 1952 10659
rect 1986 10656 1998 10659
rect 2222 10656 2228 10668
rect 1986 10628 2228 10656
rect 1986 10625 1998 10628
rect 1940 10619 1998 10625
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 4080 10665 4108 10696
rect 4614 10684 4620 10696
rect 4672 10724 4678 10736
rect 4798 10724 4804 10736
rect 4672 10696 4804 10724
rect 4672 10684 4678 10696
rect 4798 10684 4804 10696
rect 4856 10684 4862 10736
rect 6457 10727 6515 10733
rect 6457 10693 6469 10727
rect 6503 10724 6515 10727
rect 6638 10724 6644 10736
rect 6503 10696 6644 10724
rect 6503 10693 6515 10696
rect 6457 10687 6515 10693
rect 6638 10684 6644 10696
rect 6696 10684 6702 10736
rect 8573 10727 8631 10733
rect 8573 10724 8585 10727
rect 6748 10696 8585 10724
rect 6748 10668 6776 10696
rect 8573 10693 8585 10696
rect 8619 10693 8631 10727
rect 8573 10687 8631 10693
rect 9861 10727 9919 10733
rect 9861 10693 9873 10727
rect 9907 10724 9919 10727
rect 13449 10727 13507 10733
rect 9907 10696 12434 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 4338 10665 4344 10668
rect 3513 10659 3571 10665
rect 3513 10625 3525 10659
rect 3559 10656 3571 10659
rect 4065 10659 4123 10665
rect 3559 10628 4016 10656
rect 3559 10625 3571 10628
rect 3513 10619 3571 10625
rect 3988 10452 4016 10628
rect 4065 10625 4077 10659
rect 4111 10625 4123 10659
rect 4332 10656 4344 10665
rect 4299 10628 4344 10656
rect 4065 10619 4123 10625
rect 4332 10619 4344 10628
rect 4338 10616 4344 10619
rect 4396 10616 4402 10668
rect 6730 10616 6736 10668
rect 6788 10616 6794 10668
rect 7742 10656 7748 10668
rect 7703 10628 7748 10656
rect 7742 10616 7748 10628
rect 7800 10616 7806 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9732 10628 9781 10656
rect 9732 10616 9738 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 9769 10619 9827 10625
rect 10413 10659 10471 10665
rect 10413 10625 10425 10659
rect 10459 10625 10471 10659
rect 10413 10619 10471 10625
rect 5074 10548 5080 10600
rect 5132 10588 5138 10600
rect 5721 10591 5779 10597
rect 5721 10588 5733 10591
rect 5132 10560 5733 10588
rect 5132 10548 5138 10560
rect 5721 10557 5733 10560
rect 5767 10557 5779 10591
rect 7190 10588 7196 10600
rect 7151 10560 7196 10588
rect 5721 10551 5779 10557
rect 7190 10548 7196 10560
rect 7248 10548 7254 10600
rect 7377 10591 7435 10597
rect 7377 10557 7389 10591
rect 7423 10588 7435 10591
rect 8386 10588 8392 10600
rect 7423 10560 8392 10588
rect 7423 10557 7435 10560
rect 7377 10551 7435 10557
rect 8386 10548 8392 10560
rect 8444 10548 8450 10600
rect 8662 10588 8668 10600
rect 8623 10560 8668 10588
rect 8662 10548 8668 10560
rect 8720 10548 8726 10600
rect 8757 10591 8815 10597
rect 8757 10557 8769 10591
rect 8803 10557 8815 10591
rect 8757 10551 8815 10557
rect 6546 10520 6552 10532
rect 5000 10492 6552 10520
rect 5000 10452 5028 10492
rect 6546 10480 6552 10492
rect 6604 10480 6610 10532
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 8772 10520 8800 10551
rect 9122 10548 9128 10600
rect 9180 10588 9186 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9180 10560 9965 10588
rect 9180 10548 9186 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 8536 10492 8800 10520
rect 8536 10480 8542 10492
rect 9582 10480 9588 10532
rect 9640 10520 9646 10532
rect 10428 10520 10456 10619
rect 11698 10588 11704 10600
rect 11659 10560 11704 10588
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 12406 10588 12434 10696
rect 13449 10693 13461 10727
rect 13495 10724 13507 10727
rect 17954 10724 17960 10736
rect 13495 10696 17960 10724
rect 13495 10693 13507 10696
rect 13449 10687 13507 10693
rect 17954 10684 17960 10696
rect 18012 10684 18018 10736
rect 12802 10616 12808 10668
rect 12860 10656 12866 10668
rect 13722 10656 13728 10668
rect 12860 10628 13728 10656
rect 12860 10616 12866 10628
rect 13722 10616 13728 10628
rect 13780 10616 13786 10668
rect 14366 10656 14372 10668
rect 14327 10628 14372 10656
rect 14366 10616 14372 10628
rect 14424 10656 14430 10668
rect 14645 10659 14703 10665
rect 14645 10656 14657 10659
rect 14424 10628 14657 10656
rect 14424 10616 14430 10628
rect 14645 10625 14657 10628
rect 14691 10625 14703 10659
rect 18322 10656 18328 10668
rect 18283 10628 18328 10656
rect 14645 10619 14703 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 16114 10588 16120 10600
rect 12406 10560 16120 10588
rect 16114 10548 16120 10560
rect 16172 10548 16178 10600
rect 9640 10492 10456 10520
rect 13909 10523 13967 10529
rect 9640 10480 9646 10492
rect 13909 10489 13921 10523
rect 13955 10520 13967 10523
rect 14642 10520 14648 10532
rect 13955 10492 14648 10520
rect 13955 10489 13967 10492
rect 13909 10483 13967 10489
rect 14642 10480 14648 10492
rect 14700 10480 14706 10532
rect 15746 10520 15752 10532
rect 15707 10492 15752 10520
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 7926 10452 7932 10464
rect 3988 10424 5028 10452
rect 7887 10424 7932 10452
rect 7926 10412 7932 10424
rect 7984 10412 7990 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 11057 10455 11115 10461
rect 11057 10452 11069 10455
rect 8352 10424 11069 10452
rect 8352 10412 8358 10424
rect 11057 10421 11069 10424
rect 11103 10421 11115 10455
rect 11057 10415 11115 10421
rect 11330 10412 11336 10464
rect 11388 10452 11394 10464
rect 11790 10452 11796 10464
rect 11388 10424 11796 10452
rect 11388 10412 11394 10424
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 13170 10412 13176 10464
rect 13228 10452 13234 10464
rect 14185 10455 14243 10461
rect 14185 10452 14197 10455
rect 13228 10424 14197 10452
rect 13228 10412 13234 10424
rect 14185 10421 14197 10424
rect 14231 10421 14243 10455
rect 15378 10452 15384 10464
rect 15339 10424 15384 10452
rect 14185 10415 14243 10421
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 18509 10455 18567 10461
rect 18509 10421 18521 10455
rect 18555 10452 18567 10455
rect 20070 10452 20076 10464
rect 18555 10424 20076 10452
rect 18555 10421 18567 10424
rect 18509 10415 18567 10421
rect 20070 10412 20076 10424
rect 20128 10412 20134 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 2590 10248 2596 10260
rect 2551 10220 2596 10248
rect 2590 10208 2596 10220
rect 2648 10208 2654 10260
rect 3326 10208 3332 10260
rect 3384 10248 3390 10260
rect 4982 10248 4988 10260
rect 3384 10220 4988 10248
rect 3384 10208 3390 10220
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5166 10248 5172 10260
rect 5127 10220 5172 10248
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5276 10220 11192 10248
rect 2317 10183 2375 10189
rect 2317 10149 2329 10183
rect 2363 10149 2375 10183
rect 2317 10143 2375 10149
rect 1765 10115 1823 10121
rect 1765 10081 1777 10115
rect 1811 10112 1823 10115
rect 1854 10112 1860 10124
rect 1811 10084 1860 10112
rect 1811 10081 1823 10084
rect 1765 10075 1823 10081
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 2332 10044 2360 10143
rect 2682 10140 2688 10192
rect 2740 10180 2746 10192
rect 3786 10180 3792 10192
rect 2740 10152 3792 10180
rect 2740 10140 2746 10152
rect 3786 10140 3792 10152
rect 3844 10140 3850 10192
rect 4062 10140 4068 10192
rect 4120 10180 4126 10192
rect 5276 10180 5304 10220
rect 4120 10152 5304 10180
rect 4120 10140 4126 10152
rect 8938 10140 8944 10192
rect 8996 10180 9002 10192
rect 9582 10180 9588 10192
rect 8996 10152 9588 10180
rect 8996 10140 9002 10152
rect 9582 10140 9588 10152
rect 9640 10180 9646 10192
rect 9769 10183 9827 10189
rect 9769 10180 9781 10183
rect 9640 10152 9781 10180
rect 9640 10140 9646 10152
rect 9769 10149 9781 10152
rect 9815 10149 9827 10183
rect 11164 10180 11192 10220
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 14093 10251 14151 10257
rect 14093 10248 14105 10251
rect 11296 10220 14105 10248
rect 11296 10208 11302 10220
rect 14093 10217 14105 10220
rect 14139 10217 14151 10251
rect 14093 10211 14151 10217
rect 15194 10208 15200 10260
rect 15252 10248 15258 10260
rect 15749 10251 15807 10257
rect 15749 10248 15761 10251
rect 15252 10220 15761 10248
rect 15252 10208 15258 10220
rect 15749 10217 15761 10220
rect 15795 10217 15807 10251
rect 15749 10211 15807 10217
rect 11164 10152 11744 10180
rect 9769 10143 9827 10149
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3145 10115 3203 10121
rect 3145 10112 3157 10115
rect 3108 10084 3157 10112
rect 3108 10072 3114 10084
rect 3145 10081 3157 10084
rect 3191 10081 3203 10115
rect 4246 10112 4252 10124
rect 4207 10084 4252 10112
rect 3145 10075 3203 10081
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4356 10084 4936 10112
rect 2332 10016 4016 10044
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 2866 9976 2872 9988
rect 1903 9948 2872 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 2866 9936 2872 9948
rect 2924 9936 2930 9988
rect 1949 9911 2007 9917
rect 1949 9877 1961 9911
rect 1995 9908 2007 9911
rect 2222 9908 2228 9920
rect 1995 9880 2228 9908
rect 1995 9877 2007 9880
rect 1949 9871 2007 9877
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 2498 9868 2504 9920
rect 2556 9908 2562 9920
rect 2961 9911 3019 9917
rect 2961 9908 2973 9911
rect 2556 9880 2973 9908
rect 2556 9868 2562 9880
rect 2961 9877 2973 9880
rect 3007 9877 3019 9911
rect 2961 9871 3019 9877
rect 3050 9868 3056 9920
rect 3108 9908 3114 9920
rect 3108 9880 3153 9908
rect 3108 9868 3114 9880
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3789 9911 3847 9917
rect 3789 9908 3801 9911
rect 3384 9880 3801 9908
rect 3384 9868 3390 9880
rect 3789 9877 3801 9880
rect 3835 9877 3847 9911
rect 3988 9908 4016 10016
rect 4062 10004 4068 10056
rect 4120 10044 4126 10056
rect 4356 10044 4384 10084
rect 4120 10016 4384 10044
rect 4433 10047 4491 10053
rect 4120 10004 4126 10016
rect 4433 10013 4445 10047
rect 4479 10044 4491 10047
rect 4522 10044 4528 10056
rect 4479 10016 4528 10044
rect 4479 10013 4491 10016
rect 4433 10007 4491 10013
rect 4522 10004 4528 10016
rect 4580 10004 4586 10056
rect 4908 10044 4936 10084
rect 5626 10072 5632 10124
rect 5684 10112 5690 10124
rect 5813 10115 5871 10121
rect 5813 10112 5825 10115
rect 5684 10084 5825 10112
rect 5684 10072 5690 10084
rect 5813 10081 5825 10084
rect 5859 10112 5871 10115
rect 5994 10112 6000 10124
rect 5859 10084 6000 10112
rect 5859 10081 5871 10084
rect 5813 10075 5871 10081
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6822 10112 6828 10124
rect 6783 10084 6828 10112
rect 6822 10072 6828 10084
rect 6880 10072 6886 10124
rect 11072 10084 11560 10112
rect 4908 10016 5764 10044
rect 4154 9936 4160 9988
rect 4212 9976 4218 9988
rect 5629 9979 5687 9985
rect 5629 9976 5641 9979
rect 4212 9948 5641 9976
rect 4212 9936 4218 9948
rect 5629 9945 5641 9948
rect 5675 9945 5687 9979
rect 5736 9976 5764 10016
rect 6086 10004 6092 10056
rect 6144 10044 6150 10056
rect 6181 10047 6239 10053
rect 6181 10044 6193 10047
rect 6144 10016 6193 10044
rect 6144 10004 6150 10016
rect 6181 10013 6193 10016
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 7092 10047 7150 10053
rect 7092 10013 7104 10047
rect 7138 10044 7150 10047
rect 8294 10044 8300 10056
rect 7138 10016 8300 10044
rect 7138 10013 7150 10016
rect 7092 10007 7150 10013
rect 8294 10004 8300 10016
rect 8352 10004 8358 10056
rect 8570 10044 8576 10056
rect 8483 10016 8576 10044
rect 8570 10004 8576 10016
rect 8628 10044 8634 10056
rect 8846 10044 8852 10056
rect 8628 10016 8852 10044
rect 8628 10004 8634 10016
rect 8846 10004 8852 10016
rect 8904 10004 8910 10056
rect 11072 10044 11100 10084
rect 11532 10060 11560 10084
rect 9416 10016 11100 10044
rect 8754 9976 8760 9988
rect 5736 9948 8760 9976
rect 5629 9939 5687 9945
rect 8754 9936 8760 9948
rect 8812 9936 8818 9988
rect 4246 9908 4252 9920
rect 3988 9880 4252 9908
rect 3789 9871 3847 9877
rect 4246 9868 4252 9880
rect 4304 9868 4310 9920
rect 4525 9911 4583 9917
rect 4525 9877 4537 9911
rect 4571 9908 4583 9911
rect 4614 9908 4620 9920
rect 4571 9880 4620 9908
rect 4571 9877 4583 9880
rect 4525 9871 4583 9877
rect 4614 9868 4620 9880
rect 4672 9868 4678 9920
rect 4890 9908 4896 9920
rect 4851 9880 4896 9908
rect 4890 9868 4896 9880
rect 4948 9868 4954 9920
rect 5166 9868 5172 9920
rect 5224 9908 5230 9920
rect 5537 9911 5595 9917
rect 5537 9908 5549 9911
rect 5224 9880 5549 9908
rect 5224 9868 5230 9880
rect 5537 9877 5549 9880
rect 5583 9877 5595 9911
rect 5537 9871 5595 9877
rect 6365 9911 6423 9917
rect 6365 9877 6377 9911
rect 6411 9908 6423 9911
rect 7834 9908 7840 9920
rect 6411 9880 7840 9908
rect 6411 9877 6423 9880
rect 6365 9871 6423 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9908 8263 9911
rect 8386 9908 8392 9920
rect 8251 9880 8392 9908
rect 8251 9877 8263 9880
rect 8205 9871 8263 9877
rect 8386 9868 8392 9880
rect 8444 9868 8450 9920
rect 8570 9868 8576 9920
rect 8628 9908 8634 9920
rect 8941 9911 8999 9917
rect 8941 9908 8953 9911
rect 8628 9880 8953 9908
rect 8628 9868 8634 9880
rect 8941 9877 8953 9880
rect 8987 9877 8999 9911
rect 8941 9871 8999 9877
rect 9214 9868 9220 9920
rect 9272 9908 9278 9920
rect 9416 9917 9444 10016
rect 11146 10004 11152 10056
rect 11204 10044 11210 10056
rect 11532 10049 11652 10060
rect 11204 10016 11249 10044
rect 11532 10043 11667 10049
rect 11532 10032 11621 10043
rect 11204 10004 11210 10016
rect 11609 10009 11621 10032
rect 11655 10009 11667 10043
rect 11716 10044 11744 10152
rect 11790 10140 11796 10192
rect 11848 10180 11854 10192
rect 11885 10183 11943 10189
rect 11885 10180 11897 10183
rect 11848 10152 11897 10180
rect 11848 10140 11854 10152
rect 11885 10149 11897 10152
rect 11931 10149 11943 10183
rect 11885 10143 11943 10149
rect 13188 10084 14320 10112
rect 13188 10044 13216 10084
rect 11716 10016 13216 10044
rect 13265 10047 13323 10053
rect 11609 10003 11667 10009
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 13630 10044 13636 10056
rect 13311 10016 13636 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 14292 10053 14320 10084
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10044 14335 10047
rect 15013 10047 15071 10053
rect 15013 10044 15025 10047
rect 14323 10016 15025 10044
rect 14323 10013 14335 10016
rect 14277 10007 14335 10013
rect 15013 10013 15025 10016
rect 15059 10013 15071 10047
rect 15013 10007 15071 10013
rect 10042 9936 10048 9988
rect 10100 9976 10106 9988
rect 10904 9979 10962 9985
rect 10904 9976 10916 9979
rect 10100 9948 10916 9976
rect 10100 9936 10106 9948
rect 10904 9945 10916 9948
rect 10950 9976 10962 9979
rect 11330 9976 11336 9988
rect 10950 9948 11336 9976
rect 10950 9945 10962 9948
rect 10904 9939 10962 9945
rect 11330 9936 11336 9948
rect 11388 9936 11394 9988
rect 13020 9979 13078 9985
rect 13020 9945 13032 9979
rect 13066 9976 13078 9979
rect 13814 9976 13820 9988
rect 13066 9948 13820 9976
rect 13066 9945 13078 9948
rect 13020 9939 13078 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 14550 9976 14556 9988
rect 14511 9948 14556 9976
rect 14550 9936 14556 9948
rect 14608 9936 14614 9988
rect 15194 9936 15200 9988
rect 15252 9976 15258 9988
rect 16117 9979 16175 9985
rect 16117 9976 16129 9979
rect 15252 9948 16129 9976
rect 15252 9936 15258 9948
rect 16117 9945 16129 9948
rect 16163 9945 16175 9979
rect 16117 9939 16175 9945
rect 9401 9911 9459 9917
rect 9401 9908 9413 9911
rect 9272 9880 9413 9908
rect 9272 9868 9278 9880
rect 9401 9877 9413 9880
rect 9447 9877 9459 9911
rect 9401 9871 9459 9877
rect 9858 9868 9864 9920
rect 9916 9908 9922 9920
rect 11425 9911 11483 9917
rect 11425 9908 11437 9911
rect 9916 9880 11437 9908
rect 9916 9868 9922 9880
rect 11425 9877 11437 9880
rect 11471 9877 11483 9911
rect 11425 9871 11483 9877
rect 11974 9868 11980 9920
rect 12032 9908 12038 9920
rect 13541 9911 13599 9917
rect 13541 9908 13553 9911
rect 12032 9880 13553 9908
rect 12032 9868 12038 9880
rect 13541 9877 13553 9880
rect 13587 9877 13599 9911
rect 13541 9871 13599 9877
rect 15102 9868 15108 9920
rect 15160 9908 15166 9920
rect 15381 9911 15439 9917
rect 15381 9908 15393 9911
rect 15160 9880 15393 9908
rect 15160 9868 15166 9880
rect 15381 9877 15393 9880
rect 15427 9877 15439 9911
rect 15381 9871 15439 9877
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 3605 9707 3663 9713
rect 3605 9704 3617 9707
rect 3445 9676 3617 9704
rect 2314 9528 2320 9580
rect 2372 9568 2378 9580
rect 2613 9571 2671 9577
rect 2613 9568 2625 9571
rect 2372 9540 2625 9568
rect 2372 9528 2378 9540
rect 2613 9537 2625 9540
rect 2659 9568 2671 9571
rect 2869 9571 2927 9577
rect 2659 9540 2820 9568
rect 2659 9537 2671 9540
rect 2613 9531 2671 9537
rect 2792 9500 2820 9540
rect 2869 9537 2881 9571
rect 2915 9568 2927 9571
rect 3142 9568 3148 9580
rect 2915 9540 3148 9568
rect 2915 9537 2927 9540
rect 2869 9531 2927 9537
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 3326 9528 3332 9580
rect 3384 9568 3390 9580
rect 3445 9568 3473 9676
rect 3605 9673 3617 9676
rect 3651 9673 3663 9707
rect 3605 9667 3663 9673
rect 4709 9707 4767 9713
rect 4709 9673 4721 9707
rect 4755 9704 4767 9707
rect 4890 9704 4896 9716
rect 4755 9676 4896 9704
rect 4755 9673 4767 9676
rect 4709 9667 4767 9673
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5166 9664 5172 9716
rect 5224 9704 5230 9716
rect 8389 9707 8447 9713
rect 5224 9676 8340 9704
rect 5224 9664 5230 9676
rect 5902 9596 5908 9648
rect 5960 9636 5966 9648
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 5960 9608 6009 9636
rect 5960 9596 5966 9608
rect 5997 9605 6009 9608
rect 6043 9605 6055 9639
rect 7558 9636 7564 9648
rect 7519 9608 7564 9636
rect 5997 9599 6055 9605
rect 7558 9596 7564 9608
rect 7616 9596 7622 9648
rect 8312 9636 8340 9676
rect 8389 9673 8401 9707
rect 8435 9704 8447 9707
rect 8662 9704 8668 9716
rect 8435 9676 8668 9704
rect 8435 9673 8447 9676
rect 8389 9667 8447 9673
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 8754 9664 8760 9716
rect 8812 9704 8818 9716
rect 15102 9704 15108 9716
rect 8812 9676 15108 9704
rect 8812 9664 8818 9676
rect 15102 9664 15108 9676
rect 15160 9664 15166 9716
rect 9674 9636 9680 9648
rect 8312 9608 9680 9636
rect 9674 9596 9680 9608
rect 9732 9636 9738 9648
rect 9861 9639 9919 9645
rect 9861 9636 9873 9639
rect 9732 9608 9873 9636
rect 9732 9596 9738 9608
rect 9861 9605 9873 9608
rect 9907 9605 9919 9639
rect 9861 9599 9919 9605
rect 10781 9639 10839 9645
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11238 9636 11244 9648
rect 10827 9608 11244 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11238 9596 11244 9608
rect 11296 9596 11302 9648
rect 11784 9639 11842 9645
rect 11784 9605 11796 9639
rect 11830 9636 11842 9639
rect 13814 9636 13820 9648
rect 11830 9608 13676 9636
rect 13775 9608 13820 9636
rect 11830 9605 11842 9608
rect 11784 9599 11842 9605
rect 3384 9540 3473 9568
rect 3513 9571 3571 9577
rect 3384 9528 3390 9540
rect 3513 9537 3525 9571
rect 3559 9568 3571 9571
rect 4338 9568 4344 9580
rect 3559 9540 4344 9568
rect 3559 9537 3571 9540
rect 3513 9531 3571 9537
rect 4338 9528 4344 9540
rect 4396 9528 4402 9580
rect 4617 9571 4675 9577
rect 4617 9537 4629 9571
rect 4663 9568 4675 9571
rect 5074 9568 5080 9580
rect 4663 9540 5080 9568
rect 4663 9537 4675 9540
rect 4617 9531 4675 9537
rect 5074 9528 5080 9540
rect 5132 9528 5138 9580
rect 5353 9571 5411 9577
rect 5353 9537 5365 9571
rect 5399 9568 5411 9571
rect 5626 9568 5632 9580
rect 5399 9540 5632 9568
rect 5399 9537 5411 9540
rect 5353 9531 5411 9537
rect 5626 9528 5632 9540
rect 5684 9528 5690 9580
rect 6178 9528 6184 9580
rect 6236 9568 6242 9580
rect 8662 9568 8668 9580
rect 6236 9540 8668 9568
rect 6236 9528 6242 9540
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8757 9571 8815 9577
rect 8757 9537 8769 9571
rect 8803 9568 8815 9571
rect 8803 9540 9444 9568
rect 8803 9537 8815 9540
rect 8757 9531 8815 9537
rect 2792 9472 3556 9500
rect 3528 9444 3556 9472
rect 3694 9460 3700 9512
rect 3752 9500 3758 9512
rect 3752 9472 3797 9500
rect 3752 9460 3758 9472
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 4801 9503 4859 9509
rect 4801 9500 4813 9503
rect 4764 9472 4813 9500
rect 4764 9460 4770 9472
rect 4801 9469 4813 9472
rect 4847 9469 4859 9503
rect 4801 9463 4859 9469
rect 6917 9503 6975 9509
rect 6917 9469 6929 9503
rect 6963 9500 6975 9503
rect 7374 9500 7380 9512
rect 6963 9472 7380 9500
rect 6963 9469 6975 9472
rect 6917 9463 6975 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 7837 9503 7895 9509
rect 7699 9469 7716 9500
rect 7653 9463 7716 9469
rect 7837 9469 7849 9503
rect 7883 9500 7895 9503
rect 8018 9500 8024 9512
rect 7883 9472 8024 9500
rect 7883 9469 7895 9472
rect 7837 9463 7895 9469
rect 1486 9432 1492 9444
rect 1447 9404 1492 9432
rect 1486 9392 1492 9404
rect 1544 9392 1550 9444
rect 3510 9392 3516 9444
rect 3568 9392 3574 9444
rect 3786 9392 3792 9444
rect 3844 9432 3850 9444
rect 4249 9435 4307 9441
rect 4249 9432 4261 9435
rect 3844 9404 4261 9432
rect 3844 9392 3850 9404
rect 4249 9401 4261 9404
rect 4295 9401 4307 9435
rect 7558 9432 7564 9444
rect 4249 9395 4307 9401
rect 5828 9404 7564 9432
rect 3142 9324 3148 9376
rect 3200 9364 3206 9376
rect 3200 9336 3245 9364
rect 3200 9324 3206 9336
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 5828 9364 5856 9404
rect 7558 9392 7564 9404
rect 7616 9392 7622 9444
rect 7688 9432 7716 9463
rect 8018 9460 8024 9472
rect 8076 9460 8082 9512
rect 8849 9503 8907 9509
rect 8849 9469 8861 9503
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 7688 9404 7972 9432
rect 4672 9336 5856 9364
rect 4672 9324 4678 9336
rect 5902 9324 5908 9376
rect 5960 9364 5966 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5960 9336 6377 9364
rect 5960 9324 5966 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 6365 9327 6423 9333
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 7944 9364 7972 9404
rect 8110 9392 8116 9444
rect 8168 9432 8174 9444
rect 8754 9432 8760 9444
rect 8168 9404 8760 9432
rect 8168 9392 8174 9404
rect 8754 9392 8760 9404
rect 8812 9392 8818 9444
rect 8864 9432 8892 9463
rect 8938 9460 8944 9512
rect 8996 9500 9002 9512
rect 8996 9472 9041 9500
rect 8996 9460 9002 9472
rect 9306 9432 9312 9444
rect 8864 9404 9312 9432
rect 9306 9392 9312 9404
rect 9364 9392 9370 9444
rect 9416 9441 9444 9540
rect 9582 9528 9588 9580
rect 9640 9568 9646 9580
rect 9769 9571 9827 9577
rect 9769 9568 9781 9571
rect 9640 9540 9781 9568
rect 9640 9528 9646 9540
rect 9769 9537 9781 9540
rect 9815 9537 9827 9571
rect 9769 9531 9827 9537
rect 9401 9435 9459 9441
rect 9401 9401 9413 9435
rect 9447 9401 9459 9435
rect 9784 9432 9812 9531
rect 11146 9528 11152 9580
rect 11204 9568 11210 9580
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 11204 9540 11529 9568
rect 11204 9528 11210 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 11517 9531 11575 9537
rect 11624 9540 12848 9568
rect 10042 9500 10048 9512
rect 10003 9472 10048 9500
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 10689 9503 10747 9509
rect 10689 9469 10701 9503
rect 10735 9500 10747 9503
rect 10778 9500 10784 9512
rect 10735 9472 10784 9500
rect 10735 9469 10747 9472
rect 10689 9463 10747 9469
rect 10778 9460 10784 9472
rect 10836 9460 10842 9512
rect 11624 9500 11652 9540
rect 11532 9472 11652 9500
rect 12820 9500 12848 9540
rect 12894 9528 12900 9580
rect 12952 9568 12958 9580
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12952 9540 13185 9568
rect 12952 9528 12958 9540
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 13173 9531 13231 9537
rect 13648 9500 13676 9608
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14185 9571 14243 9577
rect 14185 9537 14197 9571
rect 14231 9568 14243 9571
rect 14274 9568 14280 9580
rect 14231 9540 14280 9568
rect 14231 9537 14243 9540
rect 14185 9531 14243 9537
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 15120 9577 15148 9664
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15746 9568 15752 9580
rect 15707 9540 15752 9568
rect 15105 9531 15163 9537
rect 15746 9528 15752 9540
rect 15804 9568 15810 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15804 9540 16037 9568
rect 15804 9528 15810 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 14829 9503 14887 9509
rect 14829 9500 14841 9503
rect 12820 9472 13032 9500
rect 13648 9472 14841 9500
rect 11532 9432 11560 9472
rect 9784 9404 11560 9432
rect 9401 9395 9459 9401
rect 11054 9364 11060 9376
rect 7944 9336 11060 9364
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 11149 9367 11207 9373
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 11790 9364 11796 9376
rect 11195 9336 11796 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 11790 9324 11796 9336
rect 11848 9324 11854 9376
rect 11882 9324 11888 9376
rect 11940 9364 11946 9376
rect 12618 9364 12624 9376
rect 11940 9336 12624 9364
rect 11940 9324 11946 9336
rect 12618 9324 12624 9336
rect 12676 9324 12682 9376
rect 12894 9364 12900 9376
rect 12855 9336 12900 9364
rect 12894 9324 12900 9336
rect 12952 9324 12958 9376
rect 13004 9364 13032 9472
rect 14829 9469 14841 9472
rect 14875 9469 14887 9503
rect 14829 9463 14887 9469
rect 14918 9460 14924 9512
rect 14976 9500 14982 9512
rect 16669 9503 16727 9509
rect 16669 9500 16681 9503
rect 14976 9472 16681 9500
rect 14976 9460 14982 9472
rect 16669 9469 16681 9472
rect 16715 9469 16727 9503
rect 16669 9463 16727 9469
rect 15289 9435 15347 9441
rect 15289 9401 15301 9435
rect 15335 9432 15347 9435
rect 17126 9432 17132 9444
rect 15335 9404 17132 9432
rect 15335 9401 15347 9404
rect 15289 9395 15347 9401
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 15470 9364 15476 9376
rect 13004 9336 15476 9364
rect 15470 9324 15476 9336
rect 15528 9324 15534 9376
rect 15565 9367 15623 9373
rect 15565 9333 15577 9367
rect 15611 9364 15623 9367
rect 15654 9364 15660 9376
rect 15611 9336 15660 9364
rect 15611 9333 15623 9336
rect 15565 9327 15623 9333
rect 15654 9324 15660 9336
rect 15712 9324 15718 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1578 9160 1584 9172
rect 1539 9132 1584 9160
rect 1578 9120 1584 9132
rect 1636 9120 1642 9172
rect 1946 9160 1952 9172
rect 1907 9132 1952 9160
rect 1946 9120 1952 9132
rect 2004 9120 2010 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4120 9132 8524 9160
rect 4120 9120 4126 9132
rect 1302 9052 1308 9104
rect 1360 9092 1366 9104
rect 5442 9092 5448 9104
rect 1360 9064 5448 9092
rect 1360 9052 1366 9064
rect 5442 9052 5448 9064
rect 5500 9052 5506 9104
rect 6730 9052 6736 9104
rect 6788 9092 6794 9104
rect 6825 9095 6883 9101
rect 6825 9092 6837 9095
rect 6788 9064 6837 9092
rect 6788 9052 6794 9064
rect 6825 9061 6837 9064
rect 6871 9061 6883 9095
rect 8496 9092 8524 9132
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9677 9163 9735 9169
rect 9677 9160 9689 9163
rect 9364 9132 9689 9160
rect 9364 9120 9370 9132
rect 9677 9129 9689 9132
rect 9723 9129 9735 9163
rect 12802 9160 12808 9172
rect 9677 9123 9735 9129
rect 9784 9132 12808 9160
rect 9784 9092 9812 9132
rect 12802 9120 12808 9132
rect 12860 9120 12866 9172
rect 12897 9163 12955 9169
rect 12897 9129 12909 9163
rect 12943 9160 12955 9163
rect 12943 9132 17080 9160
rect 12943 9129 12955 9132
rect 12897 9123 12955 9129
rect 8496 9064 9812 9092
rect 6825 9055 6883 9061
rect 10042 9052 10048 9104
rect 10100 9092 10106 9104
rect 10100 9064 10272 9092
rect 10100 9052 10106 9064
rect 1486 8984 1492 9036
rect 1544 9024 1550 9036
rect 2501 9027 2559 9033
rect 2501 9024 2513 9027
rect 1544 8996 2513 9024
rect 1544 8984 1550 8996
rect 2501 8993 2513 8996
rect 2547 8993 2559 9027
rect 2501 8987 2559 8993
rect 2682 8984 2688 9036
rect 2740 9024 2746 9036
rect 4709 9027 4767 9033
rect 2740 8996 3280 9024
rect 2740 8984 2746 8996
rect 1210 8916 1216 8968
rect 1268 8956 1274 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 1268 8928 1409 8956
rect 1268 8916 1274 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 2317 8959 2375 8965
rect 2317 8925 2329 8959
rect 2363 8956 2375 8959
rect 3142 8956 3148 8968
rect 2363 8928 3148 8956
rect 2363 8925 2375 8928
rect 2317 8919 2375 8925
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 3252 8965 3280 8996
rect 4709 8993 4721 9027
rect 4755 8993 4767 9027
rect 4709 8987 4767 8993
rect 3237 8959 3295 8965
rect 3237 8925 3249 8959
rect 3283 8925 3295 8959
rect 4724 8956 4752 8987
rect 4798 8984 4804 9036
rect 4856 9024 4862 9036
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 4856 8996 5641 9024
rect 4856 8984 4862 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 6270 9024 6276 9036
rect 6231 8996 6276 9024
rect 5629 8987 5687 8993
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 8662 8984 8668 9036
rect 8720 9024 8726 9036
rect 9582 9024 9588 9036
rect 8720 8996 9588 9024
rect 8720 8984 8726 8996
rect 9582 8984 9588 8996
rect 9640 8984 9646 9036
rect 10244 9033 10272 9064
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 14093 9095 14151 9101
rect 14093 9092 14105 9095
rect 10652 9064 14105 9092
rect 10652 9052 10658 9064
rect 14093 9061 14105 9064
rect 14139 9092 14151 9095
rect 14274 9092 14280 9104
rect 14139 9064 14280 9092
rect 14139 9061 14151 9064
rect 14093 9055 14151 9061
rect 14274 9052 14280 9064
rect 14332 9052 14338 9104
rect 15562 9052 15568 9104
rect 15620 9092 15626 9104
rect 15620 9064 16528 9092
rect 15620 9052 15626 9064
rect 10229 9027 10287 9033
rect 10229 8993 10241 9027
rect 10275 8993 10287 9027
rect 10229 8987 10287 8993
rect 12345 9027 12403 9033
rect 12345 8993 12357 9027
rect 12391 9024 12403 9027
rect 12894 9024 12900 9036
rect 12391 8996 12900 9024
rect 12391 8993 12403 8996
rect 12345 8987 12403 8993
rect 12894 8984 12900 8996
rect 12952 8984 12958 9036
rect 15473 9027 15531 9033
rect 15473 8993 15485 9027
rect 15519 9024 15531 9027
rect 16298 9024 16304 9036
rect 15519 8996 16304 9024
rect 15519 8993 15531 8996
rect 15473 8987 15531 8993
rect 16298 8984 16304 8996
rect 16356 8984 16362 9036
rect 5442 8956 5448 8968
rect 4724 8928 5448 8956
rect 3237 8919 3295 8925
rect 5442 8916 5448 8928
rect 5500 8916 5506 8968
rect 6457 8959 6515 8965
rect 6457 8925 6469 8959
rect 6503 8956 6515 8959
rect 6503 8928 8340 8956
rect 6503 8925 6515 8928
rect 6457 8919 6515 8925
rect 2774 8848 2780 8900
rect 2832 8888 2838 8900
rect 3786 8888 3792 8900
rect 2832 8860 3792 8888
rect 2832 8848 2838 8860
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 4982 8848 4988 8900
rect 5040 8888 5046 8900
rect 5537 8891 5595 8897
rect 5537 8888 5549 8891
rect 5040 8860 5549 8888
rect 5040 8848 5046 8860
rect 5537 8857 5549 8860
rect 5583 8857 5595 8891
rect 5537 8851 5595 8857
rect 6365 8891 6423 8897
rect 6365 8857 6377 8891
rect 6411 8888 6423 8891
rect 6411 8860 8064 8888
rect 6411 8857 6423 8860
rect 6365 8851 6423 8857
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 2464 8792 2509 8820
rect 2464 8780 2470 8792
rect 3234 8780 3240 8832
rect 3292 8820 3298 8832
rect 3421 8823 3479 8829
rect 3421 8820 3433 8823
rect 3292 8792 3433 8820
rect 3292 8780 3298 8792
rect 3421 8789 3433 8792
rect 3467 8789 3479 8823
rect 3421 8783 3479 8789
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 4028 8792 4077 8820
rect 4028 8780 4034 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 4430 8820 4436 8832
rect 4391 8792 4436 8820
rect 4065 8783 4123 8789
rect 4430 8780 4436 8792
rect 4488 8780 4494 8832
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8820 4583 8823
rect 5077 8823 5135 8829
rect 5077 8820 5089 8823
rect 4571 8792 5089 8820
rect 4571 8789 4583 8792
rect 4525 8783 4583 8789
rect 5077 8789 5089 8792
rect 5123 8789 5135 8823
rect 5077 8783 5135 8789
rect 5445 8823 5503 8829
rect 5445 8789 5457 8823
rect 5491 8820 5503 8823
rect 5994 8820 6000 8832
rect 5491 8792 6000 8820
rect 5491 8789 5503 8792
rect 5445 8783 5503 8789
rect 5994 8780 6000 8792
rect 6052 8780 6058 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7101 8823 7159 8829
rect 7101 8820 7113 8823
rect 6972 8792 7113 8820
rect 6972 8780 6978 8792
rect 7101 8789 7113 8792
rect 7147 8789 7159 8823
rect 8036 8820 8064 8860
rect 8110 8848 8116 8900
rect 8168 8888 8174 8900
rect 8214 8891 8272 8897
rect 8214 8888 8226 8891
rect 8168 8860 8226 8888
rect 8168 8848 8174 8860
rect 8214 8857 8226 8860
rect 8260 8857 8272 8891
rect 8312 8888 8340 8928
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8481 8959 8539 8965
rect 8481 8956 8493 8959
rect 8444 8928 8493 8956
rect 8444 8916 8450 8928
rect 8481 8925 8493 8928
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 10689 8959 10747 8965
rect 10689 8956 10701 8959
rect 10100 8928 10701 8956
rect 10100 8916 10106 8928
rect 10689 8925 10701 8928
rect 10735 8925 10747 8959
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 10689 8919 10747 8925
rect 11164 8928 11805 8956
rect 8570 8888 8576 8900
rect 8312 8860 8576 8888
rect 8214 8851 8272 8857
rect 8570 8848 8576 8860
rect 8628 8848 8634 8900
rect 10134 8888 10140 8900
rect 10095 8860 10140 8888
rect 10134 8848 10140 8860
rect 10192 8848 10198 8900
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 11164 8888 11192 8928
rect 11793 8925 11805 8928
rect 11839 8956 11851 8959
rect 13633 8959 13691 8965
rect 13633 8956 13645 8959
rect 11839 8928 13645 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 13633 8925 13645 8928
rect 13679 8925 13691 8959
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 13633 8919 13691 8925
rect 15028 8928 15761 8956
rect 15028 8900 15056 8928
rect 15749 8925 15761 8928
rect 15795 8925 15807 8959
rect 15749 8919 15807 8925
rect 10468 8860 11192 8888
rect 11333 8891 11391 8897
rect 10468 8848 10474 8860
rect 11333 8857 11345 8891
rect 11379 8888 11391 8891
rect 12342 8888 12348 8900
rect 11379 8860 12348 8888
rect 11379 8857 11391 8860
rect 11333 8851 11391 8857
rect 12342 8848 12348 8860
rect 12400 8848 12406 8900
rect 12529 8891 12587 8897
rect 12529 8857 12541 8891
rect 12575 8888 12587 8891
rect 13173 8891 13231 8897
rect 13173 8888 13185 8891
rect 12575 8860 13185 8888
rect 12575 8857 12587 8860
rect 12529 8851 12587 8857
rect 13173 8857 13185 8860
rect 13219 8857 13231 8891
rect 13173 8851 13231 8857
rect 15010 8848 15016 8900
rect 15068 8848 15074 8900
rect 15228 8891 15286 8897
rect 15228 8857 15240 8891
rect 15274 8888 15286 8891
rect 16393 8891 16451 8897
rect 16393 8888 16405 8891
rect 15274 8860 16405 8888
rect 15274 8857 15286 8860
rect 15228 8851 15286 8857
rect 16393 8857 16405 8860
rect 16439 8857 16451 8891
rect 16500 8888 16528 9064
rect 17052 8965 17080 9132
rect 17221 9095 17279 9101
rect 17221 9061 17233 9095
rect 17267 9092 17279 9095
rect 19886 9092 19892 9104
rect 17267 9064 19892 9092
rect 17267 9061 17279 9064
rect 17221 9055 17279 9061
rect 19886 9052 19892 9064
rect 19944 9052 19950 9104
rect 17037 8959 17095 8965
rect 17037 8925 17049 8959
rect 17083 8925 17095 8959
rect 17037 8919 17095 8925
rect 17497 8891 17555 8897
rect 17497 8888 17509 8891
rect 16500 8860 17509 8888
rect 16393 8851 16451 8857
rect 17497 8857 17509 8860
rect 17543 8857 17555 8891
rect 17497 8851 17555 8857
rect 8938 8820 8944 8832
rect 8036 8792 8944 8820
rect 7101 8783 7159 8789
rect 8938 8780 8944 8792
rect 8996 8780 9002 8832
rect 9122 8820 9128 8832
rect 9083 8792 9128 8820
rect 9122 8780 9128 8792
rect 9180 8780 9186 8832
rect 10045 8823 10103 8829
rect 10045 8789 10057 8823
rect 10091 8820 10103 8823
rect 10226 8820 10232 8832
rect 10091 8792 10232 8820
rect 10091 8789 10103 8792
rect 10045 8783 10103 8789
rect 10226 8780 10232 8792
rect 10284 8780 10290 8832
rect 11054 8780 11060 8832
rect 11112 8820 11118 8832
rect 11609 8823 11667 8829
rect 11609 8820 11621 8823
rect 11112 8792 11621 8820
rect 11112 8780 11118 8792
rect 11609 8789 11621 8792
rect 11655 8789 11667 8823
rect 11609 8783 11667 8789
rect 11790 8780 11796 8832
rect 11848 8820 11854 8832
rect 12437 8823 12495 8829
rect 12437 8820 12449 8823
rect 11848 8792 12449 8820
rect 11848 8780 11854 8792
rect 12437 8789 12449 8792
rect 12483 8789 12495 8823
rect 12437 8783 12495 8789
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 16669 8823 16727 8829
rect 16669 8820 16681 8823
rect 12676 8792 16681 8820
rect 12676 8780 12682 8792
rect 16669 8789 16681 8792
rect 16715 8789 16727 8823
rect 16669 8783 16727 8789
rect 17957 8823 18015 8829
rect 17957 8789 17969 8823
rect 18003 8820 18015 8823
rect 18230 8820 18236 8832
rect 18003 8792 18236 8820
rect 18003 8789 18015 8792
rect 17957 8783 18015 8789
rect 18230 8780 18236 8792
rect 18288 8780 18294 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 2314 8616 2320 8628
rect 2275 8588 2320 8616
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 4798 8616 4804 8628
rect 2648 8588 4804 8616
rect 2648 8576 2654 8588
rect 4798 8576 4804 8588
rect 4856 8616 4862 8628
rect 6365 8619 6423 8625
rect 6365 8616 6377 8619
rect 4856 8588 6377 8616
rect 4856 8576 4862 8588
rect 6365 8585 6377 8588
rect 6411 8585 6423 8619
rect 8110 8616 8116 8628
rect 8071 8588 8116 8616
rect 6365 8579 6423 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8938 8576 8944 8628
rect 8996 8616 9002 8628
rect 9033 8619 9091 8625
rect 9033 8616 9045 8619
rect 8996 8588 9045 8616
rect 8996 8576 9002 8588
rect 9033 8585 9045 8588
rect 9079 8585 9091 8619
rect 9033 8579 9091 8585
rect 9401 8619 9459 8625
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 9490 8616 9496 8628
rect 9447 8588 9496 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 9490 8576 9496 8588
rect 9548 8576 9554 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 12989 8619 13047 8625
rect 12989 8616 13001 8619
rect 12768 8588 13001 8616
rect 12768 8576 12774 8588
rect 12989 8585 13001 8588
rect 13035 8585 13047 8619
rect 15010 8616 15016 8628
rect 14971 8588 15016 8616
rect 12989 8579 13047 8585
rect 15010 8576 15016 8588
rect 15068 8576 15074 8628
rect 15933 8619 15991 8625
rect 15933 8585 15945 8619
rect 15979 8616 15991 8619
rect 15979 8588 17908 8616
rect 15979 8585 15991 8588
rect 15933 8579 15991 8585
rect 1397 8551 1455 8557
rect 1397 8517 1409 8551
rect 1443 8548 1455 8551
rect 2774 8548 2780 8560
rect 1443 8520 2780 8548
rect 1443 8517 1455 8520
rect 1397 8511 1455 8517
rect 2774 8508 2780 8520
rect 2832 8508 2838 8560
rect 4890 8548 4896 8560
rect 4448 8520 4896 8548
rect 2041 8483 2099 8489
rect 2041 8449 2053 8483
rect 2087 8480 2099 8483
rect 2590 8480 2596 8492
rect 2087 8452 2596 8480
rect 2087 8449 2099 8452
rect 2041 8443 2099 8449
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 3142 8440 3148 8492
rect 3200 8480 3206 8492
rect 3441 8483 3499 8489
rect 3441 8480 3453 8483
rect 3200 8452 3453 8480
rect 3200 8440 3206 8452
rect 3441 8449 3453 8452
rect 3487 8449 3499 8483
rect 3441 8443 3499 8449
rect 3786 8440 3792 8492
rect 3844 8480 3850 8492
rect 4448 8489 4476 8520
rect 4890 8508 4896 8520
rect 4948 8548 4954 8560
rect 5534 8548 5540 8560
rect 4948 8520 5540 8548
rect 4948 8508 4954 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 7374 8508 7380 8560
rect 7432 8548 7438 8560
rect 7432 8520 7880 8548
rect 7432 8508 7438 8520
rect 4433 8483 4491 8489
rect 3844 8452 4384 8480
rect 3844 8440 3850 8452
rect 3697 8415 3755 8421
rect 3697 8381 3709 8415
rect 3743 8381 3755 8415
rect 4154 8412 4160 8424
rect 4115 8384 4160 8412
rect 3697 8375 3755 8381
rect 3712 8344 3740 8375
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 4356 8412 4384 8452
rect 4433 8449 4445 8483
rect 4479 8449 4491 8483
rect 4689 8483 4747 8489
rect 4689 8480 4701 8483
rect 4433 8443 4491 8449
rect 4540 8452 4701 8480
rect 4540 8412 4568 8452
rect 4689 8449 4701 8452
rect 4735 8449 4747 8483
rect 4689 8443 4747 8449
rect 6914 8440 6920 8492
rect 6972 8480 6978 8492
rect 7478 8483 7536 8489
rect 7478 8480 7490 8483
rect 6972 8452 7490 8480
rect 6972 8440 6978 8452
rect 7478 8449 7490 8452
rect 7524 8449 7536 8483
rect 7852 8480 7880 8520
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 9214 8548 9220 8560
rect 8076 8520 9220 8548
rect 8076 8508 8082 8520
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 12158 8548 12164 8560
rect 9324 8520 12164 8548
rect 8202 8480 8208 8492
rect 7852 8452 8208 8480
rect 7478 8443 7536 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 8478 8440 8484 8492
rect 8536 8480 8542 8492
rect 8757 8483 8815 8489
rect 8757 8480 8769 8483
rect 8536 8452 8769 8480
rect 8536 8440 8542 8452
rect 8757 8449 8769 8452
rect 8803 8449 8815 8483
rect 8757 8443 8815 8449
rect 4356 8384 4568 8412
rect 7745 8415 7803 8421
rect 7745 8381 7757 8415
rect 7791 8412 7803 8415
rect 8386 8412 8392 8424
rect 7791 8384 8392 8412
rect 7791 8381 7803 8384
rect 7745 8375 7803 8381
rect 8386 8372 8392 8384
rect 8444 8372 8450 8424
rect 3712 8316 4476 8344
rect 4448 8276 4476 8316
rect 5442 8304 5448 8356
rect 5500 8344 5506 8356
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5500 8316 5825 8344
rect 5500 8304 5506 8316
rect 5813 8313 5825 8316
rect 5859 8344 5871 8347
rect 9324 8344 9352 8520
rect 12158 8508 12164 8520
rect 12216 8508 12222 8560
rect 13900 8551 13958 8557
rect 13900 8517 13912 8551
rect 13946 8548 13958 8551
rect 16942 8548 16948 8560
rect 13946 8520 16948 8548
rect 13946 8517 13958 8520
rect 13900 8511 13958 8517
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17880 8548 17908 8588
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 20714 8616 20720 8628
rect 18012 8588 20720 8616
rect 18012 8576 18018 8588
rect 20714 8576 20720 8588
rect 20772 8576 20778 8628
rect 18598 8548 18604 8560
rect 17880 8520 18604 8548
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 10318 8480 10324 8492
rect 10279 8452 10324 8480
rect 10318 8440 10324 8452
rect 10376 8440 10382 8492
rect 11054 8440 11060 8492
rect 11112 8480 11118 8492
rect 11885 8483 11943 8489
rect 11885 8480 11897 8483
rect 11112 8452 11897 8480
rect 11112 8440 11118 8452
rect 11885 8449 11897 8452
rect 11931 8449 11943 8483
rect 15654 8480 15660 8492
rect 11885 8443 11943 8449
rect 12820 8452 15660 8480
rect 9490 8412 9496 8424
rect 9451 8384 9496 8412
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 9950 8412 9956 8424
rect 9723 8384 9956 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 9950 8372 9956 8384
rect 10008 8372 10014 8424
rect 11238 8372 11244 8424
rect 11296 8412 11302 8424
rect 11609 8415 11667 8421
rect 11609 8412 11621 8415
rect 11296 8384 11621 8412
rect 11296 8372 11302 8384
rect 11609 8381 11621 8384
rect 11655 8381 11667 8415
rect 11790 8412 11796 8424
rect 11751 8384 11796 8412
rect 11609 8375 11667 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 12820 8421 12848 8452
rect 15654 8440 15660 8452
rect 15712 8440 15718 8492
rect 15746 8440 15752 8492
rect 15804 8480 15810 8492
rect 15804 8452 15849 8480
rect 15804 8440 15810 8452
rect 15930 8440 15936 8492
rect 15988 8480 15994 8492
rect 16669 8483 16727 8489
rect 16669 8480 16681 8483
rect 15988 8452 16681 8480
rect 15988 8440 15994 8452
rect 16669 8449 16681 8452
rect 16715 8449 16727 8483
rect 17310 8480 17316 8492
rect 17271 8452 17316 8480
rect 16669 8443 16727 8449
rect 17310 8440 17316 8452
rect 17368 8480 17374 8492
rect 17589 8483 17647 8489
rect 17589 8480 17601 8483
rect 17368 8452 17601 8480
rect 17368 8440 17374 8452
rect 17589 8449 17601 8452
rect 17635 8449 17647 8483
rect 17589 8443 17647 8449
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 12897 8415 12955 8421
rect 12897 8381 12909 8415
rect 12943 8412 12955 8415
rect 13262 8412 13268 8424
rect 12943 8384 13268 8412
rect 12943 8381 12955 8384
rect 12897 8375 12955 8381
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 13630 8412 13636 8424
rect 13591 8384 13636 8412
rect 13630 8372 13636 8384
rect 13688 8372 13694 8424
rect 14918 8372 14924 8424
rect 14976 8412 14982 8424
rect 15289 8415 15347 8421
rect 15289 8412 15301 8415
rect 14976 8384 15301 8412
rect 14976 8372 14982 8384
rect 15289 8381 15301 8384
rect 15335 8381 15347 8415
rect 16206 8412 16212 8424
rect 16167 8384 16212 8412
rect 15289 8375 15347 8381
rect 16206 8372 16212 8384
rect 16264 8372 16270 8424
rect 10962 8344 10968 8356
rect 5859 8316 6868 8344
rect 5859 8313 5871 8316
rect 5813 8307 5871 8313
rect 5718 8276 5724 8288
rect 4448 8248 5724 8276
rect 5718 8236 5724 8248
rect 5776 8236 5782 8288
rect 6840 8276 6868 8316
rect 7760 8316 9352 8344
rect 10923 8316 10968 8344
rect 7760 8276 7788 8316
rect 10962 8304 10968 8316
rect 11020 8304 11026 8356
rect 17129 8347 17187 8353
rect 17129 8344 17141 8347
rect 14568 8316 17141 8344
rect 12250 8276 12256 8288
rect 6840 8248 7788 8276
rect 12211 8248 12256 8276
rect 12250 8236 12256 8248
rect 12308 8236 12314 8288
rect 13354 8276 13360 8288
rect 13315 8248 13360 8276
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 14568 8276 14596 8316
rect 17129 8313 17141 8316
rect 17175 8313 17187 8347
rect 17954 8344 17960 8356
rect 17915 8316 17960 8344
rect 17129 8307 17187 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 18322 8344 18328 8356
rect 18283 8316 18328 8344
rect 18322 8304 18328 8316
rect 18380 8304 18386 8356
rect 18782 8344 18788 8356
rect 18743 8316 18788 8344
rect 18782 8304 18788 8316
rect 18840 8304 18846 8356
rect 13596 8248 14596 8276
rect 13596 8236 13602 8248
rect 15562 8236 15568 8288
rect 15620 8276 15626 8288
rect 20254 8276 20260 8288
rect 15620 8248 20260 8276
rect 15620 8236 15626 8248
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2406 8072 2412 8084
rect 2367 8044 2412 8072
rect 2406 8032 2412 8044
rect 2464 8032 2470 8084
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 3108 8044 3801 8072
rect 3108 8032 3114 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 4982 8072 4988 8084
rect 4943 8044 4988 8072
rect 3789 8035 3847 8041
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5718 8072 5724 8084
rect 5679 8044 5724 8072
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6604 8044 7144 8072
rect 6604 8032 6610 8044
rect 3418 7964 3424 8016
rect 3476 8004 3482 8016
rect 6730 8004 6736 8016
rect 3476 7976 6736 8004
rect 3476 7964 3482 7976
rect 6730 7964 6736 7976
rect 6788 7964 6794 8016
rect 1857 7939 1915 7945
rect 1857 7905 1869 7939
rect 1903 7936 1915 7939
rect 2314 7936 2320 7948
rect 1903 7908 2320 7936
rect 1903 7905 1915 7908
rect 1857 7899 1915 7905
rect 2314 7896 2320 7908
rect 2372 7896 2378 7948
rect 3142 7896 3148 7948
rect 3200 7936 3206 7948
rect 3237 7939 3295 7945
rect 3237 7936 3249 7939
rect 3200 7908 3249 7936
rect 3200 7896 3206 7908
rect 3237 7905 3249 7908
rect 3283 7905 3295 7939
rect 3237 7899 3295 7905
rect 4433 7939 4491 7945
rect 4433 7905 4445 7939
rect 4479 7936 4491 7939
rect 6914 7936 6920 7948
rect 4479 7908 6920 7936
rect 4479 7905 4491 7908
rect 4433 7899 4491 7905
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 3973 7871 4031 7877
rect 2556 7840 3096 7868
rect 2556 7828 2562 7840
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7800 2007 7803
rect 2590 7800 2596 7812
rect 1995 7772 2596 7800
rect 1995 7769 2007 7772
rect 1949 7763 2007 7769
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 3068 7809 3096 7840
rect 3973 7837 3985 7871
rect 4019 7868 4031 7871
rect 4062 7868 4068 7880
rect 4019 7840 4068 7868
rect 4019 7837 4031 7840
rect 3973 7831 4031 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 6638 7868 6644 7880
rect 4448 7840 6644 7868
rect 3053 7803 3111 7809
rect 3053 7769 3065 7803
rect 3099 7800 3111 7803
rect 4448 7800 4476 7840
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7006 7868 7012 7880
rect 6967 7840 7012 7868
rect 7006 7828 7012 7840
rect 7064 7828 7070 7880
rect 7116 7868 7144 8044
rect 7742 8032 7748 8084
rect 7800 8072 7806 8084
rect 8021 8075 8079 8081
rect 8021 8072 8033 8075
rect 7800 8044 8033 8072
rect 7800 8032 7806 8044
rect 8021 8041 8033 8044
rect 8067 8041 8079 8075
rect 8021 8035 8079 8041
rect 8481 8075 8539 8081
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 15562 8072 15568 8084
rect 8527 8044 15568 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 15654 8032 15660 8084
rect 15712 8072 15718 8084
rect 16390 8072 16396 8084
rect 15712 8044 16396 8072
rect 15712 8032 15718 8044
rect 16390 8032 16396 8044
rect 16448 8032 16454 8084
rect 14274 7964 14280 8016
rect 14332 8004 14338 8016
rect 14332 7976 15424 8004
rect 14332 7964 14338 7976
rect 7466 7936 7472 7948
rect 7427 7908 7472 7936
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7936 11023 7939
rect 11054 7936 11060 7948
rect 11011 7908 11060 7936
rect 11011 7905 11023 7908
rect 10965 7899 11023 7905
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 14461 7939 14519 7945
rect 14461 7905 14473 7939
rect 14507 7936 14519 7939
rect 15010 7936 15016 7948
rect 14507 7908 15016 7936
rect 14507 7905 14519 7908
rect 14461 7899 14519 7905
rect 15010 7896 15016 7908
rect 15068 7896 15074 7948
rect 15102 7896 15108 7948
rect 15160 7936 15166 7948
rect 15289 7939 15347 7945
rect 15289 7936 15301 7939
rect 15160 7908 15301 7936
rect 15160 7896 15166 7908
rect 15289 7905 15301 7908
rect 15335 7905 15347 7939
rect 15289 7899 15347 7905
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 7116 7840 8309 7868
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 8938 7868 8944 7880
rect 8444 7840 8944 7868
rect 8444 7828 8450 7840
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 9208 7871 9266 7877
rect 9208 7837 9220 7871
rect 9254 7868 9266 7871
rect 10594 7868 10600 7880
rect 9254 7840 10600 7868
rect 9254 7837 9266 7840
rect 9208 7831 9266 7837
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 12621 7871 12679 7877
rect 11940 7840 12572 7868
rect 11940 7828 11946 7840
rect 3099 7772 4476 7800
rect 4525 7803 4583 7809
rect 3099 7769 3111 7772
rect 3053 7763 3111 7769
rect 4525 7769 4537 7803
rect 4571 7800 4583 7803
rect 4571 7772 9260 7800
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 2041 7735 2099 7741
rect 2041 7701 2053 7735
rect 2087 7732 2099 7735
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2087 7704 2697 7732
rect 2087 7701 2099 7704
rect 2041 7695 2099 7701
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 4062 7732 4068 7744
rect 3191 7704 4068 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4614 7732 4620 7744
rect 4575 7704 4620 7732
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 5442 7692 5448 7744
rect 5500 7732 5506 7744
rect 7098 7732 7104 7744
rect 5500 7704 7104 7732
rect 5500 7692 5506 7704
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7558 7732 7564 7744
rect 7519 7704 7564 7732
rect 7558 7692 7564 7704
rect 7616 7692 7622 7744
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 8386 7732 8392 7744
rect 7699 7704 8392 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 9232 7732 9260 7772
rect 9306 7760 9312 7812
rect 9364 7800 9370 7812
rect 12434 7809 12440 7812
rect 12376 7803 12440 7809
rect 12376 7800 12388 7803
rect 9364 7772 11376 7800
rect 12347 7772 12388 7800
rect 9364 7760 9370 7772
rect 10134 7732 10140 7744
rect 9232 7704 10140 7732
rect 10134 7692 10140 7704
rect 10192 7692 10198 7744
rect 10318 7732 10324 7744
rect 10279 7704 10324 7732
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11241 7735 11299 7741
rect 11241 7732 11253 7735
rect 11112 7704 11253 7732
rect 11112 7692 11118 7704
rect 11241 7701 11253 7704
rect 11287 7701 11299 7735
rect 11348 7732 11376 7772
rect 12376 7769 12388 7772
rect 12422 7769 12440 7803
rect 12376 7763 12440 7769
rect 12434 7760 12440 7763
rect 12492 7760 12498 7812
rect 12544 7800 12572 7840
rect 12621 7837 12633 7871
rect 12667 7868 12679 7871
rect 12802 7868 12808 7880
rect 12667 7840 12808 7868
rect 12667 7837 12679 7840
rect 12621 7831 12679 7837
rect 12802 7828 12808 7840
rect 12860 7828 12866 7880
rect 12897 7871 12955 7877
rect 12897 7837 12909 7871
rect 12943 7837 12955 7871
rect 12897 7831 12955 7837
rect 12912 7800 12940 7831
rect 13354 7828 13360 7880
rect 13412 7868 13418 7880
rect 14553 7871 14611 7877
rect 14553 7868 14565 7871
rect 13412 7840 14565 7868
rect 13412 7828 13418 7840
rect 14553 7837 14565 7840
rect 14599 7837 14611 7871
rect 14553 7831 14611 7837
rect 14645 7871 14703 7877
rect 14645 7837 14657 7871
rect 14691 7868 14703 7871
rect 14918 7868 14924 7880
rect 14691 7840 14924 7868
rect 14691 7837 14703 7840
rect 14645 7831 14703 7837
rect 14918 7828 14924 7840
rect 14976 7828 14982 7880
rect 15396 7868 15424 7976
rect 15933 7871 15991 7877
rect 15933 7868 15945 7871
rect 15396 7840 15945 7868
rect 15933 7837 15945 7840
rect 15979 7837 15991 7871
rect 15933 7831 15991 7837
rect 16298 7828 16304 7880
rect 16356 7868 16362 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 16356 7840 17785 7868
rect 16356 7828 16362 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 18230 7868 18236 7880
rect 18191 7840 18236 7868
rect 17773 7831 17831 7837
rect 18230 7828 18236 7840
rect 18288 7868 18294 7880
rect 18509 7871 18567 7877
rect 18509 7868 18521 7871
rect 18288 7840 18521 7868
rect 18288 7828 18294 7840
rect 18509 7837 18521 7840
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 12544 7772 12940 7800
rect 13906 7760 13912 7812
rect 13964 7800 13970 7812
rect 15746 7800 15752 7812
rect 13964 7772 15752 7800
rect 13964 7760 13970 7772
rect 15746 7760 15752 7772
rect 15804 7760 15810 7812
rect 17528 7803 17586 7809
rect 17528 7769 17540 7803
rect 17574 7800 17586 7803
rect 18414 7800 18420 7812
rect 17574 7772 18420 7800
rect 17574 7769 17586 7772
rect 17528 7763 17586 7769
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 20993 7803 21051 7809
rect 20993 7769 21005 7803
rect 21039 7800 21051 7803
rect 21542 7800 21548 7812
rect 21039 7772 21548 7800
rect 21039 7769 21051 7772
rect 20993 7763 21051 7769
rect 21542 7760 21548 7772
rect 21600 7760 21606 7812
rect 13541 7735 13599 7741
rect 13541 7732 13553 7735
rect 11348 7704 13553 7732
rect 11241 7695 11299 7701
rect 13541 7701 13553 7704
rect 13587 7701 13599 7735
rect 13541 7695 13599 7701
rect 15013 7735 15071 7741
rect 15013 7701 15025 7735
rect 15059 7732 15071 7735
rect 16022 7732 16028 7744
rect 15059 7704 16028 7732
rect 15059 7701 15071 7704
rect 15013 7695 15071 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 16114 7692 16120 7744
rect 16172 7732 16178 7744
rect 18049 7735 18107 7741
rect 18049 7732 18061 7735
rect 16172 7704 18061 7732
rect 16172 7692 16178 7704
rect 18049 7701 18061 7704
rect 18095 7701 18107 7735
rect 18049 7695 18107 7701
rect 18966 7692 18972 7744
rect 19024 7732 19030 7744
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 19024 7704 19257 7732
rect 19024 7692 19030 7704
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 21358 7732 21364 7744
rect 21319 7704 21364 7732
rect 19245 7695 19303 7701
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 2682 7488 2688 7540
rect 2740 7528 2746 7540
rect 2774 7528 2780 7540
rect 2740 7500 2780 7528
rect 2740 7488 2746 7500
rect 2774 7488 2780 7500
rect 2832 7488 2838 7540
rect 4249 7531 4307 7537
rect 4249 7497 4261 7531
rect 4295 7528 4307 7531
rect 4430 7528 4436 7540
rect 4295 7500 4436 7528
rect 4295 7497 4307 7500
rect 4249 7491 4307 7497
rect 4430 7488 4436 7500
rect 4488 7488 4494 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 5537 7531 5595 7537
rect 5537 7528 5549 7531
rect 5500 7500 5549 7528
rect 5500 7488 5506 7500
rect 5537 7497 5549 7500
rect 5583 7497 5595 7531
rect 5537 7491 5595 7497
rect 5994 7488 6000 7540
rect 6052 7528 6058 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 6052 7500 6377 7528
rect 6052 7488 6058 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6638 7488 6644 7540
rect 6696 7528 6702 7540
rect 6733 7531 6791 7537
rect 6733 7528 6745 7531
rect 6696 7500 6745 7528
rect 6696 7488 6702 7500
rect 6733 7497 6745 7500
rect 6779 7497 6791 7531
rect 6733 7491 6791 7497
rect 7098 7488 7104 7540
rect 7156 7528 7162 7540
rect 8478 7528 8484 7540
rect 7156 7500 8484 7528
rect 7156 7488 7162 7500
rect 8478 7488 8484 7500
rect 8536 7488 8542 7540
rect 9122 7488 9128 7540
rect 9180 7528 9186 7540
rect 9861 7531 9919 7537
rect 9861 7528 9873 7531
rect 9180 7500 9873 7528
rect 9180 7488 9186 7500
rect 9861 7497 9873 7500
rect 9907 7497 9919 7531
rect 9861 7491 9919 7497
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7497 10287 7531
rect 10229 7491 10287 7497
rect 1394 7420 1400 7472
rect 1452 7460 1458 7472
rect 2010 7463 2068 7469
rect 2010 7460 2022 7463
rect 1452 7432 2022 7460
rect 1452 7420 1458 7432
rect 2010 7429 2022 7432
rect 2056 7429 2068 7463
rect 2010 7423 2068 7429
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4617 7463 4675 7469
rect 4617 7460 4629 7463
rect 4212 7432 4629 7460
rect 4212 7420 4218 7432
rect 4617 7429 4629 7432
rect 4663 7429 4675 7463
rect 4617 7423 4675 7429
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 7190 7460 7196 7472
rect 5675 7432 7196 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 7190 7420 7196 7432
rect 7248 7420 7254 7472
rect 10244 7460 10272 7491
rect 11238 7488 11244 7540
rect 11296 7528 11302 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11296 7500 11529 7528
rect 11296 7488 11302 7500
rect 11517 7497 11529 7500
rect 11563 7528 11575 7531
rect 11974 7528 11980 7540
rect 11563 7500 11980 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 13906 7528 13912 7540
rect 12406 7500 13912 7528
rect 12406 7460 12434 7500
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 16942 7528 16948 7540
rect 16715 7500 16948 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17773 7531 17831 7537
rect 17773 7497 17785 7531
rect 17819 7497 17831 7531
rect 17773 7491 17831 7497
rect 10244 7432 12434 7460
rect 12652 7463 12710 7469
rect 12652 7429 12664 7463
rect 12698 7460 12710 7463
rect 15102 7460 15108 7472
rect 12698 7432 15108 7460
rect 12698 7429 12710 7432
rect 12652 7423 12710 7429
rect 15102 7420 15108 7432
rect 15160 7420 15166 7472
rect 15390 7463 15448 7469
rect 15390 7429 15402 7463
rect 15436 7460 15448 7463
rect 15654 7460 15660 7472
rect 15436 7432 15660 7460
rect 15436 7429 15448 7432
rect 15390 7423 15448 7429
rect 15654 7420 15660 7432
rect 15712 7420 15718 7472
rect 16022 7420 16028 7472
rect 16080 7460 16086 7472
rect 17788 7460 17816 7491
rect 18874 7488 18880 7540
rect 18932 7528 18938 7540
rect 18969 7531 19027 7537
rect 18969 7528 18981 7531
rect 18932 7500 18981 7528
rect 18932 7488 18938 7500
rect 18969 7497 18981 7500
rect 19015 7497 19027 7531
rect 18969 7491 19027 7497
rect 21266 7460 21272 7472
rect 16080 7432 17632 7460
rect 17788 7432 21272 7460
rect 16080 7420 16086 7432
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 3326 7392 3332 7404
rect 2464 7364 3332 7392
rect 2464 7352 2470 7364
rect 3326 7352 3332 7364
rect 3384 7392 3390 7404
rect 4709 7395 4767 7401
rect 4709 7392 4721 7395
rect 3384 7364 4721 7392
rect 3384 7352 3390 7364
rect 4709 7361 4721 7364
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 7561 7395 7619 7401
rect 7561 7392 7573 7395
rect 5224 7364 7573 7392
rect 5224 7352 5230 7364
rect 7561 7361 7573 7364
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 8104 7395 8162 7401
rect 8104 7361 8116 7395
rect 8150 7392 8162 7395
rect 9306 7392 9312 7404
rect 8150 7364 9312 7392
rect 8150 7361 8162 7364
rect 8104 7355 8162 7361
rect 9306 7352 9312 7364
rect 9364 7352 9370 7404
rect 9490 7352 9496 7404
rect 9548 7392 9554 7404
rect 10505 7395 10563 7401
rect 10505 7392 10517 7395
rect 9548 7364 10517 7392
rect 9548 7352 9554 7364
rect 10505 7361 10517 7364
rect 10551 7361 10563 7395
rect 10505 7355 10563 7361
rect 11054 7352 11060 7404
rect 11112 7392 11118 7404
rect 11422 7392 11428 7404
rect 11112 7364 11428 7392
rect 11112 7352 11118 7364
rect 11422 7352 11428 7364
rect 11480 7392 11486 7404
rect 11882 7392 11888 7404
rect 11480 7364 11888 7392
rect 11480 7352 11486 7364
rect 11882 7352 11888 7364
rect 11940 7352 11946 7404
rect 12802 7352 12808 7404
rect 12860 7392 12866 7404
rect 12860 7364 12940 7392
rect 12860 7352 12866 7364
rect 1762 7324 1768 7336
rect 1723 7296 1768 7324
rect 1762 7284 1768 7296
rect 1820 7284 1826 7336
rect 3973 7327 4031 7333
rect 3973 7293 3985 7327
rect 4019 7293 4031 7327
rect 4798 7324 4804 7336
rect 4759 7296 4804 7324
rect 3973 7287 4031 7293
rect 3988 7256 4016 7287
rect 4798 7284 4804 7296
rect 4856 7284 4862 7336
rect 5445 7327 5503 7333
rect 5445 7293 5457 7327
rect 5491 7324 5503 7327
rect 6638 7324 6644 7336
rect 5491 7296 6644 7324
rect 5491 7293 5503 7296
rect 5445 7287 5503 7293
rect 6638 7284 6644 7296
rect 6696 7284 6702 7336
rect 6730 7284 6736 7336
rect 6788 7324 6794 7336
rect 6825 7327 6883 7333
rect 6825 7324 6837 7327
rect 6788 7296 6837 7324
rect 6788 7284 6794 7296
rect 6825 7293 6837 7296
rect 6871 7293 6883 7327
rect 6825 7287 6883 7293
rect 6914 7284 6920 7336
rect 6972 7324 6978 7336
rect 7837 7327 7895 7333
rect 6972 7296 7017 7324
rect 6972 7284 6978 7296
rect 7837 7293 7849 7327
rect 7883 7293 7895 7327
rect 7837 7287 7895 7293
rect 9585 7327 9643 7333
rect 9585 7293 9597 7327
rect 9631 7293 9643 7327
rect 9766 7324 9772 7336
rect 9727 7296 9772 7324
rect 9585 7287 9643 7293
rect 7098 7256 7104 7268
rect 3988 7228 7104 7256
rect 7098 7216 7104 7228
rect 7156 7216 7162 7268
rect 1489 7191 1547 7197
rect 1489 7157 1501 7191
rect 1535 7188 1547 7191
rect 1578 7188 1584 7200
rect 1535 7160 1584 7188
rect 1535 7157 1547 7160
rect 1489 7151 1547 7157
rect 1578 7148 1584 7160
rect 1636 7148 1642 7200
rect 3142 7188 3148 7200
rect 3103 7160 3148 7188
rect 3142 7148 3148 7160
rect 3200 7148 3206 7200
rect 3513 7191 3571 7197
rect 3513 7157 3525 7191
rect 3559 7188 3571 7191
rect 4246 7188 4252 7200
rect 3559 7160 4252 7188
rect 3559 7157 3571 7160
rect 3513 7151 3571 7157
rect 4246 7148 4252 7160
rect 4304 7188 4310 7200
rect 5166 7188 5172 7200
rect 4304 7160 5172 7188
rect 4304 7148 4310 7160
rect 5166 7148 5172 7160
rect 5224 7148 5230 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 5997 7191 6055 7197
rect 5997 7188 6009 7191
rect 5684 7160 6009 7188
rect 5684 7148 5690 7160
rect 5997 7157 6009 7160
rect 6043 7157 6055 7191
rect 7374 7188 7380 7200
rect 7335 7160 7380 7188
rect 5997 7151 6055 7157
rect 7374 7148 7380 7160
rect 7432 7148 7438 7200
rect 7852 7188 7880 7287
rect 8938 7216 8944 7268
rect 8996 7216 9002 7268
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7256 9275 7259
rect 9600 7256 9628 7287
rect 9766 7284 9772 7296
rect 9824 7284 9830 7336
rect 12912 7333 12940 7364
rect 13078 7352 13084 7404
rect 13136 7392 13142 7404
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13136 7364 13369 7392
rect 13136 7352 13142 7364
rect 13357 7361 13369 7364
rect 13403 7361 13415 7395
rect 15933 7395 15991 7401
rect 15933 7392 15945 7395
rect 13357 7355 13415 7361
rect 13924 7364 15945 7392
rect 12897 7327 12955 7333
rect 12897 7293 12909 7327
rect 12943 7324 12955 7327
rect 13630 7324 13636 7336
rect 12943 7296 13636 7324
rect 12943 7293 12955 7296
rect 12897 7287 12955 7293
rect 13630 7284 13636 7296
rect 13688 7284 13694 7336
rect 9950 7256 9956 7268
rect 9263 7228 9956 7256
rect 9263 7225 9275 7228
rect 9217 7219 9275 7225
rect 9950 7216 9956 7228
rect 10008 7216 10014 7268
rect 10134 7216 10140 7268
rect 10192 7256 10198 7268
rect 11882 7256 11888 7268
rect 10192 7228 11888 7256
rect 10192 7216 10198 7228
rect 11882 7216 11888 7228
rect 11940 7216 11946 7268
rect 8018 7188 8024 7200
rect 7852 7160 8024 7188
rect 8018 7148 8024 7160
rect 8076 7188 8082 7200
rect 8956 7188 8984 7216
rect 8076 7160 8984 7188
rect 8076 7148 8082 7160
rect 11054 7148 11060 7200
rect 11112 7188 11118 7200
rect 11149 7191 11207 7197
rect 11149 7188 11161 7191
rect 11112 7160 11161 7188
rect 11112 7148 11118 7160
rect 11149 7157 11161 7160
rect 11195 7157 11207 7191
rect 11149 7151 11207 7157
rect 12250 7148 12256 7200
rect 12308 7188 12314 7200
rect 13924 7188 13952 7364
rect 15933 7361 15945 7364
rect 15979 7361 15991 7395
rect 15933 7355 15991 7361
rect 16390 7352 16396 7404
rect 16448 7392 16454 7404
rect 17604 7401 17632 7432
rect 21266 7420 21272 7432
rect 21324 7420 21330 7472
rect 17313 7395 17371 7401
rect 17313 7392 17325 7395
rect 16448 7364 17325 7392
rect 16448 7352 16454 7364
rect 17313 7361 17325 7364
rect 17359 7361 17371 7395
rect 17313 7355 17371 7361
rect 17589 7395 17647 7401
rect 17589 7361 17601 7395
rect 17635 7361 17647 7395
rect 18690 7392 18696 7404
rect 18651 7364 18696 7392
rect 17589 7355 17647 7361
rect 18690 7352 18696 7364
rect 18748 7352 18754 7404
rect 18966 7352 18972 7404
rect 19024 7392 19030 7404
rect 19153 7395 19211 7401
rect 19153 7392 19165 7395
rect 19024 7364 19165 7392
rect 19024 7352 19030 7364
rect 19153 7361 19165 7364
rect 19199 7361 19211 7395
rect 19886 7392 19892 7404
rect 19847 7364 19892 7392
rect 19153 7355 19211 7361
rect 19886 7352 19892 7364
rect 19944 7352 19950 7404
rect 15657 7327 15715 7333
rect 15657 7293 15669 7327
rect 15703 7324 15715 7327
rect 16298 7324 16304 7336
rect 15703 7296 16304 7324
rect 15703 7293 15715 7296
rect 15657 7287 15715 7293
rect 16298 7284 16304 7296
rect 16356 7284 16362 7336
rect 17034 7284 17040 7336
rect 17092 7324 17098 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17092 7296 18061 7324
rect 17092 7284 17098 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 14001 7259 14059 7265
rect 14001 7225 14013 7259
rect 14047 7256 14059 7259
rect 14366 7256 14372 7268
rect 14047 7228 14372 7256
rect 14047 7225 14059 7228
rect 14001 7219 14059 7225
rect 14366 7216 14372 7228
rect 14424 7216 14430 7268
rect 16117 7259 16175 7265
rect 16117 7225 16129 7259
rect 16163 7256 16175 7259
rect 18506 7256 18512 7268
rect 16163 7228 18368 7256
rect 18467 7228 18512 7256
rect 16163 7225 16175 7228
rect 16117 7219 16175 7225
rect 14274 7188 14280 7200
rect 12308 7160 13952 7188
rect 14235 7160 14280 7188
rect 12308 7148 12314 7160
rect 14274 7148 14280 7160
rect 14332 7148 14338 7200
rect 18340 7188 18368 7228
rect 18506 7216 18512 7228
rect 18564 7216 18570 7268
rect 19518 7216 19524 7268
rect 19576 7256 19582 7268
rect 20165 7259 20223 7265
rect 20165 7256 20177 7259
rect 19576 7228 20177 7256
rect 19576 7216 19582 7228
rect 20165 7225 20177 7228
rect 20211 7225 20223 7259
rect 20165 7219 20223 7225
rect 18874 7188 18880 7200
rect 18340 7160 18880 7188
rect 18874 7148 18880 7160
rect 18932 7148 18938 7200
rect 19705 7191 19763 7197
rect 19705 7157 19717 7191
rect 19751 7188 19763 7191
rect 19794 7188 19800 7200
rect 19751 7160 19800 7188
rect 19751 7157 19763 7160
rect 19705 7151 19763 7157
rect 19794 7148 19800 7160
rect 19852 7148 19858 7200
rect 20438 7148 20444 7200
rect 20496 7188 20502 7200
rect 20533 7191 20591 7197
rect 20533 7188 20545 7191
rect 20496 7160 20545 7188
rect 20496 7148 20502 7160
rect 20533 7157 20545 7160
rect 20579 7157 20591 7191
rect 20990 7188 20996 7200
rect 20951 7160 20996 7188
rect 20533 7151 20591 7157
rect 20990 7148 20996 7160
rect 21048 7148 21054 7200
rect 21361 7191 21419 7197
rect 21361 7157 21373 7191
rect 21407 7188 21419 7191
rect 21450 7188 21456 7200
rect 21407 7160 21456 7188
rect 21407 7157 21419 7160
rect 21361 7151 21419 7157
rect 21450 7148 21456 7160
rect 21508 7148 21514 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 1394 6944 1400 6996
rect 1452 6984 1458 6996
rect 2038 6984 2044 6996
rect 1452 6956 2044 6984
rect 1452 6944 1458 6956
rect 2038 6944 2044 6956
rect 2096 6944 2102 6996
rect 2590 6944 2596 6996
rect 2648 6984 2654 6996
rect 3789 6987 3847 6993
rect 3789 6984 3801 6987
rect 2648 6956 3801 6984
rect 2648 6944 2654 6956
rect 3789 6953 3801 6956
rect 3835 6953 3847 6987
rect 3789 6947 3847 6953
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 5258 6984 5264 6996
rect 4120 6956 5264 6984
rect 4120 6944 4126 6956
rect 5258 6944 5264 6956
rect 5316 6984 5322 6996
rect 5534 6984 5540 6996
rect 5316 6956 5396 6984
rect 5495 6956 5540 6984
rect 5316 6944 5322 6956
rect 3142 6876 3148 6928
rect 3200 6916 3206 6928
rect 4801 6919 4859 6925
rect 3200 6888 4384 6916
rect 3200 6876 3206 6888
rect 4356 6857 4384 6888
rect 4801 6885 4813 6919
rect 4847 6885 4859 6919
rect 5368 6916 5396 6956
rect 5534 6944 5540 6956
rect 5592 6944 5598 6996
rect 8386 6944 8392 6996
rect 8444 6984 8450 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8444 6956 8953 6984
rect 8444 6944 8450 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 18690 6944 18696 6996
rect 18748 6984 18754 6996
rect 18785 6987 18843 6993
rect 18785 6984 18797 6987
rect 18748 6956 18797 6984
rect 18748 6944 18754 6956
rect 18785 6953 18797 6956
rect 18831 6953 18843 6987
rect 18785 6947 18843 6953
rect 6730 6916 6736 6928
rect 5368 6888 6736 6916
rect 4801 6879 4859 6885
rect 4341 6851 4399 6857
rect 4341 6817 4353 6851
rect 4387 6817 4399 6851
rect 4341 6811 4399 6817
rect 4522 6808 4528 6860
rect 4580 6848 4586 6860
rect 4816 6848 4844 6879
rect 6730 6876 6736 6888
rect 6788 6876 6794 6928
rect 7576 6888 7788 6916
rect 7576 6848 7604 6888
rect 4580 6820 4844 6848
rect 4908 6820 7604 6848
rect 7653 6851 7711 6857
rect 4580 6808 4586 6820
rect 1397 6783 1455 6789
rect 1397 6749 1409 6783
rect 1443 6780 1455 6783
rect 3237 6783 3295 6789
rect 1443 6752 1808 6780
rect 1443 6749 1455 6752
rect 1397 6743 1455 6749
rect 1780 6724 1808 6752
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 3970 6780 3976 6792
rect 3283 6752 3976 6780
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6780 4307 6783
rect 4908 6780 4936 6820
rect 7653 6817 7665 6851
rect 7699 6817 7711 6851
rect 7760 6848 7788 6888
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8481 6919 8539 6925
rect 8481 6916 8493 6919
rect 8352 6888 8493 6916
rect 8352 6876 8358 6888
rect 8481 6885 8493 6888
rect 8527 6916 8539 6919
rect 8570 6916 8576 6928
rect 8527 6888 8576 6916
rect 8527 6885 8539 6888
rect 8481 6879 8539 6885
rect 8570 6876 8576 6888
rect 8628 6876 8634 6928
rect 11422 6916 11428 6928
rect 10980 6888 11428 6916
rect 8662 6848 8668 6860
rect 7760 6820 8668 6848
rect 7653 6811 7711 6817
rect 4295 6752 4936 6780
rect 4985 6783 5043 6789
rect 4295 6749 4307 6752
rect 4249 6743 4307 6749
rect 4985 6749 4997 6783
rect 5031 6780 5043 6783
rect 5258 6780 5264 6792
rect 5031 6752 5264 6780
rect 5031 6749 5043 6752
rect 4985 6743 5043 6749
rect 5258 6740 5264 6752
rect 5316 6780 5322 6792
rect 6730 6780 6736 6792
rect 5316 6752 6736 6780
rect 5316 6740 5322 6752
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7006 6780 7012 6792
rect 6967 6752 7012 6780
rect 7006 6740 7012 6752
rect 7064 6740 7070 6792
rect 7668 6780 7696 6811
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 9306 6808 9312 6860
rect 9364 6848 9370 6860
rect 9493 6851 9551 6857
rect 9493 6848 9505 6851
rect 9364 6820 9505 6848
rect 9364 6808 9370 6820
rect 9493 6817 9505 6820
rect 9539 6817 9551 6851
rect 10594 6848 10600 6860
rect 9493 6811 9551 6817
rect 9784 6820 10456 6848
rect 10555 6820 10600 6848
rect 9784 6780 9812 6820
rect 9950 6780 9956 6792
rect 7668 6752 9812 6780
rect 9911 6752 9956 6780
rect 9950 6740 9956 6752
rect 10008 6740 10014 6792
rect 10428 6780 10456 6820
rect 10594 6808 10600 6820
rect 10652 6808 10658 6860
rect 10980 6780 11008 6888
rect 11422 6876 11428 6888
rect 11480 6876 11486 6928
rect 11057 6851 11115 6857
rect 11057 6817 11069 6851
rect 11103 6817 11115 6851
rect 11057 6811 11115 6817
rect 10428 6752 11008 6780
rect 11072 6780 11100 6811
rect 12434 6808 12440 6860
rect 12492 6848 12498 6860
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 12492 6820 12633 6848
rect 12492 6808 12498 6820
rect 12621 6817 12633 6820
rect 12667 6817 12679 6851
rect 13078 6848 13084 6860
rect 13039 6820 13084 6848
rect 12621 6811 12679 6817
rect 13078 6808 13084 6820
rect 13136 6808 13142 6860
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 18509 6851 18567 6857
rect 18509 6848 18521 6851
rect 18472 6820 18521 6848
rect 18472 6808 18478 6820
rect 18509 6817 18521 6820
rect 18555 6817 18567 6851
rect 20625 6851 20683 6857
rect 20625 6848 20637 6851
rect 18509 6811 18567 6817
rect 19444 6820 20637 6848
rect 19444 6792 19472 6820
rect 20625 6817 20637 6820
rect 20671 6817 20683 6851
rect 20625 6811 20683 6817
rect 11330 6780 11336 6792
rect 11072 6752 11192 6780
rect 11291 6752 11336 6780
rect 1664 6715 1722 6721
rect 1664 6681 1676 6715
rect 1710 6681 1722 6715
rect 1664 6675 1722 6681
rect 1688 6644 1716 6675
rect 1762 6672 1768 6724
rect 1820 6672 1826 6724
rect 3436 6684 7144 6712
rect 1854 6644 1860 6656
rect 1688 6616 1860 6644
rect 1854 6604 1860 6616
rect 1912 6604 1918 6656
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2682 6644 2688 6656
rect 2188 6616 2688 6644
rect 2188 6604 2194 6616
rect 2682 6604 2688 6616
rect 2740 6644 2746 6656
rect 3436 6653 3464 6684
rect 2777 6647 2835 6653
rect 2777 6644 2789 6647
rect 2740 6616 2789 6644
rect 2740 6604 2746 6616
rect 2777 6613 2789 6616
rect 2823 6613 2835 6647
rect 2777 6607 2835 6613
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6613 3479 6647
rect 3421 6607 3479 6613
rect 4157 6647 4215 6653
rect 4157 6613 4169 6647
rect 4203 6644 4215 6647
rect 4430 6644 4436 6656
rect 4203 6616 4436 6644
rect 4203 6613 4215 6616
rect 4157 6607 4215 6613
rect 4430 6604 4436 6616
rect 4488 6604 4494 6656
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 5166 6644 5172 6656
rect 4856 6616 5172 6644
rect 4856 6604 4862 6616
rect 5166 6604 5172 6616
rect 5224 6644 5230 6656
rect 5718 6644 5724 6656
rect 5224 6616 5724 6644
rect 5224 6604 5230 6616
rect 5718 6604 5724 6616
rect 5776 6604 5782 6656
rect 7116 6644 7144 6684
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 7745 6715 7803 6721
rect 7745 6712 7757 6715
rect 7248 6684 7757 6712
rect 7248 6672 7254 6684
rect 7745 6681 7757 6684
rect 7791 6712 7803 6715
rect 8110 6712 8116 6724
rect 7791 6684 8116 6712
rect 7791 6681 7803 6684
rect 7745 6675 7803 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 9766 6712 9772 6724
rect 8220 6684 9772 6712
rect 7466 6644 7472 6656
rect 7116 6616 7472 6644
rect 7466 6604 7472 6616
rect 7524 6604 7530 6656
rect 7834 6604 7840 6656
rect 7892 6644 7898 6656
rect 8220 6653 8248 6684
rect 9766 6672 9772 6684
rect 9824 6672 9830 6724
rect 11164 6712 11192 6752
rect 11330 6740 11336 6752
rect 11388 6740 11394 6792
rect 11974 6780 11980 6792
rect 11935 6752 11980 6780
rect 11974 6740 11980 6752
rect 12032 6740 12038 6792
rect 13357 6783 13415 6789
rect 13357 6749 13369 6783
rect 13403 6780 13415 6783
rect 13538 6780 13544 6792
rect 13403 6752 13544 6780
rect 13403 6749 13415 6752
rect 13357 6743 13415 6749
rect 13538 6740 13544 6752
rect 13596 6740 13602 6792
rect 13630 6740 13636 6792
rect 13688 6780 13694 6792
rect 14366 6789 14372 6792
rect 14093 6783 14151 6789
rect 14093 6780 14105 6783
rect 13688 6752 14105 6780
rect 13688 6740 13694 6752
rect 14093 6749 14105 6752
rect 14139 6749 14151 6783
rect 14360 6780 14372 6789
rect 14327 6752 14372 6780
rect 14093 6743 14151 6749
rect 14360 6743 14372 6752
rect 14366 6740 14372 6743
rect 14424 6740 14430 6792
rect 16209 6783 16267 6789
rect 16209 6749 16221 6783
rect 16255 6780 16267 6783
rect 16298 6780 16304 6792
rect 16255 6752 16304 6780
rect 16255 6749 16267 6752
rect 16209 6743 16267 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 17865 6783 17923 6789
rect 17865 6780 17877 6783
rect 17604 6752 17877 6780
rect 14274 6712 14280 6724
rect 11164 6684 14280 6712
rect 14274 6672 14280 6684
rect 14332 6672 14338 6724
rect 16476 6715 16534 6721
rect 16476 6681 16488 6715
rect 16522 6712 16534 6715
rect 16942 6712 16948 6724
rect 16522 6684 16948 6712
rect 16522 6681 16534 6684
rect 16476 6675 16534 6681
rect 16942 6672 16948 6684
rect 17000 6672 17006 6724
rect 8205 6647 8263 6653
rect 7892 6616 7937 6644
rect 7892 6604 7898 6616
rect 8205 6613 8217 6647
rect 8251 6613 8263 6647
rect 8205 6607 8263 6613
rect 8294 6604 8300 6656
rect 8352 6644 8358 6656
rect 9309 6647 9367 6653
rect 9309 6644 9321 6647
rect 8352 6616 9321 6644
rect 8352 6604 8358 6616
rect 9309 6613 9321 6616
rect 9355 6613 9367 6647
rect 9309 6607 9367 6613
rect 9398 6604 9404 6656
rect 9456 6644 9462 6656
rect 9456 6616 9501 6644
rect 9456 6604 9462 6616
rect 10778 6604 10784 6656
rect 10836 6644 10842 6656
rect 11238 6644 11244 6656
rect 10836 6616 11244 6644
rect 10836 6604 10842 6616
rect 11238 6604 11244 6616
rect 11296 6604 11302 6656
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6644 11759 6647
rect 11790 6644 11796 6656
rect 11747 6616 11796 6644
rect 11747 6613 11759 6616
rect 11701 6607 11759 6613
rect 11790 6604 11796 6616
rect 11848 6604 11854 6656
rect 13262 6644 13268 6656
rect 13223 6616 13268 6644
rect 13262 6604 13268 6616
rect 13320 6604 13326 6656
rect 13725 6647 13783 6653
rect 13725 6613 13737 6647
rect 13771 6644 13783 6647
rect 14458 6644 14464 6656
rect 13771 6616 14464 6644
rect 13771 6613 13783 6616
rect 13725 6607 13783 6613
rect 14458 6604 14464 6616
rect 14516 6604 14522 6656
rect 15470 6644 15476 6656
rect 15431 6616 15476 6644
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 15746 6644 15752 6656
rect 15707 6616 15752 6644
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16390 6604 16396 6656
rect 16448 6644 16454 6656
rect 17604 6653 17632 6752
rect 17865 6749 17877 6752
rect 17911 6749 17923 6783
rect 19426 6780 19432 6792
rect 19387 6752 19432 6780
rect 17865 6743 17923 6749
rect 19426 6740 19432 6752
rect 19484 6740 19490 6792
rect 19886 6780 19892 6792
rect 19847 6752 19892 6780
rect 19886 6740 19892 6752
rect 19944 6740 19950 6792
rect 20165 6783 20223 6789
rect 20165 6749 20177 6783
rect 20211 6780 20223 6783
rect 20254 6780 20260 6792
rect 20211 6752 20260 6780
rect 20211 6749 20223 6752
rect 20165 6743 20223 6749
rect 20254 6740 20260 6752
rect 20312 6740 20318 6792
rect 20898 6712 20904 6724
rect 20364 6684 20904 6712
rect 17589 6647 17647 6653
rect 17589 6644 17601 6647
rect 16448 6616 17601 6644
rect 16448 6604 16454 6616
rect 17589 6613 17601 6616
rect 17635 6613 17647 6647
rect 17589 6607 17647 6613
rect 17678 6604 17684 6656
rect 17736 6644 17742 6656
rect 19245 6647 19303 6653
rect 19245 6644 19257 6647
rect 17736 6616 19257 6644
rect 17736 6604 17742 6616
rect 19245 6613 19257 6616
rect 19291 6613 19303 6647
rect 19702 6644 19708 6656
rect 19663 6616 19708 6644
rect 19245 6607 19303 6613
rect 19702 6604 19708 6616
rect 19760 6604 19766 6656
rect 20364 6653 20392 6684
rect 20898 6672 20904 6684
rect 20956 6672 20962 6724
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6613 20407 6647
rect 20349 6607 20407 6613
rect 20806 6604 20812 6656
rect 20864 6644 20870 6656
rect 20993 6647 21051 6653
rect 20993 6644 21005 6647
rect 20864 6616 21005 6644
rect 20864 6604 20870 6616
rect 20993 6613 21005 6616
rect 21039 6613 21051 6647
rect 20993 6607 21051 6613
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 1670 6440 1676 6452
rect 1631 6412 1676 6440
rect 1670 6400 1676 6412
rect 1728 6400 1734 6452
rect 2314 6440 2320 6452
rect 2275 6412 2320 6440
rect 2314 6400 2320 6412
rect 2372 6400 2378 6452
rect 7374 6440 7380 6452
rect 2746 6412 7380 6440
rect 2225 6375 2283 6381
rect 2225 6341 2237 6375
rect 2271 6372 2283 6375
rect 2746 6372 2774 6412
rect 7374 6400 7380 6412
rect 7432 6400 7438 6452
rect 8202 6440 8208 6452
rect 7484 6412 8208 6440
rect 2271 6344 2774 6372
rect 2271 6341 2283 6344
rect 2225 6335 2283 6341
rect 3418 6332 3424 6384
rect 3476 6332 3482 6384
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 7484 6372 7512 6412
rect 8202 6400 8208 6412
rect 8260 6400 8266 6452
rect 9674 6400 9680 6452
rect 9732 6440 9738 6452
rect 9769 6443 9827 6449
rect 9769 6440 9781 6443
rect 9732 6412 9781 6440
rect 9732 6400 9738 6412
rect 9769 6409 9781 6412
rect 9815 6440 9827 6443
rect 10042 6440 10048 6452
rect 9815 6412 10048 6440
rect 9815 6409 9827 6412
rect 9769 6403 9827 6409
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 11057 6443 11115 6449
rect 11057 6409 11069 6443
rect 11103 6409 11115 6443
rect 11057 6403 11115 6409
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6440 12311 6443
rect 13078 6440 13084 6452
rect 12299 6412 13084 6440
rect 12299 6409 12311 6412
rect 12253 6403 12311 6409
rect 6788 6344 7512 6372
rect 6788 6332 6794 6344
rect 7834 6332 7840 6384
rect 7892 6372 7898 6384
rect 11072 6372 11100 6403
rect 13078 6400 13084 6412
rect 13136 6400 13142 6452
rect 14458 6440 14464 6452
rect 14419 6412 14464 6440
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 14553 6443 14611 6449
rect 14553 6409 14565 6443
rect 14599 6440 14611 6443
rect 15746 6440 15752 6452
rect 14599 6412 15752 6440
rect 14599 6409 14611 6412
rect 14553 6403 14611 6409
rect 15746 6400 15752 6412
rect 15804 6400 15810 6452
rect 15933 6443 15991 6449
rect 15933 6409 15945 6443
rect 15979 6440 15991 6443
rect 16669 6443 16727 6449
rect 16669 6440 16681 6443
rect 15979 6412 16681 6440
rect 15979 6409 15991 6412
rect 15933 6403 15991 6409
rect 16669 6409 16681 6412
rect 16715 6409 16727 6443
rect 17034 6440 17040 6452
rect 16995 6412 17040 6440
rect 16669 6403 16727 6409
rect 17034 6400 17040 6412
rect 17092 6400 17098 6452
rect 17126 6400 17132 6452
rect 17184 6440 17190 6452
rect 17865 6443 17923 6449
rect 17184 6412 17229 6440
rect 17184 6400 17190 6412
rect 17865 6409 17877 6443
rect 17911 6409 17923 6443
rect 18138 6440 18144 6452
rect 18099 6412 18144 6440
rect 17865 6403 17923 6409
rect 17770 6372 17776 6384
rect 7892 6344 10824 6372
rect 11072 6344 17776 6372
rect 7892 6332 7898 6344
rect 1486 6304 1492 6316
rect 1447 6276 1492 6304
rect 1486 6264 1492 6276
rect 1544 6264 1550 6316
rect 3436 6304 3464 6332
rect 4074 6307 4132 6313
rect 4074 6304 4086 6307
rect 2148 6276 4086 6304
rect 2148 6245 2176 6276
rect 4074 6273 4086 6276
rect 4120 6304 4132 6307
rect 4341 6307 4399 6313
rect 4120 6276 4292 6304
rect 4120 6273 4132 6276
rect 4074 6267 4132 6273
rect 2133 6239 2191 6245
rect 2133 6205 2145 6239
rect 2179 6205 2191 6239
rect 2133 6199 2191 6205
rect 2682 6196 2688 6248
rect 2740 6236 2746 6248
rect 3326 6236 3332 6248
rect 2740 6208 3332 6236
rect 2740 6196 2746 6208
rect 3326 6196 3332 6208
rect 3384 6196 3390 6248
rect 4264 6236 4292 6276
rect 4341 6273 4353 6307
rect 4387 6304 4399 6307
rect 4798 6304 4804 6316
rect 4387 6276 4804 6304
rect 4387 6273 4399 6276
rect 4341 6267 4399 6273
rect 4798 6264 4804 6276
rect 4856 6264 4862 6316
rect 5741 6307 5799 6313
rect 5741 6273 5753 6307
rect 5787 6304 5799 6307
rect 6362 6304 6368 6316
rect 5787 6276 6368 6304
rect 5787 6273 5799 6276
rect 5741 6267 5799 6273
rect 6362 6264 6368 6276
rect 6420 6264 6426 6316
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6989 6307 7047 6313
rect 6989 6304 7001 6307
rect 6604 6276 7001 6304
rect 6604 6264 6610 6276
rect 6989 6273 7001 6276
rect 7035 6273 7047 6307
rect 6989 6267 7047 6273
rect 7282 6264 7288 6316
rect 7340 6304 7346 6316
rect 8645 6307 8703 6313
rect 8645 6304 8657 6307
rect 7340 6276 8657 6304
rect 7340 6264 7346 6276
rect 8645 6273 8657 6276
rect 8691 6273 8703 6307
rect 8645 6267 8703 6273
rect 9122 6264 9128 6316
rect 9180 6304 9186 6316
rect 10689 6307 10747 6313
rect 10689 6304 10701 6307
rect 9180 6276 10701 6304
rect 9180 6264 9186 6276
rect 10689 6273 10701 6276
rect 10735 6273 10747 6307
rect 10796 6304 10824 6344
rect 17770 6332 17776 6344
rect 17828 6332 17834 6384
rect 17880 6372 17908 6403
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 18230 6400 18236 6452
rect 18288 6440 18294 6452
rect 19061 6443 19119 6449
rect 19061 6440 19073 6443
rect 18288 6412 19073 6440
rect 18288 6400 18294 6412
rect 19061 6409 19073 6412
rect 19107 6409 19119 6443
rect 19061 6403 19119 6409
rect 19150 6400 19156 6452
rect 19208 6440 19214 6452
rect 19978 6440 19984 6452
rect 19208 6412 19840 6440
rect 19939 6412 19984 6440
rect 19208 6400 19214 6412
rect 17880 6344 19748 6372
rect 13078 6304 13084 6316
rect 10796 6276 13084 6304
rect 10689 6267 10747 6273
rect 13078 6264 13084 6276
rect 13136 6264 13142 6316
rect 13377 6307 13435 6313
rect 13377 6273 13389 6307
rect 13423 6304 13435 6307
rect 14734 6304 14740 6316
rect 13423 6276 14740 6304
rect 13423 6273 13435 6276
rect 13377 6267 13435 6273
rect 14734 6264 14740 6276
rect 14792 6264 14798 6316
rect 16390 6304 16396 6316
rect 15764 6276 16396 6304
rect 5994 6236 6000 6248
rect 4264 6208 4660 6236
rect 5955 6208 6000 6236
rect 1854 6128 1860 6180
rect 1912 6168 1918 6180
rect 2590 6168 2596 6180
rect 1912 6140 2596 6168
rect 1912 6128 1918 6140
rect 2590 6128 2596 6140
rect 2648 6168 2654 6180
rect 4632 6177 4660 6208
rect 5994 6196 6000 6208
rect 6052 6236 6058 6248
rect 6733 6239 6791 6245
rect 6733 6236 6745 6239
rect 6052 6208 6745 6236
rect 6052 6196 6058 6208
rect 6733 6205 6745 6208
rect 6779 6205 6791 6239
rect 8018 6236 8024 6248
rect 6733 6199 6791 6205
rect 7760 6208 8024 6236
rect 2961 6171 3019 6177
rect 2961 6168 2973 6171
rect 2648 6140 2973 6168
rect 2648 6128 2654 6140
rect 2961 6137 2973 6140
rect 3007 6137 3019 6171
rect 2961 6131 3019 6137
rect 4617 6171 4675 6177
rect 4617 6137 4629 6171
rect 4663 6137 4675 6171
rect 4617 6131 4675 6137
rect 2682 6100 2688 6112
rect 2643 6072 2688 6100
rect 2682 6060 2688 6072
rect 2740 6060 2746 6112
rect 3142 6060 3148 6112
rect 3200 6100 3206 6112
rect 5350 6100 5356 6112
rect 3200 6072 5356 6100
rect 3200 6060 3206 6072
rect 5350 6060 5356 6072
rect 5408 6060 5414 6112
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 5776 6072 6377 6100
rect 5776 6060 5782 6072
rect 6365 6069 6377 6072
rect 6411 6100 6423 6103
rect 6454 6100 6460 6112
rect 6411 6072 6460 6100
rect 6411 6069 6423 6072
rect 6365 6063 6423 6069
rect 6454 6060 6460 6072
rect 6512 6060 6518 6112
rect 6748 6100 6776 6199
rect 7760 6100 7788 6208
rect 8018 6196 8024 6208
rect 8076 6236 8082 6248
rect 8389 6239 8447 6245
rect 8389 6236 8401 6239
rect 8076 6208 8401 6236
rect 8076 6196 8082 6208
rect 8389 6205 8401 6208
rect 8435 6205 8447 6239
rect 8389 6199 8447 6205
rect 9490 6196 9496 6248
rect 9548 6236 9554 6248
rect 10413 6239 10471 6245
rect 10413 6236 10425 6239
rect 9548 6208 10425 6236
rect 9548 6196 9554 6208
rect 10413 6205 10425 6208
rect 10459 6205 10471 6239
rect 10413 6199 10471 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6205 10655 6239
rect 10597 6199 10655 6205
rect 11977 6239 12035 6245
rect 11977 6205 11989 6239
rect 12023 6236 12035 6239
rect 12342 6236 12348 6248
rect 12023 6208 12348 6236
rect 12023 6205 12035 6208
rect 11977 6199 12035 6205
rect 10134 6128 10140 6180
rect 10192 6168 10198 6180
rect 10612 6168 10640 6199
rect 12342 6196 12348 6208
rect 12400 6196 12406 6248
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14369 6239 14427 6245
rect 13688 6208 13781 6236
rect 13688 6196 13694 6208
rect 14369 6205 14381 6239
rect 14415 6236 14427 6239
rect 15470 6236 15476 6248
rect 14415 6208 15476 6236
rect 14415 6205 14427 6208
rect 14369 6199 14427 6205
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 15764 6245 15792 6276
rect 16390 6264 16396 6276
rect 16448 6264 16454 6316
rect 16850 6264 16856 6316
rect 16908 6304 16914 6316
rect 16908 6276 17264 6304
rect 16908 6264 16914 6276
rect 17236 6248 17264 6276
rect 17310 6264 17316 6316
rect 17368 6304 17374 6316
rect 17681 6307 17739 6313
rect 17681 6304 17693 6307
rect 17368 6276 17693 6304
rect 17368 6264 17374 6276
rect 17681 6273 17693 6276
rect 17727 6273 17739 6307
rect 17681 6267 17739 6273
rect 17862 6264 17868 6316
rect 17920 6304 17926 6316
rect 18325 6307 18383 6313
rect 18325 6304 18337 6307
rect 17920 6276 18337 6304
rect 17920 6264 17926 6276
rect 18325 6273 18337 6276
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 18414 6264 18420 6316
rect 18472 6304 18478 6316
rect 19720 6313 19748 6344
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18472 6276 18613 6304
rect 18472 6264 18478 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 18601 6267 18659 6273
rect 19245 6307 19303 6313
rect 19245 6273 19257 6307
rect 19291 6304 19303 6307
rect 19705 6307 19763 6313
rect 19291 6276 19380 6304
rect 19291 6273 19303 6276
rect 19245 6267 19303 6273
rect 15749 6239 15807 6245
rect 15749 6205 15761 6239
rect 15795 6205 15807 6239
rect 15749 6199 15807 6205
rect 15841 6239 15899 6245
rect 15841 6205 15853 6239
rect 15887 6236 15899 6239
rect 16942 6236 16948 6248
rect 15887 6208 16948 6236
rect 15887 6205 15899 6208
rect 15841 6199 15899 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17218 6196 17224 6248
rect 17276 6236 17282 6248
rect 17276 6208 17369 6236
rect 17276 6196 17282 6208
rect 18506 6196 18512 6248
rect 18564 6236 18570 6248
rect 19150 6236 19156 6248
rect 18564 6208 19156 6236
rect 18564 6196 18570 6208
rect 19150 6196 19156 6208
rect 19208 6196 19214 6248
rect 10192 6140 10640 6168
rect 10192 6128 10198 6140
rect 6748 6072 7788 6100
rect 7834 6060 7840 6112
rect 7892 6100 7898 6112
rect 8113 6103 8171 6109
rect 8113 6100 8125 6103
rect 7892 6072 8125 6100
rect 7892 6060 7898 6072
rect 8113 6069 8125 6072
rect 8159 6069 8171 6103
rect 8113 6063 8171 6069
rect 8662 6060 8668 6112
rect 8720 6100 8726 6112
rect 11790 6100 11796 6112
rect 8720 6072 11796 6100
rect 8720 6060 8726 6072
rect 11790 6060 11796 6072
rect 11848 6060 11854 6112
rect 12710 6060 12716 6112
rect 12768 6100 12774 6112
rect 13648 6100 13676 6196
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 15197 6171 15255 6177
rect 15197 6168 15209 6171
rect 13780 6140 15209 6168
rect 13780 6128 13786 6140
rect 15197 6137 15209 6140
rect 15243 6137 15255 6171
rect 15197 6131 15255 6137
rect 15286 6128 15292 6180
rect 15344 6168 15350 6180
rect 19352 6168 19380 6276
rect 19705 6273 19717 6307
rect 19751 6273 19763 6307
rect 19812 6304 19840 6412
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 20165 6307 20223 6313
rect 20165 6304 20177 6307
rect 19812 6276 20177 6304
rect 19705 6267 19763 6273
rect 20165 6273 20177 6276
rect 20211 6304 20223 6307
rect 20806 6304 20812 6316
rect 20211 6276 20812 6304
rect 20211 6273 20223 6276
rect 20165 6267 20223 6273
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 20901 6307 20959 6313
rect 20901 6273 20913 6307
rect 20947 6304 20959 6307
rect 21082 6304 21088 6316
rect 20947 6276 21088 6304
rect 20947 6273 20959 6276
rect 20901 6267 20959 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 21361 6307 21419 6313
rect 21361 6273 21373 6307
rect 21407 6304 21419 6307
rect 21450 6304 21456 6316
rect 21407 6276 21456 6304
rect 21407 6273 21419 6276
rect 21361 6267 21419 6273
rect 21450 6264 21456 6276
rect 21508 6264 21514 6316
rect 15344 6140 19380 6168
rect 15344 6128 15350 6140
rect 12768 6072 13676 6100
rect 14921 6103 14979 6109
rect 12768 6060 12774 6072
rect 14921 6069 14933 6103
rect 14967 6100 14979 6103
rect 15010 6100 15016 6112
rect 14967 6072 15016 6100
rect 14967 6069 14979 6072
rect 14921 6063 14979 6069
rect 15010 6060 15016 6072
rect 15068 6060 15074 6112
rect 16301 6103 16359 6109
rect 16301 6069 16313 6103
rect 16347 6100 16359 6103
rect 18690 6100 18696 6112
rect 16347 6072 18696 6100
rect 16347 6069 16359 6072
rect 16301 6063 16359 6069
rect 18690 6060 18696 6072
rect 18748 6060 18754 6112
rect 18785 6103 18843 6109
rect 18785 6069 18797 6103
rect 18831 6100 18843 6103
rect 18966 6100 18972 6112
rect 18831 6072 18972 6100
rect 18831 6069 18843 6072
rect 18785 6063 18843 6069
rect 18966 6060 18972 6072
rect 19024 6060 19030 6112
rect 19521 6103 19579 6109
rect 19521 6069 19533 6103
rect 19567 6100 19579 6103
rect 19978 6100 19984 6112
rect 19567 6072 19984 6100
rect 19567 6069 19579 6072
rect 19521 6063 19579 6069
rect 19978 6060 19984 6072
rect 20036 6060 20042 6112
rect 20717 6103 20775 6109
rect 20717 6069 20729 6103
rect 20763 6100 20775 6103
rect 20806 6100 20812 6112
rect 20763 6072 20812 6100
rect 20763 6069 20775 6072
rect 20717 6063 20775 6069
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 21174 6100 21180 6112
rect 21135 6072 21180 6100
rect 21174 6060 21180 6072
rect 21232 6060 21238 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 3142 5896 3148 5908
rect 2455 5868 3148 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3789 5899 3847 5905
rect 3789 5865 3801 5899
rect 3835 5896 3847 5899
rect 3878 5896 3884 5908
rect 3835 5868 3884 5896
rect 3835 5865 3847 5868
rect 3789 5859 3847 5865
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 4338 5856 4344 5908
rect 4396 5856 4402 5908
rect 5721 5899 5779 5905
rect 5721 5865 5733 5899
rect 5767 5896 5779 5899
rect 5994 5896 6000 5908
rect 5767 5868 6000 5896
rect 5767 5865 5779 5868
rect 5721 5859 5779 5865
rect 5994 5856 6000 5868
rect 6052 5856 6058 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7650 5896 7656 5908
rect 6972 5868 7656 5896
rect 6972 5856 6978 5868
rect 7650 5856 7656 5868
rect 7708 5856 7714 5908
rect 9125 5899 9183 5905
rect 9125 5865 9137 5899
rect 9171 5896 9183 5899
rect 10594 5896 10600 5908
rect 9171 5868 10600 5896
rect 9171 5865 9183 5868
rect 9125 5859 9183 5865
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 11882 5856 11888 5908
rect 11940 5896 11946 5908
rect 13357 5899 13415 5905
rect 13357 5896 13369 5899
rect 11940 5868 13369 5896
rect 11940 5856 11946 5868
rect 13357 5865 13369 5868
rect 13403 5865 13415 5899
rect 14734 5896 14740 5908
rect 14695 5868 14740 5896
rect 13357 5859 13415 5865
rect 14734 5856 14740 5868
rect 14792 5856 14798 5908
rect 15197 5899 15255 5905
rect 15197 5865 15209 5899
rect 15243 5896 15255 5899
rect 15286 5896 15292 5908
rect 15243 5868 15292 5896
rect 15243 5865 15255 5868
rect 15197 5859 15255 5865
rect 15286 5856 15292 5868
rect 15344 5856 15350 5908
rect 15654 5856 15660 5908
rect 15712 5896 15718 5908
rect 16117 5899 16175 5905
rect 16117 5896 16129 5899
rect 15712 5868 16129 5896
rect 15712 5856 15718 5868
rect 16117 5865 16129 5868
rect 16163 5865 16175 5899
rect 16117 5859 16175 5865
rect 16669 5899 16727 5905
rect 16669 5865 16681 5899
rect 16715 5896 16727 5899
rect 16850 5896 16856 5908
rect 16715 5868 16856 5896
rect 16715 5865 16727 5868
rect 16669 5859 16727 5865
rect 16850 5856 16856 5868
rect 16908 5856 16914 5908
rect 17402 5896 17408 5908
rect 16960 5868 17408 5896
rect 2682 5788 2688 5840
rect 2740 5828 2746 5840
rect 2740 5800 3004 5828
rect 2740 5788 2746 5800
rect 1854 5760 1860 5772
rect 1815 5732 1860 5760
rect 1854 5720 1860 5732
rect 1912 5720 1918 5772
rect 2590 5720 2596 5772
rect 2648 5760 2654 5772
rect 2976 5769 3004 5800
rect 3510 5788 3516 5840
rect 3568 5828 3574 5840
rect 4356 5828 4384 5856
rect 3568 5800 4384 5828
rect 3568 5788 3574 5800
rect 5902 5788 5908 5840
rect 5960 5828 5966 5840
rect 5960 5800 8064 5828
rect 5960 5788 5966 5800
rect 2777 5763 2835 5769
rect 2777 5760 2789 5763
rect 2648 5732 2789 5760
rect 2648 5720 2654 5732
rect 2777 5729 2789 5732
rect 2823 5729 2835 5763
rect 2777 5723 2835 5729
rect 2961 5763 3019 5769
rect 2961 5729 2973 5763
rect 3007 5729 3019 5763
rect 2961 5723 3019 5729
rect 3326 5720 3332 5772
rect 3384 5760 3390 5772
rect 4341 5763 4399 5769
rect 4341 5760 4353 5763
rect 3384 5732 4353 5760
rect 3384 5720 3390 5732
rect 4341 5729 4353 5732
rect 4387 5729 4399 5763
rect 7834 5760 7840 5772
rect 4341 5723 4399 5729
rect 4448 5732 7512 5760
rect 7795 5732 7840 5760
rect 2038 5692 2044 5704
rect 1999 5664 2044 5692
rect 2038 5652 2044 5664
rect 2096 5652 2102 5704
rect 3970 5692 3976 5704
rect 3344 5664 3976 5692
rect 1949 5627 2007 5633
rect 1949 5593 1961 5627
rect 1995 5624 2007 5627
rect 3344 5624 3372 5664
rect 3970 5652 3976 5664
rect 4028 5652 4034 5704
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4448 5692 4476 5732
rect 4798 5692 4804 5704
rect 4120 5664 4476 5692
rect 4759 5664 4804 5692
rect 4120 5652 4126 5664
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 7006 5692 7012 5704
rect 6967 5664 7012 5692
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 7484 5701 7512 5732
rect 7834 5720 7840 5732
rect 7892 5720 7898 5772
rect 8036 5769 8064 5800
rect 9950 5788 9956 5840
rect 10008 5828 10014 5840
rect 16960 5828 16988 5868
rect 17402 5856 17408 5868
rect 17460 5856 17466 5908
rect 17678 5856 17684 5908
rect 17736 5896 17742 5908
rect 17736 5868 19380 5896
rect 17736 5856 17742 5868
rect 10008 5800 16988 5828
rect 10008 5788 10014 5800
rect 18230 5788 18236 5840
rect 18288 5828 18294 5840
rect 19245 5831 19303 5837
rect 19245 5828 19257 5831
rect 18288 5800 19257 5828
rect 18288 5788 18294 5800
rect 19245 5797 19257 5800
rect 19291 5797 19303 5831
rect 19352 5828 19380 5868
rect 19886 5856 19892 5908
rect 19944 5896 19950 5908
rect 20165 5899 20223 5905
rect 20165 5896 20177 5899
rect 19944 5868 20177 5896
rect 19944 5856 19950 5868
rect 20165 5865 20177 5868
rect 20211 5865 20223 5899
rect 21082 5896 21088 5908
rect 21043 5868 21088 5896
rect 20165 5859 20223 5865
rect 21082 5856 21088 5868
rect 21140 5856 21146 5908
rect 19352 5800 20392 5828
rect 19245 5791 19303 5797
rect 8021 5763 8079 5769
rect 8021 5729 8033 5763
rect 8067 5729 8079 5763
rect 8021 5723 8079 5729
rect 8202 5720 8208 5772
rect 8260 5760 8266 5772
rect 9585 5763 9643 5769
rect 8260 5732 9076 5760
rect 8260 5720 8266 5732
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 8294 5652 8300 5704
rect 8352 5692 8358 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8352 5664 8953 5692
rect 8352 5652 8358 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 9048 5692 9076 5732
rect 9585 5729 9597 5763
rect 9631 5760 9643 5763
rect 9674 5760 9680 5772
rect 9631 5732 9680 5760
rect 9631 5729 9643 5732
rect 9585 5723 9643 5729
rect 9674 5720 9680 5732
rect 9732 5720 9738 5772
rect 16206 5760 16212 5772
rect 9876 5732 16212 5760
rect 9876 5692 9904 5732
rect 16206 5720 16212 5732
rect 16264 5720 16270 5772
rect 18046 5720 18052 5772
rect 18104 5760 18110 5772
rect 18104 5732 18149 5760
rect 18104 5720 18110 5732
rect 18690 5720 18696 5772
rect 18748 5760 18754 5772
rect 18748 5732 19748 5760
rect 18748 5720 18754 5732
rect 9048 5664 9904 5692
rect 8941 5655 8999 5661
rect 11882 5652 11888 5704
rect 11940 5692 11946 5704
rect 12437 5695 12495 5701
rect 12437 5692 12449 5695
rect 11940 5664 12449 5692
rect 11940 5652 11946 5664
rect 12437 5661 12449 5664
rect 12483 5661 12495 5695
rect 13538 5692 13544 5704
rect 13499 5664 13544 5692
rect 12437 5655 12495 5661
rect 13538 5652 13544 5664
rect 13596 5652 13602 5704
rect 13630 5652 13636 5704
rect 13688 5692 13694 5704
rect 14093 5695 14151 5701
rect 14093 5692 14105 5695
rect 13688 5664 14105 5692
rect 13688 5652 13694 5664
rect 14093 5661 14105 5664
rect 14139 5661 14151 5695
rect 15010 5692 15016 5704
rect 14971 5664 15016 5692
rect 14093 5655 14151 5661
rect 15010 5652 15016 5664
rect 15068 5652 15074 5704
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 18138 5692 18144 5704
rect 16172 5664 18144 5692
rect 16172 5652 16178 5664
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18509 5695 18567 5701
rect 18509 5661 18521 5695
rect 18555 5692 18567 5695
rect 18598 5692 18604 5704
rect 18555 5664 18604 5692
rect 18555 5661 18567 5664
rect 18509 5655 18567 5661
rect 18598 5652 18604 5664
rect 18656 5652 18662 5704
rect 18874 5652 18880 5704
rect 18932 5692 18938 5704
rect 19720 5701 19748 5732
rect 20364 5701 20392 5800
rect 21266 5788 21272 5840
rect 21324 5788 21330 5840
rect 21284 5760 21312 5788
rect 20824 5732 21312 5760
rect 20824 5701 20852 5732
rect 19429 5695 19487 5701
rect 19429 5692 19441 5695
rect 18932 5664 19441 5692
rect 18932 5652 18938 5664
rect 19429 5661 19441 5664
rect 19475 5661 19487 5695
rect 19429 5655 19487 5661
rect 19705 5695 19763 5701
rect 19705 5661 19717 5695
rect 19751 5661 19763 5695
rect 19705 5655 19763 5661
rect 20349 5695 20407 5701
rect 20349 5661 20361 5695
rect 20395 5661 20407 5695
rect 20349 5655 20407 5661
rect 20809 5695 20867 5701
rect 20809 5661 20821 5695
rect 20855 5661 20867 5695
rect 20809 5655 20867 5661
rect 20990 5652 20996 5704
rect 21048 5692 21054 5704
rect 21269 5695 21327 5701
rect 21269 5692 21281 5695
rect 21048 5664 21281 5692
rect 21048 5652 21054 5664
rect 21269 5661 21281 5664
rect 21315 5692 21327 5695
rect 21818 5692 21824 5704
rect 21315 5664 21824 5692
rect 21315 5661 21327 5664
rect 21269 5655 21327 5661
rect 21818 5652 21824 5664
rect 21876 5652 21882 5704
rect 4249 5627 4307 5633
rect 4249 5624 4261 5627
rect 1995 5596 3372 5624
rect 3436 5596 4261 5624
rect 1995 5593 2007 5596
rect 1949 5587 2007 5593
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 3436 5565 3464 5596
rect 4249 5593 4261 5596
rect 4295 5593 4307 5627
rect 7024 5624 7052 5652
rect 10413 5627 10471 5633
rect 10413 5624 10425 5627
rect 7024 5596 10425 5624
rect 4249 5587 4307 5593
rect 10413 5593 10425 5596
rect 10459 5624 10471 5627
rect 11698 5624 11704 5636
rect 10459 5596 11704 5624
rect 10459 5593 10471 5596
rect 10413 5587 10471 5593
rect 11698 5584 11704 5596
rect 11756 5584 11762 5636
rect 12161 5627 12219 5633
rect 12161 5593 12173 5627
rect 12207 5624 12219 5627
rect 12710 5624 12716 5636
rect 12207 5596 12716 5624
rect 12207 5593 12219 5596
rect 12161 5587 12219 5593
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 17804 5627 17862 5633
rect 17804 5593 17816 5627
rect 17850 5624 17862 5627
rect 18690 5624 18696 5636
rect 17850 5596 18696 5624
rect 17850 5593 17862 5596
rect 17804 5587 17862 5593
rect 18690 5584 18696 5596
rect 18748 5584 18754 5636
rect 3421 5559 3479 5565
rect 3108 5528 3153 5556
rect 3108 5516 3114 5528
rect 3421 5525 3433 5559
rect 3467 5525 3479 5559
rect 4154 5556 4160 5568
rect 4115 5528 4160 5556
rect 3421 5519 3479 5525
rect 4154 5516 4160 5528
rect 4212 5516 4218 5568
rect 4985 5559 5043 5565
rect 4985 5525 4997 5559
rect 5031 5556 5043 5559
rect 6822 5556 6828 5568
rect 5031 5528 6828 5556
rect 5031 5525 5043 5528
rect 4985 5519 5043 5525
rect 6822 5516 6828 5528
rect 6880 5516 6886 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7285 5559 7343 5565
rect 7285 5556 7297 5559
rect 6972 5528 7297 5556
rect 6972 5516 6978 5528
rect 7285 5525 7297 5528
rect 7331 5525 7343 5559
rect 7285 5519 7343 5525
rect 7374 5516 7380 5568
rect 7432 5556 7438 5568
rect 8113 5559 8171 5565
rect 8113 5556 8125 5559
rect 7432 5528 8125 5556
rect 7432 5516 7438 5528
rect 8113 5525 8125 5528
rect 8159 5525 8171 5559
rect 8113 5519 8171 5525
rect 8481 5559 8539 5565
rect 8481 5525 8493 5559
rect 8527 5556 8539 5559
rect 8662 5556 8668 5568
rect 8527 5528 8668 5556
rect 8527 5525 8539 5528
rect 8481 5519 8539 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 9674 5556 9680 5568
rect 9635 5528 9680 5556
rect 9674 5516 9680 5528
rect 9732 5516 9738 5568
rect 9769 5559 9827 5565
rect 9769 5525 9781 5559
rect 9815 5556 9827 5559
rect 9950 5556 9956 5568
rect 9815 5528 9956 5556
rect 9815 5525 9827 5528
rect 9769 5519 9827 5525
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10137 5559 10195 5565
rect 10137 5525 10149 5559
rect 10183 5556 10195 5559
rect 12250 5556 12256 5568
rect 10183 5528 12256 5556
rect 10183 5525 10195 5528
rect 10137 5519 10195 5525
rect 12250 5516 12256 5528
rect 12308 5516 12314 5568
rect 13078 5556 13084 5568
rect 13039 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 17494 5516 17500 5568
rect 17552 5556 17558 5568
rect 18325 5559 18383 5565
rect 18325 5556 18337 5559
rect 17552 5528 18337 5556
rect 17552 5516 17558 5528
rect 18325 5525 18337 5528
rect 18371 5525 18383 5559
rect 18325 5519 18383 5525
rect 18506 5516 18512 5568
rect 18564 5556 18570 5568
rect 18785 5559 18843 5565
rect 18785 5556 18797 5559
rect 18564 5528 18797 5556
rect 18564 5516 18570 5528
rect 18785 5525 18797 5528
rect 18831 5525 18843 5559
rect 19886 5556 19892 5568
rect 19847 5528 19892 5556
rect 18785 5519 18843 5525
rect 19886 5516 19892 5528
rect 19944 5516 19950 5568
rect 20622 5556 20628 5568
rect 20583 5528 20628 5556
rect 20622 5516 20628 5528
rect 20680 5516 20686 5568
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 2866 5352 2872 5364
rect 2827 5324 2872 5352
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3881 5355 3939 5361
rect 3881 5352 3893 5355
rect 3108 5324 3893 5352
rect 3108 5312 3114 5324
rect 3881 5321 3893 5324
rect 3927 5321 3939 5355
rect 3881 5315 3939 5321
rect 4249 5355 4307 5361
rect 4249 5321 4261 5355
rect 4295 5352 4307 5355
rect 4706 5352 4712 5364
rect 4295 5324 4712 5352
rect 4295 5321 4307 5324
rect 4249 5315 4307 5321
rect 4706 5312 4712 5324
rect 4764 5312 4770 5364
rect 5353 5355 5411 5361
rect 5353 5321 5365 5355
rect 5399 5352 5411 5355
rect 8021 5355 8079 5361
rect 8021 5352 8033 5355
rect 5399 5324 8033 5352
rect 5399 5321 5411 5324
rect 5353 5315 5411 5321
rect 8021 5321 8033 5324
rect 8067 5321 8079 5355
rect 8021 5315 8079 5321
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8168 5324 8401 5352
rect 8168 5312 8174 5324
rect 8389 5321 8401 5324
rect 8435 5352 8447 5355
rect 9217 5355 9275 5361
rect 8435 5324 8708 5352
rect 8435 5321 8447 5324
rect 8389 5315 8447 5321
rect 1670 5244 1676 5296
rect 1728 5284 1734 5296
rect 3237 5287 3295 5293
rect 3237 5284 3249 5287
rect 1728 5256 3249 5284
rect 1728 5244 1734 5256
rect 3237 5253 3249 5256
rect 3283 5284 3295 5287
rect 3510 5284 3516 5296
rect 3283 5256 3516 5284
rect 3283 5253 3295 5256
rect 3237 5247 3295 5253
rect 3510 5244 3516 5256
rect 3568 5244 3574 5296
rect 7500 5287 7558 5293
rect 4172 5256 7420 5284
rect 1949 5219 2007 5225
rect 1949 5185 1961 5219
rect 1995 5216 2007 5219
rect 2498 5216 2504 5228
rect 1995 5188 2504 5216
rect 1995 5185 2007 5188
rect 1949 5179 2007 5185
rect 2498 5176 2504 5188
rect 2556 5176 2562 5228
rect 4172 5216 4200 5256
rect 3344 5188 4200 5216
rect 4341 5219 4399 5225
rect 3344 5160 3372 5188
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4522 5216 4528 5228
rect 4387 5188 4528 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4522 5176 4528 5188
rect 4580 5216 4586 5228
rect 4982 5216 4988 5228
rect 4580 5188 4988 5216
rect 4580 5176 4586 5188
rect 4982 5176 4988 5188
rect 5040 5176 5046 5228
rect 5442 5216 5448 5228
rect 5403 5188 5448 5216
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 7392 5216 7420 5256
rect 7500 5253 7512 5287
rect 7546 5284 7558 5287
rect 8680 5284 8708 5324
rect 9217 5321 9229 5355
rect 9263 5352 9275 5355
rect 9398 5352 9404 5364
rect 9263 5324 9404 5352
rect 9263 5321 9275 5324
rect 9217 5315 9275 5321
rect 9398 5312 9404 5324
rect 9456 5312 9462 5364
rect 9490 5312 9496 5364
rect 9548 5352 9554 5364
rect 16669 5355 16727 5361
rect 9548 5324 9593 5352
rect 9692 5324 16436 5352
rect 9548 5312 9554 5324
rect 9692 5284 9720 5324
rect 7546 5256 8616 5284
rect 8680 5256 9720 5284
rect 10628 5287 10686 5293
rect 7546 5253 7558 5256
rect 7500 5247 7558 5253
rect 7745 5219 7803 5225
rect 7392 5188 7696 5216
rect 2130 5108 2136 5160
rect 2188 5148 2194 5160
rect 2225 5151 2283 5157
rect 2225 5148 2237 5151
rect 2188 5120 2237 5148
rect 2188 5108 2194 5120
rect 2225 5117 2237 5120
rect 2271 5117 2283 5151
rect 3326 5148 3332 5160
rect 3287 5120 3332 5148
rect 2225 5111 2283 5117
rect 3326 5108 3332 5120
rect 3384 5108 3390 5160
rect 3418 5108 3424 5160
rect 3476 5148 3482 5160
rect 4433 5151 4491 5157
rect 3476 5120 3521 5148
rect 3476 5108 3482 5120
rect 4433 5117 4445 5151
rect 4479 5117 4491 5151
rect 4433 5111 4491 5117
rect 5261 5151 5319 5157
rect 5261 5117 5273 5151
rect 5307 5148 5319 5151
rect 7668 5148 7696 5188
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 8018 5216 8024 5228
rect 7791 5188 8024 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 8018 5176 8024 5188
rect 8076 5176 8082 5228
rect 8478 5216 8484 5228
rect 8439 5188 8484 5216
rect 8478 5176 8484 5188
rect 8536 5176 8542 5228
rect 8588 5160 8616 5256
rect 10628 5253 10640 5287
rect 10674 5284 10686 5287
rect 10962 5284 10968 5296
rect 10674 5256 10968 5284
rect 10674 5253 10686 5256
rect 10628 5247 10686 5253
rect 10962 5244 10968 5256
rect 11020 5244 11026 5296
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 12158 5284 12164 5296
rect 11756 5256 12164 5284
rect 11756 5244 11762 5256
rect 12158 5244 12164 5256
rect 12216 5284 12222 5296
rect 12989 5287 13047 5293
rect 12989 5284 13001 5287
rect 12216 5256 13001 5284
rect 12216 5244 12222 5256
rect 12989 5253 13001 5256
rect 13035 5253 13047 5287
rect 12989 5247 13047 5253
rect 14366 5244 14372 5296
rect 14424 5284 14430 5296
rect 14737 5287 14795 5293
rect 14737 5284 14749 5287
rect 14424 5256 14749 5284
rect 14424 5244 14430 5256
rect 14737 5253 14749 5256
rect 14783 5284 14795 5287
rect 16298 5284 16304 5296
rect 14783 5256 16304 5284
rect 14783 5253 14795 5256
rect 14737 5247 14795 5253
rect 16298 5244 16304 5256
rect 16356 5244 16362 5296
rect 16408 5284 16436 5324
rect 16669 5321 16681 5355
rect 16715 5352 16727 5355
rect 16942 5352 16948 5364
rect 16715 5324 16948 5352
rect 16715 5321 16727 5324
rect 16669 5315 16727 5321
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17681 5355 17739 5361
rect 17681 5321 17693 5355
rect 17727 5321 17739 5355
rect 17681 5315 17739 5321
rect 17696 5284 17724 5315
rect 17770 5312 17776 5364
rect 17828 5352 17834 5364
rect 18601 5355 18659 5361
rect 17828 5324 18184 5352
rect 17828 5312 17834 5324
rect 16408 5256 17724 5284
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 10873 5219 10931 5225
rect 10100 5188 10824 5216
rect 10100 5176 10106 5188
rect 8386 5148 8392 5160
rect 5307 5120 6408 5148
rect 7668 5120 8392 5148
rect 5307 5117 5319 5120
rect 5261 5111 5319 5117
rect 3436 5080 3464 5108
rect 4448 5080 4476 5111
rect 2746 5052 3004 5080
rect 3436 5052 4476 5080
rect 5813 5083 5871 5089
rect 2314 4972 2320 5024
rect 2372 5012 2378 5024
rect 2501 5015 2559 5021
rect 2501 5012 2513 5015
rect 2372 4984 2513 5012
rect 2372 4972 2378 4984
rect 2501 4981 2513 4984
rect 2547 5012 2559 5015
rect 2746 5012 2774 5052
rect 2547 4984 2774 5012
rect 2976 5012 3004 5052
rect 5813 5049 5825 5083
rect 5859 5080 5871 5083
rect 5902 5080 5908 5092
rect 5859 5052 5908 5080
rect 5859 5049 5871 5052
rect 5813 5043 5871 5049
rect 5902 5040 5908 5052
rect 5960 5040 5966 5092
rect 6380 5089 6408 5120
rect 8386 5108 8392 5120
rect 8444 5108 8450 5160
rect 8570 5108 8576 5160
rect 8628 5148 8634 5160
rect 10796 5148 10824 5188
rect 10873 5185 10885 5219
rect 10919 5216 10931 5219
rect 11146 5216 11152 5228
rect 10919 5188 11152 5216
rect 10919 5185 10931 5188
rect 10873 5179 10931 5185
rect 11146 5176 11152 5188
rect 11204 5176 11210 5228
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 12342 5216 12348 5228
rect 12303 5188 12348 5216
rect 11517 5179 11575 5185
rect 11532 5148 11560 5179
rect 12342 5176 12348 5188
rect 12400 5176 12406 5228
rect 15013 5219 15071 5225
rect 15013 5216 15025 5219
rect 12728 5188 15025 5216
rect 8628 5120 8673 5148
rect 10796 5120 11560 5148
rect 12161 5151 12219 5157
rect 8628 5108 8634 5120
rect 12161 5117 12173 5151
rect 12207 5117 12219 5151
rect 12161 5111 12219 5117
rect 6365 5083 6423 5089
rect 6365 5049 6377 5083
rect 6411 5080 6423 5083
rect 6546 5080 6552 5092
rect 6411 5052 6552 5080
rect 6411 5049 6423 5052
rect 6365 5043 6423 5049
rect 6546 5040 6552 5052
rect 6604 5040 6610 5092
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 12176 5080 12204 5111
rect 12250 5108 12256 5160
rect 12308 5148 12314 5160
rect 12308 5120 12353 5148
rect 12308 5108 12314 5120
rect 12728 5089 12756 5188
rect 15013 5185 15025 5188
rect 15059 5185 15071 5219
rect 15838 5216 15844 5228
rect 15799 5188 15844 5216
rect 15013 5179 15071 5185
rect 15838 5176 15844 5188
rect 15896 5176 15902 5228
rect 15930 5176 15936 5228
rect 15988 5216 15994 5228
rect 17037 5219 17095 5225
rect 17037 5216 17049 5219
rect 15988 5188 17049 5216
rect 15988 5176 15994 5188
rect 17037 5185 17049 5188
rect 17083 5185 17095 5219
rect 17037 5179 17095 5185
rect 17402 5176 17408 5228
rect 17460 5216 17466 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17460 5188 17877 5216
rect 17460 5176 17466 5188
rect 17865 5185 17877 5188
rect 17911 5216 17923 5219
rect 17954 5216 17960 5228
rect 17911 5188 17960 5216
rect 17911 5185 17923 5188
rect 17865 5179 17923 5185
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 18156 5225 18184 5324
rect 18601 5321 18613 5355
rect 18647 5352 18659 5355
rect 19058 5352 19064 5364
rect 18647 5324 19064 5352
rect 18647 5321 18659 5324
rect 18601 5315 18659 5321
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 20346 5312 20352 5364
rect 20404 5352 20410 5364
rect 20441 5355 20499 5361
rect 20441 5352 20453 5355
rect 20404 5324 20453 5352
rect 20404 5312 20410 5324
rect 20441 5321 20453 5324
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 18966 5244 18972 5296
rect 19024 5284 19030 5296
rect 19024 5256 21128 5284
rect 19024 5244 19030 5256
rect 18141 5219 18199 5225
rect 18141 5185 18153 5219
rect 18187 5185 18199 5219
rect 18141 5179 18199 5185
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 18785 5219 18843 5225
rect 18785 5216 18797 5219
rect 18656 5188 18797 5216
rect 18656 5176 18662 5188
rect 18785 5185 18797 5188
rect 18831 5216 18843 5219
rect 19150 5216 19156 5228
rect 18831 5188 19156 5216
rect 18831 5185 18843 5188
rect 18785 5179 18843 5185
rect 19150 5176 19156 5188
rect 19208 5176 19214 5228
rect 19245 5219 19303 5225
rect 19245 5185 19257 5219
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 15562 5148 15568 5160
rect 15523 5120 15568 5148
rect 15562 5108 15568 5120
rect 15620 5108 15626 5160
rect 15746 5148 15752 5160
rect 15707 5120 15752 5148
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 17126 5148 17132 5160
rect 17087 5120 17132 5148
rect 17126 5108 17132 5120
rect 17184 5108 17190 5160
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 19260 5148 19288 5179
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20165 5219 20223 5225
rect 20165 5216 20177 5219
rect 19944 5188 20177 5216
rect 19944 5176 19950 5188
rect 20165 5185 20177 5188
rect 20211 5185 20223 5219
rect 20165 5179 20223 5185
rect 20438 5176 20444 5228
rect 20496 5216 20502 5228
rect 21100 5225 21128 5256
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20496 5188 20637 5216
rect 20496 5176 20502 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 21085 5219 21143 5225
rect 21085 5185 21097 5219
rect 21131 5185 21143 5219
rect 21085 5179 21143 5185
rect 19518 5148 19524 5160
rect 17276 5120 17321 5148
rect 18340 5120 19288 5148
rect 19479 5120 19524 5148
rect 17276 5108 17282 5120
rect 12713 5083 12771 5089
rect 8260 5052 8432 5080
rect 12176 5052 12434 5080
rect 8260 5040 8266 5052
rect 8294 5012 8300 5024
rect 2976 4984 8300 5012
rect 2547 4981 2559 4984
rect 2501 4975 2559 4981
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 8404 5012 8432 5052
rect 11698 5012 11704 5024
rect 8404 4984 11704 5012
rect 11698 4972 11704 4984
rect 11756 4972 11762 5024
rect 12406 5012 12434 5052
rect 12713 5049 12725 5083
rect 12759 5049 12771 5083
rect 12713 5043 12771 5049
rect 16209 5083 16267 5089
rect 16209 5049 16221 5083
rect 16255 5080 16267 5083
rect 17034 5080 17040 5092
rect 16255 5052 17040 5080
rect 16255 5049 16267 5052
rect 16209 5043 16267 5049
rect 17034 5040 17040 5052
rect 17092 5040 17098 5092
rect 18340 5089 18368 5120
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 18325 5083 18383 5089
rect 18325 5049 18337 5083
rect 18371 5049 18383 5083
rect 18325 5043 18383 5049
rect 18874 5040 18880 5092
rect 18932 5080 18938 5092
rect 19981 5083 20039 5089
rect 19981 5080 19993 5083
rect 18932 5052 19993 5080
rect 18932 5040 18938 5052
rect 19981 5049 19993 5052
rect 20027 5049 20039 5083
rect 19981 5043 20039 5049
rect 13630 5012 13636 5024
rect 12406 4984 13636 5012
rect 13630 4972 13636 4984
rect 13688 4972 13694 5024
rect 15197 5015 15255 5021
rect 15197 4981 15209 5015
rect 15243 5012 15255 5015
rect 17954 5012 17960 5024
rect 15243 4984 17960 5012
rect 15243 4981 15255 4984
rect 15197 4975 15255 4981
rect 17954 4972 17960 4984
rect 18012 4972 18018 5024
rect 18138 4972 18144 5024
rect 18196 5012 18202 5024
rect 19061 5015 19119 5021
rect 19061 5012 19073 5015
rect 18196 4984 19073 5012
rect 18196 4972 18202 4984
rect 19061 4981 19073 4984
rect 19107 4981 19119 5015
rect 20898 5012 20904 5024
rect 20859 4984 20904 5012
rect 19061 4975 19119 4981
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 3970 4808 3976 4820
rect 3375 4780 3976 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 5442 4768 5448 4820
rect 5500 4808 5506 4820
rect 7745 4811 7803 4817
rect 7745 4808 7757 4811
rect 5500 4780 7757 4808
rect 5500 4768 5506 4780
rect 7745 4777 7757 4780
rect 7791 4777 7803 4811
rect 10134 4808 10140 4820
rect 10095 4780 10140 4808
rect 7745 4771 7803 4777
rect 10134 4768 10140 4780
rect 10192 4768 10198 4820
rect 11882 4808 11888 4820
rect 10520 4780 11744 4808
rect 11843 4780 11888 4808
rect 1670 4740 1676 4752
rect 1631 4712 1676 4740
rect 1670 4700 1676 4712
rect 1728 4700 1734 4752
rect 7469 4743 7527 4749
rect 7469 4709 7481 4743
rect 7515 4709 7527 4743
rect 10520 4740 10548 4780
rect 7469 4703 7527 4709
rect 9508 4712 10548 4740
rect 11716 4740 11744 4780
rect 11882 4768 11888 4780
rect 11940 4768 11946 4820
rect 15746 4808 15752 4820
rect 11992 4780 15752 4808
rect 11992 4740 12020 4780
rect 15746 4768 15752 4780
rect 15804 4768 15810 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16080 4780 19288 4808
rect 16080 4768 16086 4780
rect 13630 4740 13636 4752
rect 11716 4712 12020 4740
rect 13591 4712 13636 4740
rect 1762 4632 1768 4684
rect 1820 4672 1826 4684
rect 1949 4675 2007 4681
rect 1949 4672 1961 4675
rect 1820 4644 1961 4672
rect 1820 4632 1826 4644
rect 1949 4641 1961 4644
rect 1995 4641 2007 4675
rect 5166 4672 5172 4684
rect 5127 4644 5172 4672
rect 1949 4635 2007 4641
rect 1964 4604 1992 4635
rect 5166 4632 5172 4644
rect 5224 4672 5230 4684
rect 6089 4675 6147 4681
rect 6089 4672 6101 4675
rect 5224 4644 6101 4672
rect 5224 4632 5230 4644
rect 6089 4641 6101 4644
rect 6135 4641 6147 4675
rect 7484 4672 7512 4703
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 7484 4644 8401 4672
rect 6089 4635 6147 4641
rect 8389 4641 8401 4644
rect 8435 4672 8447 4675
rect 8570 4672 8576 4684
rect 8435 4644 8576 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 8570 4632 8576 4644
rect 8628 4632 8634 4684
rect 9122 4672 9128 4684
rect 9083 4644 9128 4672
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 2682 4604 2688 4616
rect 1964 4576 2688 4604
rect 2682 4564 2688 4576
rect 2740 4604 2746 4616
rect 5184 4604 5212 4632
rect 2740 4576 5212 4604
rect 2740 4564 2746 4576
rect 7926 4564 7932 4616
rect 7984 4604 7990 4616
rect 8113 4607 8171 4613
rect 8113 4604 8125 4607
rect 7984 4576 8125 4604
rect 7984 4564 7990 4576
rect 8113 4573 8125 4576
rect 8159 4604 8171 4607
rect 9508 4604 9536 4712
rect 13630 4700 13636 4712
rect 13688 4700 13694 4752
rect 9585 4675 9643 4681
rect 9585 4641 9597 4675
rect 9631 4672 9643 4675
rect 10318 4672 10324 4684
rect 9631 4644 10324 4672
rect 9631 4641 9643 4644
rect 9585 4635 9643 4641
rect 10318 4632 10324 4644
rect 10376 4632 10382 4684
rect 18046 4632 18052 4684
rect 18104 4672 18110 4684
rect 19260 4681 19288 4780
rect 19245 4675 19303 4681
rect 18104 4644 18644 4672
rect 18104 4632 18110 4644
rect 8159 4576 9536 4604
rect 9769 4607 9827 4613
rect 8159 4573 8171 4576
rect 8113 4567 8171 4573
rect 9769 4573 9781 4607
rect 9815 4604 9827 4607
rect 9858 4604 9864 4616
rect 9815 4576 9864 4604
rect 9815 4573 9827 4576
rect 9769 4567 9827 4573
rect 9858 4564 9864 4576
rect 9916 4564 9922 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 11146 4604 11152 4616
rect 10551 4576 11152 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 11146 4564 11152 4576
rect 11204 4604 11210 4616
rect 12526 4613 12532 4616
rect 12253 4607 12311 4613
rect 12253 4604 12265 4607
rect 11204 4576 12265 4604
rect 11204 4564 11210 4576
rect 12253 4573 12265 4576
rect 12299 4573 12311 4607
rect 12253 4567 12311 4573
rect 12520 4567 12532 4613
rect 12584 4604 12590 4616
rect 14090 4604 14096 4616
rect 12584 4576 12620 4604
rect 14051 4576 14096 4604
rect 12526 4564 12532 4567
rect 12584 4564 12590 4576
rect 14090 4564 14096 4576
rect 14148 4564 14154 4616
rect 16298 4564 16304 4616
rect 16356 4604 16362 4616
rect 16393 4607 16451 4613
rect 16393 4604 16405 4607
rect 16356 4576 16405 4604
rect 16356 4564 16362 4576
rect 16393 4573 16405 4576
rect 16439 4604 16451 4607
rect 18064 4604 18092 4632
rect 18506 4604 18512 4616
rect 16439 4576 18092 4604
rect 18467 4576 18512 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 18506 4564 18512 4576
rect 18564 4564 18570 4616
rect 18616 4604 18644 4644
rect 19245 4641 19257 4675
rect 19291 4641 19303 4675
rect 19245 4635 19303 4641
rect 21094 4607 21152 4613
rect 18616 4576 20116 4604
rect 1489 4539 1547 4545
rect 1489 4505 1501 4539
rect 1535 4505 1547 4539
rect 1489 4499 1547 4505
rect 1504 4468 1532 4499
rect 1578 4496 1584 4548
rect 1636 4536 1642 4548
rect 2194 4539 2252 4545
rect 2194 4536 2206 4539
rect 1636 4508 2206 4536
rect 1636 4496 1642 4508
rect 2194 4505 2206 4508
rect 2240 4505 2252 4539
rect 2194 4499 2252 4505
rect 4924 4539 4982 4545
rect 4924 4505 4936 4539
rect 4970 4536 4982 4539
rect 5442 4536 5448 4548
rect 4970 4508 5448 4536
rect 4970 4505 4982 4508
rect 4924 4499 4982 4505
rect 5442 4496 5448 4508
rect 5500 4496 5506 4548
rect 6356 4539 6414 4545
rect 6356 4505 6368 4539
rect 6402 4536 6414 4539
rect 6638 4536 6644 4548
rect 6402 4508 6644 4536
rect 6402 4505 6414 4508
rect 6356 4499 6414 4505
rect 6638 4496 6644 4508
rect 6696 4496 6702 4548
rect 9677 4539 9735 4545
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 9950 4536 9956 4548
rect 9723 4508 9956 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 10318 4496 10324 4548
rect 10376 4536 10382 4548
rect 10772 4539 10830 4545
rect 10376 4508 10548 4536
rect 10376 4496 10382 4508
rect 3050 4468 3056 4480
rect 1504 4440 3056 4468
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3789 4471 3847 4477
rect 3789 4437 3801 4471
rect 3835 4468 3847 4471
rect 4798 4468 4804 4480
rect 3835 4440 4804 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4798 4428 4804 4440
rect 4856 4428 4862 4480
rect 5813 4471 5871 4477
rect 5813 4437 5825 4471
rect 5859 4468 5871 4471
rect 7926 4468 7932 4480
rect 5859 4440 7932 4468
rect 5859 4437 5871 4440
rect 5813 4431 5871 4437
rect 7926 4428 7932 4440
rect 7984 4428 7990 4480
rect 8202 4468 8208 4480
rect 8163 4440 8208 4468
rect 8202 4428 8208 4440
rect 8260 4428 8266 4480
rect 9490 4428 9496 4480
rect 9548 4468 9554 4480
rect 10410 4468 10416 4480
rect 9548 4440 10416 4468
rect 9548 4428 9554 4440
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10520 4468 10548 4508
rect 10772 4505 10784 4539
rect 10818 4536 10830 4539
rect 11054 4536 11060 4548
rect 10818 4508 11060 4536
rect 10818 4505 10830 4508
rect 10772 4499 10830 4505
rect 11054 4496 11060 4508
rect 11112 4496 11118 4548
rect 15930 4536 15936 4548
rect 11164 4508 15936 4536
rect 11164 4468 11192 4508
rect 15930 4496 15936 4508
rect 15988 4496 15994 4548
rect 16148 4539 16206 4545
rect 16148 4505 16160 4539
rect 16194 4536 16206 4539
rect 17034 4536 17040 4548
rect 16194 4508 17040 4536
rect 16194 4505 16206 4508
rect 16148 4499 16206 4505
rect 17034 4496 17040 4508
rect 17092 4496 17098 4548
rect 17678 4496 17684 4548
rect 17736 4536 17742 4548
rect 17782 4539 17840 4545
rect 17782 4536 17794 4539
rect 17736 4508 17794 4536
rect 17736 4496 17742 4508
rect 17782 4505 17794 4508
rect 17828 4505 17840 4539
rect 18785 4539 18843 4545
rect 18785 4536 18797 4539
rect 17782 4499 17840 4505
rect 17880 4508 18797 4536
rect 17880 4480 17908 4508
rect 18785 4505 18797 4508
rect 18831 4505 18843 4539
rect 18785 4499 18843 4505
rect 14734 4468 14740 4480
rect 10520 4440 11192 4468
rect 14695 4440 14740 4468
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15013 4471 15071 4477
rect 15013 4437 15025 4471
rect 15059 4468 15071 4471
rect 15562 4468 15568 4480
rect 15059 4440 15568 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 15562 4428 15568 4440
rect 15620 4468 15626 4480
rect 16390 4468 16396 4480
rect 15620 4440 16396 4468
rect 15620 4428 15626 4440
rect 16390 4428 16396 4440
rect 16448 4428 16454 4480
rect 16669 4471 16727 4477
rect 16669 4437 16681 4471
rect 16715 4468 16727 4471
rect 16942 4468 16948 4480
rect 16715 4440 16948 4468
rect 16715 4437 16727 4440
rect 16669 4431 16727 4437
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17862 4428 17868 4480
rect 17920 4428 17926 4480
rect 18046 4428 18052 4480
rect 18104 4468 18110 4480
rect 18325 4471 18383 4477
rect 18325 4468 18337 4471
rect 18104 4440 18337 4468
rect 18104 4428 18110 4440
rect 18325 4437 18337 4440
rect 18371 4437 18383 4471
rect 18325 4431 18383 4437
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 19981 4471 20039 4477
rect 19981 4468 19993 4471
rect 19024 4440 19993 4468
rect 19024 4428 19030 4440
rect 19981 4437 19993 4440
rect 20027 4437 20039 4471
rect 20088 4468 20116 4576
rect 21094 4573 21106 4607
rect 21140 4573 21152 4607
rect 21094 4567 21152 4573
rect 21361 4607 21419 4613
rect 21361 4573 21373 4607
rect 21407 4573 21419 4607
rect 21361 4567 21419 4573
rect 21100 4536 21128 4567
rect 21174 4536 21180 4548
rect 21100 4508 21180 4536
rect 21174 4496 21180 4508
rect 21232 4496 21238 4548
rect 21376 4468 21404 4567
rect 20088 4440 21404 4468
rect 19981 4431 20039 4437
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 4617 4267 4675 4273
rect 4617 4264 4629 4267
rect 3292 4236 4629 4264
rect 3292 4224 3298 4236
rect 4617 4233 4629 4236
rect 4663 4233 4675 4267
rect 4617 4227 4675 4233
rect 5350 4224 5356 4276
rect 5408 4264 5414 4276
rect 5629 4267 5687 4273
rect 5629 4264 5641 4267
rect 5408 4236 5641 4264
rect 5408 4224 5414 4236
rect 5629 4233 5641 4236
rect 5675 4233 5687 4267
rect 5994 4264 6000 4276
rect 5955 4236 6000 4264
rect 5629 4227 5687 4233
rect 5994 4224 6000 4236
rect 6052 4224 6058 4276
rect 7009 4267 7067 4273
rect 7009 4233 7021 4267
rect 7055 4264 7067 4267
rect 7098 4264 7104 4276
rect 7055 4236 7104 4264
rect 7055 4233 7067 4236
rect 7009 4227 7067 4233
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 7929 4267 7987 4273
rect 7929 4233 7941 4267
rect 7975 4264 7987 4267
rect 8202 4264 8208 4276
rect 7975 4236 8208 4264
rect 7975 4233 7987 4236
rect 7929 4227 7987 4233
rect 8202 4224 8208 4236
rect 8260 4224 8266 4276
rect 9125 4267 9183 4273
rect 9125 4233 9137 4267
rect 9171 4264 9183 4267
rect 9214 4264 9220 4276
rect 9171 4236 9220 4264
rect 9171 4233 9183 4236
rect 9125 4227 9183 4233
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 10318 4264 10324 4276
rect 9968 4236 10324 4264
rect 3712 4168 4016 4196
rect 2866 4088 2872 4140
rect 2924 4128 2930 4140
rect 3329 4131 3387 4137
rect 3329 4128 3341 4131
rect 2924 4100 3341 4128
rect 2924 4088 2930 4100
rect 3329 4097 3341 4100
rect 3375 4097 3387 4131
rect 3712 4128 3740 4168
rect 3329 4091 3387 4097
rect 3620 4100 3740 4128
rect 3789 4131 3847 4137
rect 1949 4063 2007 4069
rect 1949 4029 1961 4063
rect 1995 4029 2007 4063
rect 2222 4060 2228 4072
rect 2135 4032 2228 4060
rect 1949 4023 2007 4029
rect 1964 3924 1992 4023
rect 2222 4020 2228 4032
rect 2280 4060 2286 4072
rect 2958 4060 2964 4072
rect 2280 4032 2964 4060
rect 2280 4020 2286 4032
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3053 4063 3111 4069
rect 3053 4029 3065 4063
rect 3099 4060 3111 4063
rect 3142 4060 3148 4072
rect 3099 4032 3148 4060
rect 3099 4029 3111 4032
rect 3053 4023 3111 4029
rect 3142 4020 3148 4032
rect 3200 4020 3206 4072
rect 3620 3992 3648 4100
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 3988 4128 4016 4168
rect 6472 4168 7052 4196
rect 4430 4128 4436 4140
rect 3988 4100 4436 4128
rect 3789 4091 3847 4097
rect 2746 3964 3648 3992
rect 2746 3924 2774 3964
rect 1964 3896 2774 3924
rect 3804 3924 3832 4091
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4709 4131 4767 4137
rect 4709 4097 4721 4131
rect 4755 4128 4767 4131
rect 4890 4128 4896 4140
rect 4755 4100 4896 4128
rect 4755 4097 4767 4100
rect 4709 4091 4767 4097
rect 4890 4088 4896 4100
rect 4948 4128 4954 4140
rect 6472 4128 6500 4168
rect 4948 4100 6500 4128
rect 4948 4088 4954 4100
rect 6546 4088 6552 4140
rect 6604 4088 6610 4140
rect 6914 4128 6920 4140
rect 6875 4100 6920 4128
rect 6914 4088 6920 4100
rect 6972 4088 6978 4140
rect 7024 4128 7052 4168
rect 7466 4156 7472 4208
rect 7524 4196 7530 4208
rect 9858 4196 9864 4208
rect 7524 4168 9864 4196
rect 7524 4156 7530 4168
rect 9858 4156 9864 4168
rect 9916 4156 9922 4208
rect 8018 4128 8024 4140
rect 7024 4100 7880 4128
rect 7979 4100 8024 4128
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5258 4060 5264 4072
rect 4856 4032 5264 4060
rect 4856 4020 4862 4032
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5353 4063 5411 4069
rect 5353 4029 5365 4063
rect 5399 4029 5411 4063
rect 5534 4060 5540 4072
rect 5495 4032 5540 4060
rect 5353 4023 5411 4029
rect 3970 3992 3976 4004
rect 3931 3964 3976 3992
rect 3970 3952 3976 3964
rect 4028 3952 4034 4004
rect 4062 3952 4068 4004
rect 4120 3992 4126 4004
rect 4249 3995 4307 4001
rect 4249 3992 4261 3995
rect 4120 3964 4261 3992
rect 4120 3952 4126 3964
rect 4249 3961 4261 3964
rect 4295 3961 4307 3995
rect 5368 3992 5396 4023
rect 5534 4020 5540 4032
rect 5592 4020 5598 4072
rect 5902 4020 5908 4072
rect 5960 4060 5966 4072
rect 6454 4060 6460 4072
rect 5960 4032 6460 4060
rect 5960 4020 5966 4032
rect 6454 4020 6460 4032
rect 6512 4020 6518 4072
rect 6564 4060 6592 4088
rect 6733 4063 6791 4069
rect 6733 4060 6745 4063
rect 6564 4032 6745 4060
rect 6733 4029 6745 4032
rect 6779 4029 6791 4063
rect 6733 4023 6791 4029
rect 6822 4020 6828 4072
rect 6880 4060 6886 4072
rect 7745 4063 7803 4069
rect 6880 4032 7512 4060
rect 6880 4020 6886 4032
rect 6546 3992 6552 4004
rect 5368 3964 6552 3992
rect 4249 3955 4307 3961
rect 6546 3952 6552 3964
rect 6604 3952 6610 4004
rect 7374 3992 7380 4004
rect 7335 3964 7380 3992
rect 7374 3952 7380 3964
rect 7432 3952 7438 4004
rect 7484 3992 7512 4032
rect 7745 4029 7757 4063
rect 7791 4029 7803 4063
rect 7852 4060 7880 4100
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 9217 4063 9275 4069
rect 9217 4060 9229 4063
rect 7852 4032 9229 4060
rect 7745 4023 7803 4029
rect 9217 4029 9229 4032
rect 9263 4029 9275 4063
rect 9217 4023 9275 4029
rect 9401 4063 9459 4069
rect 9401 4029 9413 4063
rect 9447 4060 9459 4063
rect 9674 4060 9680 4072
rect 9447 4032 9680 4060
rect 9447 4029 9459 4032
rect 9401 4023 9459 4029
rect 7760 3992 7788 4023
rect 8570 3992 8576 4004
rect 7484 3964 7788 3992
rect 8220 3964 8576 3992
rect 8220 3924 8248 3964
rect 8570 3952 8576 3964
rect 8628 3992 8634 4004
rect 9232 3992 9260 4023
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 9858 4060 9864 4072
rect 9819 4032 9864 4060
rect 9858 4020 9864 4032
rect 9916 4020 9922 4072
rect 9968 3992 9996 4236
rect 10318 4224 10324 4236
rect 10376 4224 10382 4276
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10560 4236 10605 4264
rect 10560 4224 10566 4236
rect 11698 4224 11704 4276
rect 11756 4264 11762 4276
rect 11793 4267 11851 4273
rect 11793 4264 11805 4267
rect 11756 4236 11805 4264
rect 11756 4224 11762 4236
rect 11793 4233 11805 4236
rect 11839 4233 11851 4267
rect 11793 4227 11851 4233
rect 13814 4224 13820 4276
rect 13872 4224 13878 4276
rect 14090 4264 14096 4276
rect 14051 4236 14096 4264
rect 14090 4224 14096 4236
rect 14148 4224 14154 4276
rect 17037 4267 17095 4273
rect 17037 4233 17049 4267
rect 17083 4264 17095 4267
rect 19518 4264 19524 4276
rect 17083 4236 19524 4264
rect 17083 4233 17095 4236
rect 17037 4227 17095 4233
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 10134 4196 10140 4208
rect 10095 4168 10140 4196
rect 10134 4156 10140 4168
rect 10192 4156 10198 4208
rect 10410 4156 10416 4208
rect 10468 4196 10474 4208
rect 11885 4199 11943 4205
rect 11885 4196 11897 4199
rect 10468 4168 11897 4196
rect 10468 4156 10474 4168
rect 11885 4165 11897 4168
rect 11931 4165 11943 4199
rect 13832 4196 13860 4224
rect 11885 4159 11943 4165
rect 11992 4168 13860 4196
rect 14636 4199 14694 4205
rect 10318 4088 10324 4140
rect 10376 4128 10382 4140
rect 11149 4131 11207 4137
rect 11149 4128 11161 4131
rect 10376 4100 11161 4128
rect 10376 4088 10382 4100
rect 11149 4097 11161 4100
rect 11195 4097 11207 4131
rect 11992 4128 12020 4168
rect 14636 4165 14648 4199
rect 14682 4196 14694 4199
rect 14734 4196 14740 4208
rect 14682 4168 14740 4196
rect 14682 4165 14694 4168
rect 14636 4159 14694 4165
rect 14734 4156 14740 4168
rect 14792 4156 14798 4208
rect 16942 4156 16948 4208
rect 17000 4196 17006 4208
rect 17773 4199 17831 4205
rect 17000 4168 17172 4196
rect 17000 4156 17006 4168
rect 12710 4128 12716 4140
rect 11149 4091 11207 4097
rect 11256 4100 12020 4128
rect 12671 4100 12716 4128
rect 10045 4063 10103 4069
rect 10045 4029 10057 4063
rect 10091 4029 10103 4063
rect 11256 4060 11284 4100
rect 12710 4088 12716 4100
rect 12768 4088 12774 4140
rect 12980 4131 13038 4137
rect 12980 4097 12992 4131
rect 13026 4128 13038 4131
rect 13814 4128 13820 4140
rect 13026 4100 13820 4128
rect 13026 4097 13038 4100
rect 12980 4091 13038 4097
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14366 4128 14372 4140
rect 14327 4100 14372 4128
rect 14366 4088 14372 4100
rect 14424 4088 14430 4140
rect 16206 4128 16212 4140
rect 14476 4100 15424 4128
rect 16167 4100 16212 4128
rect 10045 4023 10103 4029
rect 10520 4032 11284 4060
rect 11701 4063 11759 4069
rect 8628 3964 9168 3992
rect 9232 3964 9996 3992
rect 10060 3992 10088 4023
rect 10410 3992 10416 4004
rect 10060 3964 10416 3992
rect 8628 3952 8634 3964
rect 3804 3896 8248 3924
rect 8294 3884 8300 3936
rect 8352 3924 8358 3936
rect 8389 3927 8447 3933
rect 8389 3924 8401 3927
rect 8352 3896 8401 3924
rect 8352 3884 8358 3896
rect 8389 3893 8401 3896
rect 8435 3893 8447 3927
rect 8389 3887 8447 3893
rect 8478 3884 8484 3936
rect 8536 3924 8542 3936
rect 8757 3927 8815 3933
rect 8757 3924 8769 3927
rect 8536 3896 8769 3924
rect 8536 3884 8542 3896
rect 8757 3893 8769 3896
rect 8803 3893 8815 3927
rect 9140 3924 9168 3964
rect 10410 3952 10416 3964
rect 10468 3952 10474 4004
rect 10520 3924 10548 4032
rect 11701 4029 11713 4063
rect 11747 4029 11759 4063
rect 14476 4060 14504 4100
rect 11701 4023 11759 4029
rect 13740 4032 14504 4060
rect 10686 3952 10692 4004
rect 10744 3992 10750 4004
rect 10965 3995 11023 4001
rect 10965 3992 10977 3995
rect 10744 3964 10977 3992
rect 10744 3952 10750 3964
rect 10965 3961 10977 3964
rect 11011 3961 11023 3995
rect 11716 3992 11744 4023
rect 11882 3992 11888 4004
rect 11716 3964 11888 3992
rect 10965 3955 11023 3961
rect 11882 3952 11888 3964
rect 11940 3952 11946 4004
rect 13740 3992 13768 4032
rect 13648 3964 13768 3992
rect 15396 3992 15424 4100
rect 16206 4088 16212 4100
rect 16264 4088 16270 4140
rect 17144 4128 17172 4168
rect 17773 4165 17785 4199
rect 17819 4196 17831 4199
rect 17862 4196 17868 4208
rect 17819 4168 17868 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 17862 4156 17868 4168
rect 17920 4156 17926 4208
rect 17954 4156 17960 4208
rect 18012 4196 18018 4208
rect 18012 4168 19288 4196
rect 18012 4156 18018 4168
rect 18049 4131 18107 4137
rect 18049 4128 18061 4131
rect 17144 4100 18061 4128
rect 18049 4097 18061 4100
rect 18095 4097 18107 4131
rect 18690 4128 18696 4140
rect 18651 4100 18696 4128
rect 18049 4091 18107 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4097 19211 4131
rect 19260 4128 19288 4168
rect 19613 4131 19671 4137
rect 19613 4128 19625 4131
rect 19260 4100 19625 4128
rect 19153 4091 19211 4097
rect 19613 4097 19625 4100
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 20073 4131 20131 4137
rect 20073 4097 20085 4131
rect 20119 4097 20131 4131
rect 20073 4091 20131 4097
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4128 20775 4131
rect 20806 4128 20812 4140
rect 20763 4100 20812 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 16850 4060 16856 4072
rect 16811 4032 16856 4060
rect 16850 4020 16856 4032
rect 16908 4020 16914 4072
rect 16945 4063 17003 4069
rect 16945 4029 16957 4063
rect 16991 4060 17003 4063
rect 17126 4060 17132 4072
rect 16991 4032 17132 4060
rect 16991 4029 17003 4032
rect 16945 4023 17003 4029
rect 17126 4020 17132 4032
rect 17184 4020 17190 4072
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 19168 4060 19196 4091
rect 17828 4032 19196 4060
rect 17828 4020 17834 4032
rect 19242 4020 19248 4072
rect 19300 4060 19306 4072
rect 20088 4060 20116 4091
rect 20806 4088 20812 4100
rect 20864 4088 20870 4140
rect 20990 4128 20996 4140
rect 20951 4100 20996 4128
rect 20990 4088 20996 4100
rect 21048 4088 21054 4140
rect 19300 4032 20116 4060
rect 19300 4020 19306 4032
rect 15396 3964 17264 3992
rect 9140 3896 10548 3924
rect 12253 3927 12311 3933
rect 8757 3887 8815 3893
rect 12253 3893 12265 3927
rect 12299 3924 12311 3927
rect 12894 3924 12900 3936
rect 12299 3896 12900 3924
rect 12299 3893 12311 3896
rect 12253 3887 12311 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13354 3884 13360 3936
rect 13412 3924 13418 3936
rect 13648 3924 13676 3964
rect 17236 3936 17264 3964
rect 17310 3952 17316 4004
rect 17368 3992 17374 4004
rect 19429 3995 19487 4001
rect 19429 3992 19441 3995
rect 17368 3964 19441 3992
rect 17368 3952 17374 3964
rect 19429 3961 19441 3964
rect 19475 3961 19487 3995
rect 19886 3992 19892 4004
rect 19847 3964 19892 3992
rect 19429 3955 19487 3961
rect 19886 3952 19892 3964
rect 19944 3952 19950 4004
rect 20533 3995 20591 4001
rect 20533 3961 20545 3995
rect 20579 3992 20591 3995
rect 22278 3992 22284 4004
rect 20579 3964 22284 3992
rect 20579 3961 20591 3964
rect 20533 3955 20591 3961
rect 22278 3952 22284 3964
rect 22336 3952 22342 4004
rect 13412 3896 13676 3924
rect 13412 3884 13418 3896
rect 13722 3884 13728 3936
rect 13780 3924 13786 3936
rect 14550 3924 14556 3936
rect 13780 3896 14556 3924
rect 13780 3884 13786 3896
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 15746 3924 15752 3936
rect 15707 3896 15752 3924
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 15838 3884 15844 3936
rect 15896 3924 15902 3936
rect 16025 3927 16083 3933
rect 16025 3924 16037 3927
rect 15896 3896 16037 3924
rect 15896 3884 15902 3896
rect 16025 3893 16037 3896
rect 16071 3893 16083 3927
rect 16025 3887 16083 3893
rect 17218 3884 17224 3936
rect 17276 3884 17282 3936
rect 17405 3927 17463 3933
rect 17405 3893 17417 3927
rect 17451 3924 17463 3927
rect 17586 3924 17592 3936
rect 17451 3896 17592 3924
rect 17451 3893 17463 3896
rect 17405 3887 17463 3893
rect 17586 3884 17592 3896
rect 17644 3884 17650 3936
rect 17770 3884 17776 3936
rect 17828 3924 17834 3936
rect 18969 3927 19027 3933
rect 18969 3924 18981 3927
rect 17828 3896 18981 3924
rect 17828 3884 17834 3896
rect 18969 3893 18981 3896
rect 19015 3893 19027 3927
rect 18969 3887 19027 3893
rect 20990 3884 20996 3936
rect 21048 3924 21054 3936
rect 21177 3927 21235 3933
rect 21177 3924 21189 3927
rect 21048 3896 21189 3924
rect 21048 3884 21054 3896
rect 21177 3893 21189 3896
rect 21223 3893 21235 3927
rect 21177 3887 21235 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 3142 3680 3148 3732
rect 3200 3720 3206 3732
rect 3200 3692 3832 3720
rect 3200 3680 3206 3692
rect 3326 3652 3332 3664
rect 3287 3624 3332 3652
rect 3326 3612 3332 3624
rect 3384 3612 3390 3664
rect 3804 3652 3832 3692
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 4387 3723 4445 3729
rect 4387 3720 4399 3723
rect 3936 3692 4399 3720
rect 3936 3680 3942 3692
rect 4387 3689 4399 3692
rect 4433 3689 4445 3723
rect 4387 3683 4445 3689
rect 5534 3680 5540 3732
rect 5592 3720 5598 3732
rect 6825 3723 6883 3729
rect 6825 3720 6837 3723
rect 5592 3692 6837 3720
rect 5592 3680 5598 3692
rect 6825 3689 6837 3692
rect 6871 3689 6883 3723
rect 6825 3683 6883 3689
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 10873 3723 10931 3729
rect 7156 3692 9536 3720
rect 7156 3680 7162 3692
rect 4522 3652 4528 3664
rect 3804 3624 4528 3652
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 6546 3652 6552 3664
rect 6507 3624 6552 3652
rect 6546 3612 6552 3624
rect 6604 3652 6610 3664
rect 7006 3652 7012 3664
rect 6604 3624 7012 3652
rect 6604 3612 6610 3624
rect 7006 3612 7012 3624
rect 7064 3612 7070 3664
rect 7466 3612 7472 3664
rect 7524 3652 7530 3664
rect 7650 3652 7656 3664
rect 7524 3624 7656 3652
rect 7524 3612 7530 3624
rect 7650 3612 7656 3624
rect 7708 3612 7714 3664
rect 8941 3655 8999 3661
rect 8941 3652 8953 3655
rect 7852 3624 8953 3652
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 2832 3556 2877 3584
rect 2832 3544 2838 3556
rect 3418 3544 3424 3596
rect 3476 3584 3482 3596
rect 5166 3584 5172 3596
rect 3476 3556 5028 3584
rect 5127 3556 5172 3584
rect 3476 3544 3482 3556
rect 2746 3488 4108 3516
rect 2746 3460 2774 3488
rect 2532 3451 2590 3457
rect 2532 3417 2544 3451
rect 2578 3448 2590 3451
rect 2746 3448 2780 3460
rect 2578 3420 2780 3448
rect 2578 3417 2590 3420
rect 2532 3411 2590 3417
rect 2774 3408 2780 3420
rect 2832 3408 2838 3460
rect 3142 3448 3148 3460
rect 3103 3420 3148 3448
rect 3142 3408 3148 3420
rect 3200 3408 3206 3460
rect 1397 3383 1455 3389
rect 1397 3349 1409 3383
rect 1443 3380 1455 3383
rect 1578 3380 1584 3392
rect 1443 3352 1584 3380
rect 1443 3349 1455 3352
rect 1397 3343 1455 3349
rect 1578 3340 1584 3352
rect 1636 3340 1642 3392
rect 4080 3380 4108 3488
rect 4522 3476 4528 3528
rect 4580 3516 4586 3528
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 4580 3488 4629 3516
rect 4580 3476 4586 3488
rect 4617 3485 4629 3488
rect 4663 3485 4675 3519
rect 5000 3516 5028 3556
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 7377 3587 7435 3593
rect 7377 3584 7389 3587
rect 6196 3556 7389 3584
rect 5718 3516 5724 3528
rect 5000 3488 5724 3516
rect 4617 3479 4675 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 4430 3408 4436 3460
rect 4488 3448 4494 3460
rect 5414 3451 5472 3457
rect 5414 3448 5426 3451
rect 4488 3420 5426 3448
rect 4488 3408 4494 3420
rect 5414 3417 5426 3420
rect 5460 3448 5472 3451
rect 6196 3448 6224 3556
rect 7377 3553 7389 3556
rect 7423 3553 7435 3587
rect 7377 3547 7435 3553
rect 5460 3420 6224 3448
rect 7285 3451 7343 3457
rect 5460 3417 5472 3420
rect 5414 3411 5472 3417
rect 7285 3417 7297 3451
rect 7331 3448 7343 3451
rect 7852 3448 7880 3624
rect 8941 3621 8953 3624
rect 8987 3621 8999 3655
rect 8941 3615 8999 3621
rect 8018 3584 8024 3596
rect 7979 3556 8024 3584
rect 8018 3544 8024 3556
rect 8076 3544 8082 3596
rect 8113 3587 8171 3593
rect 8113 3553 8125 3587
rect 8159 3584 8171 3587
rect 8478 3584 8484 3596
rect 8159 3556 8484 3584
rect 8159 3553 8171 3556
rect 8113 3547 8171 3553
rect 8478 3544 8484 3556
rect 8536 3544 8542 3596
rect 9508 3593 9536 3692
rect 10873 3689 10885 3723
rect 10919 3720 10931 3723
rect 11146 3720 11152 3732
rect 10919 3692 11152 3720
rect 10919 3689 10931 3692
rect 10873 3683 10931 3689
rect 11146 3680 11152 3692
rect 11204 3680 11210 3732
rect 16761 3723 16819 3729
rect 16761 3689 16773 3723
rect 16807 3720 16819 3723
rect 17034 3720 17040 3732
rect 16807 3692 17040 3720
rect 16807 3689 16819 3692
rect 16761 3683 16819 3689
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 17954 3680 17960 3732
rect 18012 3720 18018 3732
rect 18230 3720 18236 3732
rect 18012 3692 18236 3720
rect 18012 3680 18018 3692
rect 18230 3680 18236 3692
rect 18288 3680 18294 3732
rect 10137 3655 10195 3661
rect 10137 3621 10149 3655
rect 10183 3652 10195 3655
rect 11054 3652 11060 3664
rect 10183 3624 11060 3652
rect 10183 3621 10195 3624
rect 10137 3615 10195 3621
rect 11054 3612 11060 3624
rect 11112 3612 11118 3664
rect 12066 3652 12072 3664
rect 11348 3624 12072 3652
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 11238 3584 11244 3596
rect 9493 3547 9551 3553
rect 9646 3556 11244 3584
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8205 3519 8263 3525
rect 8205 3516 8217 3519
rect 7984 3488 8217 3516
rect 7984 3476 7990 3488
rect 8205 3485 8217 3488
rect 8251 3485 8263 3519
rect 8205 3479 8263 3485
rect 8312 3488 9076 3516
rect 7331 3420 7880 3448
rect 7331 3417 7343 3420
rect 7285 3411 7343 3417
rect 6822 3380 6828 3392
rect 4080 3352 6828 3380
rect 6822 3340 6828 3352
rect 6880 3340 6886 3392
rect 7190 3380 7196 3392
rect 7151 3352 7196 3380
rect 7190 3340 7196 3352
rect 7248 3340 7254 3392
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 8312 3380 8340 3488
rect 8570 3380 8576 3392
rect 7432 3352 8340 3380
rect 8531 3352 8576 3380
rect 7432 3340 7438 3352
rect 8570 3340 8576 3352
rect 8628 3340 8634 3392
rect 9048 3380 9076 3488
rect 9214 3476 9220 3528
rect 9272 3516 9278 3528
rect 9309 3519 9367 3525
rect 9309 3516 9321 3519
rect 9272 3488 9321 3516
rect 9272 3476 9278 3488
rect 9309 3485 9321 3488
rect 9355 3516 9367 3519
rect 9646 3516 9674 3556
rect 11238 3544 11244 3556
rect 11296 3544 11302 3596
rect 9355 3488 9674 3516
rect 9953 3519 10011 3525
rect 9355 3485 9367 3488
rect 9309 3479 9367 3485
rect 9953 3485 9965 3519
rect 9999 3516 10011 3519
rect 10870 3516 10876 3528
rect 9999 3488 10876 3516
rect 9999 3485 10011 3488
rect 9953 3479 10011 3485
rect 10870 3476 10876 3488
rect 10928 3476 10934 3528
rect 11054 3476 11060 3528
rect 11112 3516 11118 3528
rect 11348 3516 11376 3624
rect 12066 3612 12072 3624
rect 12124 3652 12130 3664
rect 17862 3652 17868 3664
rect 12124 3624 17868 3652
rect 12124 3612 12130 3624
rect 17862 3612 17868 3624
rect 17920 3612 17926 3664
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 19797 3655 19855 3661
rect 19797 3652 19809 3655
rect 19116 3624 19809 3652
rect 19116 3612 19122 3624
rect 19797 3621 19809 3624
rect 19843 3621 19855 3655
rect 19797 3615 19855 3621
rect 12805 3587 12863 3593
rect 12805 3553 12817 3587
rect 12851 3584 12863 3587
rect 13630 3584 13636 3596
rect 12851 3556 13636 3584
rect 12851 3553 12863 3556
rect 12805 3547 12863 3553
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 14274 3584 14280 3596
rect 14235 3556 14280 3584
rect 14274 3544 14280 3556
rect 14332 3544 14338 3596
rect 15289 3587 15347 3593
rect 15289 3553 15301 3587
rect 15335 3553 15347 3587
rect 15289 3547 15347 3553
rect 12158 3516 12164 3528
rect 11112 3488 11376 3516
rect 12119 3488 12164 3516
rect 11112 3476 11118 3488
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12894 3516 12900 3528
rect 12855 3488 12900 3516
rect 12894 3476 12900 3488
rect 12952 3476 12958 3528
rect 12989 3519 13047 3525
rect 12989 3485 13001 3519
rect 13035 3516 13047 3519
rect 15304 3516 15332 3547
rect 15470 3544 15476 3596
rect 15528 3584 15534 3596
rect 16022 3584 16028 3596
rect 15528 3556 16028 3584
rect 15528 3544 15534 3556
rect 16022 3544 16028 3556
rect 16080 3544 16086 3596
rect 20070 3584 20076 3596
rect 19628 3556 20076 3584
rect 15746 3516 15752 3528
rect 13035 3488 15271 3516
rect 15304 3488 15752 3516
rect 13035 3485 13047 3488
rect 12989 3479 13047 3485
rect 9401 3451 9459 3457
rect 9401 3417 9413 3451
rect 9447 3448 9459 3451
rect 10594 3448 10600 3460
rect 9447 3420 10600 3448
rect 9447 3417 9459 3420
rect 9401 3411 9459 3417
rect 10594 3408 10600 3420
rect 10652 3408 10658 3460
rect 13633 3451 13691 3457
rect 13633 3448 13645 3451
rect 12406 3420 13645 3448
rect 10226 3380 10232 3392
rect 9048 3352 10232 3380
rect 10226 3340 10232 3352
rect 10284 3340 10290 3392
rect 10318 3340 10324 3392
rect 10376 3380 10382 3392
rect 12406 3380 12434 3420
rect 13633 3417 13645 3420
rect 13679 3417 13691 3451
rect 13633 3411 13691 3417
rect 14461 3451 14519 3457
rect 14461 3417 14473 3451
rect 14507 3448 14519 3451
rect 14642 3448 14648 3460
rect 14507 3420 14648 3448
rect 14507 3417 14519 3420
rect 14461 3411 14519 3417
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 15243 3448 15271 3488
rect 15746 3476 15752 3488
rect 15804 3516 15810 3528
rect 16117 3519 16175 3525
rect 16117 3516 16129 3519
rect 15804 3488 16129 3516
rect 15804 3476 15810 3488
rect 16117 3485 16129 3488
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 16574 3476 16580 3528
rect 16632 3516 16638 3528
rect 17037 3519 17095 3525
rect 17037 3516 17049 3519
rect 16632 3488 17049 3516
rect 16632 3476 16638 3488
rect 17037 3485 17049 3488
rect 17083 3485 17095 3519
rect 17678 3516 17684 3528
rect 17639 3488 17684 3516
rect 17037 3479 17095 3485
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 18598 3516 18604 3528
rect 18559 3488 18604 3516
rect 18598 3476 18604 3488
rect 18656 3476 18662 3528
rect 19628 3525 19656 3556
rect 20070 3544 20076 3556
rect 20128 3544 20134 3596
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3485 19671 3519
rect 20162 3516 20168 3528
rect 20123 3488 20168 3516
rect 19613 3479 19671 3485
rect 20162 3476 20168 3488
rect 20220 3476 20226 3528
rect 20530 3476 20536 3528
rect 20588 3516 20594 3528
rect 20717 3519 20775 3525
rect 20717 3516 20729 3519
rect 20588 3488 20729 3516
rect 20588 3476 20594 3488
rect 20717 3485 20729 3488
rect 20763 3485 20775 3519
rect 20717 3479 20775 3485
rect 17957 3451 18015 3457
rect 17957 3448 17969 3451
rect 15243 3420 16068 3448
rect 13354 3380 13360 3392
rect 10376 3352 12434 3380
rect 13315 3352 13360 3380
rect 10376 3340 10382 3352
rect 13354 3340 13360 3352
rect 13412 3340 13418 3392
rect 14366 3380 14372 3392
rect 14327 3352 14372 3380
rect 14366 3340 14372 3352
rect 14424 3340 14430 3392
rect 14829 3383 14887 3389
rect 14829 3349 14841 3383
rect 14875 3380 14887 3383
rect 15381 3383 15439 3389
rect 15381 3380 15393 3383
rect 14875 3352 15393 3380
rect 14875 3349 14887 3352
rect 14829 3343 14887 3349
rect 15381 3349 15393 3352
rect 15427 3349 15439 3383
rect 15381 3343 15439 3349
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 15841 3383 15899 3389
rect 15528 3352 15573 3380
rect 15528 3340 15534 3352
rect 15841 3349 15853 3383
rect 15887 3380 15899 3383
rect 15930 3380 15936 3392
rect 15887 3352 15936 3380
rect 15887 3349 15899 3352
rect 15841 3343 15899 3349
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16040 3380 16068 3420
rect 16316 3420 17969 3448
rect 16316 3380 16344 3420
rect 17957 3417 17969 3420
rect 18003 3417 18015 3451
rect 17957 3411 18015 3417
rect 18690 3408 18696 3460
rect 18748 3448 18754 3460
rect 21269 3451 21327 3457
rect 21269 3448 21281 3451
rect 18748 3420 21281 3448
rect 18748 3408 18754 3420
rect 21269 3417 21281 3420
rect 21315 3417 21327 3451
rect 21269 3411 21327 3417
rect 16040 3352 16344 3380
rect 16942 3340 16948 3392
rect 17000 3380 17006 3392
rect 18417 3383 18475 3389
rect 18417 3380 18429 3383
rect 17000 3352 18429 3380
rect 17000 3340 17006 3352
rect 18417 3349 18429 3352
rect 18463 3349 18475 3383
rect 18417 3343 18475 3349
rect 18506 3340 18512 3392
rect 18564 3380 18570 3392
rect 19245 3383 19303 3389
rect 19245 3380 19257 3383
rect 18564 3352 19257 3380
rect 18564 3340 18570 3352
rect 19245 3349 19257 3352
rect 19291 3349 19303 3383
rect 19245 3343 19303 3349
rect 20070 3340 20076 3392
rect 20128 3380 20134 3392
rect 20349 3383 20407 3389
rect 20349 3380 20361 3383
rect 20128 3352 20361 3380
rect 20128 3340 20134 3352
rect 20349 3349 20361 3352
rect 20395 3349 20407 3383
rect 20349 3343 20407 3349
rect 20530 3340 20536 3392
rect 20588 3380 20594 3392
rect 20901 3383 20959 3389
rect 20901 3380 20913 3383
rect 20588 3352 20913 3380
rect 20588 3340 20594 3352
rect 20901 3349 20913 3352
rect 20947 3349 20959 3383
rect 20901 3343 20959 3349
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 2682 3176 2688 3188
rect 2643 3148 2688 3176
rect 2682 3136 2688 3148
rect 2740 3136 2746 3188
rect 2774 3136 2780 3188
rect 2832 3176 2838 3188
rect 2961 3179 3019 3185
rect 2961 3176 2973 3179
rect 2832 3148 2973 3176
rect 2832 3136 2838 3148
rect 2961 3145 2973 3148
rect 3007 3145 3019 3179
rect 2961 3139 3019 3145
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3145 4675 3179
rect 4617 3139 4675 3145
rect 1854 3068 1860 3120
rect 1912 3108 1918 3120
rect 4430 3108 4436 3120
rect 1912 3080 4436 3108
rect 1912 3068 1918 3080
rect 4430 3068 4436 3080
rect 4488 3108 4494 3120
rect 4632 3108 4660 3139
rect 4706 3136 4712 3188
rect 4764 3176 4770 3188
rect 6365 3179 6423 3185
rect 4764 3148 6132 3176
rect 4764 3136 4770 3148
rect 6104 3108 6132 3148
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 7282 3176 7288 3188
rect 6411 3148 7288 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 7282 3136 7288 3148
rect 7340 3136 7346 3188
rect 8941 3179 8999 3185
rect 8941 3176 8953 3179
rect 8588 3148 8953 3176
rect 4488 3080 4660 3108
rect 5184 3080 6040 3108
rect 6104 3080 7972 3108
rect 4488 3068 4494 3080
rect 5184 3052 5212 3080
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3040 2007 3043
rect 2406 3040 2412 3052
rect 1995 3012 2412 3040
rect 1995 3009 2007 3012
rect 1949 3003 2007 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 2498 3000 2504 3052
rect 2556 3040 2562 3052
rect 4085 3043 4143 3049
rect 2556 3012 2601 3040
rect 2556 3000 2562 3012
rect 4085 3009 4097 3043
rect 4131 3040 4143 3043
rect 4341 3043 4399 3049
rect 4131 3012 4292 3040
rect 4131 3009 4143 3012
rect 4085 3003 4143 3009
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2774 2972 2780 2984
rect 2271 2944 2780 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2774 2932 2780 2944
rect 2832 2932 2838 2984
rect 4264 2972 4292 3012
rect 4341 3009 4353 3043
rect 4387 3040 4399 3043
rect 5166 3040 5172 3052
rect 4387 3012 5172 3040
rect 4387 3009 4399 3012
rect 4341 3003 4399 3009
rect 5166 3000 5172 3012
rect 5224 3000 5230 3052
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 6012 3049 6040 3080
rect 5730 3043 5788 3049
rect 5730 3040 5742 3043
rect 5316 3012 5742 3040
rect 5316 3000 5322 3012
rect 5730 3009 5742 3012
rect 5776 3040 5788 3043
rect 5997 3043 6055 3049
rect 5776 3012 5948 3040
rect 5776 3009 5788 3012
rect 5730 3003 5788 3009
rect 4430 2972 4436 2984
rect 4264 2944 4436 2972
rect 4430 2932 4436 2944
rect 4488 2932 4494 2984
rect 4706 2932 4712 2984
rect 4764 2972 4770 2984
rect 4890 2972 4896 2984
rect 4764 2944 4896 2972
rect 4764 2932 4770 2944
rect 4890 2932 4896 2944
rect 4948 2932 4954 2984
rect 5920 2972 5948 3012
rect 5997 3009 6009 3043
rect 6043 3009 6055 3043
rect 5997 3003 6055 3009
rect 7009 3043 7067 3049
rect 7009 3009 7021 3043
rect 7055 3040 7067 3043
rect 7834 3040 7840 3052
rect 7055 3012 7840 3040
rect 7055 3009 7067 3012
rect 7009 3003 7067 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 7944 3040 7972 3080
rect 8018 3068 8024 3120
rect 8076 3108 8082 3120
rect 8420 3111 8478 3117
rect 8420 3108 8432 3111
rect 8076 3080 8432 3108
rect 8076 3068 8082 3080
rect 8420 3077 8432 3080
rect 8466 3108 8478 3111
rect 8588 3108 8616 3148
rect 8941 3145 8953 3148
rect 8987 3176 8999 3179
rect 9858 3176 9864 3188
rect 8987 3148 9864 3176
rect 8987 3145 8999 3148
rect 8941 3139 8999 3145
rect 9858 3136 9864 3148
rect 9916 3136 9922 3188
rect 10042 3136 10048 3188
rect 10100 3176 10106 3188
rect 10100 3148 10456 3176
rect 10100 3136 10106 3148
rect 10428 3108 10456 3148
rect 11790 3136 11796 3188
rect 11848 3176 11854 3188
rect 12526 3176 12532 3188
rect 11848 3148 12532 3176
rect 11848 3136 11854 3148
rect 12526 3136 12532 3148
rect 12584 3136 12590 3188
rect 13630 3176 13636 3188
rect 13591 3148 13636 3176
rect 13630 3136 13636 3148
rect 13688 3136 13694 3188
rect 13814 3136 13820 3188
rect 13872 3176 13878 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 13872 3148 14565 3176
rect 13872 3136 13878 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 15473 3179 15531 3185
rect 15473 3176 15485 3179
rect 15436 3148 15485 3176
rect 15436 3136 15442 3148
rect 15473 3145 15485 3148
rect 15519 3145 15531 3179
rect 15473 3139 15531 3145
rect 15654 3136 15660 3188
rect 15712 3176 15718 3188
rect 17313 3179 17371 3185
rect 17313 3176 17325 3179
rect 15712 3148 17325 3176
rect 15712 3136 15718 3148
rect 17313 3145 17325 3148
rect 17359 3145 17371 3179
rect 17313 3139 17371 3145
rect 17862 3136 17868 3188
rect 17920 3176 17926 3188
rect 18417 3179 18475 3185
rect 18417 3176 18429 3179
rect 17920 3148 18429 3176
rect 17920 3136 17926 3148
rect 18417 3145 18429 3148
rect 18463 3145 18475 3179
rect 18417 3139 18475 3145
rect 10597 3111 10655 3117
rect 10597 3108 10609 3111
rect 8466 3080 8616 3108
rect 8680 3080 10364 3108
rect 10428 3080 10609 3108
rect 8466 3077 8478 3080
rect 8420 3071 8478 3077
rect 8680 3049 8708 3080
rect 8665 3043 8723 3049
rect 7944 3012 8616 3040
rect 7098 2972 7104 2984
rect 5920 2944 7104 2972
rect 7098 2932 7104 2944
rect 7156 2932 7162 2984
rect 8588 2972 8616 3012
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 9122 3000 9128 3052
rect 9180 3040 9186 3052
rect 9490 3040 9496 3052
rect 9180 3012 9496 3040
rect 9180 3000 9186 3012
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10336 3049 10364 3080
rect 10597 3077 10609 3080
rect 10643 3077 10655 3111
rect 10597 3071 10655 3077
rect 11238 3068 11244 3120
rect 11296 3108 11302 3120
rect 12342 3108 12348 3120
rect 11296 3080 12348 3108
rect 11296 3068 11302 3080
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 13078 3108 13084 3120
rect 12535 3080 13084 3108
rect 10054 3043 10112 3049
rect 10054 3040 10066 3043
rect 9732 3012 10066 3040
rect 9732 3000 9738 3012
rect 10054 3009 10066 3012
rect 10100 3009 10112 3043
rect 10054 3003 10112 3009
rect 10321 3044 10379 3049
rect 10321 3043 10456 3044
rect 10321 3009 10333 3043
rect 10367 3040 10456 3043
rect 10965 3043 11023 3049
rect 10367 3016 10916 3040
rect 10367 3009 10379 3016
rect 10428 3012 10916 3016
rect 10321 3003 10379 3009
rect 10888 2972 10916 3012
rect 10965 3009 10977 3043
rect 11011 3040 11023 3043
rect 11698 3040 11704 3052
rect 11011 3012 11704 3040
rect 11011 3009 11023 3012
rect 10965 3003 11023 3009
rect 11698 3000 11704 3012
rect 11756 3000 11762 3052
rect 11977 3043 12035 3049
rect 11977 3009 11989 3043
rect 12023 3040 12035 3043
rect 12066 3040 12072 3052
rect 12023 3012 12072 3040
rect 12023 3009 12035 3012
rect 11977 3003 12035 3009
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 12535 3049 12563 3080
rect 13078 3068 13084 3080
rect 13136 3068 13142 3120
rect 12520 3043 12578 3049
rect 12520 3009 12532 3043
rect 12566 3009 12578 3043
rect 13648 3040 13676 3136
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 18966 3108 18972 3120
rect 13780 3080 18972 3108
rect 13780 3068 13786 3080
rect 18966 3068 18972 3080
rect 19024 3068 19030 3120
rect 19794 3108 19800 3120
rect 19168 3080 19800 3108
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13648 3012 13921 3040
rect 12520 3003 12578 3009
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 14550 3000 14556 3052
rect 14608 3040 14614 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14608 3012 14841 3040
rect 14608 3000 14614 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 14829 3003 14887 3009
rect 16025 3043 16083 3049
rect 16025 3009 16037 3043
rect 16071 3040 16083 3043
rect 16114 3040 16120 3052
rect 16071 3012 16120 3040
rect 16071 3009 16083 3012
rect 16025 3003 16083 3009
rect 16114 3000 16120 3012
rect 16172 3000 16178 3052
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17310 3040 17316 3052
rect 16991 3012 17316 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17494 3040 17500 3052
rect 17455 3012 17500 3040
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3009 18107 3043
rect 18049 3003 18107 3009
rect 18601 3043 18659 3049
rect 18601 3009 18613 3043
rect 18647 3040 18659 3043
rect 18874 3040 18880 3052
rect 18647 3012 18880 3040
rect 18647 3009 18659 3012
rect 18601 3003 18659 3009
rect 11146 2972 11152 2984
rect 8588 2944 8708 2972
rect 10888 2944 11152 2972
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 3326 2904 3332 2916
rect 624 2876 3332 2904
rect 624 2864 630 2876
rect 3326 2864 3332 2876
rect 3384 2864 3390 2916
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1302 2836 1308 2848
rect 256 2808 1308 2836
rect 256 2796 262 2808
rect 1302 2796 1308 2808
rect 1360 2836 1366 2848
rect 2222 2836 2228 2848
rect 1360 2808 2228 2836
rect 1360 2796 1366 2808
rect 2222 2796 2228 2808
rect 2280 2796 2286 2848
rect 2774 2796 2780 2848
rect 2832 2836 2838 2848
rect 6546 2836 6552 2848
rect 2832 2808 6552 2836
rect 2832 2796 2838 2808
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2836 7343 2839
rect 8018 2836 8024 2848
rect 7331 2808 8024 2836
rect 7331 2805 7343 2808
rect 7285 2799 7343 2805
rect 8018 2796 8024 2808
rect 8076 2796 8082 2848
rect 8680 2836 8708 2944
rect 11146 2932 11152 2944
rect 11204 2972 11210 2984
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11204 2944 12265 2972
rect 11204 2932 11210 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12253 2935 12311 2941
rect 14274 2932 14280 2984
rect 14332 2972 14338 2984
rect 18064 2972 18092 3003
rect 18874 3000 18880 3012
rect 18932 3000 18938 3052
rect 19168 3049 19196 3080
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 19610 3000 19616 3052
rect 19668 3040 19674 3052
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 19668 3012 19717 3040
rect 19668 3000 19674 3012
rect 19705 3009 19717 3012
rect 19751 3009 19763 3043
rect 21358 3040 21364 3052
rect 21319 3012 21364 3040
rect 19705 3003 19763 3009
rect 21358 3000 21364 3012
rect 21416 3040 21422 3052
rect 22738 3040 22744 3052
rect 21416 3012 22744 3040
rect 21416 3000 21422 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 19978 2972 19984 2984
rect 14332 2944 15976 2972
rect 18064 2944 19984 2972
rect 14332 2932 14338 2944
rect 12158 2904 12164 2916
rect 11164 2876 12164 2904
rect 11054 2836 11060 2848
rect 8680 2808 11060 2836
rect 11054 2796 11060 2808
rect 11112 2796 11118 2848
rect 11164 2845 11192 2876
rect 12158 2864 12164 2876
rect 12216 2864 12222 2916
rect 14734 2864 14740 2916
rect 14792 2904 14798 2916
rect 15841 2907 15899 2913
rect 15841 2904 15853 2907
rect 14792 2876 15853 2904
rect 14792 2864 14798 2876
rect 15841 2873 15853 2876
rect 15887 2873 15899 2907
rect 15841 2867 15899 2873
rect 11149 2839 11207 2845
rect 11149 2805 11161 2839
rect 11195 2805 11207 2839
rect 11149 2799 11207 2805
rect 11793 2839 11851 2845
rect 11793 2805 11805 2839
rect 11839 2836 11851 2839
rect 11882 2836 11888 2848
rect 11839 2808 11888 2836
rect 11839 2805 11851 2808
rect 11793 2799 11851 2805
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 15286 2836 15292 2848
rect 12124 2808 15292 2836
rect 12124 2796 12130 2808
rect 15286 2796 15292 2808
rect 15344 2796 15350 2848
rect 15948 2836 15976 2944
rect 19978 2932 19984 2944
rect 20036 2932 20042 2984
rect 20714 2972 20720 2984
rect 20675 2944 20720 2972
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 16390 2864 16396 2916
rect 16448 2904 16454 2916
rect 17865 2907 17923 2913
rect 17865 2904 17877 2907
rect 16448 2876 17877 2904
rect 16448 2864 16454 2876
rect 17865 2873 17877 2876
rect 17911 2873 17923 2907
rect 17865 2867 17923 2873
rect 16761 2839 16819 2845
rect 16761 2836 16773 2839
rect 15948 2808 16773 2836
rect 16761 2805 16773 2808
rect 16807 2805 16819 2839
rect 16761 2799 16819 2805
rect 18690 2796 18696 2848
rect 18748 2836 18754 2848
rect 18969 2839 19027 2845
rect 18969 2836 18981 2839
rect 18748 2808 18981 2836
rect 18748 2796 18754 2808
rect 18969 2805 18981 2808
rect 19015 2805 19027 2839
rect 18969 2799 19027 2805
rect 19610 2796 19616 2848
rect 19668 2836 19674 2848
rect 19889 2839 19947 2845
rect 19889 2836 19901 2839
rect 19668 2808 19901 2836
rect 19668 2796 19674 2808
rect 19889 2805 19901 2808
rect 19935 2805 19947 2839
rect 19889 2799 19947 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7377 2635 7435 2641
rect 7377 2632 7389 2635
rect 7248 2604 7389 2632
rect 7248 2592 7254 2604
rect 7377 2601 7389 2604
rect 7423 2601 7435 2635
rect 7377 2595 7435 2601
rect 7558 2592 7564 2644
rect 7616 2632 7622 2644
rect 7837 2635 7895 2641
rect 7837 2632 7849 2635
rect 7616 2604 7849 2632
rect 7616 2592 7622 2604
rect 7837 2601 7849 2604
rect 7883 2601 7895 2635
rect 7837 2595 7895 2601
rect 8018 2592 8024 2644
rect 8076 2632 8082 2644
rect 10134 2632 10140 2644
rect 8076 2604 9996 2632
rect 10095 2604 10140 2632
rect 8076 2592 8082 2604
rect 5258 2564 5264 2576
rect 1964 2536 5264 2564
rect 1964 2505 1992 2536
rect 5258 2524 5264 2536
rect 5316 2524 5322 2576
rect 6638 2524 6644 2576
rect 6696 2564 6702 2576
rect 8202 2564 8208 2576
rect 6696 2536 8208 2564
rect 6696 2524 6702 2536
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 9674 2524 9680 2576
rect 9732 2524 9738 2576
rect 9968 2564 9996 2604
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 10410 2632 10416 2644
rect 10371 2604 10416 2632
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10870 2592 10876 2644
rect 10928 2632 10934 2644
rect 11517 2635 11575 2641
rect 11517 2632 11529 2635
rect 10928 2604 11529 2632
rect 10928 2592 10934 2604
rect 11517 2601 11529 2604
rect 11563 2601 11575 2635
rect 11517 2595 11575 2601
rect 13446 2592 13452 2644
rect 13504 2632 13510 2644
rect 15749 2635 15807 2641
rect 15749 2632 15761 2635
rect 13504 2604 15761 2632
rect 13504 2592 13510 2604
rect 15749 2601 15761 2604
rect 15795 2601 15807 2635
rect 15749 2595 15807 2601
rect 16114 2592 16120 2644
rect 16172 2632 16178 2644
rect 16172 2604 17448 2632
rect 16172 2592 16178 2604
rect 9968 2536 12112 2564
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 2222 2496 2228 2508
rect 2183 2468 2228 2496
rect 1949 2459 2007 2465
rect 2222 2456 2228 2468
rect 2280 2456 2286 2508
rect 3326 2496 3332 2508
rect 3287 2468 3332 2496
rect 3326 2456 3332 2468
rect 3384 2456 3390 2508
rect 4341 2499 4399 2505
rect 4341 2465 4353 2499
rect 4387 2496 4399 2499
rect 4706 2496 4712 2508
rect 4387 2468 4712 2496
rect 4387 2465 4399 2468
rect 4341 2459 4399 2465
rect 4706 2456 4712 2468
rect 4764 2456 4770 2508
rect 4798 2456 4804 2508
rect 4856 2496 4862 2508
rect 5445 2499 5503 2505
rect 5445 2496 5457 2499
rect 4856 2468 5457 2496
rect 4856 2456 4862 2468
rect 5445 2465 5457 2468
rect 5491 2465 5503 2499
rect 5445 2459 5503 2465
rect 6825 2499 6883 2505
rect 6825 2465 6837 2499
rect 6871 2496 6883 2499
rect 7098 2496 7104 2508
rect 6871 2468 7104 2496
rect 6871 2465 6883 2468
rect 6825 2459 6883 2465
rect 7098 2456 7104 2468
rect 7156 2456 7162 2508
rect 8481 2499 8539 2505
rect 8481 2465 8493 2499
rect 8527 2496 8539 2499
rect 9306 2496 9312 2508
rect 8527 2468 9312 2496
rect 8527 2465 8539 2468
rect 8481 2459 8539 2465
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3234 2388 3240 2440
rect 3292 2428 3298 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 3292 2400 4629 2428
rect 3292 2388 3298 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 5810 2428 5816 2440
rect 5767 2400 5816 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 4062 2320 4068 2372
rect 4120 2360 4126 2372
rect 5736 2360 5764 2391
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 8205 2431 8263 2437
rect 6963 2400 8156 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 8128 2360 8156 2400
rect 8205 2397 8217 2431
rect 8251 2428 8263 2431
rect 8294 2428 8300 2440
rect 8251 2400 8300 2428
rect 8251 2397 8263 2400
rect 8205 2391 8263 2397
rect 8294 2388 8300 2400
rect 8352 2388 8358 2440
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 8496 2428 8524 2459
rect 9306 2456 9312 2468
rect 9364 2456 9370 2508
rect 9585 2499 9643 2505
rect 9585 2465 9597 2499
rect 9631 2496 9643 2499
rect 9692 2496 9720 2524
rect 10962 2496 10968 2508
rect 9631 2468 9720 2496
rect 10923 2468 10968 2496
rect 9631 2465 9643 2468
rect 9585 2459 9643 2465
rect 10962 2456 10968 2468
rect 11020 2456 11026 2508
rect 12084 2505 12112 2536
rect 12526 2524 12532 2576
rect 12584 2564 12590 2576
rect 13541 2567 13599 2573
rect 13541 2564 13553 2567
rect 12584 2536 13553 2564
rect 12584 2524 12590 2536
rect 13541 2533 13553 2536
rect 13587 2533 13599 2567
rect 13541 2527 13599 2533
rect 13630 2524 13636 2576
rect 13688 2564 13694 2576
rect 13688 2536 16160 2564
rect 13688 2524 13694 2536
rect 12069 2499 12127 2505
rect 12069 2465 12081 2499
rect 12115 2465 12127 2499
rect 12069 2459 12127 2465
rect 8444 2400 8524 2428
rect 8444 2388 8450 2400
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8720 2400 8953 2428
rect 8720 2388 8726 2400
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 9674 2428 9680 2440
rect 8941 2391 8999 2397
rect 9048 2400 9680 2428
rect 9048 2360 9076 2400
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 9950 2428 9956 2440
rect 9732 2400 9956 2428
rect 9732 2388 9738 2400
rect 9950 2388 9956 2400
rect 10008 2388 10014 2440
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 10560 2400 11989 2428
rect 10560 2388 10566 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 12084 2428 12112 2459
rect 12158 2456 12164 2508
rect 12216 2496 12222 2508
rect 12216 2468 15608 2496
rect 12216 2456 12222 2468
rect 12529 2431 12587 2437
rect 12529 2428 12541 2431
rect 12084 2400 12541 2428
rect 11977 2391 12035 2397
rect 12529 2397 12541 2400
rect 12575 2397 12587 2431
rect 13630 2428 13636 2440
rect 12529 2391 12587 2397
rect 12636 2400 13636 2428
rect 12636 2360 12664 2400
rect 13630 2388 13636 2400
rect 13688 2388 13694 2440
rect 13725 2431 13783 2437
rect 13725 2397 13737 2431
rect 13771 2428 13783 2431
rect 13814 2428 13820 2440
rect 13771 2400 13820 2428
rect 13771 2397 13783 2400
rect 13725 2391 13783 2397
rect 13814 2388 13820 2400
rect 13872 2388 13878 2440
rect 14090 2428 14096 2440
rect 14051 2400 14096 2428
rect 14090 2388 14096 2400
rect 14148 2388 14154 2440
rect 15286 2428 15292 2440
rect 15247 2400 15292 2428
rect 15286 2388 15292 2400
rect 15344 2388 15350 2440
rect 15580 2437 15608 2468
rect 16132 2437 16160 2536
rect 16206 2524 16212 2576
rect 16264 2564 16270 2576
rect 16853 2567 16911 2573
rect 16853 2564 16865 2567
rect 16264 2536 16865 2564
rect 16264 2524 16270 2536
rect 16853 2533 16865 2536
rect 16899 2533 16911 2567
rect 16853 2527 16911 2533
rect 17313 2567 17371 2573
rect 17313 2533 17325 2567
rect 17359 2533 17371 2567
rect 17420 2564 17448 2604
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 19337 2635 19395 2641
rect 19337 2632 19349 2635
rect 17552 2604 19349 2632
rect 17552 2592 17558 2604
rect 19337 2601 19349 2604
rect 19383 2601 19395 2635
rect 19337 2595 19395 2601
rect 17865 2567 17923 2573
rect 17865 2564 17877 2567
rect 17420 2536 17877 2564
rect 17313 2527 17371 2533
rect 17865 2533 17877 2536
rect 17911 2533 17923 2567
rect 17865 2527 17923 2533
rect 17328 2496 17356 2527
rect 18322 2524 18328 2576
rect 18380 2564 18386 2576
rect 19889 2567 19947 2573
rect 19889 2564 19901 2567
rect 18380 2536 19901 2564
rect 18380 2524 18386 2536
rect 19889 2533 19901 2536
rect 19935 2533 19947 2567
rect 19889 2527 19947 2533
rect 19978 2524 19984 2576
rect 20036 2564 20042 2576
rect 20036 2536 21128 2564
rect 20036 2524 20042 2536
rect 20806 2496 20812 2508
rect 16224 2468 17356 2496
rect 18616 2468 20812 2496
rect 15565 2431 15623 2437
rect 15565 2397 15577 2431
rect 15611 2397 15623 2431
rect 15565 2391 15623 2397
rect 16117 2431 16175 2437
rect 16117 2397 16129 2431
rect 16163 2397 16175 2431
rect 16117 2391 16175 2397
rect 4120 2332 5764 2360
rect 6886 2332 7972 2360
rect 8128 2332 9076 2360
rect 9140 2332 12664 2360
rect 4120 2320 4126 2332
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 6886 2292 6914 2332
rect 5776 2264 6914 2292
rect 7009 2295 7067 2301
rect 5776 2252 5782 2264
rect 7009 2261 7021 2295
rect 7055 2292 7067 2295
rect 7282 2292 7288 2304
rect 7055 2264 7288 2292
rect 7055 2261 7067 2264
rect 7009 2255 7067 2261
rect 7282 2252 7288 2264
rect 7340 2252 7346 2304
rect 7944 2292 7972 2332
rect 9140 2301 9168 2332
rect 12986 2320 12992 2372
rect 13044 2360 13050 2372
rect 13044 2332 15148 2360
rect 13044 2320 13050 2332
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 7944 2264 8309 2292
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8297 2255 8355 2261
rect 9125 2295 9183 2301
rect 9125 2261 9137 2295
rect 9171 2261 9183 2295
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9125 2255 9183 2261
rect 9766 2252 9772 2264
rect 9824 2252 9830 2304
rect 10134 2252 10140 2304
rect 10192 2292 10198 2304
rect 10781 2295 10839 2301
rect 10781 2292 10793 2295
rect 10192 2264 10793 2292
rect 10192 2252 10198 2264
rect 10781 2261 10793 2264
rect 10827 2261 10839 2295
rect 10781 2255 10839 2261
rect 10873 2295 10931 2301
rect 10873 2261 10885 2295
rect 10919 2292 10931 2295
rect 10962 2292 10968 2304
rect 10919 2264 10968 2292
rect 10919 2261 10931 2264
rect 10873 2255 10931 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11882 2292 11888 2304
rect 11843 2264 11888 2292
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 13170 2292 13176 2304
rect 13131 2264 13176 2292
rect 13170 2252 13176 2264
rect 13228 2252 13234 2304
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 15120 2301 15148 2332
rect 15194 2320 15200 2372
rect 15252 2360 15258 2372
rect 16224 2360 16252 2468
rect 16669 2431 16727 2437
rect 16669 2428 16681 2431
rect 15252 2332 16252 2360
rect 16546 2400 16681 2428
rect 15252 2320 15258 2332
rect 14737 2295 14795 2301
rect 14737 2292 14749 2295
rect 13320 2264 14749 2292
rect 13320 2252 13326 2264
rect 14737 2261 14749 2264
rect 14783 2261 14795 2295
rect 14737 2255 14795 2261
rect 15105 2295 15163 2301
rect 15105 2261 15117 2295
rect 15151 2261 15163 2295
rect 15105 2255 15163 2261
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2292 16359 2295
rect 16546 2292 16574 2400
rect 16669 2397 16681 2400
rect 16715 2397 16727 2431
rect 16669 2391 16727 2397
rect 17497 2431 17555 2437
rect 17497 2397 17509 2431
rect 17543 2428 17555 2431
rect 17954 2428 17960 2440
rect 17543 2400 17960 2428
rect 17543 2397 17555 2400
rect 17497 2391 17555 2397
rect 17954 2388 17960 2400
rect 18012 2388 18018 2440
rect 18049 2431 18107 2437
rect 18049 2397 18061 2431
rect 18095 2428 18107 2431
rect 18138 2428 18144 2440
rect 18095 2400 18144 2428
rect 18095 2397 18107 2400
rect 18049 2391 18107 2397
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 18616 2437 18644 2468
rect 20806 2456 20812 2468
rect 20864 2456 20870 2508
rect 21100 2505 21128 2536
rect 21085 2499 21143 2505
rect 21085 2465 21097 2499
rect 21131 2465 21143 2499
rect 21085 2459 21143 2465
rect 21361 2499 21419 2505
rect 21361 2465 21373 2499
rect 21407 2496 21419 2499
rect 21450 2496 21456 2508
rect 21407 2468 21456 2496
rect 21407 2465 21419 2468
rect 21361 2459 21419 2465
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 18601 2431 18659 2437
rect 18601 2397 18613 2431
rect 18647 2397 18659 2431
rect 18601 2391 18659 2397
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 19702 2428 19708 2440
rect 19567 2400 19708 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 19702 2388 19708 2400
rect 19760 2388 19766 2440
rect 20073 2431 20131 2437
rect 20073 2397 20085 2431
rect 20119 2428 20131 2431
rect 20622 2428 20628 2440
rect 20119 2400 20628 2428
rect 20119 2397 20131 2400
rect 20073 2391 20131 2397
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 16942 2320 16948 2372
rect 17000 2360 17006 2372
rect 17000 2332 18460 2360
rect 17000 2320 17006 2332
rect 18432 2301 18460 2332
rect 16347 2264 16574 2292
rect 18417 2295 18475 2301
rect 16347 2261 16359 2264
rect 16301 2255 16359 2261
rect 18417 2261 18429 2295
rect 18463 2261 18475 2295
rect 18417 2255 18475 2261
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
rect 8570 2048 8576 2100
rect 8628 2088 8634 2100
rect 11882 2088 11888 2100
rect 8628 2060 11888 2088
rect 8628 2048 8634 2060
rect 11882 2048 11888 2060
rect 11940 2048 11946 2100
rect 15286 2048 15292 2100
rect 15344 2088 15350 2100
rect 18046 2088 18052 2100
rect 15344 2060 18052 2088
rect 15344 2048 15350 2060
rect 18046 2048 18052 2060
rect 18104 2048 18110 2100
rect 8202 1980 8208 2032
rect 8260 2020 8266 2032
rect 13262 2020 13268 2032
rect 8260 1992 13268 2020
rect 8260 1980 8266 1992
rect 13262 1980 13268 1992
rect 13320 1980 13326 2032
rect 13906 1980 13912 2032
rect 13964 2020 13970 2032
rect 16206 2020 16212 2032
rect 13964 1992 16212 2020
rect 13964 1980 13970 1992
rect 16206 1980 16212 1992
rect 16264 1980 16270 2032
rect 4430 1912 4436 1964
rect 4488 1952 4494 1964
rect 13170 1952 13176 1964
rect 4488 1924 13176 1952
rect 4488 1912 4494 1924
rect 13170 1912 13176 1924
rect 13228 1912 13234 1964
rect 13814 1912 13820 1964
rect 13872 1952 13878 1964
rect 17770 1952 17776 1964
rect 13872 1924 17776 1952
rect 13872 1912 13878 1924
rect 17770 1912 17776 1924
rect 17828 1912 17834 1964
rect 3050 1844 3056 1896
rect 3108 1884 3114 1896
rect 3108 1856 6914 1884
rect 3108 1844 3114 1856
rect 6886 1816 6914 1856
rect 7006 1844 7012 1896
rect 7064 1884 7070 1896
rect 14090 1884 14096 1896
rect 7064 1856 14096 1884
rect 7064 1844 7070 1856
rect 14090 1844 14096 1856
rect 14148 1844 14154 1896
rect 6886 1788 7144 1816
rect 1578 1708 1584 1760
rect 1636 1748 1642 1760
rect 1636 1720 6914 1748
rect 1636 1708 1642 1720
rect 6886 1612 6914 1720
rect 7116 1680 7144 1788
rect 9674 1776 9680 1828
rect 9732 1816 9738 1828
rect 15838 1816 15844 1828
rect 9732 1788 15844 1816
rect 9732 1776 9738 1788
rect 15838 1776 15844 1788
rect 15896 1776 15902 1828
rect 7282 1708 7288 1760
rect 7340 1748 7346 1760
rect 9766 1748 9772 1760
rect 7340 1720 9772 1748
rect 7340 1708 7346 1720
rect 9766 1708 9772 1720
rect 9824 1748 9830 1760
rect 10686 1748 10692 1760
rect 9824 1720 10692 1748
rect 9824 1708 9830 1720
rect 10686 1708 10692 1720
rect 10744 1748 10750 1760
rect 14366 1748 14372 1760
rect 10744 1720 14372 1748
rect 10744 1708 10750 1720
rect 14366 1708 14372 1720
rect 14424 1708 14430 1760
rect 9214 1680 9220 1692
rect 7116 1652 9220 1680
rect 9214 1640 9220 1652
rect 9272 1680 9278 1692
rect 10134 1680 10140 1692
rect 9272 1652 10140 1680
rect 9272 1640 9278 1652
rect 10134 1640 10140 1652
rect 10192 1640 10198 1692
rect 8386 1612 8392 1624
rect 6886 1584 8392 1612
rect 8386 1572 8392 1584
rect 8444 1572 8450 1624
rect 2866 1300 2872 1352
rect 2924 1340 2930 1352
rect 18414 1340 18420 1352
rect 2924 1312 18420 1340
rect 2924 1300 2930 1312
rect 18414 1300 18420 1312
rect 18472 1300 18478 1352
<< via1 >>
rect 1492 20748 1544 20800
rect 4712 20748 4764 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 2780 20544 2832 20596
rect 3148 20587 3200 20596
rect 3148 20553 3157 20587
rect 3157 20553 3191 20587
rect 3191 20553 3200 20587
rect 3148 20544 3200 20553
rect 4712 20587 4764 20596
rect 4712 20553 4721 20587
rect 4721 20553 4755 20587
rect 4755 20553 4764 20587
rect 4712 20544 4764 20553
rect 1492 20519 1544 20528
rect 1492 20485 1501 20519
rect 1501 20485 1535 20519
rect 1535 20485 1544 20519
rect 1492 20476 1544 20485
rect 2228 20451 2280 20460
rect 2228 20417 2237 20451
rect 2237 20417 2271 20451
rect 2271 20417 2280 20451
rect 2228 20408 2280 20417
rect 8208 20476 8260 20528
rect 3976 20451 4028 20460
rect 3976 20417 3985 20451
rect 3985 20417 4019 20451
rect 4019 20417 4028 20451
rect 3976 20408 4028 20417
rect 8668 20408 8720 20460
rect 4160 20340 4212 20392
rect 1860 20272 1912 20324
rect 2044 20315 2096 20324
rect 2044 20281 2053 20315
rect 2053 20281 2087 20315
rect 2087 20281 2096 20315
rect 2044 20272 2096 20281
rect 2320 20272 2372 20324
rect 4436 20247 4488 20256
rect 4436 20213 4445 20247
rect 4445 20213 4479 20247
rect 4479 20213 4488 20247
rect 4436 20204 4488 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2596 20043 2648 20052
rect 2596 20009 2605 20043
rect 2605 20009 2639 20043
rect 2639 20009 2648 20043
rect 2596 20000 2648 20009
rect 3976 20000 4028 20052
rect 4160 20000 4212 20052
rect 2228 19932 2280 19984
rect 2964 19864 3016 19916
rect 6552 19864 6604 19916
rect 3608 19796 3660 19848
rect 4436 19839 4488 19848
rect 4436 19805 4445 19839
rect 4445 19805 4479 19839
rect 4479 19805 4488 19839
rect 4436 19796 4488 19805
rect 4528 19796 4580 19848
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 2044 19703 2096 19712
rect 2044 19669 2053 19703
rect 2053 19669 2087 19703
rect 2087 19669 2096 19703
rect 2044 19660 2096 19669
rect 3884 19660 3936 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 1952 19456 2004 19508
rect 3608 19499 3660 19508
rect 3608 19465 3617 19499
rect 3617 19465 3651 19499
rect 3651 19465 3660 19499
rect 3608 19456 3660 19465
rect 3884 19499 3936 19508
rect 3884 19465 3893 19499
rect 3893 19465 3927 19499
rect 3927 19465 3936 19499
rect 3884 19456 3936 19465
rect 4528 19499 4580 19508
rect 4528 19465 4537 19499
rect 4537 19465 4571 19499
rect 4571 19465 4580 19499
rect 4528 19456 4580 19465
rect 2320 19320 2372 19372
rect 2688 19320 2740 19372
rect 3332 19252 3384 19304
rect 5908 19388 5960 19440
rect 9680 19320 9732 19372
rect 2688 19184 2740 19236
rect 8484 19184 8536 19236
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 2044 19116 2096 19168
rect 6000 19116 6052 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 8208 18912 8260 18964
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 2228 18708 2280 18760
rect 5632 18844 5684 18896
rect 3148 18776 3200 18828
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 1676 18572 1728 18624
rect 2596 18615 2648 18624
rect 2596 18581 2605 18615
rect 2605 18581 2639 18615
rect 2639 18581 2648 18615
rect 2596 18572 2648 18581
rect 10692 18751 10744 18760
rect 3148 18640 3200 18692
rect 10692 18717 10701 18751
rect 10701 18717 10735 18751
rect 10735 18717 10744 18751
rect 10692 18708 10744 18717
rect 3240 18572 3292 18624
rect 4712 18615 4764 18624
rect 4712 18581 4721 18615
rect 4721 18581 4755 18615
rect 4755 18581 4764 18615
rect 4712 18572 4764 18581
rect 5816 18615 5868 18624
rect 5816 18581 5825 18615
rect 5825 18581 5859 18615
rect 5859 18581 5868 18615
rect 5816 18572 5868 18581
rect 6920 18615 6972 18624
rect 6920 18581 6929 18615
rect 6929 18581 6963 18615
rect 6963 18581 6972 18615
rect 6920 18572 6972 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 2136 18368 2188 18420
rect 2596 18368 2648 18420
rect 9680 18411 9732 18420
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 3240 18300 3292 18352
rect 9680 18377 9689 18411
rect 9689 18377 9723 18411
rect 9723 18377 9732 18411
rect 9680 18368 9732 18377
rect 10692 18368 10744 18420
rect 3884 18275 3936 18284
rect 3884 18241 3893 18275
rect 3893 18241 3927 18275
rect 3927 18241 3936 18275
rect 3884 18232 3936 18241
rect 4528 18232 4580 18284
rect 5724 18232 5776 18284
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 6828 18207 6880 18216
rect 4712 18096 4764 18148
rect 6828 18173 6837 18207
rect 6837 18173 6871 18207
rect 6871 18173 6880 18207
rect 6828 18164 6880 18173
rect 11704 18275 11756 18284
rect 11704 18241 11713 18275
rect 11713 18241 11747 18275
rect 11747 18241 11756 18275
rect 11704 18232 11756 18241
rect 6644 18096 6696 18148
rect 8208 18164 8260 18216
rect 10140 18207 10192 18216
rect 10140 18173 10149 18207
rect 10149 18173 10183 18207
rect 10183 18173 10192 18207
rect 10140 18164 10192 18173
rect 11060 18164 11112 18216
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2964 18028 3016 18080
rect 3148 18071 3200 18080
rect 3148 18037 3157 18071
rect 3157 18037 3191 18071
rect 3191 18037 3200 18071
rect 3148 18028 3200 18037
rect 3332 18028 3384 18080
rect 4620 18028 4672 18080
rect 5356 18071 5408 18080
rect 5356 18037 5365 18071
rect 5365 18037 5399 18071
rect 5399 18037 5408 18071
rect 5356 18028 5408 18037
rect 7012 18028 7064 18080
rect 9496 18028 9548 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 6828 17824 6880 17876
rect 10140 17824 10192 17876
rect 3148 17756 3200 17808
rect 6920 17756 6972 17808
rect 5724 17688 5776 17740
rect 15752 17756 15804 17808
rect 1676 17663 1728 17672
rect 1676 17629 1685 17663
rect 1685 17629 1719 17663
rect 1719 17629 1728 17663
rect 1676 17620 1728 17629
rect 2412 17663 2464 17672
rect 2412 17629 2421 17663
rect 2421 17629 2455 17663
rect 2455 17629 2464 17663
rect 2412 17620 2464 17629
rect 2780 17620 2832 17672
rect 4528 17620 4580 17672
rect 6920 17620 6972 17672
rect 7288 17620 7340 17672
rect 7748 17620 7800 17672
rect 9404 17688 9456 17740
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 12900 17663 12952 17672
rect 12900 17629 12909 17663
rect 12909 17629 12943 17663
rect 12943 17629 12952 17663
rect 12900 17620 12952 17629
rect 13268 17620 13320 17672
rect 2320 17552 2372 17604
rect 3424 17552 3476 17604
rect 6736 17552 6788 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 1676 17484 1728 17536
rect 2872 17527 2924 17536
rect 2872 17493 2881 17527
rect 2881 17493 2915 17527
rect 2915 17493 2924 17527
rect 2872 17484 2924 17493
rect 3884 17484 3936 17536
rect 5816 17484 5868 17536
rect 9496 17552 9548 17604
rect 12532 17595 12584 17604
rect 12532 17561 12541 17595
rect 12541 17561 12575 17595
rect 12575 17561 12584 17595
rect 12532 17552 12584 17561
rect 7472 17484 7524 17536
rect 8576 17527 8628 17536
rect 8576 17493 8585 17527
rect 8585 17493 8619 17527
rect 8619 17493 8628 17527
rect 8576 17484 8628 17493
rect 9772 17484 9824 17536
rect 11796 17484 11848 17536
rect 11980 17527 12032 17536
rect 11980 17493 11989 17527
rect 11989 17493 12023 17527
rect 12023 17493 12032 17527
rect 11980 17484 12032 17493
rect 13544 17527 13596 17536
rect 13544 17493 13553 17527
rect 13553 17493 13587 17527
rect 13587 17493 13596 17527
rect 13544 17484 13596 17493
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 5724 17323 5776 17332
rect 5724 17289 5733 17323
rect 5733 17289 5767 17323
rect 5767 17289 5776 17323
rect 5724 17280 5776 17289
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 4252 17144 4304 17196
rect 4620 17187 4672 17196
rect 4620 17153 4654 17187
rect 4654 17153 4672 17187
rect 4620 17144 4672 17153
rect 6920 17212 6972 17264
rect 7932 17212 7984 17264
rect 7012 17144 7064 17196
rect 8300 17187 8352 17196
rect 8300 17153 8334 17187
rect 8334 17153 8352 17187
rect 11060 17212 11112 17264
rect 8300 17144 8352 17153
rect 9772 17144 9824 17196
rect 11796 17187 11848 17196
rect 11796 17153 11830 17187
rect 11830 17153 11848 17187
rect 11796 17144 11848 17153
rect 2964 17076 3016 17128
rect 4160 17076 4212 17128
rect 1492 17051 1544 17060
rect 1492 17017 1501 17051
rect 1501 17017 1535 17051
rect 1535 17017 1544 17051
rect 1492 17008 1544 17017
rect 1768 17008 1820 17060
rect 11152 17008 11204 17060
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 7748 16983 7800 16992
rect 7748 16949 7757 16983
rect 7757 16949 7791 16983
rect 7791 16949 7800 16983
rect 7748 16940 7800 16949
rect 12900 16983 12952 16992
rect 12900 16949 12909 16983
rect 12909 16949 12943 16983
rect 12943 16949 12952 16983
rect 12900 16940 12952 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 2780 16736 2832 16788
rect 2964 16779 3016 16788
rect 2964 16745 2973 16779
rect 2973 16745 3007 16779
rect 3007 16745 3016 16779
rect 2964 16736 3016 16745
rect 3884 16600 3936 16652
rect 6920 16736 6972 16788
rect 13268 16779 13320 16788
rect 6644 16711 6696 16720
rect 6644 16677 6653 16711
rect 6653 16677 6687 16711
rect 6687 16677 6696 16711
rect 6644 16668 6696 16677
rect 13268 16745 13277 16779
rect 13277 16745 13311 16779
rect 13311 16745 13320 16779
rect 13268 16736 13320 16745
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 2688 16532 2740 16584
rect 3148 16575 3200 16584
rect 3148 16541 3157 16575
rect 3157 16541 3191 16575
rect 3191 16541 3200 16575
rect 3148 16532 3200 16541
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 5356 16532 5408 16584
rect 7840 16600 7892 16652
rect 9404 16600 9456 16652
rect 8208 16575 8260 16584
rect 8208 16541 8217 16575
rect 8217 16541 8251 16575
rect 8251 16541 8260 16575
rect 8208 16532 8260 16541
rect 8300 16532 8352 16584
rect 2872 16464 2924 16516
rect 11060 16600 11112 16652
rect 11152 16532 11204 16584
rect 11980 16532 12032 16584
rect 13544 16532 13596 16584
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2044 16439 2096 16448
rect 2044 16405 2053 16439
rect 2053 16405 2087 16439
rect 2087 16405 2096 16439
rect 2044 16396 2096 16405
rect 3240 16396 3292 16448
rect 4252 16439 4304 16448
rect 4252 16405 4261 16439
rect 4261 16405 4295 16439
rect 4295 16405 4304 16439
rect 4252 16396 4304 16405
rect 5724 16396 5776 16448
rect 6552 16396 6604 16448
rect 9312 16439 9364 16448
rect 9312 16405 9321 16439
rect 9321 16405 9355 16439
rect 9355 16405 9364 16439
rect 9312 16396 9364 16405
rect 11152 16439 11204 16448
rect 11152 16405 11161 16439
rect 11161 16405 11195 16439
rect 11195 16405 11204 16439
rect 11152 16396 11204 16405
rect 11704 16396 11756 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 2596 16235 2648 16244
rect 2596 16201 2605 16235
rect 2605 16201 2639 16235
rect 2639 16201 2648 16235
rect 2596 16192 2648 16201
rect 4252 16192 4304 16244
rect 6000 16192 6052 16244
rect 7840 16235 7892 16244
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 4528 16124 4580 16176
rect 6644 16124 6696 16176
rect 9312 16192 9364 16244
rect 11152 16192 11204 16244
rect 1768 16056 1820 16108
rect 2136 16056 2188 16108
rect 2596 16056 2648 16108
rect 2872 16056 2924 16108
rect 9312 16056 9364 16108
rect 11152 16056 11204 16108
rect 7196 16031 7248 16040
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4344 15963 4396 15972
rect 4344 15929 4353 15963
rect 4353 15929 4387 15963
rect 4387 15929 4396 15963
rect 7196 15997 7205 16031
rect 7205 15997 7239 16031
rect 7239 15997 7248 16031
rect 7196 15988 7248 15997
rect 7288 16031 7340 16040
rect 7288 15997 7297 16031
rect 7297 15997 7331 16031
rect 7331 15997 7340 16031
rect 9220 16031 9272 16040
rect 7288 15988 7340 15997
rect 9220 15997 9229 16031
rect 9229 15997 9263 16031
rect 9263 15997 9272 16031
rect 9220 15988 9272 15997
rect 10416 16031 10468 16040
rect 10416 15997 10425 16031
rect 10425 15997 10459 16031
rect 10459 15997 10468 16031
rect 10416 15988 10468 15997
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 12900 15988 12952 16040
rect 4344 15920 4396 15929
rect 8024 15920 8076 15972
rect 3884 15852 3936 15904
rect 6552 15852 6604 15904
rect 11152 15895 11204 15904
rect 11152 15861 11161 15895
rect 11161 15861 11195 15895
rect 11195 15861 11204 15895
rect 11152 15852 11204 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 2412 15648 2464 15700
rect 2780 15648 2832 15700
rect 7288 15648 7340 15700
rect 9312 15648 9364 15700
rect 1952 15512 2004 15564
rect 8024 15580 8076 15632
rect 11704 15648 11756 15700
rect 3332 15555 3384 15564
rect 3332 15521 3341 15555
rect 3341 15521 3375 15555
rect 3375 15521 3384 15555
rect 3332 15512 3384 15521
rect 4896 15555 4948 15564
rect 4896 15521 4905 15555
rect 4905 15521 4939 15555
rect 4939 15521 4948 15555
rect 4896 15512 4948 15521
rect 5908 15555 5960 15564
rect 5908 15521 5917 15555
rect 5917 15521 5951 15555
rect 5951 15521 5960 15555
rect 5908 15512 5960 15521
rect 7932 15555 7984 15564
rect 7932 15521 7941 15555
rect 7941 15521 7975 15555
rect 7975 15521 7984 15555
rect 7932 15512 7984 15521
rect 1860 15444 1912 15496
rect 8576 15444 8628 15496
rect 9220 15444 9272 15496
rect 10968 15444 11020 15496
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 1676 15308 1728 15360
rect 4160 15308 4212 15360
rect 4712 15351 4764 15360
rect 4712 15317 4721 15351
rect 4721 15317 4755 15351
rect 4755 15317 4764 15351
rect 5724 15351 5776 15360
rect 4712 15308 4764 15317
rect 5724 15317 5733 15351
rect 5733 15317 5767 15351
rect 5767 15317 5776 15351
rect 5724 15308 5776 15317
rect 10784 15376 10836 15428
rect 12440 15308 12492 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 2320 15147 2372 15156
rect 2320 15113 2329 15147
rect 2329 15113 2363 15147
rect 2363 15113 2372 15147
rect 2320 15104 2372 15113
rect 2872 15104 2924 15156
rect 1676 15011 1728 15020
rect 1676 14977 1685 15011
rect 1685 14977 1719 15011
rect 1719 14977 1728 15011
rect 1676 14968 1728 14977
rect 3332 14968 3384 15020
rect 7196 15147 7248 15156
rect 7196 15113 7205 15147
rect 7205 15113 7239 15147
rect 7239 15113 7248 15147
rect 7196 15104 7248 15113
rect 5908 14968 5960 15020
rect 6920 15036 6972 15088
rect 7932 15036 7984 15088
rect 8668 15104 8720 15156
rect 10416 15104 10468 15156
rect 11152 15104 11204 15156
rect 6460 14968 6512 15020
rect 4252 14900 4304 14952
rect 6552 14875 6604 14884
rect 6552 14841 6561 14875
rect 6561 14841 6595 14875
rect 6595 14841 6604 14875
rect 6552 14832 6604 14841
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1768 14764 1820 14816
rect 2320 14764 2372 14816
rect 5080 14764 5132 14816
rect 11796 15036 11848 15088
rect 10876 15011 10928 15020
rect 10876 14977 10894 15011
rect 10894 14977 10928 15011
rect 10876 14968 10928 14977
rect 11060 14968 11112 15020
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 7748 14943 7800 14952
rect 7748 14909 7757 14943
rect 7757 14909 7791 14943
rect 7791 14909 7800 14943
rect 9220 14943 9272 14952
rect 7748 14900 7800 14909
rect 9220 14909 9229 14943
rect 9229 14909 9263 14943
rect 9263 14909 9272 14943
rect 9220 14900 9272 14909
rect 7288 14764 7340 14816
rect 10784 14764 10836 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 2412 14356 2464 14408
rect 4988 14560 5040 14612
rect 5908 14560 5960 14612
rect 6000 14560 6052 14612
rect 10876 14560 10928 14612
rect 8760 14492 8812 14544
rect 4160 14424 4212 14476
rect 3884 14356 3936 14408
rect 5540 14424 5592 14476
rect 6920 14467 6972 14476
rect 6920 14433 6929 14467
rect 6929 14433 6963 14467
rect 6963 14433 6972 14467
rect 6920 14424 6972 14433
rect 7012 14356 7064 14408
rect 7472 14356 7524 14408
rect 5724 14288 5776 14340
rect 9312 14288 9364 14340
rect 9588 14288 9640 14340
rect 11060 14356 11112 14408
rect 11704 14424 11756 14476
rect 19984 14424 20036 14476
rect 12256 14288 12308 14340
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 6920 14220 6972 14272
rect 8024 14220 8076 14272
rect 10324 14220 10376 14272
rect 11244 14220 11296 14272
rect 18144 14220 18196 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 2412 14059 2464 14068
rect 2412 14025 2421 14059
rect 2421 14025 2455 14059
rect 2455 14025 2464 14059
rect 2412 14016 2464 14025
rect 4896 14016 4948 14068
rect 8668 14016 8720 14068
rect 8760 14059 8812 14068
rect 8760 14025 8769 14059
rect 8769 14025 8803 14059
rect 8803 14025 8812 14059
rect 8760 14016 8812 14025
rect 9220 14016 9272 14068
rect 2320 13948 2372 14000
rect 5908 13948 5960 14000
rect 2136 13923 2188 13932
rect 2136 13889 2145 13923
rect 2145 13889 2179 13923
rect 2179 13889 2188 13923
rect 2136 13880 2188 13889
rect 2964 13923 3016 13932
rect 1400 13812 1452 13864
rect 2964 13889 2973 13923
rect 2973 13889 3007 13923
rect 3007 13889 3016 13923
rect 2964 13880 3016 13889
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 4160 13923 4212 13932
rect 4160 13889 4194 13923
rect 4194 13889 4212 13923
rect 4160 13880 4212 13889
rect 4436 13880 4488 13932
rect 6000 13880 6052 13932
rect 2872 13812 2924 13864
rect 8576 13948 8628 14000
rect 8024 13923 8076 13932
rect 8024 13889 8042 13923
rect 8042 13889 8076 13923
rect 8024 13880 8076 13889
rect 9864 13880 9916 13932
rect 9220 13744 9272 13796
rect 9588 13812 9640 13864
rect 10692 13880 10744 13932
rect 10324 13855 10376 13864
rect 10324 13821 10333 13855
rect 10333 13821 10367 13855
rect 10367 13821 10376 13855
rect 10324 13812 10376 13821
rect 11980 13812 12032 13864
rect 19064 13812 19116 13864
rect 9956 13744 10008 13796
rect 3240 13676 3292 13728
rect 7012 13676 7064 13728
rect 7380 13676 7432 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 4160 13472 4212 13524
rect 5540 13515 5592 13524
rect 5540 13481 5549 13515
rect 5549 13481 5583 13515
rect 5583 13481 5592 13515
rect 5540 13472 5592 13481
rect 9956 13515 10008 13524
rect 9956 13481 9965 13515
rect 9965 13481 9999 13515
rect 9999 13481 10008 13515
rect 12256 13515 12308 13524
rect 9956 13472 10008 13481
rect 3792 13404 3844 13456
rect 4436 13404 4488 13456
rect 5264 13404 5316 13456
rect 10232 13404 10284 13456
rect 4804 13379 4856 13388
rect 4804 13345 4813 13379
rect 4813 13345 4847 13379
rect 4847 13345 4856 13379
rect 4804 13336 4856 13345
rect 5908 13336 5960 13388
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 5448 13268 5500 13320
rect 7288 13311 7340 13320
rect 7288 13277 7297 13311
rect 7297 13277 7331 13311
rect 7331 13277 7340 13311
rect 7288 13268 7340 13277
rect 8024 13336 8076 13388
rect 8576 13336 8628 13388
rect 8760 13268 8812 13320
rect 9128 13268 9180 13320
rect 9680 13268 9732 13320
rect 7012 13243 7064 13252
rect 7012 13209 7021 13243
rect 7021 13209 7055 13243
rect 7055 13209 7064 13243
rect 7012 13200 7064 13209
rect 2228 13175 2280 13184
rect 2228 13141 2237 13175
rect 2237 13141 2271 13175
rect 2271 13141 2280 13175
rect 2228 13132 2280 13141
rect 4252 13132 4304 13184
rect 4528 13175 4580 13184
rect 4528 13141 4537 13175
rect 4537 13141 4571 13175
rect 4571 13141 4580 13175
rect 4528 13132 4580 13141
rect 5172 13132 5224 13184
rect 7564 13132 7616 13184
rect 8208 13175 8260 13184
rect 8208 13141 8217 13175
rect 8217 13141 8251 13175
rect 8251 13141 8260 13175
rect 9680 13175 9732 13184
rect 8208 13132 8260 13141
rect 9680 13141 9689 13175
rect 9689 13141 9723 13175
rect 9723 13141 9732 13175
rect 9680 13132 9732 13141
rect 11244 13268 11296 13320
rect 12256 13481 12265 13515
rect 12265 13481 12299 13515
rect 12299 13481 12308 13515
rect 12256 13472 12308 13481
rect 12072 13200 12124 13252
rect 15292 13132 15344 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 1492 12971 1544 12980
rect 1492 12937 1501 12971
rect 1501 12937 1535 12971
rect 1535 12937 1544 12971
rect 1492 12928 1544 12937
rect 4344 12928 4396 12980
rect 4528 12928 4580 12980
rect 5816 12928 5868 12980
rect 9864 12971 9916 12980
rect 4620 12860 4672 12912
rect 5908 12860 5960 12912
rect 7012 12860 7064 12912
rect 3148 12724 3200 12776
rect 3884 12792 3936 12844
rect 4160 12792 4212 12844
rect 9864 12937 9873 12971
rect 9873 12937 9907 12971
rect 9907 12937 9916 12971
rect 9864 12928 9916 12937
rect 10232 12903 10284 12912
rect 10232 12869 10241 12903
rect 10241 12869 10275 12903
rect 10275 12869 10284 12903
rect 10232 12860 10284 12869
rect 18880 12860 18932 12912
rect 3976 12724 4028 12776
rect 4068 12656 4120 12708
rect 5448 12699 5500 12708
rect 5448 12665 5457 12699
rect 5457 12665 5491 12699
rect 5491 12665 5500 12699
rect 5448 12656 5500 12665
rect 7748 12724 7800 12776
rect 10416 12767 10468 12776
rect 8024 12656 8076 12708
rect 4436 12588 4488 12640
rect 7472 12631 7524 12640
rect 7472 12597 7481 12631
rect 7481 12597 7515 12631
rect 7515 12597 7524 12631
rect 7472 12588 7524 12597
rect 9220 12588 9272 12640
rect 10416 12733 10425 12767
rect 10425 12733 10459 12767
rect 10459 12733 10468 12767
rect 10416 12724 10468 12733
rect 11520 12631 11572 12640
rect 11520 12597 11529 12631
rect 11529 12597 11563 12631
rect 11563 12597 11572 12631
rect 11520 12588 11572 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1860 12427 1912 12436
rect 1860 12393 1869 12427
rect 1869 12393 1903 12427
rect 1903 12393 1912 12427
rect 1860 12384 1912 12393
rect 2044 12384 2096 12436
rect 2872 12384 2924 12436
rect 4160 12384 4212 12436
rect 4804 12427 4856 12436
rect 4804 12393 4813 12427
rect 4813 12393 4847 12427
rect 4847 12393 4856 12427
rect 4804 12384 4856 12393
rect 3056 12316 3108 12368
rect 10416 12384 10468 12436
rect 12072 12427 12124 12436
rect 9036 12316 9088 12368
rect 9220 12316 9272 12368
rect 2780 12291 2832 12300
rect 2780 12257 2789 12291
rect 2789 12257 2823 12291
rect 2823 12257 2832 12291
rect 2780 12248 2832 12257
rect 7748 12248 7800 12300
rect 9588 12248 9640 12300
rect 1860 12180 1912 12232
rect 3884 12180 3936 12232
rect 4804 12180 4856 12232
rect 5540 12180 5592 12232
rect 6644 12223 6696 12232
rect 6644 12189 6653 12223
rect 6653 12189 6687 12223
rect 6687 12189 6696 12223
rect 6644 12180 6696 12189
rect 6920 12223 6972 12232
rect 6920 12189 6954 12223
rect 6954 12189 6972 12223
rect 6920 12180 6972 12189
rect 7840 12180 7892 12232
rect 10416 12180 10468 12232
rect 11060 12180 11112 12232
rect 12072 12393 12081 12427
rect 12081 12393 12115 12427
rect 12115 12393 12124 12427
rect 12072 12384 12124 12393
rect 19708 12223 19760 12232
rect 19708 12189 19717 12223
rect 19717 12189 19751 12223
rect 19751 12189 19760 12223
rect 19708 12180 19760 12189
rect 2320 12112 2372 12164
rect 5724 12112 5776 12164
rect 5908 12155 5960 12164
rect 5908 12121 5926 12155
rect 5926 12121 5960 12155
rect 5908 12112 5960 12121
rect 7104 12112 7156 12164
rect 8668 12112 8720 12164
rect 2504 12087 2556 12096
rect 2504 12053 2513 12087
rect 2513 12053 2547 12087
rect 2547 12053 2556 12087
rect 2504 12044 2556 12053
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 4068 12044 4120 12096
rect 6000 12044 6052 12096
rect 6920 12044 6972 12096
rect 7748 12044 7800 12096
rect 8024 12087 8076 12096
rect 8024 12053 8033 12087
rect 8033 12053 8067 12087
rect 8067 12053 8076 12087
rect 8024 12044 8076 12053
rect 8576 12044 8628 12096
rect 9312 12044 9364 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 12164 12112 12216 12164
rect 10232 12044 10284 12096
rect 12992 12044 13044 12096
rect 13452 12044 13504 12096
rect 20536 12044 20588 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 1676 11883 1728 11892
rect 1676 11849 1685 11883
rect 1685 11849 1719 11883
rect 1719 11849 1728 11883
rect 1676 11840 1728 11849
rect 2504 11840 2556 11892
rect 1584 11704 1636 11756
rect 2872 11704 2924 11756
rect 3976 11772 4028 11824
rect 4252 11840 4304 11892
rect 4620 11840 4672 11892
rect 4804 11883 4856 11892
rect 4804 11849 4813 11883
rect 4813 11849 4847 11883
rect 4847 11849 4856 11883
rect 4804 11840 4856 11849
rect 4528 11772 4580 11824
rect 3240 11747 3292 11756
rect 3240 11713 3274 11747
rect 3274 11713 3292 11747
rect 3240 11704 3292 11713
rect 4068 11704 4120 11756
rect 5264 11704 5316 11756
rect 5724 11840 5776 11892
rect 7472 11840 7524 11892
rect 12164 11883 12216 11892
rect 6000 11772 6052 11824
rect 6644 11772 6696 11824
rect 6920 11704 6972 11756
rect 7564 11704 7616 11756
rect 1952 11636 2004 11688
rect 2044 11500 2096 11552
rect 5356 11636 5408 11688
rect 7380 11679 7432 11688
rect 4712 11568 4764 11620
rect 5448 11568 5500 11620
rect 7380 11645 7389 11679
rect 7389 11645 7423 11679
rect 7423 11645 7432 11679
rect 7380 11636 7432 11645
rect 9680 11815 9732 11824
rect 9680 11781 9714 11815
rect 9714 11781 9732 11815
rect 9680 11772 9732 11781
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 12440 11883 12492 11892
rect 12440 11849 12449 11883
rect 12449 11849 12483 11883
rect 12483 11849 12492 11883
rect 12440 11840 12492 11849
rect 6644 11500 6696 11552
rect 9312 11636 9364 11688
rect 9036 11568 9088 11620
rect 10600 11704 10652 11756
rect 12624 11747 12676 11756
rect 12624 11713 12633 11747
rect 12633 11713 12667 11747
rect 12667 11713 12676 11747
rect 12624 11704 12676 11713
rect 19248 11747 19300 11756
rect 19248 11713 19257 11747
rect 19257 11713 19291 11747
rect 19291 11713 19300 11747
rect 19248 11704 19300 11713
rect 9128 11543 9180 11552
rect 9128 11509 9137 11543
rect 9137 11509 9171 11543
rect 9171 11509 9180 11543
rect 9128 11500 9180 11509
rect 10784 11543 10836 11552
rect 10784 11509 10793 11543
rect 10793 11509 10827 11543
rect 10827 11509 10836 11543
rect 10784 11500 10836 11509
rect 11060 11543 11112 11552
rect 11060 11509 11069 11543
rect 11069 11509 11103 11543
rect 11103 11509 11112 11543
rect 11060 11500 11112 11509
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 14280 11500 14332 11552
rect 20168 11500 20220 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1584 11339 1636 11348
rect 1584 11305 1593 11339
rect 1593 11305 1627 11339
rect 1627 11305 1636 11339
rect 1584 11296 1636 11305
rect 2780 11296 2832 11348
rect 3424 11296 3476 11348
rect 7196 11296 7248 11348
rect 8484 11296 8536 11348
rect 10600 11296 10652 11348
rect 8668 11228 8720 11280
rect 9036 11228 9088 11280
rect 15844 11228 15896 11280
rect 19616 11228 19668 11280
rect 2872 11160 2924 11212
rect 8024 11160 8076 11212
rect 1768 11092 1820 11144
rect 1952 11092 2004 11144
rect 3056 11092 3108 11144
rect 3240 11092 3292 11144
rect 4068 11092 4120 11144
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 4712 11092 4764 11144
rect 6644 11092 6696 11144
rect 3976 11024 4028 11076
rect 4436 11024 4488 11076
rect 3424 10956 3476 11008
rect 6460 11024 6512 11076
rect 6828 11092 6880 11144
rect 8852 11092 8904 11144
rect 9496 11092 9548 11144
rect 10784 11160 10836 11212
rect 14832 11203 14884 11212
rect 10416 11092 10468 11144
rect 12164 11135 12216 11144
rect 8208 11024 8260 11076
rect 6000 10999 6052 11008
rect 6000 10965 6009 10999
rect 6009 10965 6043 10999
rect 6043 10965 6052 10999
rect 6000 10956 6052 10965
rect 6552 10999 6604 11008
rect 6552 10965 6561 10999
rect 6561 10965 6595 10999
rect 6595 10965 6604 10999
rect 6552 10956 6604 10965
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 9404 11024 9456 11076
rect 12164 11101 12173 11135
rect 12173 11101 12207 11135
rect 12207 11101 12216 11135
rect 12164 11092 12216 11101
rect 12256 11092 12308 11144
rect 14832 11169 14841 11203
rect 14841 11169 14875 11203
rect 14875 11169 14884 11203
rect 14832 11160 14884 11169
rect 15200 11092 15252 11144
rect 15292 11092 15344 11144
rect 12072 11024 12124 11076
rect 13728 11024 13780 11076
rect 14464 11067 14516 11076
rect 14464 11033 14473 11067
rect 14473 11033 14507 11067
rect 14507 11033 14516 11067
rect 14464 11024 14516 11033
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 3056 10795 3108 10804
rect 3056 10761 3065 10795
rect 3065 10761 3099 10795
rect 3099 10761 3108 10795
rect 3056 10752 3108 10761
rect 3148 10752 3200 10804
rect 4160 10752 4212 10804
rect 4712 10752 4764 10804
rect 5632 10752 5684 10804
rect 7104 10795 7156 10804
rect 7104 10761 7113 10795
rect 7113 10761 7147 10795
rect 7147 10761 7156 10795
rect 7104 10752 7156 10761
rect 8208 10795 8260 10804
rect 8208 10761 8217 10795
rect 8217 10761 8251 10795
rect 8251 10761 8260 10795
rect 8208 10752 8260 10761
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 13820 10752 13872 10804
rect 1768 10684 1820 10736
rect 2228 10616 2280 10668
rect 4620 10684 4672 10736
rect 4804 10684 4856 10736
rect 6644 10684 6696 10736
rect 4344 10659 4396 10668
rect 4344 10625 4378 10659
rect 4378 10625 4396 10659
rect 4344 10616 4396 10625
rect 6736 10616 6788 10668
rect 7748 10659 7800 10668
rect 7748 10625 7757 10659
rect 7757 10625 7791 10659
rect 7791 10625 7800 10659
rect 7748 10616 7800 10625
rect 9680 10616 9732 10668
rect 5080 10548 5132 10600
rect 7196 10591 7248 10600
rect 7196 10557 7205 10591
rect 7205 10557 7239 10591
rect 7239 10557 7248 10591
rect 7196 10548 7248 10557
rect 8392 10548 8444 10600
rect 8668 10591 8720 10600
rect 8668 10557 8677 10591
rect 8677 10557 8711 10591
rect 8711 10557 8720 10591
rect 8668 10548 8720 10557
rect 6552 10480 6604 10532
rect 8484 10480 8536 10532
rect 9128 10548 9180 10600
rect 9588 10480 9640 10532
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 17960 10684 18012 10736
rect 12808 10616 12860 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 14372 10616 14424 10625
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 16120 10548 16172 10600
rect 14648 10480 14700 10532
rect 15752 10523 15804 10532
rect 15752 10489 15761 10523
rect 15761 10489 15795 10523
rect 15795 10489 15804 10523
rect 15752 10480 15804 10489
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 8300 10412 8352 10464
rect 11336 10412 11388 10464
rect 11796 10412 11848 10464
rect 13176 10412 13228 10464
rect 15384 10455 15436 10464
rect 15384 10421 15393 10455
rect 15393 10421 15427 10455
rect 15427 10421 15436 10455
rect 15384 10412 15436 10421
rect 20076 10412 20128 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 2596 10251 2648 10260
rect 2596 10217 2605 10251
rect 2605 10217 2639 10251
rect 2639 10217 2648 10251
rect 2596 10208 2648 10217
rect 3332 10208 3384 10260
rect 4988 10208 5040 10260
rect 5172 10251 5224 10260
rect 5172 10217 5181 10251
rect 5181 10217 5215 10251
rect 5215 10217 5224 10251
rect 5172 10208 5224 10217
rect 1860 10072 1912 10124
rect 2688 10140 2740 10192
rect 3792 10140 3844 10192
rect 4068 10140 4120 10192
rect 8944 10140 8996 10192
rect 9588 10140 9640 10192
rect 11244 10208 11296 10260
rect 15200 10208 15252 10260
rect 3056 10072 3108 10124
rect 4252 10115 4304 10124
rect 4252 10081 4261 10115
rect 4261 10081 4295 10115
rect 4295 10081 4304 10115
rect 4252 10072 4304 10081
rect 2872 9936 2924 9988
rect 2228 9868 2280 9920
rect 2504 9868 2556 9920
rect 3056 9911 3108 9920
rect 3056 9877 3065 9911
rect 3065 9877 3099 9911
rect 3099 9877 3108 9911
rect 3056 9868 3108 9877
rect 3332 9868 3384 9920
rect 4068 10004 4120 10056
rect 4528 10004 4580 10056
rect 5632 10072 5684 10124
rect 6000 10072 6052 10124
rect 6828 10115 6880 10124
rect 6828 10081 6837 10115
rect 6837 10081 6871 10115
rect 6871 10081 6880 10115
rect 6828 10072 6880 10081
rect 4160 9936 4212 9988
rect 6092 10004 6144 10056
rect 8300 10004 8352 10056
rect 8576 10047 8628 10056
rect 8576 10013 8585 10047
rect 8585 10013 8619 10047
rect 8619 10013 8628 10047
rect 8576 10004 8628 10013
rect 8852 10004 8904 10056
rect 8760 9936 8812 9988
rect 4252 9868 4304 9920
rect 4620 9868 4672 9920
rect 4896 9911 4948 9920
rect 4896 9877 4905 9911
rect 4905 9877 4939 9911
rect 4939 9877 4948 9911
rect 4896 9868 4948 9877
rect 5172 9868 5224 9920
rect 7840 9868 7892 9920
rect 8392 9868 8444 9920
rect 8576 9868 8628 9920
rect 9220 9868 9272 9920
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 11796 10140 11848 10192
rect 13636 10004 13688 10056
rect 10048 9936 10100 9988
rect 11336 9936 11388 9988
rect 13820 9936 13872 9988
rect 14556 9979 14608 9988
rect 14556 9945 14565 9979
rect 14565 9945 14599 9979
rect 14599 9945 14608 9979
rect 14556 9936 14608 9945
rect 15200 9936 15252 9988
rect 9864 9868 9916 9920
rect 11980 9868 12032 9920
rect 15108 9868 15160 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 2320 9528 2372 9580
rect 3148 9528 3200 9580
rect 3332 9528 3384 9580
rect 4896 9664 4948 9716
rect 5172 9664 5224 9716
rect 5908 9596 5960 9648
rect 7564 9639 7616 9648
rect 7564 9605 7573 9639
rect 7573 9605 7607 9639
rect 7607 9605 7616 9639
rect 7564 9596 7616 9605
rect 8668 9664 8720 9716
rect 8760 9664 8812 9716
rect 15108 9664 15160 9716
rect 9680 9596 9732 9648
rect 11244 9596 11296 9648
rect 13820 9639 13872 9648
rect 4344 9528 4396 9580
rect 5080 9528 5132 9580
rect 5632 9528 5684 9580
rect 6184 9528 6236 9580
rect 8668 9528 8720 9580
rect 3700 9503 3752 9512
rect 3700 9469 3709 9503
rect 3709 9469 3743 9503
rect 3743 9469 3752 9503
rect 3700 9460 3752 9469
rect 4712 9460 4764 9512
rect 7380 9460 7432 9512
rect 1492 9435 1544 9444
rect 1492 9401 1501 9435
rect 1501 9401 1535 9435
rect 1535 9401 1544 9435
rect 1492 9392 1544 9401
rect 3516 9392 3568 9444
rect 3792 9392 3844 9444
rect 3148 9367 3200 9376
rect 3148 9333 3157 9367
rect 3157 9333 3191 9367
rect 3191 9333 3200 9367
rect 3148 9324 3200 9333
rect 4620 9324 4672 9376
rect 7564 9392 7616 9444
rect 8024 9460 8076 9512
rect 5908 9324 5960 9376
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 8116 9392 8168 9444
rect 8760 9392 8812 9444
rect 8944 9503 8996 9512
rect 8944 9469 8953 9503
rect 8953 9469 8987 9503
rect 8987 9469 8996 9503
rect 8944 9460 8996 9469
rect 9312 9392 9364 9444
rect 9588 9528 9640 9580
rect 11152 9528 11204 9580
rect 10048 9503 10100 9512
rect 10048 9469 10057 9503
rect 10057 9469 10091 9503
rect 10091 9469 10100 9503
rect 10048 9460 10100 9469
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 10784 9460 10836 9512
rect 12900 9528 12952 9580
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14280 9528 14332 9580
rect 15752 9571 15804 9580
rect 15752 9537 15761 9571
rect 15761 9537 15795 9571
rect 15795 9537 15804 9571
rect 15752 9528 15804 9537
rect 11060 9324 11112 9376
rect 11796 9324 11848 9376
rect 11888 9324 11940 9376
rect 12624 9324 12676 9376
rect 12900 9367 12952 9376
rect 12900 9333 12909 9367
rect 12909 9333 12943 9367
rect 12943 9333 12952 9367
rect 12900 9324 12952 9333
rect 14924 9460 14976 9512
rect 17132 9392 17184 9444
rect 15476 9324 15528 9376
rect 15660 9324 15712 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1584 9163 1636 9172
rect 1584 9129 1593 9163
rect 1593 9129 1627 9163
rect 1627 9129 1636 9163
rect 1584 9120 1636 9129
rect 1952 9163 2004 9172
rect 1952 9129 1961 9163
rect 1961 9129 1995 9163
rect 1995 9129 2004 9163
rect 1952 9120 2004 9129
rect 4068 9120 4120 9172
rect 1308 9052 1360 9104
rect 5448 9052 5500 9104
rect 6736 9052 6788 9104
rect 9312 9120 9364 9172
rect 12808 9120 12860 9172
rect 10048 9052 10100 9104
rect 1492 8984 1544 9036
rect 2688 8984 2740 9036
rect 1216 8916 1268 8968
rect 3148 8916 3200 8968
rect 4804 8984 4856 9036
rect 6276 9027 6328 9036
rect 6276 8993 6285 9027
rect 6285 8993 6319 9027
rect 6319 8993 6328 9027
rect 6276 8984 6328 8993
rect 8668 8984 8720 9036
rect 9588 8984 9640 9036
rect 10600 9052 10652 9104
rect 14280 9052 14332 9104
rect 15568 9052 15620 9104
rect 12900 8984 12952 9036
rect 16304 8984 16356 9036
rect 5448 8916 5500 8968
rect 2780 8848 2832 8900
rect 3792 8848 3844 8900
rect 4988 8848 5040 8900
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 3240 8780 3292 8832
rect 3976 8780 4028 8832
rect 4436 8823 4488 8832
rect 4436 8789 4445 8823
rect 4445 8789 4479 8823
rect 4479 8789 4488 8823
rect 4436 8780 4488 8789
rect 6000 8780 6052 8832
rect 6920 8780 6972 8832
rect 8116 8848 8168 8900
rect 8392 8916 8444 8968
rect 10048 8916 10100 8968
rect 8576 8848 8628 8900
rect 10140 8891 10192 8900
rect 10140 8857 10149 8891
rect 10149 8857 10183 8891
rect 10183 8857 10192 8891
rect 10140 8848 10192 8857
rect 10416 8848 10468 8900
rect 12348 8848 12400 8900
rect 15016 8848 15068 8900
rect 19892 9052 19944 9104
rect 8944 8780 8996 8832
rect 9128 8823 9180 8832
rect 9128 8789 9137 8823
rect 9137 8789 9171 8823
rect 9171 8789 9180 8823
rect 9128 8780 9180 8789
rect 10232 8780 10284 8832
rect 11060 8780 11112 8832
rect 11796 8780 11848 8832
rect 12624 8780 12676 8832
rect 18236 8780 18288 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 2320 8619 2372 8628
rect 2320 8585 2329 8619
rect 2329 8585 2363 8619
rect 2363 8585 2372 8619
rect 2320 8576 2372 8585
rect 2596 8576 2648 8628
rect 4804 8576 4856 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8944 8576 8996 8628
rect 9496 8576 9548 8628
rect 12716 8576 12768 8628
rect 15016 8619 15068 8628
rect 15016 8585 15025 8619
rect 15025 8585 15059 8619
rect 15059 8585 15068 8619
rect 15016 8576 15068 8585
rect 2780 8508 2832 8560
rect 2596 8440 2648 8492
rect 3148 8440 3200 8492
rect 3792 8440 3844 8492
rect 4896 8508 4948 8560
rect 5540 8508 5592 8560
rect 7380 8508 7432 8560
rect 4160 8415 4212 8424
rect 4160 8381 4169 8415
rect 4169 8381 4203 8415
rect 4203 8381 4212 8415
rect 4160 8372 4212 8381
rect 6920 8440 6972 8492
rect 8024 8508 8076 8560
rect 9220 8508 9272 8560
rect 8208 8440 8260 8492
rect 8484 8440 8536 8492
rect 8392 8372 8444 8424
rect 5448 8304 5500 8356
rect 12164 8508 12216 8560
rect 16948 8508 17000 8560
rect 17960 8576 18012 8628
rect 20720 8576 20772 8628
rect 18604 8508 18656 8560
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 11060 8440 11112 8492
rect 9496 8415 9548 8424
rect 9496 8381 9505 8415
rect 9505 8381 9539 8415
rect 9539 8381 9548 8415
rect 9496 8372 9548 8381
rect 9956 8372 10008 8424
rect 11244 8372 11296 8424
rect 11796 8415 11848 8424
rect 11796 8381 11805 8415
rect 11805 8381 11839 8415
rect 11839 8381 11848 8415
rect 11796 8372 11848 8381
rect 15660 8440 15712 8492
rect 15752 8483 15804 8492
rect 15752 8449 15761 8483
rect 15761 8449 15795 8483
rect 15795 8449 15804 8483
rect 15752 8440 15804 8449
rect 15936 8440 15988 8492
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 13268 8372 13320 8424
rect 13636 8415 13688 8424
rect 13636 8381 13645 8415
rect 13645 8381 13679 8415
rect 13679 8381 13688 8415
rect 13636 8372 13688 8381
rect 14924 8372 14976 8424
rect 16212 8415 16264 8424
rect 16212 8381 16221 8415
rect 16221 8381 16255 8415
rect 16255 8381 16264 8415
rect 16212 8372 16264 8381
rect 10968 8347 11020 8356
rect 5724 8236 5776 8288
rect 10968 8313 10977 8347
rect 10977 8313 11011 8347
rect 11011 8313 11020 8347
rect 10968 8304 11020 8313
rect 12256 8279 12308 8288
rect 12256 8245 12265 8279
rect 12265 8245 12299 8279
rect 12299 8245 12308 8279
rect 12256 8236 12308 8245
rect 13360 8279 13412 8288
rect 13360 8245 13369 8279
rect 13369 8245 13403 8279
rect 13403 8245 13412 8279
rect 13360 8236 13412 8245
rect 13544 8236 13596 8288
rect 17960 8347 18012 8356
rect 17960 8313 17969 8347
rect 17969 8313 18003 8347
rect 18003 8313 18012 8347
rect 17960 8304 18012 8313
rect 18328 8347 18380 8356
rect 18328 8313 18337 8347
rect 18337 8313 18371 8347
rect 18371 8313 18380 8347
rect 18328 8304 18380 8313
rect 18788 8347 18840 8356
rect 18788 8313 18797 8347
rect 18797 8313 18831 8347
rect 18831 8313 18840 8347
rect 18788 8304 18840 8313
rect 15568 8236 15620 8288
rect 20260 8236 20312 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2412 8075 2464 8084
rect 2412 8041 2421 8075
rect 2421 8041 2455 8075
rect 2455 8041 2464 8075
rect 2412 8032 2464 8041
rect 3056 8032 3108 8084
rect 4988 8075 5040 8084
rect 4988 8041 4997 8075
rect 4997 8041 5031 8075
rect 5031 8041 5040 8075
rect 4988 8032 5040 8041
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6552 8032 6604 8084
rect 3424 7964 3476 8016
rect 6736 7964 6788 8016
rect 2320 7896 2372 7948
rect 3148 7896 3200 7948
rect 6920 7896 6972 7948
rect 2504 7828 2556 7880
rect 2596 7760 2648 7812
rect 4068 7828 4120 7880
rect 6644 7828 6696 7880
rect 7012 7871 7064 7880
rect 7012 7837 7021 7871
rect 7021 7837 7055 7871
rect 7055 7837 7064 7871
rect 7012 7828 7064 7837
rect 7748 8032 7800 8084
rect 15568 8032 15620 8084
rect 15660 8032 15712 8084
rect 16396 8075 16448 8084
rect 16396 8041 16405 8075
rect 16405 8041 16439 8075
rect 16439 8041 16448 8075
rect 16396 8032 16448 8041
rect 14280 7964 14332 8016
rect 7472 7939 7524 7948
rect 7472 7905 7481 7939
rect 7481 7905 7515 7939
rect 7515 7905 7524 7939
rect 7472 7896 7524 7905
rect 11060 7896 11112 7948
rect 15016 7896 15068 7948
rect 15108 7896 15160 7948
rect 8392 7828 8444 7880
rect 8944 7871 8996 7880
rect 8944 7837 8953 7871
rect 8953 7837 8987 7871
rect 8987 7837 8996 7871
rect 8944 7828 8996 7837
rect 10600 7828 10652 7880
rect 11888 7828 11940 7880
rect 4068 7692 4120 7744
rect 4620 7735 4672 7744
rect 4620 7701 4629 7735
rect 4629 7701 4663 7735
rect 4663 7701 4672 7735
rect 4620 7692 4672 7701
rect 5448 7692 5500 7744
rect 7104 7692 7156 7744
rect 7564 7735 7616 7744
rect 7564 7701 7573 7735
rect 7573 7701 7607 7735
rect 7607 7701 7616 7735
rect 7564 7692 7616 7701
rect 8392 7692 8444 7744
rect 9312 7760 9364 7812
rect 10140 7692 10192 7744
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 11060 7692 11112 7744
rect 12440 7760 12492 7812
rect 12808 7828 12860 7880
rect 13360 7828 13412 7880
rect 14924 7828 14976 7880
rect 16304 7828 16356 7880
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 13912 7760 13964 7812
rect 15752 7760 15804 7812
rect 18420 7760 18472 7812
rect 21548 7760 21600 7812
rect 16028 7692 16080 7744
rect 16120 7692 16172 7744
rect 18972 7692 19024 7744
rect 21364 7735 21416 7744
rect 21364 7701 21373 7735
rect 21373 7701 21407 7735
rect 21407 7701 21416 7735
rect 21364 7692 21416 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 2688 7488 2740 7540
rect 2780 7488 2832 7540
rect 4436 7488 4488 7540
rect 5448 7488 5500 7540
rect 6000 7488 6052 7540
rect 6644 7488 6696 7540
rect 7104 7488 7156 7540
rect 8484 7488 8536 7540
rect 9128 7488 9180 7540
rect 1400 7420 1452 7472
rect 4160 7420 4212 7472
rect 7196 7420 7248 7472
rect 11244 7488 11296 7540
rect 11980 7488 12032 7540
rect 13912 7488 13964 7540
rect 16948 7488 17000 7540
rect 15108 7420 15160 7472
rect 15660 7420 15712 7472
rect 16028 7420 16080 7472
rect 18880 7488 18932 7540
rect 2412 7352 2464 7404
rect 3332 7352 3384 7404
rect 5172 7352 5224 7404
rect 9312 7352 9364 7404
rect 9496 7352 9548 7404
rect 11060 7352 11112 7404
rect 11428 7352 11480 7404
rect 11888 7352 11940 7404
rect 12808 7352 12860 7404
rect 1768 7327 1820 7336
rect 1768 7293 1777 7327
rect 1777 7293 1811 7327
rect 1811 7293 1820 7327
rect 1768 7284 1820 7293
rect 4804 7327 4856 7336
rect 4804 7293 4813 7327
rect 4813 7293 4847 7327
rect 4847 7293 4856 7327
rect 4804 7284 4856 7293
rect 6644 7284 6696 7336
rect 6736 7284 6788 7336
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 9772 7327 9824 7336
rect 7104 7216 7156 7268
rect 1584 7148 1636 7200
rect 3148 7191 3200 7200
rect 3148 7157 3157 7191
rect 3157 7157 3191 7191
rect 3191 7157 3200 7191
rect 3148 7148 3200 7157
rect 4252 7148 4304 7200
rect 5172 7148 5224 7200
rect 5632 7148 5684 7200
rect 7380 7191 7432 7200
rect 7380 7157 7389 7191
rect 7389 7157 7423 7191
rect 7423 7157 7432 7191
rect 7380 7148 7432 7157
rect 8944 7216 8996 7268
rect 9772 7293 9781 7327
rect 9781 7293 9815 7327
rect 9815 7293 9824 7327
rect 9772 7284 9824 7293
rect 13084 7352 13136 7404
rect 13636 7284 13688 7336
rect 9956 7216 10008 7268
rect 10140 7216 10192 7268
rect 11888 7216 11940 7268
rect 8024 7148 8076 7200
rect 11060 7148 11112 7200
rect 12256 7148 12308 7200
rect 16396 7352 16448 7404
rect 21272 7420 21324 7472
rect 18696 7395 18748 7404
rect 18696 7361 18705 7395
rect 18705 7361 18739 7395
rect 18739 7361 18748 7395
rect 18696 7352 18748 7361
rect 18972 7352 19024 7404
rect 19892 7395 19944 7404
rect 19892 7361 19901 7395
rect 19901 7361 19935 7395
rect 19935 7361 19944 7395
rect 19892 7352 19944 7361
rect 16304 7284 16356 7336
rect 17040 7284 17092 7336
rect 14372 7216 14424 7268
rect 18512 7259 18564 7268
rect 14280 7191 14332 7200
rect 14280 7157 14289 7191
rect 14289 7157 14323 7191
rect 14323 7157 14332 7191
rect 14280 7148 14332 7157
rect 18512 7225 18521 7259
rect 18521 7225 18555 7259
rect 18555 7225 18564 7259
rect 18512 7216 18564 7225
rect 19524 7216 19576 7268
rect 18880 7148 18932 7200
rect 19800 7148 19852 7200
rect 20444 7148 20496 7200
rect 20996 7191 21048 7200
rect 20996 7157 21005 7191
rect 21005 7157 21039 7191
rect 21039 7157 21048 7191
rect 20996 7148 21048 7157
rect 21456 7148 21508 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 1400 6944 1452 6996
rect 2044 6944 2096 6996
rect 2596 6944 2648 6996
rect 4068 6944 4120 6996
rect 5264 6944 5316 6996
rect 5540 6987 5592 6996
rect 3148 6876 3200 6928
rect 5540 6953 5549 6987
rect 5549 6953 5583 6987
rect 5583 6953 5592 6987
rect 5540 6944 5592 6953
rect 8392 6944 8444 6996
rect 18696 6944 18748 6996
rect 4528 6808 4580 6860
rect 6736 6876 6788 6928
rect 3976 6740 4028 6792
rect 8300 6876 8352 6928
rect 8576 6876 8628 6928
rect 5264 6740 5316 6792
rect 6736 6740 6788 6792
rect 7012 6783 7064 6792
rect 7012 6749 7021 6783
rect 7021 6749 7055 6783
rect 7055 6749 7064 6783
rect 7012 6740 7064 6749
rect 8668 6808 8720 6860
rect 9312 6808 9364 6860
rect 10600 6851 10652 6860
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10600 6817 10609 6851
rect 10609 6817 10643 6851
rect 10643 6817 10652 6851
rect 10600 6808 10652 6817
rect 11428 6876 11480 6928
rect 12440 6808 12492 6860
rect 13084 6851 13136 6860
rect 13084 6817 13093 6851
rect 13093 6817 13127 6851
rect 13127 6817 13136 6851
rect 13084 6808 13136 6817
rect 18420 6808 18472 6860
rect 11336 6783 11388 6792
rect 1768 6672 1820 6724
rect 1860 6604 1912 6656
rect 2136 6604 2188 6656
rect 2688 6604 2740 6656
rect 4436 6604 4488 6656
rect 4804 6604 4856 6656
rect 5172 6604 5224 6656
rect 5724 6604 5776 6656
rect 7196 6672 7248 6724
rect 8116 6672 8168 6724
rect 7472 6604 7524 6656
rect 7840 6647 7892 6656
rect 7840 6613 7849 6647
rect 7849 6613 7883 6647
rect 7883 6613 7892 6647
rect 9772 6672 9824 6724
rect 11336 6749 11345 6783
rect 11345 6749 11379 6783
rect 11379 6749 11388 6783
rect 11336 6740 11388 6749
rect 11980 6783 12032 6792
rect 11980 6749 11989 6783
rect 11989 6749 12023 6783
rect 12023 6749 12032 6783
rect 11980 6740 12032 6749
rect 13544 6740 13596 6792
rect 13636 6740 13688 6792
rect 14372 6783 14424 6792
rect 14372 6749 14406 6783
rect 14406 6749 14424 6783
rect 14372 6740 14424 6749
rect 16304 6740 16356 6792
rect 14280 6672 14332 6724
rect 16948 6672 17000 6724
rect 7840 6604 7892 6613
rect 8300 6604 8352 6656
rect 9404 6647 9456 6656
rect 9404 6613 9413 6647
rect 9413 6613 9447 6647
rect 9447 6613 9456 6647
rect 9404 6604 9456 6613
rect 10784 6604 10836 6656
rect 11244 6647 11296 6656
rect 11244 6613 11253 6647
rect 11253 6613 11287 6647
rect 11287 6613 11296 6647
rect 11244 6604 11296 6613
rect 11796 6604 11848 6656
rect 13268 6647 13320 6656
rect 13268 6613 13277 6647
rect 13277 6613 13311 6647
rect 13311 6613 13320 6647
rect 13268 6604 13320 6613
rect 14464 6604 14516 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16396 6604 16448 6656
rect 19432 6783 19484 6792
rect 19432 6749 19441 6783
rect 19441 6749 19475 6783
rect 19475 6749 19484 6783
rect 19432 6740 19484 6749
rect 19892 6783 19944 6792
rect 19892 6749 19901 6783
rect 19901 6749 19935 6783
rect 19935 6749 19944 6783
rect 19892 6740 19944 6749
rect 20260 6740 20312 6792
rect 17684 6604 17736 6656
rect 19708 6647 19760 6656
rect 19708 6613 19717 6647
rect 19717 6613 19751 6647
rect 19751 6613 19760 6647
rect 19708 6604 19760 6613
rect 20904 6672 20956 6724
rect 20812 6604 20864 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 2320 6443 2372 6452
rect 2320 6409 2329 6443
rect 2329 6409 2363 6443
rect 2363 6409 2372 6443
rect 2320 6400 2372 6409
rect 7380 6400 7432 6452
rect 3424 6332 3476 6384
rect 6736 6332 6788 6384
rect 8208 6400 8260 6452
rect 9680 6400 9732 6452
rect 10048 6400 10100 6452
rect 7840 6332 7892 6384
rect 13084 6400 13136 6452
rect 14464 6443 14516 6452
rect 14464 6409 14473 6443
rect 14473 6409 14507 6443
rect 14507 6409 14516 6443
rect 14464 6400 14516 6409
rect 15752 6400 15804 6452
rect 17040 6443 17092 6452
rect 17040 6409 17049 6443
rect 17049 6409 17083 6443
rect 17083 6409 17092 6443
rect 17040 6400 17092 6409
rect 17132 6443 17184 6452
rect 17132 6409 17141 6443
rect 17141 6409 17175 6443
rect 17175 6409 17184 6443
rect 17132 6400 17184 6409
rect 18144 6443 18196 6452
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 2688 6196 2740 6248
rect 3332 6196 3384 6248
rect 4804 6264 4856 6316
rect 6368 6264 6420 6316
rect 6552 6264 6604 6316
rect 7288 6264 7340 6316
rect 9128 6264 9180 6316
rect 17776 6332 17828 6384
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 18236 6400 18288 6452
rect 19156 6400 19208 6452
rect 19984 6443 20036 6452
rect 13084 6264 13136 6316
rect 14740 6264 14792 6316
rect 6000 6239 6052 6248
rect 1860 6128 1912 6180
rect 2596 6128 2648 6180
rect 6000 6205 6009 6239
rect 6009 6205 6043 6239
rect 6043 6205 6052 6239
rect 6000 6196 6052 6205
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3148 6060 3200 6112
rect 5356 6060 5408 6112
rect 5724 6060 5776 6112
rect 6460 6060 6512 6112
rect 8024 6196 8076 6248
rect 9496 6196 9548 6248
rect 10140 6128 10192 6180
rect 12348 6196 12400 6248
rect 13636 6239 13688 6248
rect 13636 6205 13645 6239
rect 13645 6205 13679 6239
rect 13679 6205 13688 6239
rect 13636 6196 13688 6205
rect 15476 6196 15528 6248
rect 16396 6264 16448 6316
rect 16856 6264 16908 6316
rect 17316 6264 17368 6316
rect 17868 6264 17920 6316
rect 18420 6264 18472 6316
rect 16948 6196 17000 6248
rect 17224 6239 17276 6248
rect 17224 6205 17233 6239
rect 17233 6205 17267 6239
rect 17267 6205 17276 6239
rect 17224 6196 17276 6205
rect 18512 6196 18564 6248
rect 19156 6196 19208 6248
rect 7840 6060 7892 6112
rect 8668 6060 8720 6112
rect 11796 6060 11848 6112
rect 12716 6060 12768 6112
rect 13728 6128 13780 6180
rect 15292 6128 15344 6180
rect 19984 6409 19993 6443
rect 19993 6409 20027 6443
rect 20027 6409 20036 6443
rect 19984 6400 20036 6409
rect 20812 6264 20864 6316
rect 21088 6264 21140 6316
rect 21456 6264 21508 6316
rect 15016 6060 15068 6112
rect 18696 6060 18748 6112
rect 18972 6060 19024 6112
rect 19984 6060 20036 6112
rect 20812 6060 20864 6112
rect 21180 6103 21232 6112
rect 21180 6069 21189 6103
rect 21189 6069 21223 6103
rect 21223 6069 21232 6103
rect 21180 6060 21232 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 3148 5856 3200 5908
rect 3884 5856 3936 5908
rect 4344 5856 4396 5908
rect 6000 5856 6052 5908
rect 6920 5856 6972 5908
rect 7656 5856 7708 5908
rect 10600 5856 10652 5908
rect 11888 5856 11940 5908
rect 14740 5899 14792 5908
rect 14740 5865 14749 5899
rect 14749 5865 14783 5899
rect 14783 5865 14792 5899
rect 14740 5856 14792 5865
rect 15292 5856 15344 5908
rect 15660 5856 15712 5908
rect 16856 5856 16908 5908
rect 2688 5788 2740 5840
rect 1860 5763 1912 5772
rect 1860 5729 1869 5763
rect 1869 5729 1903 5763
rect 1903 5729 1912 5763
rect 1860 5720 1912 5729
rect 2596 5720 2648 5772
rect 3516 5788 3568 5840
rect 5908 5788 5960 5840
rect 3332 5720 3384 5772
rect 7840 5763 7892 5772
rect 2044 5695 2096 5704
rect 2044 5661 2053 5695
rect 2053 5661 2087 5695
rect 2087 5661 2096 5695
rect 2044 5652 2096 5661
rect 3976 5652 4028 5704
rect 4068 5652 4120 5704
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 7840 5729 7849 5763
rect 7849 5729 7883 5763
rect 7883 5729 7892 5763
rect 7840 5720 7892 5729
rect 9956 5788 10008 5840
rect 17408 5856 17460 5908
rect 17684 5856 17736 5908
rect 18236 5788 18288 5840
rect 19892 5856 19944 5908
rect 21088 5899 21140 5908
rect 21088 5865 21097 5899
rect 21097 5865 21131 5899
rect 21131 5865 21140 5899
rect 21088 5856 21140 5865
rect 8208 5720 8260 5772
rect 8300 5652 8352 5704
rect 9680 5720 9732 5772
rect 16212 5720 16264 5772
rect 18052 5763 18104 5772
rect 18052 5729 18061 5763
rect 18061 5729 18095 5763
rect 18095 5729 18104 5763
rect 18052 5720 18104 5729
rect 18696 5720 18748 5772
rect 11888 5652 11940 5704
rect 13544 5695 13596 5704
rect 13544 5661 13553 5695
rect 13553 5661 13587 5695
rect 13587 5661 13596 5695
rect 13544 5652 13596 5661
rect 13636 5652 13688 5704
rect 15016 5695 15068 5704
rect 15016 5661 15025 5695
rect 15025 5661 15059 5695
rect 15059 5661 15068 5695
rect 15016 5652 15068 5661
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 16120 5652 16172 5704
rect 18144 5652 18196 5704
rect 18604 5652 18656 5704
rect 18880 5652 18932 5704
rect 21272 5788 21324 5840
rect 20996 5652 21048 5704
rect 21824 5652 21876 5704
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 11704 5584 11756 5636
rect 12716 5584 12768 5636
rect 18696 5584 18748 5636
rect 3056 5516 3108 5525
rect 4160 5559 4212 5568
rect 4160 5525 4169 5559
rect 4169 5525 4203 5559
rect 4203 5525 4212 5559
rect 4160 5516 4212 5525
rect 6828 5516 6880 5568
rect 6920 5516 6972 5568
rect 7380 5516 7432 5568
rect 8668 5516 8720 5568
rect 9680 5559 9732 5568
rect 9680 5525 9689 5559
rect 9689 5525 9723 5559
rect 9723 5525 9732 5559
rect 9680 5516 9732 5525
rect 9956 5516 10008 5568
rect 12256 5516 12308 5568
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 17500 5516 17552 5568
rect 18512 5516 18564 5568
rect 19892 5559 19944 5568
rect 19892 5525 19901 5559
rect 19901 5525 19935 5559
rect 19935 5525 19944 5559
rect 19892 5516 19944 5525
rect 20628 5559 20680 5568
rect 20628 5525 20637 5559
rect 20637 5525 20671 5559
rect 20671 5525 20680 5559
rect 20628 5516 20680 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 2872 5355 2924 5364
rect 2872 5321 2881 5355
rect 2881 5321 2915 5355
rect 2915 5321 2924 5355
rect 2872 5312 2924 5321
rect 3056 5312 3108 5364
rect 4712 5312 4764 5364
rect 8116 5312 8168 5364
rect 1676 5244 1728 5296
rect 3516 5244 3568 5296
rect 2504 5176 2556 5228
rect 4528 5176 4580 5228
rect 4988 5176 5040 5228
rect 5448 5219 5500 5228
rect 5448 5185 5457 5219
rect 5457 5185 5491 5219
rect 5491 5185 5500 5219
rect 5448 5176 5500 5185
rect 9404 5312 9456 5364
rect 9496 5355 9548 5364
rect 9496 5321 9505 5355
rect 9505 5321 9539 5355
rect 9539 5321 9548 5355
rect 9496 5312 9548 5321
rect 2136 5108 2188 5160
rect 3332 5151 3384 5160
rect 3332 5117 3341 5151
rect 3341 5117 3375 5151
rect 3375 5117 3384 5151
rect 3332 5108 3384 5117
rect 3424 5151 3476 5160
rect 3424 5117 3433 5151
rect 3433 5117 3467 5151
rect 3467 5117 3476 5151
rect 3424 5108 3476 5117
rect 8024 5176 8076 5228
rect 8484 5219 8536 5228
rect 8484 5185 8493 5219
rect 8493 5185 8527 5219
rect 8527 5185 8536 5219
rect 8484 5176 8536 5185
rect 10968 5244 11020 5296
rect 11704 5244 11756 5296
rect 12164 5244 12216 5296
rect 14372 5244 14424 5296
rect 16304 5244 16356 5296
rect 16948 5312 17000 5364
rect 17776 5312 17828 5364
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 10048 5176 10100 5228
rect 2320 4972 2372 5024
rect 5908 5040 5960 5092
rect 8392 5108 8444 5160
rect 8576 5151 8628 5160
rect 8576 5117 8585 5151
rect 8585 5117 8619 5151
rect 8619 5117 8628 5151
rect 11152 5176 11204 5228
rect 12348 5219 12400 5228
rect 12348 5185 12357 5219
rect 12357 5185 12391 5219
rect 12391 5185 12400 5219
rect 12348 5176 12400 5185
rect 8576 5108 8628 5117
rect 6552 5040 6604 5092
rect 8208 5040 8260 5092
rect 12256 5151 12308 5160
rect 12256 5117 12265 5151
rect 12265 5117 12299 5151
rect 12299 5117 12308 5151
rect 12256 5108 12308 5117
rect 15844 5219 15896 5228
rect 15844 5185 15853 5219
rect 15853 5185 15887 5219
rect 15887 5185 15896 5219
rect 15844 5176 15896 5185
rect 15936 5176 15988 5228
rect 17408 5176 17460 5228
rect 17960 5176 18012 5228
rect 19064 5312 19116 5364
rect 20352 5312 20404 5364
rect 18972 5244 19024 5296
rect 18604 5176 18656 5228
rect 19156 5176 19208 5228
rect 15568 5151 15620 5160
rect 15568 5117 15577 5151
rect 15577 5117 15611 5151
rect 15611 5117 15620 5151
rect 15568 5108 15620 5117
rect 15752 5151 15804 5160
rect 15752 5117 15761 5151
rect 15761 5117 15795 5151
rect 15795 5117 15804 5151
rect 15752 5108 15804 5117
rect 17132 5151 17184 5160
rect 17132 5117 17141 5151
rect 17141 5117 17175 5151
rect 17175 5117 17184 5151
rect 17132 5108 17184 5117
rect 17224 5151 17276 5160
rect 17224 5117 17233 5151
rect 17233 5117 17267 5151
rect 17267 5117 17276 5151
rect 19892 5176 19944 5228
rect 20444 5176 20496 5228
rect 19524 5151 19576 5160
rect 17224 5108 17276 5117
rect 8300 4972 8352 5024
rect 11704 5015 11756 5024
rect 11704 4981 11713 5015
rect 11713 4981 11747 5015
rect 11747 4981 11756 5015
rect 11704 4972 11756 4981
rect 17040 5040 17092 5092
rect 19524 5117 19533 5151
rect 19533 5117 19567 5151
rect 19567 5117 19576 5151
rect 19524 5108 19576 5117
rect 18880 5040 18932 5092
rect 13636 4972 13688 5024
rect 17960 4972 18012 5024
rect 18144 4972 18196 5024
rect 20904 5015 20956 5024
rect 20904 4981 20913 5015
rect 20913 4981 20947 5015
rect 20947 4981 20956 5015
rect 20904 4972 20956 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 3976 4768 4028 4820
rect 5448 4768 5500 4820
rect 10140 4811 10192 4820
rect 10140 4777 10149 4811
rect 10149 4777 10183 4811
rect 10183 4777 10192 4811
rect 10140 4768 10192 4777
rect 11888 4811 11940 4820
rect 1676 4743 1728 4752
rect 1676 4709 1685 4743
rect 1685 4709 1719 4743
rect 1719 4709 1728 4743
rect 1676 4700 1728 4709
rect 11888 4777 11897 4811
rect 11897 4777 11931 4811
rect 11931 4777 11940 4811
rect 11888 4768 11940 4777
rect 15752 4768 15804 4820
rect 16028 4768 16080 4820
rect 13636 4743 13688 4752
rect 1768 4632 1820 4684
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 8576 4632 8628 4684
rect 9128 4675 9180 4684
rect 9128 4641 9137 4675
rect 9137 4641 9171 4675
rect 9171 4641 9180 4675
rect 9128 4632 9180 4641
rect 2688 4564 2740 4616
rect 7932 4564 7984 4616
rect 13636 4709 13645 4743
rect 13645 4709 13679 4743
rect 13679 4709 13688 4743
rect 13636 4700 13688 4709
rect 10324 4632 10376 4684
rect 18052 4675 18104 4684
rect 18052 4641 18061 4675
rect 18061 4641 18095 4675
rect 18095 4641 18104 4675
rect 18052 4632 18104 4641
rect 9864 4564 9916 4616
rect 11152 4564 11204 4616
rect 12532 4607 12584 4616
rect 12532 4573 12566 4607
rect 12566 4573 12584 4607
rect 14096 4607 14148 4616
rect 12532 4564 12584 4573
rect 14096 4573 14105 4607
rect 14105 4573 14139 4607
rect 14139 4573 14148 4607
rect 14096 4564 14148 4573
rect 16304 4564 16356 4616
rect 18512 4607 18564 4616
rect 18512 4573 18521 4607
rect 18521 4573 18555 4607
rect 18555 4573 18564 4607
rect 18512 4564 18564 4573
rect 1584 4496 1636 4548
rect 5448 4496 5500 4548
rect 6644 4496 6696 4548
rect 9956 4496 10008 4548
rect 10324 4496 10376 4548
rect 3056 4428 3108 4480
rect 4804 4428 4856 4480
rect 7932 4428 7984 4480
rect 8208 4471 8260 4480
rect 8208 4437 8217 4471
rect 8217 4437 8251 4471
rect 8251 4437 8260 4471
rect 8208 4428 8260 4437
rect 9496 4428 9548 4480
rect 10416 4428 10468 4480
rect 11060 4496 11112 4548
rect 15936 4496 15988 4548
rect 17040 4496 17092 4548
rect 17684 4496 17736 4548
rect 14740 4471 14792 4480
rect 14740 4437 14749 4471
rect 14749 4437 14783 4471
rect 14783 4437 14792 4471
rect 14740 4428 14792 4437
rect 15568 4428 15620 4480
rect 16396 4428 16448 4480
rect 16948 4428 17000 4480
rect 17868 4428 17920 4480
rect 18052 4428 18104 4480
rect 18972 4428 19024 4480
rect 21180 4496 21232 4548
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 3240 4224 3292 4276
rect 5356 4224 5408 4276
rect 6000 4267 6052 4276
rect 6000 4233 6009 4267
rect 6009 4233 6043 4267
rect 6043 4233 6052 4267
rect 6000 4224 6052 4233
rect 7104 4224 7156 4276
rect 8208 4224 8260 4276
rect 9220 4224 9272 4276
rect 2872 4088 2924 4140
rect 2228 4063 2280 4072
rect 2228 4029 2237 4063
rect 2237 4029 2271 4063
rect 2271 4029 2280 4063
rect 2228 4020 2280 4029
rect 2964 4020 3016 4072
rect 3148 4020 3200 4072
rect 4436 4088 4488 4140
rect 4896 4088 4948 4140
rect 6552 4088 6604 4140
rect 6920 4131 6972 4140
rect 6920 4097 6929 4131
rect 6929 4097 6963 4131
rect 6963 4097 6972 4131
rect 6920 4088 6972 4097
rect 7472 4156 7524 4208
rect 9864 4156 9916 4208
rect 8024 4131 8076 4140
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 5264 4020 5316 4072
rect 5540 4063 5592 4072
rect 3976 3995 4028 4004
rect 3976 3961 3985 3995
rect 3985 3961 4019 3995
rect 4019 3961 4028 3995
rect 3976 3952 4028 3961
rect 4068 3952 4120 4004
rect 5540 4029 5549 4063
rect 5549 4029 5583 4063
rect 5583 4029 5592 4063
rect 5540 4020 5592 4029
rect 5908 4020 5960 4072
rect 6460 4020 6512 4072
rect 6828 4020 6880 4072
rect 6552 3952 6604 4004
rect 7380 3995 7432 4004
rect 7380 3961 7389 3995
rect 7389 3961 7423 3995
rect 7423 3961 7432 3995
rect 7380 3952 7432 3961
rect 8024 4097 8033 4131
rect 8033 4097 8067 4131
rect 8067 4097 8076 4131
rect 8024 4088 8076 4097
rect 8576 3952 8628 4004
rect 9680 4020 9732 4072
rect 9864 4063 9916 4072
rect 9864 4029 9873 4063
rect 9873 4029 9907 4063
rect 9907 4029 9916 4063
rect 9864 4020 9916 4029
rect 10324 4224 10376 4276
rect 10508 4267 10560 4276
rect 10508 4233 10517 4267
rect 10517 4233 10551 4267
rect 10551 4233 10560 4267
rect 10508 4224 10560 4233
rect 11704 4224 11756 4276
rect 13820 4224 13872 4276
rect 14096 4267 14148 4276
rect 14096 4233 14105 4267
rect 14105 4233 14139 4267
rect 14139 4233 14148 4267
rect 14096 4224 14148 4233
rect 19524 4224 19576 4276
rect 10140 4199 10192 4208
rect 10140 4165 10149 4199
rect 10149 4165 10183 4199
rect 10183 4165 10192 4199
rect 10140 4156 10192 4165
rect 10416 4156 10468 4208
rect 10324 4088 10376 4140
rect 14740 4156 14792 4208
rect 16948 4156 17000 4208
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 13820 4088 13872 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 16212 4131 16264 4140
rect 8300 3884 8352 3936
rect 8484 3884 8536 3936
rect 10416 3952 10468 4004
rect 10692 3952 10744 4004
rect 11888 3952 11940 4004
rect 16212 4097 16221 4131
rect 16221 4097 16255 4131
rect 16255 4097 16264 4131
rect 16212 4088 16264 4097
rect 17868 4156 17920 4208
rect 17960 4156 18012 4208
rect 18696 4131 18748 4140
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 16856 4063 16908 4072
rect 16856 4029 16865 4063
rect 16865 4029 16899 4063
rect 16899 4029 16908 4063
rect 16856 4020 16908 4029
rect 17132 4020 17184 4072
rect 17776 4020 17828 4072
rect 19248 4020 19300 4072
rect 20812 4088 20864 4140
rect 20996 4131 21048 4140
rect 20996 4097 21005 4131
rect 21005 4097 21039 4131
rect 21039 4097 21048 4131
rect 20996 4088 21048 4097
rect 12900 3884 12952 3936
rect 13360 3884 13412 3936
rect 17316 3952 17368 4004
rect 19892 3995 19944 4004
rect 19892 3961 19901 3995
rect 19901 3961 19935 3995
rect 19935 3961 19944 3995
rect 19892 3952 19944 3961
rect 22284 3952 22336 4004
rect 13728 3884 13780 3936
rect 14556 3884 14608 3936
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 15844 3884 15896 3936
rect 17224 3884 17276 3936
rect 17592 3884 17644 3936
rect 17776 3884 17828 3936
rect 20996 3884 21048 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 3148 3680 3200 3732
rect 3332 3655 3384 3664
rect 3332 3621 3341 3655
rect 3341 3621 3375 3655
rect 3375 3621 3384 3655
rect 3332 3612 3384 3621
rect 3884 3680 3936 3732
rect 5540 3680 5592 3732
rect 7104 3680 7156 3732
rect 4528 3612 4580 3664
rect 6552 3655 6604 3664
rect 6552 3621 6561 3655
rect 6561 3621 6595 3655
rect 6595 3621 6604 3655
rect 6552 3612 6604 3621
rect 7012 3612 7064 3664
rect 7472 3612 7524 3664
rect 7656 3612 7708 3664
rect 2780 3587 2832 3596
rect 2780 3553 2789 3587
rect 2789 3553 2823 3587
rect 2823 3553 2832 3587
rect 2780 3544 2832 3553
rect 3424 3544 3476 3596
rect 5172 3587 5224 3596
rect 2780 3408 2832 3460
rect 3148 3451 3200 3460
rect 3148 3417 3157 3451
rect 3157 3417 3191 3451
rect 3191 3417 3200 3451
rect 3148 3408 3200 3417
rect 1584 3340 1636 3392
rect 4528 3476 4580 3528
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5724 3476 5776 3528
rect 4436 3408 4488 3460
rect 8024 3587 8076 3596
rect 8024 3553 8033 3587
rect 8033 3553 8067 3587
rect 8067 3553 8076 3587
rect 8024 3544 8076 3553
rect 8484 3544 8536 3596
rect 11152 3680 11204 3732
rect 17040 3680 17092 3732
rect 17960 3680 18012 3732
rect 18236 3680 18288 3732
rect 11060 3612 11112 3664
rect 7932 3476 7984 3528
rect 6828 3340 6880 3392
rect 7196 3383 7248 3392
rect 7196 3349 7205 3383
rect 7205 3349 7239 3383
rect 7239 3349 7248 3383
rect 7196 3340 7248 3349
rect 7380 3340 7432 3392
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9220 3476 9272 3528
rect 11244 3544 11296 3596
rect 10876 3476 10928 3528
rect 11060 3476 11112 3528
rect 12072 3612 12124 3664
rect 17868 3612 17920 3664
rect 19064 3612 19116 3664
rect 13636 3544 13688 3596
rect 14280 3587 14332 3596
rect 14280 3553 14289 3587
rect 14289 3553 14323 3587
rect 14323 3553 14332 3587
rect 14280 3544 14332 3553
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 12900 3519 12952 3528
rect 12900 3485 12909 3519
rect 12909 3485 12943 3519
rect 12943 3485 12952 3519
rect 12900 3476 12952 3485
rect 15476 3544 15528 3596
rect 16028 3544 16080 3596
rect 10600 3408 10652 3460
rect 10232 3340 10284 3392
rect 10324 3340 10376 3392
rect 14648 3408 14700 3460
rect 15752 3476 15804 3528
rect 16580 3476 16632 3528
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 20076 3544 20128 3596
rect 20168 3519 20220 3528
rect 20168 3485 20177 3519
rect 20177 3485 20211 3519
rect 20211 3485 20220 3519
rect 20168 3476 20220 3485
rect 20536 3476 20588 3528
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 14372 3383 14424 3392
rect 14372 3349 14381 3383
rect 14381 3349 14415 3383
rect 14415 3349 14424 3383
rect 14372 3340 14424 3349
rect 15476 3383 15528 3392
rect 15476 3349 15485 3383
rect 15485 3349 15519 3383
rect 15519 3349 15528 3383
rect 15476 3340 15528 3349
rect 15936 3340 15988 3392
rect 18696 3408 18748 3460
rect 16948 3340 17000 3392
rect 18512 3340 18564 3392
rect 20076 3340 20128 3392
rect 20536 3340 20588 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 2688 3179 2740 3188
rect 2688 3145 2697 3179
rect 2697 3145 2731 3179
rect 2731 3145 2740 3179
rect 2688 3136 2740 3145
rect 2780 3136 2832 3188
rect 1860 3068 1912 3120
rect 4436 3068 4488 3120
rect 4712 3136 4764 3188
rect 7288 3136 7340 3188
rect 2412 3000 2464 3052
rect 2504 3043 2556 3052
rect 2504 3009 2513 3043
rect 2513 3009 2547 3043
rect 2547 3009 2556 3043
rect 2504 3000 2556 3009
rect 2780 2932 2832 2984
rect 5172 3000 5224 3052
rect 5264 3000 5316 3052
rect 4436 2932 4488 2984
rect 4712 2932 4764 2984
rect 4896 2932 4948 2984
rect 7840 3000 7892 3052
rect 8024 3068 8076 3120
rect 9864 3136 9916 3188
rect 10048 3136 10100 3188
rect 11796 3136 11848 3188
rect 12532 3136 12584 3188
rect 13636 3179 13688 3188
rect 13636 3145 13645 3179
rect 13645 3145 13679 3179
rect 13679 3145 13688 3179
rect 13636 3136 13688 3145
rect 13820 3136 13872 3188
rect 15384 3136 15436 3188
rect 15660 3136 15712 3188
rect 17868 3136 17920 3188
rect 7104 2932 7156 2984
rect 9128 3000 9180 3052
rect 9496 3000 9548 3052
rect 9680 3000 9732 3052
rect 11244 3068 11296 3120
rect 12348 3068 12400 3120
rect 11704 3000 11756 3052
rect 12072 3000 12124 3052
rect 13084 3068 13136 3120
rect 13728 3068 13780 3120
rect 18972 3068 19024 3120
rect 14556 3000 14608 3052
rect 16120 3000 16172 3052
rect 17316 3000 17368 3052
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 572 2864 624 2916
rect 3332 2864 3384 2916
rect 204 2796 256 2848
rect 1308 2796 1360 2848
rect 2228 2796 2280 2848
rect 2780 2796 2832 2848
rect 6552 2796 6604 2848
rect 8024 2796 8076 2848
rect 11152 2932 11204 2984
rect 14280 2932 14332 2984
rect 18880 3000 18932 3052
rect 19800 3068 19852 3120
rect 19616 3000 19668 3052
rect 21364 3043 21416 3052
rect 21364 3009 21373 3043
rect 21373 3009 21407 3043
rect 21407 3009 21416 3043
rect 21364 3000 21416 3009
rect 22744 3000 22796 3052
rect 11060 2796 11112 2848
rect 12164 2864 12216 2916
rect 14740 2864 14792 2916
rect 11888 2796 11940 2848
rect 12072 2796 12124 2848
rect 15292 2796 15344 2848
rect 19984 2932 20036 2984
rect 20720 2975 20772 2984
rect 20720 2941 20729 2975
rect 20729 2941 20763 2975
rect 20763 2941 20772 2975
rect 20720 2932 20772 2941
rect 16396 2864 16448 2916
rect 18696 2796 18748 2848
rect 19616 2796 19668 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 7196 2592 7248 2644
rect 7564 2592 7616 2644
rect 8024 2592 8076 2644
rect 10140 2635 10192 2644
rect 5264 2524 5316 2576
rect 6644 2524 6696 2576
rect 8208 2524 8260 2576
rect 9680 2524 9732 2576
rect 10140 2601 10149 2635
rect 10149 2601 10183 2635
rect 10183 2601 10192 2635
rect 10140 2592 10192 2601
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 10876 2592 10928 2644
rect 13452 2592 13504 2644
rect 16120 2592 16172 2644
rect 2228 2499 2280 2508
rect 2228 2465 2237 2499
rect 2237 2465 2271 2499
rect 2271 2465 2280 2499
rect 2228 2456 2280 2465
rect 3332 2499 3384 2508
rect 3332 2465 3341 2499
rect 3341 2465 3375 2499
rect 3375 2465 3384 2499
rect 3332 2456 3384 2465
rect 4712 2456 4764 2508
rect 4804 2456 4856 2508
rect 7104 2456 7156 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3240 2388 3292 2440
rect 4068 2320 4120 2372
rect 5816 2388 5868 2440
rect 8300 2388 8352 2440
rect 8392 2388 8444 2440
rect 9312 2456 9364 2508
rect 10968 2499 11020 2508
rect 10968 2465 10977 2499
rect 10977 2465 11011 2499
rect 11011 2465 11020 2499
rect 10968 2456 11020 2465
rect 12532 2524 12584 2576
rect 13636 2524 13688 2576
rect 8668 2388 8720 2440
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 9956 2388 10008 2440
rect 10508 2388 10560 2440
rect 12164 2456 12216 2508
rect 13636 2388 13688 2440
rect 13820 2388 13872 2440
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 15292 2431 15344 2440
rect 15292 2397 15301 2431
rect 15301 2397 15335 2431
rect 15335 2397 15344 2431
rect 15292 2388 15344 2397
rect 16212 2524 16264 2576
rect 17500 2592 17552 2644
rect 18328 2524 18380 2576
rect 19984 2524 20036 2576
rect 5724 2252 5776 2304
rect 7288 2252 7340 2304
rect 12992 2320 13044 2372
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 10140 2252 10192 2304
rect 10968 2252 11020 2304
rect 11888 2295 11940 2304
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 13176 2295 13228 2304
rect 13176 2261 13185 2295
rect 13185 2261 13219 2295
rect 13219 2261 13228 2295
rect 13176 2252 13228 2261
rect 13268 2252 13320 2304
rect 15200 2320 15252 2372
rect 17960 2388 18012 2440
rect 18144 2388 18196 2440
rect 20812 2456 20864 2508
rect 21456 2456 21508 2508
rect 19708 2388 19760 2440
rect 20628 2388 20680 2440
rect 16948 2320 17000 2372
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 8576 2048 8628 2100
rect 11888 2048 11940 2100
rect 15292 2048 15344 2100
rect 18052 2048 18104 2100
rect 8208 1980 8260 2032
rect 13268 1980 13320 2032
rect 13912 1980 13964 2032
rect 16212 1980 16264 2032
rect 4436 1912 4488 1964
rect 13176 1912 13228 1964
rect 13820 1912 13872 1964
rect 17776 1912 17828 1964
rect 3056 1844 3108 1896
rect 7012 1844 7064 1896
rect 14096 1844 14148 1896
rect 1584 1708 1636 1760
rect 9680 1776 9732 1828
rect 15844 1776 15896 1828
rect 7288 1708 7340 1760
rect 9772 1708 9824 1760
rect 10692 1708 10744 1760
rect 14372 1708 14424 1760
rect 9220 1640 9272 1692
rect 10140 1640 10192 1692
rect 8392 1572 8444 1624
rect 2872 1300 2924 1352
rect 18420 1300 18472 1352
<< metal2 >>
rect 1490 22672 1546 22681
rect 1490 22607 1546 22616
rect 1504 20806 1532 22607
rect 3146 22264 3202 22273
rect 3146 22199 3202 22208
rect 2594 21720 2650 21729
rect 2594 21655 2650 21664
rect 1950 21312 2006 21321
rect 1950 21247 2006 21256
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20534 1532 20742
rect 1492 20528 1544 20534
rect 1492 20470 1544 20476
rect 1860 20324 1912 20330
rect 1860 20266 1912 20272
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1490 18864 1546 18873
rect 1490 18799 1546 18808
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1676 18624 1728 18630
rect 1676 18566 1728 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1688 17678 1716 18566
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1492 17536 1544 17542
rect 1490 17504 1492 17513
rect 1676 17536 1728 17542
rect 1544 17504 1546 17513
rect 1676 17478 1728 17484
rect 1490 17439 1546 17448
rect 1490 17096 1546 17105
rect 1490 17031 1492 17040
rect 1544 17031 1546 17040
rect 1492 17002 1544 17008
rect 1688 16590 1716 17478
rect 1768 17060 1820 17066
rect 1768 17002 1820 17008
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16153 1532 16390
rect 1490 16144 1546 16153
rect 1780 16114 1808 17002
rect 1490 16079 1546 16088
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15609 1532 15846
rect 1490 15600 1546 15609
rect 1872 15586 1900 20266
rect 1964 19514 1992 21247
rect 2228 20460 2280 20466
rect 2228 20402 2280 20408
rect 2042 20360 2098 20369
rect 2042 20295 2044 20304
rect 2096 20295 2098 20304
rect 2044 20266 2096 20272
rect 2240 19990 2268 20402
rect 2320 20324 2372 20330
rect 2320 20266 2372 20272
rect 2228 19984 2280 19990
rect 2228 19926 2280 19932
rect 2042 19816 2098 19825
rect 2042 19751 2098 19760
rect 2056 19718 2084 19751
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 2332 19378 2360 20266
rect 2608 20058 2636 21655
rect 2778 20768 2834 20777
rect 2778 20703 2834 20712
rect 2792 20602 2820 20703
rect 3160 20602 3188 22199
rect 4712 20800 4764 20806
rect 4712 20742 4764 20748
rect 4724 20602 4752 20742
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 2780 20596 2832 20602
rect 2780 20538 2832 20544
rect 3148 20596 3200 20602
rect 3148 20538 3200 20544
rect 4712 20596 4764 20602
rect 4712 20538 4764 20544
rect 8208 20528 8260 20534
rect 8208 20470 8260 20476
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 3988 20058 4016 20402
rect 4160 20392 4212 20398
rect 4160 20334 4212 20340
rect 4172 20058 4200 20334
rect 4436 20256 4488 20262
rect 4436 20198 4488 20204
rect 2596 20052 2648 20058
rect 2596 19994 2648 20000
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4160 20052 4212 20058
rect 4160 19994 4212 20000
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2700 19242 2728 19314
rect 2688 19236 2740 19242
rect 2688 19178 2740 19184
rect 2044 19168 2096 19174
rect 2044 19110 2096 19116
rect 2056 18290 2084 19110
rect 2976 18986 3004 19858
rect 4448 19854 4476 20198
rect 6552 19916 6604 19922
rect 6552 19858 6604 19864
rect 3608 19848 3660 19854
rect 3608 19790 3660 19796
rect 4436 19848 4488 19854
rect 4436 19790 4488 19796
rect 4528 19848 4580 19854
rect 4528 19790 4580 19796
rect 3620 19514 3648 19790
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 3896 19514 3924 19654
rect 4540 19514 4568 19790
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 3608 19508 3660 19514
rect 3608 19450 3660 19456
rect 3884 19508 3936 19514
rect 3884 19450 3936 19456
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 5908 19440 5960 19446
rect 5908 19382 5960 19388
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 2976 18958 3280 18986
rect 3068 18834 3188 18850
rect 3068 18828 3200 18834
rect 3068 18822 3148 18828
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 2148 18426 2176 18702
rect 2136 18420 2188 18426
rect 2136 18362 2188 18368
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1490 15535 1546 15544
rect 1780 15558 1900 15586
rect 1964 15570 1992 16934
rect 2042 16552 2098 16561
rect 2042 16487 2098 16496
rect 2056 16454 2084 16487
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2148 16250 2176 17138
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2136 16108 2188 16114
rect 2136 16050 2188 16056
rect 1952 15564 2004 15570
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1676 15360 1728 15366
rect 1676 15302 1728 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 1688 15026 1716 15302
rect 1676 15020 1728 15026
rect 1676 14962 1728 14968
rect 1780 14822 1808 15558
rect 1952 15506 2004 15512
rect 1860 15496 1912 15502
rect 1860 15438 1912 15444
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1768 14816 1820 14822
rect 1768 14758 1820 14764
rect 1504 14657 1532 14758
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1400 13864 1452 13870
rect 1504 13841 1532 14214
rect 1400 13806 1452 13812
rect 1490 13832 1546 13841
rect 1214 12336 1270 12345
rect 1214 12271 1270 12280
rect 1228 8974 1256 12271
rect 1308 9104 1360 9110
rect 1308 9046 1360 9052
rect 1216 8968 1268 8974
rect 1216 8910 1268 8916
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 800 244 2790
rect 584 800 612 2858
rect 1320 2854 1348 9046
rect 1412 7478 1440 13806
rect 1490 13767 1546 13776
rect 1584 13320 1636 13326
rect 1490 13288 1546 13297
rect 1584 13262 1636 13268
rect 1490 13223 1546 13232
rect 1504 12986 1532 13223
rect 1492 12980 1544 12986
rect 1492 12922 1544 12928
rect 1596 11914 1624 13262
rect 1504 11886 1624 11914
rect 1688 11898 1716 14350
rect 1872 12442 1900 15438
rect 2044 14272 2096 14278
rect 2042 14240 2044 14249
rect 2096 14240 2098 14249
rect 2042 14175 2098 14184
rect 2148 14090 2176 16050
rect 2056 14062 2176 14090
rect 2056 12442 2084 14062
rect 2136 13932 2188 13938
rect 2136 13874 2188 13880
rect 1860 12436 1912 12442
rect 1860 12378 1912 12384
rect 2044 12436 2096 12442
rect 2044 12378 2096 12384
rect 1860 12232 1912 12238
rect 1860 12174 1912 12180
rect 1676 11892 1728 11898
rect 1504 9450 1532 11886
rect 1676 11834 1728 11840
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 11354 1624 11698
rect 1584 11348 1636 11354
rect 1584 11290 1636 11296
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1780 10742 1808 11086
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1872 10554 1900 12174
rect 1952 11688 2004 11694
rect 1952 11630 2004 11636
rect 1964 11150 1992 11630
rect 2044 11552 2096 11558
rect 2044 11494 2096 11500
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 1872 10526 1992 10554
rect 1860 10124 1912 10130
rect 1860 10066 1912 10072
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 9042 1532 9386
rect 1582 9208 1638 9217
rect 1582 9143 1584 9152
rect 1636 9143 1638 9152
rect 1584 9114 1636 9120
rect 1492 9036 1544 9042
rect 1492 8978 1544 8984
rect 1674 8800 1730 8809
rect 1674 8735 1730 8744
rect 1400 7472 1452 7478
rect 1400 7414 1452 7420
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1400 6996 1452 7002
rect 1400 6938 1452 6944
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1412 2553 1440 6938
rect 1490 6352 1546 6361
rect 1490 6287 1492 6296
rect 1544 6287 1546 6296
rect 1492 6258 1544 6264
rect 1504 3369 1532 6258
rect 1596 5681 1624 7142
rect 1688 6458 1716 8735
rect 1768 7336 1820 7342
rect 1768 7278 1820 7284
rect 1780 6730 1808 7278
rect 1768 6724 1820 6730
rect 1768 6666 1820 6672
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1582 5672 1638 5681
rect 1582 5607 1638 5616
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1688 4758 1716 5238
rect 1676 4752 1728 4758
rect 1676 4694 1728 4700
rect 1780 4690 1808 6666
rect 1872 6662 1900 10066
rect 1964 9178 1992 10526
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 2056 7002 2084 11494
rect 2044 6996 2096 7002
rect 2044 6938 2096 6944
rect 2148 6662 2176 13874
rect 2240 13274 2268 18702
rect 2596 18624 2648 18630
rect 2596 18566 2648 18572
rect 2608 18426 2636 18566
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 3068 18170 3096 18822
rect 3148 18770 3200 18776
rect 3148 18692 3200 18698
rect 3148 18634 3200 18640
rect 2976 18142 3096 18170
rect 2976 18086 3004 18142
rect 3160 18086 3188 18634
rect 3252 18630 3280 18958
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 3148 18080 3200 18086
rect 3148 18022 3200 18028
rect 3148 17808 3200 17814
rect 3148 17750 3200 17756
rect 2412 17672 2464 17678
rect 2412 17614 2464 17620
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2320 17604 2372 17610
rect 2320 17546 2372 17552
rect 2332 15162 2360 17546
rect 2424 15706 2452 17614
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2608 16250 2636 17138
rect 2792 16794 2820 17614
rect 2872 17536 2924 17542
rect 2872 17478 2924 17484
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2688 16584 2740 16590
rect 2688 16526 2740 16532
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2320 14816 2372 14822
rect 2320 14758 2372 14764
rect 2332 14006 2360 14758
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2424 14074 2452 14350
rect 2412 14068 2464 14074
rect 2412 14010 2464 14016
rect 2320 14000 2372 14006
rect 2372 13948 2452 13954
rect 2320 13942 2452 13948
rect 2332 13926 2452 13942
rect 2332 13877 2360 13926
rect 2240 13246 2360 13274
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 10674 2268 13126
rect 2332 12170 2360 13246
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2424 11778 2452 13926
rect 2608 12186 2636 16050
rect 2700 15858 2728 16526
rect 2884 16522 2912 17478
rect 2964 17128 3016 17134
rect 2964 17070 3016 17076
rect 2976 16794 3004 17070
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 3160 16590 3188 17750
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 2872 16516 2924 16522
rect 2872 16458 2924 16464
rect 3252 16454 3280 18294
rect 3344 18086 3372 19246
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 5632 18896 5684 18902
rect 5632 18838 5684 18844
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 4528 18284 4580 18290
rect 4528 18226 4580 18232
rect 3332 18080 3384 18086
rect 3332 18022 3384 18028
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3424 17604 3476 17610
rect 3424 17546 3476 17552
rect 3436 17338 3464 17546
rect 3896 17542 3924 18226
rect 4540 17678 4568 18226
rect 4724 18154 4752 18566
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 5356 18080 5408 18086
rect 5356 18022 5408 18028
rect 4528 17672 4580 17678
rect 4528 17614 4580 17620
rect 3884 17536 3936 17542
rect 3884 17478 3936 17484
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 3896 16658 3924 17478
rect 4252 17196 4304 17202
rect 4304 17156 4384 17184
rect 4252 17138 4304 17144
rect 4160 17128 4212 17134
rect 4160 17070 4212 17076
rect 3884 16652 3936 16658
rect 3884 16594 3936 16600
rect 4172 16590 4200 17070
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3240 16448 3292 16454
rect 3240 16390 3292 16396
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4264 16250 4292 16390
rect 4252 16244 4304 16250
rect 4252 16186 4304 16192
rect 2872 16108 2924 16114
rect 2872 16050 2924 16056
rect 2700 15830 2820 15858
rect 2792 15706 2820 15830
rect 2780 15700 2832 15706
rect 2780 15642 2832 15648
rect 2884 15162 2912 16050
rect 4356 15978 4384 17156
rect 4540 16182 4568 17614
rect 4632 17202 4660 18022
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 5368 16590 5396 18022
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 4528 16176 4580 16182
rect 4528 16118 4580 16124
rect 4344 15972 4396 15978
rect 4344 15914 4396 15920
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 3332 15564 3384 15570
rect 3332 15506 3384 15512
rect 2872 15156 2924 15162
rect 2872 15098 2924 15104
rect 3344 15026 3372 15506
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 3896 14414 3924 15846
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4160 15360 4212 15366
rect 4160 15302 4212 15308
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4172 14482 4200 15302
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3896 13938 3924 14350
rect 2964 13932 3016 13938
rect 2964 13874 3016 13880
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 4160 13932 4212 13938
rect 4160 13874 4212 13880
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2884 12442 2912 13806
rect 2872 12436 2924 12442
rect 2872 12378 2924 12384
rect 2976 12322 3004 13874
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 2792 12306 3004 12322
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 2780 12300 3004 12306
rect 2832 12294 3004 12300
rect 2780 12242 2832 12248
rect 2608 12158 2728 12186
rect 2504 12096 2556 12102
rect 2504 12038 2556 12044
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2516 11898 2544 12038
rect 2504 11892 2556 11898
rect 2504 11834 2556 11840
rect 2424 11750 2544 11778
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2516 9926 2544 11750
rect 2608 10266 2636 12038
rect 2596 10260 2648 10266
rect 2596 10202 2648 10208
rect 2700 10198 2728 12158
rect 2792 11354 2820 12242
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2884 11218 2912 11698
rect 3068 11234 3096 12310
rect 2872 11212 2924 11218
rect 2872 11154 2924 11160
rect 2976 11206 3096 11234
rect 2688 10192 2740 10198
rect 2976 10146 3004 11206
rect 3056 11144 3108 11150
rect 3056 11086 3108 11092
rect 3068 10810 3096 11086
rect 3160 10810 3188 12718
rect 3252 11762 3280 13670
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 3792 13456 3844 13462
rect 3792 13398 3844 13404
rect 3804 12889 3832 13398
rect 3790 12880 3846 12889
rect 3896 12850 3924 13874
rect 4172 13530 4200 13874
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4264 13190 4292 14894
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4448 13462 4476 13874
rect 4436 13456 4488 13462
rect 4436 13398 4488 13404
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4528 13184 4580 13190
rect 4528 13126 4580 13132
rect 4540 12986 4568 13126
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 4528 12980 4580 12986
rect 4528 12922 4580 12928
rect 3790 12815 3846 12824
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 4160 12844 4212 12850
rect 4160 12786 4212 12792
rect 3976 12776 4028 12782
rect 3976 12718 4028 12724
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3422 11384 3478 11393
rect 3549 11376 3857 11396
rect 3422 11319 3424 11328
rect 3476 11319 3478 11328
rect 3424 11290 3476 11296
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2688 10134 2740 10140
rect 2792 10118 3004 10146
rect 3068 10130 3096 10746
rect 3056 10124 3108 10130
rect 2228 9920 2280 9926
rect 2226 9888 2228 9897
rect 2504 9920 2556 9926
rect 2280 9888 2282 9897
rect 2504 9862 2556 9868
rect 2226 9823 2282 9832
rect 2320 9580 2372 9586
rect 2320 9522 2372 9528
rect 2332 8634 2360 9522
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2332 7954 2360 8570
rect 2424 8090 2452 8774
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2516 7970 2544 9862
rect 2792 9194 2820 10118
rect 3056 10066 3108 10072
rect 3252 10010 3280 11086
rect 3424 11008 3476 11014
rect 3424 10950 3476 10956
rect 3436 10441 3464 10950
rect 3422 10432 3478 10441
rect 3422 10367 3478 10376
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2976 9982 3280 10010
rect 2700 9166 2820 9194
rect 2700 9042 2728 9166
rect 2688 9036 2740 9042
rect 2688 8978 2740 8984
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2608 8498 2636 8570
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2320 7948 2372 7954
rect 2320 7890 2372 7896
rect 2424 7942 2544 7970
rect 2424 7834 2452 7942
rect 2332 7806 2452 7834
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1872 6186 1900 6598
rect 2332 6458 2360 7806
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2320 6452 2372 6458
rect 2320 6394 2372 6400
rect 1860 6180 1912 6186
rect 1860 6122 1912 6128
rect 2042 5808 2098 5817
rect 1860 5772 1912 5778
rect 2042 5743 2098 5752
rect 1860 5714 1912 5720
rect 1768 4684 1820 4690
rect 1768 4626 1820 4632
rect 1584 4548 1636 4554
rect 1584 4490 1636 4496
rect 1596 3398 1624 4490
rect 1584 3392 1636 3398
rect 1490 3360 1546 3369
rect 1584 3334 1636 3340
rect 1490 3295 1546 3304
rect 1398 2544 1454 2553
rect 1398 2479 1454 2488
rect 1030 2000 1086 2009
rect 1030 1935 1086 1944
rect 1044 800 1072 1935
rect 1596 1766 1624 3334
rect 1872 3126 1900 5714
rect 2056 5710 2084 5743
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2148 4185 2176 5102
rect 2320 5024 2372 5030
rect 2320 4966 2372 4972
rect 2134 4176 2190 4185
rect 2134 4111 2190 4120
rect 1860 3120 1912 3126
rect 1860 3062 1912 3068
rect 1950 2816 2006 2825
rect 1950 2751 2006 2760
rect 1584 1760 1636 1766
rect 1490 1728 1546 1737
rect 1584 1702 1636 1708
rect 1490 1663 1546 1672
rect 1504 800 1532 1663
rect 1964 800 1992 2751
rect 2148 2145 2176 4111
rect 2228 4072 2280 4078
rect 2226 4040 2228 4049
rect 2280 4040 2282 4049
rect 2226 3975 2282 3984
rect 2332 2938 2360 4966
rect 2424 3058 2452 7346
rect 2516 5234 2544 7822
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2608 7002 2636 7754
rect 2700 7546 2728 8978
rect 2780 8900 2832 8906
rect 2780 8842 2832 8848
rect 2792 8566 2820 8842
rect 2780 8560 2832 8566
rect 2780 8502 2832 8508
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2792 7721 2820 8191
rect 2778 7712 2834 7721
rect 2778 7647 2834 7656
rect 2688 7540 2740 7546
rect 2688 7482 2740 7488
rect 2780 7540 2832 7546
rect 2780 7482 2832 7488
rect 2596 6996 2648 7002
rect 2596 6938 2648 6944
rect 2688 6656 2740 6662
rect 2688 6598 2740 6604
rect 2700 6254 2728 6598
rect 2688 6248 2740 6254
rect 2688 6190 2740 6196
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2608 5778 2636 6122
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5846 2728 6054
rect 2688 5840 2740 5846
rect 2688 5782 2740 5788
rect 2596 5772 2648 5778
rect 2596 5714 2648 5720
rect 2792 5273 2820 7482
rect 2884 5370 2912 9930
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 2778 5264 2834 5273
rect 2504 5228 2556 5234
rect 2778 5199 2834 5208
rect 2504 5170 2556 5176
rect 2688 4616 2740 4622
rect 2688 4558 2740 4564
rect 2700 3618 2728 4558
rect 2976 4457 3004 9982
rect 3344 9926 3372 10202
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 3056 9920 3108 9926
rect 3056 9862 3108 9868
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3068 8090 3096 9862
rect 3146 9752 3202 9761
rect 3146 9687 3202 9696
rect 3160 9586 3188 9687
rect 3344 9586 3372 9862
rect 3422 9616 3478 9625
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3332 9580 3384 9586
rect 3422 9551 3478 9560
rect 3332 9522 3384 9528
rect 3148 9376 3200 9382
rect 3148 9318 3200 9324
rect 3160 8974 3188 9318
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3054 7984 3110 7993
rect 3160 7954 3188 8434
rect 3054 7919 3110 7928
rect 3148 7948 3200 7954
rect 3068 5658 3096 7919
rect 3148 7890 3200 7896
rect 3160 7206 3188 7890
rect 3148 7200 3200 7206
rect 3148 7142 3200 7148
rect 3160 6934 3188 7142
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3160 5914 3188 6054
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3068 5630 3188 5658
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3068 5370 3096 5510
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 4480 3108 4486
rect 2962 4448 3018 4457
rect 3056 4422 3108 4428
rect 2962 4383 3018 4392
rect 2872 4140 2924 4146
rect 2872 4082 2924 4088
rect 2700 3602 2820 3618
rect 2700 3596 2832 3602
rect 2700 3590 2780 3596
rect 2780 3538 2832 3544
rect 2780 3460 2832 3466
rect 2780 3402 2832 3408
rect 2686 3224 2742 3233
rect 2792 3194 2820 3402
rect 2686 3159 2688 3168
rect 2740 3159 2742 3168
rect 2780 3188 2832 3194
rect 2688 3130 2740 3136
rect 2780 3130 2832 3136
rect 2778 3088 2834 3097
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 2504 3052 2556 3058
rect 2778 3023 2834 3032
rect 2504 2994 2556 3000
rect 2332 2910 2452 2938
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 2240 2514 2268 2790
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2134 2136 2190 2145
rect 2134 2071 2190 2080
rect 2424 800 2452 2910
rect 2516 2417 2544 2994
rect 2792 2990 2820 3023
rect 2780 2984 2832 2990
rect 2780 2926 2832 2932
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2502 2408 2558 2417
rect 2502 2343 2558 2352
rect 2792 800 2820 2790
rect 2884 1358 2912 4082
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2872 1352 2924 1358
rect 2872 1294 2924 1300
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2778 0 2834 800
rect 2884 649 2912 1294
rect 2870 640 2926 649
rect 2870 575 2926 584
rect 2976 241 3004 4014
rect 3068 3505 3096 4422
rect 3160 4162 3188 5630
rect 3252 4282 3280 8774
rect 3344 7410 3372 9522
rect 3436 8673 3464 9551
rect 3700 9512 3752 9518
rect 3620 9472 3700 9500
rect 3620 9466 3648 9472
rect 3528 9450 3648 9466
rect 3700 9454 3752 9460
rect 3804 9450 3832 10134
rect 3516 9444 3648 9450
rect 3568 9438 3648 9444
rect 3792 9444 3844 9450
rect 3516 9386 3568 9392
rect 3792 9386 3844 9392
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3422 8664 3478 8673
rect 3422 8599 3478 8608
rect 3422 8528 3478 8537
rect 3804 8498 3832 8842
rect 3422 8463 3478 8472
rect 3792 8492 3844 8498
rect 3436 8265 3464 8463
rect 3792 8434 3844 8440
rect 3422 8256 3478 8265
rect 3422 8191 3478 8200
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3422 8120 3478 8129
rect 3549 8112 3857 8132
rect 3422 8055 3478 8064
rect 3436 8022 3464 8055
rect 3424 8016 3476 8022
rect 3424 7958 3476 7964
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3332 6248 3384 6254
rect 3332 6190 3384 6196
rect 3344 5778 3372 6190
rect 3332 5772 3384 5778
rect 3332 5714 3384 5720
rect 3436 5166 3464 6326
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3896 5914 3924 12174
rect 3988 11830 4016 12718
rect 4068 12708 4120 12714
rect 4068 12650 4120 12656
rect 4080 12322 4108 12650
rect 4172 12442 4200 12786
rect 4160 12436 4212 12442
rect 4160 12378 4212 12384
rect 4080 12294 4200 12322
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 4080 11937 4108 12038
rect 4066 11928 4122 11937
rect 4066 11863 4122 11872
rect 3976 11824 4028 11830
rect 3976 11766 4028 11772
rect 4068 11756 4120 11762
rect 4068 11698 4120 11704
rect 4080 11150 4108 11698
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 3976 11076 4028 11082
rect 3976 11018 4028 11024
rect 3988 8838 4016 11018
rect 4066 10976 4122 10985
rect 4066 10911 4122 10920
rect 4080 10198 4108 10911
rect 4172 10810 4200 12294
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4068 10192 4120 10198
rect 4068 10134 4120 10140
rect 4264 10130 4292 11834
rect 4356 10674 4384 12922
rect 4620 12912 4672 12918
rect 4620 12854 4672 12860
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 4448 11082 4476 12582
rect 4632 11898 4660 12854
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4342 10160 4398 10169
rect 4252 10124 4304 10130
rect 4540 10146 4568 11766
rect 4724 11626 4752 15302
rect 4908 14634 4936 15506
rect 5080 14816 5132 14822
rect 5080 14758 5132 14764
rect 4908 14618 5028 14634
rect 4908 14612 5040 14618
rect 4908 14606 4988 14612
rect 4908 14074 4936 14606
rect 4988 14554 5040 14560
rect 5092 14498 5120 14758
rect 5000 14470 5120 14498
rect 5540 14476 5592 14482
rect 4896 14068 4948 14074
rect 4896 14010 4948 14016
rect 4804 13388 4856 13394
rect 4804 13330 4856 13336
rect 4816 12442 4844 13330
rect 4804 12436 4856 12442
rect 4804 12378 4856 12384
rect 4816 12238 4844 12378
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11620 4764 11626
rect 4712 11562 4764 11568
rect 4816 11234 4844 11834
rect 4724 11206 4844 11234
rect 4724 11150 4752 11206
rect 4620 11144 4672 11150
rect 4618 11112 4620 11121
rect 4712 11144 4764 11150
rect 4672 11112 4674 11121
rect 4712 11086 4764 11092
rect 4618 11047 4674 11056
rect 4632 10742 4660 11047
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4620 10736 4672 10742
rect 4620 10678 4672 10684
rect 4342 10095 4398 10104
rect 4448 10118 4568 10146
rect 4252 10066 4304 10072
rect 4068 10056 4120 10062
rect 4066 10024 4068 10033
rect 4120 10024 4122 10033
rect 4066 9959 4122 9968
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 4080 9081 4108 9114
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 3976 8832 4028 8838
rect 4172 8809 4200 9930
rect 4252 9920 4304 9926
rect 4252 9862 4304 9868
rect 3976 8774 4028 8780
rect 4158 8800 4214 8809
rect 4158 8735 4214 8744
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3988 6798 4016 8599
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 4068 7880 4120 7886
rect 4066 7848 4068 7857
rect 4120 7848 4122 7857
rect 4066 7783 4122 7792
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4080 7002 4108 7686
rect 4172 7478 4200 8366
rect 4160 7472 4212 7478
rect 4160 7414 4212 7420
rect 4264 7290 4292 9862
rect 4356 9586 4384 10095
rect 4344 9580 4396 9586
rect 4344 9522 4396 9528
rect 4448 8922 4476 10118
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4172 7262 4292 7290
rect 4356 8894 4476 8922
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3516 5840 3568 5846
rect 4080 5794 4108 6938
rect 3516 5782 3568 5788
rect 3528 5302 3556 5782
rect 3896 5766 4108 5794
rect 3516 5296 3568 5302
rect 3516 5238 3568 5244
rect 3332 5160 3384 5166
rect 3332 5102 3384 5108
rect 3424 5160 3476 5166
rect 3424 5102 3476 5108
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3160 4134 3280 4162
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3160 3738 3188 4014
rect 3148 3732 3200 3738
rect 3148 3674 3200 3680
rect 3054 3496 3110 3505
rect 3054 3431 3110 3440
rect 3148 3460 3200 3466
rect 3148 3402 3200 3408
rect 3160 2553 3188 3402
rect 3146 2544 3202 2553
rect 3146 2479 3202 2488
rect 3252 2446 3280 4134
rect 3344 3670 3372 5102
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3422 3904 3478 3913
rect 3422 3839 3478 3848
rect 3332 3664 3384 3670
rect 3332 3606 3384 3612
rect 3436 3602 3464 3839
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3896 3738 3924 5766
rect 3976 5704 4028 5710
rect 4068 5704 4120 5710
rect 3976 5646 4028 5652
rect 4066 5672 4068 5681
rect 4120 5672 4122 5681
rect 3988 4978 4016 5646
rect 4066 5607 4122 5616
rect 4172 5574 4200 7262
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4160 5568 4212 5574
rect 4160 5510 4212 5516
rect 4264 5386 4292 7142
rect 4356 5914 4384 8894
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 7546 4476 8774
rect 4436 7540 4488 7546
rect 4436 7482 4488 7488
rect 4540 6866 4568 9998
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4632 9382 4660 9862
rect 4724 9518 4752 10746
rect 4804 10736 4856 10742
rect 4804 10678 4856 10684
rect 4816 9761 4844 10678
rect 5000 10266 5028 14470
rect 5540 14418 5592 14424
rect 5552 13530 5580 14418
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5264 13456 5316 13462
rect 5264 13398 5316 13404
rect 5172 13184 5224 13190
rect 5172 13126 5224 13132
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 4896 9920 4948 9926
rect 4896 9862 4948 9868
rect 4802 9752 4858 9761
rect 4908 9722 4936 9862
rect 4802 9687 4858 9696
rect 4896 9716 4948 9722
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4632 7750 4660 9318
rect 4710 9208 4766 9217
rect 4710 9143 4766 9152
rect 4816 9160 4844 9687
rect 4896 9658 4948 9664
rect 5092 9586 5120 10542
rect 5184 10266 5212 13126
rect 5276 11762 5304 13398
rect 5448 13320 5500 13326
rect 5448 13262 5500 13268
rect 5460 12714 5488 13262
rect 5448 12708 5500 12714
rect 5448 12650 5500 12656
rect 5264 11756 5316 11762
rect 5264 11698 5316 11704
rect 5172 10260 5224 10266
rect 5172 10202 5224 10208
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9722 5212 9862
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4528 6860 4580 6866
rect 4528 6802 4580 6808
rect 4436 6656 4488 6662
rect 4632 6644 4660 7686
rect 4488 6616 4660 6644
rect 4436 6598 4488 6604
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4172 5358 4292 5386
rect 3988 4950 4108 4978
rect 3974 4856 4030 4865
rect 3974 4791 3976 4800
rect 4028 4791 4030 4800
rect 3976 4762 4028 4768
rect 3974 4040 4030 4049
rect 4080 4010 4108 4950
rect 3974 3975 3976 3984
rect 4028 3975 4030 3984
rect 4068 4004 4120 4010
rect 3976 3946 4028 3952
rect 4068 3946 4120 3952
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3424 3596 3476 3602
rect 3424 3538 3476 3544
rect 3422 3224 3478 3233
rect 3422 3159 3478 3168
rect 3332 2916 3384 2922
rect 3332 2858 3384 2864
rect 3344 2553 3372 2858
rect 3436 2825 3464 3159
rect 3882 2952 3938 2961
rect 3882 2887 3938 2896
rect 3422 2816 3478 2825
rect 3422 2751 3478 2760
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 3330 2544 3386 2553
rect 3330 2479 3332 2488
rect 3384 2479 3386 2488
rect 3332 2450 3384 2456
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3068 1902 3096 2382
rect 3056 1896 3108 1902
rect 3056 1838 3108 1844
rect 3252 800 3280 2382
rect 3896 1714 3924 2887
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 3712 1686 3924 1714
rect 3712 800 3740 1686
rect 4080 1601 4108 2314
rect 4066 1592 4122 1601
rect 4066 1527 4122 1536
rect 4172 800 4200 5358
rect 4448 4146 4476 6598
rect 4724 5370 4752 9143
rect 4816 9132 4936 9160
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 4816 8634 4844 8978
rect 4804 8628 4856 8634
rect 4804 8570 4856 8576
rect 4816 7342 4844 8570
rect 4908 8566 4936 9132
rect 4988 8900 5040 8906
rect 4988 8842 5040 8848
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 5000 8090 5028 8842
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 5184 7970 5212 9658
rect 5000 7942 5212 7970
rect 4804 7336 4856 7342
rect 4804 7278 4856 7284
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4816 6322 4844 6598
rect 4804 6316 4856 6322
rect 4804 6258 4856 6264
rect 4804 5704 4856 5710
rect 4802 5672 4804 5681
rect 4856 5672 4858 5681
rect 4802 5607 4858 5616
rect 4712 5364 4764 5370
rect 4712 5306 4764 5312
rect 4528 5228 4580 5234
rect 4528 5170 4580 5176
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4540 3670 4568 5170
rect 4724 3924 4752 5306
rect 5000 5234 5028 7942
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5184 7206 5212 7346
rect 5172 7200 5224 7206
rect 5172 7142 5224 7148
rect 5276 7002 5304 11698
rect 5356 11688 5408 11694
rect 5354 11656 5356 11665
rect 5408 11656 5410 11665
rect 5460 11626 5488 12650
rect 5552 12238 5580 13466
rect 5540 12232 5592 12238
rect 5540 12174 5592 12180
rect 5354 11591 5410 11600
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5644 10810 5672 18838
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5736 17746 5764 18226
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5736 17338 5764 17682
rect 5828 17542 5856 18566
rect 5816 17536 5868 17542
rect 5816 17478 5868 17484
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5724 16448 5776 16454
rect 5724 16390 5776 16396
rect 5736 15366 5764 16390
rect 5920 15688 5948 19382
rect 6000 19168 6052 19174
rect 6000 19110 6052 19116
rect 6012 16250 6040 19110
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6564 16454 6592 19858
rect 8220 18970 8248 20470
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8484 19236 8536 19242
rect 8484 19178 8536 19184
rect 8208 18964 8260 18970
rect 8208 18906 8260 18912
rect 6920 18624 6972 18630
rect 6920 18566 6972 18572
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6644 18148 6696 18154
rect 6644 18090 6696 18096
rect 6656 16726 6684 18090
rect 6748 17610 6776 18226
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6840 17882 6868 18158
rect 6828 17876 6880 17882
rect 6828 17818 6880 17824
rect 6932 17814 6960 18566
rect 8208 18216 8260 18222
rect 8208 18158 8260 18164
rect 7012 18080 7064 18086
rect 7012 18022 7064 18028
rect 6920 17808 6972 17814
rect 6920 17750 6972 17756
rect 6920 17672 6972 17678
rect 6920 17614 6972 17620
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6932 17270 6960 17614
rect 6920 17264 6972 17270
rect 6920 17206 6972 17212
rect 6932 16794 6960 17206
rect 7024 17202 7052 18022
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 7012 17196 7064 17202
rect 7012 17138 7064 17144
rect 6920 16788 6972 16794
rect 6920 16730 6972 16736
rect 6644 16720 6696 16726
rect 6644 16662 6696 16668
rect 6552 16448 6604 16454
rect 6552 16390 6604 16396
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 6000 16244 6052 16250
rect 6000 16186 6052 16192
rect 6644 16176 6696 16182
rect 6644 16118 6696 16124
rect 6552 15904 6604 15910
rect 6552 15846 6604 15852
rect 5920 15660 6040 15688
rect 5908 15564 5960 15570
rect 5908 15506 5960 15512
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 14346 5764 15302
rect 5920 15026 5948 15506
rect 5908 15020 5960 15026
rect 5908 14962 5960 14968
rect 5920 14618 5948 14962
rect 6012 14618 6040 15660
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6564 15144 6592 15846
rect 6472 15116 6592 15144
rect 6472 15026 6500 15116
rect 6460 15020 6512 15026
rect 6460 14962 6512 14968
rect 6472 14770 6500 14962
rect 6550 14920 6606 14929
rect 6550 14855 6552 14864
rect 6604 14855 6606 14864
rect 6552 14826 6604 14832
rect 6472 14742 6592 14770
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6000 14612 6052 14618
rect 6000 14554 6052 14560
rect 5724 14340 5776 14346
rect 5724 14282 5776 14288
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 5908 14000 5960 14006
rect 5908 13942 5960 13948
rect 5920 13394 5948 13942
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5908 13388 5960 13394
rect 5908 13330 5960 13336
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11898 5764 12106
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5722 10704 5778 10713
rect 5722 10639 5778 10648
rect 5446 10568 5502 10577
rect 5446 10503 5502 10512
rect 5460 9110 5488 10503
rect 5632 10124 5684 10130
rect 5632 10066 5684 10072
rect 5644 9586 5672 10066
rect 5632 9580 5684 9586
rect 5632 9522 5684 9528
rect 5448 9104 5500 9110
rect 5448 9046 5500 9052
rect 5630 9072 5686 9081
rect 5630 9007 5686 9016
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8362 5488 8910
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5448 8356 5500 8362
rect 5448 8298 5500 8304
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 5460 7546 5488 7686
rect 5448 7540 5500 7546
rect 5368 7500 5448 7528
rect 5264 6996 5316 7002
rect 5264 6938 5316 6944
rect 5368 6882 5396 7500
rect 5448 7482 5500 7488
rect 5552 7002 5580 8502
rect 5644 7313 5672 9007
rect 5736 8537 5764 10639
rect 5722 8528 5778 8537
rect 5722 8463 5778 8472
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5736 8090 5764 8230
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5630 7304 5686 7313
rect 5630 7239 5686 7248
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5540 6996 5592 7002
rect 5540 6938 5592 6944
rect 5092 6854 5396 6882
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4804 4480 4856 4486
rect 4804 4422 4856 4428
rect 4816 4078 4844 4422
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4724 3896 4844 3924
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4448 3126 4476 3402
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4436 2984 4488 2990
rect 4436 2926 4488 2932
rect 4448 1970 4476 2926
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 4540 1057 4568 3470
rect 4712 3188 4764 3194
rect 4632 3148 4712 3176
rect 4526 1048 4582 1057
rect 4526 983 4582 992
rect 4632 800 4660 3148
rect 4712 3130 4764 3136
rect 4712 2984 4764 2990
rect 4712 2926 4764 2932
rect 4724 2514 4752 2926
rect 4816 2514 4844 3896
rect 4908 2990 4936 4082
rect 4896 2984 4948 2990
rect 4896 2926 4948 2932
rect 5092 2938 5120 6854
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5172 6656 5224 6662
rect 5172 6598 5224 6604
rect 5184 4690 5212 6598
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5184 3602 5212 4626
rect 5276 4162 5304 6734
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 5368 4282 5396 6054
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4826 5488 5170
rect 5448 4820 5500 4826
rect 5448 4762 5500 4768
rect 5446 4584 5502 4593
rect 5446 4519 5448 4528
rect 5500 4519 5502 4528
rect 5448 4490 5500 4496
rect 5356 4276 5408 4282
rect 5356 4218 5408 4224
rect 5276 4134 5488 4162
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5184 3058 5212 3538
rect 5276 3058 5304 4014
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5092 2910 5304 2938
rect 4986 2680 5042 2689
rect 4986 2615 5042 2624
rect 4712 2508 4764 2514
rect 4712 2450 4764 2456
rect 4804 2508 4856 2514
rect 4804 2450 4856 2456
rect 5000 800 5028 2615
rect 5276 2582 5304 2910
rect 5264 2576 5316 2582
rect 5264 2518 5316 2524
rect 5460 800 5488 4134
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 5552 3738 5580 4014
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5538 3360 5594 3369
rect 5538 3295 5594 3304
rect 2962 232 3018 241
rect 2962 167 3018 176
rect 3238 0 3294 800
rect 3698 0 3754 800
rect 4158 0 4214 800
rect 4618 0 4674 800
rect 4986 0 5042 800
rect 5446 0 5502 800
rect 5552 762 5580 3295
rect 5644 2774 5672 7142
rect 5736 6662 5764 8026
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5736 3534 5764 6054
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5644 2746 5764 2774
rect 5736 2310 5764 2746
rect 5828 2446 5856 12922
rect 5920 12918 5948 13330
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 5908 12164 5960 12170
rect 5908 12106 5960 12112
rect 5920 9654 5948 12106
rect 6012 12102 6040 13874
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11830 6040 12038
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6564 11098 6592 14742
rect 6656 12434 6684 16118
rect 7300 16046 7328 17614
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7196 16040 7248 16046
rect 7196 15982 7248 15988
rect 7288 16040 7340 16046
rect 7288 15982 7340 15988
rect 7208 15162 7236 15982
rect 7300 15706 7328 15982
rect 7288 15700 7340 15706
rect 7288 15642 7340 15648
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6932 14482 6960 15030
rect 7288 14816 7340 14822
rect 7288 14758 7340 14764
rect 6920 14476 6972 14482
rect 6920 14418 6972 14424
rect 7012 14408 7064 14414
rect 7012 14350 7064 14356
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6656 12406 6776 12434
rect 6644 12232 6696 12238
rect 6644 12174 6696 12180
rect 6656 11830 6684 12174
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6644 11552 6696 11558
rect 6644 11494 6696 11500
rect 6656 11150 6684 11494
rect 6472 11082 6592 11098
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 6460 11076 6592 11082
rect 6512 11070 6592 11076
rect 6460 11018 6512 11024
rect 6000 11008 6052 11014
rect 6000 10950 6052 10956
rect 6552 11008 6604 11014
rect 6552 10950 6604 10956
rect 6012 10130 6040 10950
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6564 10538 6592 10950
rect 6748 10826 6776 12406
rect 6932 12238 6960 14214
rect 7024 13734 7052 14350
rect 7012 13728 7064 13734
rect 7012 13670 7064 13676
rect 7300 13326 7328 14758
rect 7484 14414 7512 17478
rect 7760 16998 7788 17614
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7748 16992 7800 16998
rect 7748 16934 7800 16940
rect 7760 14958 7788 16934
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7852 16250 7880 16594
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7944 15570 7972 17206
rect 8220 16590 8248 18158
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 8312 16590 8340 17138
rect 8208 16584 8260 16590
rect 8208 16526 8260 16532
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8024 15972 8076 15978
rect 8024 15914 8076 15920
rect 8036 15638 8064 15914
rect 8024 15632 8076 15638
rect 8024 15574 8076 15580
rect 7932 15564 7984 15570
rect 7932 15506 7984 15512
rect 7944 15094 7972 15506
rect 7932 15088 7984 15094
rect 7932 15030 7984 15036
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7748 14952 7800 14958
rect 7748 14894 7800 14900
rect 7472 14408 7524 14414
rect 7472 14350 7524 14356
rect 7380 13728 7432 13734
rect 7380 13670 7432 13676
rect 7288 13320 7340 13326
rect 7116 13268 7288 13274
rect 7116 13262 7340 13268
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7116 13246 7328 13262
rect 7024 12918 7052 13194
rect 7012 12912 7064 12918
rect 7012 12854 7064 12860
rect 6920 12232 6972 12238
rect 6920 12174 6972 12180
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11762 6960 12038
rect 6920 11756 6972 11762
rect 6920 11698 6972 11704
rect 6828 11144 6880 11150
rect 6826 11112 6828 11121
rect 6880 11112 6882 11121
rect 6826 11047 6882 11056
rect 6656 10798 6776 10826
rect 6656 10742 6684 10798
rect 6644 10736 6696 10742
rect 6644 10678 6696 10684
rect 6552 10532 6604 10538
rect 6552 10474 6604 10480
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 6092 10056 6144 10062
rect 6012 10004 6092 10010
rect 6012 9998 6144 10004
rect 6012 9982 6132 9998
rect 5908 9648 5960 9654
rect 5908 9590 5960 9596
rect 5908 9376 5960 9382
rect 6012 9364 6040 9982
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6184 9580 6236 9586
rect 6184 9522 6236 9528
rect 5960 9336 6040 9364
rect 5908 9318 5960 9324
rect 5920 6440 5948 9318
rect 6196 9217 6224 9522
rect 6274 9344 6330 9353
rect 6274 9279 6330 9288
rect 6182 9208 6238 9217
rect 6182 9143 6238 9152
rect 6288 9042 6316 9279
rect 6276 9036 6328 9042
rect 6276 8978 6328 8984
rect 6000 8832 6052 8838
rect 6000 8774 6052 8780
rect 6012 7546 6040 8774
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 6564 6440 6592 8026
rect 6656 7886 6684 10678
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6748 9110 6776 10610
rect 6840 10130 6868 11047
rect 6828 10124 6880 10130
rect 6828 10066 6880 10072
rect 6736 9104 6788 9110
rect 6736 9046 6788 9052
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6734 8664 6790 8673
rect 6734 8599 6790 8608
rect 6748 8022 6776 8599
rect 6826 8528 6882 8537
rect 6932 8498 6960 8774
rect 6826 8463 6882 8472
rect 6920 8492 6972 8498
rect 6736 8016 6788 8022
rect 6736 7958 6788 7964
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6656 7546 6684 7822
rect 6644 7540 6696 7546
rect 6644 7482 6696 7488
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6736 7336 6788 7342
rect 6736 7278 6788 7284
rect 5920 6412 6132 6440
rect 6000 6248 6052 6254
rect 6000 6190 6052 6196
rect 6012 5914 6040 6190
rect 6000 5908 6052 5914
rect 6000 5850 6052 5856
rect 5908 5840 5960 5846
rect 6104 5794 6132 6412
rect 6472 6412 6592 6440
rect 6366 6352 6422 6361
rect 6366 6287 6368 6296
rect 6420 6287 6422 6296
rect 6368 6258 6420 6264
rect 6472 6118 6500 6412
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6460 6112 6512 6118
rect 6460 6054 6512 6060
rect 5908 5782 5960 5788
rect 5920 5098 5948 5782
rect 6012 5766 6132 5794
rect 5908 5092 5960 5098
rect 5908 5034 5960 5040
rect 6012 4978 6040 5766
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 6564 5098 6592 6258
rect 6552 5092 6604 5098
rect 6552 5034 6604 5040
rect 5920 4950 6040 4978
rect 5920 4078 5948 4950
rect 6148 4380 6456 4400
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 6000 4276 6052 4282
rect 6000 4218 6052 4224
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 6012 3641 6040 4218
rect 6564 4146 6592 5034
rect 6656 4706 6684 7278
rect 6748 6934 6776 7278
rect 6736 6928 6788 6934
rect 6840 6905 6868 8463
rect 6920 8434 6972 8440
rect 6932 7954 6960 8434
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7342 6960 7890
rect 7024 7886 7052 12854
rect 7116 12434 7144 13246
rect 7116 12406 7236 12434
rect 7104 12164 7156 12170
rect 7104 12106 7156 12112
rect 7116 10810 7144 12106
rect 7208 11354 7236 12406
rect 7286 12200 7342 12209
rect 7286 12135 7342 12144
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 7104 10804 7156 10810
rect 7104 10746 7156 10752
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7208 9382 7236 10542
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7300 8401 7328 12135
rect 7392 11694 7420 13670
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7472 12640 7524 12646
rect 7472 12582 7524 12588
rect 7484 11898 7512 12582
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7576 11762 7604 13126
rect 7564 11756 7616 11762
rect 7564 11698 7616 11704
rect 7380 11688 7432 11694
rect 7380 11630 7432 11636
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7392 8566 7420 9454
rect 7576 9450 7604 9590
rect 7564 9444 7616 9450
rect 7564 9386 7616 9392
rect 7380 8560 7432 8566
rect 7380 8502 7432 8508
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7472 7948 7524 7954
rect 7472 7890 7524 7896
rect 7012 7880 7064 7886
rect 7484 7857 7512 7890
rect 7012 7822 7064 7828
rect 7470 7848 7526 7857
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6736 6870 6788 6876
rect 6826 6896 6882 6905
rect 6826 6831 6882 6840
rect 7024 6798 7052 7822
rect 7470 7783 7526 7792
rect 7104 7744 7156 7750
rect 7104 7686 7156 7692
rect 7564 7744 7616 7750
rect 7564 7686 7616 7692
rect 7116 7546 7144 7686
rect 7104 7540 7156 7546
rect 7104 7482 7156 7488
rect 7196 7472 7248 7478
rect 7196 7414 7248 7420
rect 7104 7268 7156 7274
rect 7104 7210 7156 7216
rect 6736 6792 6788 6798
rect 6736 6734 6788 6740
rect 7012 6792 7064 6798
rect 7012 6734 7064 6740
rect 6748 6390 6776 6734
rect 6918 6488 6974 6497
rect 6918 6423 6974 6432
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6932 6225 6960 6423
rect 6918 6216 6974 6225
rect 6918 6151 6974 6160
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6932 5658 6960 5850
rect 7024 5710 7052 6734
rect 6840 5630 6960 5658
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 6840 5574 6868 5630
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6656 4678 6868 4706
rect 6644 4548 6696 4554
rect 6644 4490 6696 4496
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6460 4072 6512 4078
rect 6460 4014 6512 4020
rect 5998 3632 6054 3641
rect 5998 3567 6054 3576
rect 6472 3516 6500 4014
rect 6552 4004 6604 4010
rect 6552 3946 6604 3952
rect 6564 3670 6592 3946
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6472 3488 6592 3516
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 6564 2854 6592 3488
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6656 2582 6684 4490
rect 6840 4078 6868 4678
rect 6932 4146 6960 5510
rect 7116 4282 7144 7210
rect 7208 6730 7236 7414
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 7196 6724 7248 6730
rect 7196 6666 7248 6672
rect 7392 6458 7420 7142
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7380 6452 7432 6458
rect 7380 6394 7432 6400
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6840 3398 6868 4014
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7012 3664 7064 3670
rect 7012 3606 7064 3612
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6826 3224 6882 3233
rect 6826 3159 6882 3168
rect 6644 2576 6696 2582
rect 6644 2518 6696 2524
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 6366 1864 6422 1873
rect 6366 1799 6422 1808
rect 5828 870 5948 898
rect 5828 762 5856 870
rect 5920 800 5948 870
rect 6380 800 6408 1799
rect 6840 800 6868 3159
rect 7024 1902 7052 3606
rect 7116 2990 7144 3674
rect 7196 3392 7248 3398
rect 7196 3334 7248 3340
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7116 2514 7144 2926
rect 7208 2650 7236 3334
rect 7300 3194 7328 6258
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 4010 7420 5510
rect 7484 4214 7512 6598
rect 7472 4208 7524 4214
rect 7472 4150 7524 4156
rect 7380 4004 7432 4010
rect 7380 3946 7432 3952
rect 7472 3664 7524 3670
rect 7472 3606 7524 3612
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7288 3188 7340 3194
rect 7288 3130 7340 3136
rect 7392 2774 7420 3334
rect 7300 2746 7420 2774
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7300 2530 7328 2746
rect 7104 2508 7156 2514
rect 7104 2450 7156 2456
rect 7208 2502 7328 2530
rect 7484 2530 7512 3606
rect 7576 2650 7604 7686
rect 7668 5914 7696 14894
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 13938 8064 14214
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8036 13394 8064 13874
rect 8024 13388 8076 13394
rect 8024 13330 8076 13336
rect 7748 12776 7800 12782
rect 7748 12718 7800 12724
rect 7760 12306 7788 12718
rect 8036 12714 8064 13330
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8220 12889 8248 13126
rect 8206 12880 8262 12889
rect 8206 12815 8262 12824
rect 8024 12708 8076 12714
rect 8024 12650 8076 12656
rect 7838 12336 7894 12345
rect 7748 12300 7800 12306
rect 7838 12271 7894 12280
rect 7748 12242 7800 12248
rect 7760 12102 7788 12242
rect 7852 12238 7880 12271
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 8024 12096 8076 12102
rect 8024 12038 8076 12044
rect 8036 11218 8064 12038
rect 8496 11354 8524 19178
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8588 15502 8616 17478
rect 8576 15496 8628 15502
rect 8576 15438 8628 15444
rect 8680 15162 8708 20402
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 9680 19372 9732 19378
rect 9680 19314 9732 19320
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 9692 18426 9720 19314
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 10692 18760 10744 18766
rect 10692 18702 10744 18708
rect 10704 18426 10732 18702
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 10692 18420 10744 18426
rect 10692 18362 10744 18368
rect 11704 18284 11756 18290
rect 11704 18226 11756 18232
rect 10140 18216 10192 18222
rect 10140 18158 10192 18164
rect 11060 18216 11112 18222
rect 11060 18158 11112 18164
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 9404 17740 9456 17746
rect 9404 17682 9456 17688
rect 9416 17338 9444 17682
rect 9508 17610 9536 18022
rect 10152 17882 10180 18158
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 11072 17678 11100 18158
rect 11060 17672 11112 17678
rect 11112 17632 11192 17660
rect 11060 17614 11112 17620
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 9404 16652 9456 16658
rect 9404 16594 9456 16600
rect 9312 16448 9364 16454
rect 9312 16390 9364 16396
rect 9324 16250 9352 16390
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9312 16108 9364 16114
rect 9416 16096 9444 16594
rect 9364 16068 9444 16096
rect 9312 16050 9364 16056
rect 9220 16040 9272 16046
rect 9220 15982 9272 15988
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 9232 15502 9260 15982
rect 9324 15706 9352 16050
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8668 15156 8720 15162
rect 8668 15098 8720 15104
rect 9220 14952 9272 14958
rect 9220 14894 9272 14900
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 8760 14544 8812 14550
rect 8760 14486 8812 14492
rect 8772 14074 8800 14486
rect 9232 14074 9260 14894
rect 9312 14340 9364 14346
rect 9312 14282 9364 14288
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8760 14068 8812 14074
rect 8760 14010 8812 14016
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8588 13394 8616 13942
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8680 13297 8708 14010
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 8760 13320 8812 13326
rect 8666 13288 8722 13297
rect 8760 13262 8812 13268
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8666 13223 8722 13232
rect 8772 12730 8800 13262
rect 8680 12702 8800 12730
rect 8680 12170 8708 12702
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 9036 12368 9088 12374
rect 9036 12310 9088 12316
rect 8668 12164 8720 12170
rect 8668 12106 8720 12112
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7748 10668 7800 10674
rect 7748 10610 7800 10616
rect 7760 8090 7788 10610
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7852 6746 7880 9862
rect 7944 7313 7972 10406
rect 8036 9518 8064 11154
rect 8208 11076 8260 11082
rect 8208 11018 8260 11024
rect 8220 10810 8248 11018
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8208 10804 8260 10810
rect 8208 10746 8260 10752
rect 8404 10606 8432 10950
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8312 10062 8340 10406
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8392 9920 8444 9926
rect 8496 9908 8524 10474
rect 8588 10062 8616 12038
rect 8680 11286 8708 12106
rect 9048 11626 9076 12310
rect 9036 11620 9088 11626
rect 9036 11562 9088 11568
rect 9140 11558 9168 13262
rect 9232 12646 9260 13738
rect 9220 12640 9272 12646
rect 9220 12582 9272 12588
rect 9232 12481 9260 12582
rect 9218 12472 9274 12481
rect 9218 12407 9274 12416
rect 9232 12374 9260 12407
rect 9220 12368 9272 12374
rect 9220 12310 9272 12316
rect 9324 12102 9352 14282
rect 9508 12434 9536 17546
rect 9772 17536 9824 17542
rect 9772 17478 9824 17484
rect 9784 17202 9812 17478
rect 11060 17264 11112 17270
rect 11060 17206 11112 17212
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 11072 16658 11100 17206
rect 11164 17066 11192 17632
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11060 16652 11112 16658
rect 11060 16594 11112 16600
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10428 15162 10456 15982
rect 10968 15496 11020 15502
rect 11072 15450 11100 16594
rect 11152 16584 11204 16590
rect 11204 16544 11284 16572
rect 11152 16526 11204 16532
rect 11152 16448 11204 16454
rect 11152 16390 11204 16396
rect 11164 16250 11192 16390
rect 11152 16244 11204 16250
rect 11152 16186 11204 16192
rect 11152 16108 11204 16114
rect 11152 16050 11204 16056
rect 11164 15910 11192 16050
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11020 15444 11100 15450
rect 10968 15438 11100 15444
rect 10784 15428 10836 15434
rect 10980 15422 11100 15438
rect 10784 15370 10836 15376
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10796 14822 10824 15370
rect 11072 15026 11100 15422
rect 11164 15162 11192 15846
rect 11152 15156 11204 15162
rect 11152 15098 11204 15104
rect 10876 15020 10928 15026
rect 10876 14962 10928 14968
rect 11060 15020 11112 15026
rect 11060 14962 11112 14968
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10888 14618 10916 14962
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 11072 14414 11100 14962
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 9588 14340 9640 14346
rect 9588 14282 9640 14288
rect 9600 13870 9628 14282
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 9864 13932 9916 13938
rect 9864 13874 9916 13880
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9678 13424 9734 13433
rect 9678 13359 9734 13368
rect 9692 13326 9720 13359
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9416 12406 9536 12434
rect 9312 12096 9364 12102
rect 9312 12038 9364 12044
rect 9416 11778 9444 12406
rect 9588 12300 9640 12306
rect 9588 12242 9640 12248
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9232 11750 9444 11778
rect 9128 11552 9180 11558
rect 9128 11494 9180 11500
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 8668 11280 8720 11286
rect 9036 11280 9088 11286
rect 8668 11222 8720 11228
rect 8864 11240 9036 11268
rect 8864 11150 8892 11240
rect 9036 11222 9088 11228
rect 8852 11144 8904 11150
rect 8852 11086 8904 11092
rect 9140 10606 9168 11494
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 9128 10600 9180 10606
rect 9128 10542 9180 10548
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8444 9880 8524 9908
rect 8392 9862 8444 9868
rect 8024 9512 8076 9518
rect 8024 9454 8076 9460
rect 8116 9444 8168 9450
rect 8116 9386 8168 9392
rect 8128 9353 8156 9386
rect 8114 9344 8170 9353
rect 8114 9279 8170 9288
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8116 8900 8168 8906
rect 8116 8842 8168 8848
rect 8022 8664 8078 8673
rect 8128 8634 8156 8842
rect 8022 8599 8078 8608
rect 8116 8628 8168 8634
rect 8036 8566 8064 8599
rect 8116 8570 8168 8576
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 7930 7304 7986 7313
rect 7930 7239 7986 7248
rect 8024 7200 8076 7206
rect 8024 7142 8076 7148
rect 7852 6718 7972 6746
rect 7840 6656 7892 6662
rect 7840 6598 7892 6604
rect 7852 6390 7880 6598
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7852 5778 7880 6054
rect 7840 5772 7892 5778
rect 7840 5714 7892 5720
rect 7654 5264 7710 5273
rect 7654 5199 7710 5208
rect 7668 3670 7696 5199
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7852 3058 7880 5714
rect 7944 4622 7972 6718
rect 8036 6254 8064 7142
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 8024 6248 8076 6254
rect 8024 6190 8076 6196
rect 8036 5234 8064 6190
rect 8128 5370 8156 6666
rect 8220 6644 8248 8434
rect 8404 8430 8432 8910
rect 8496 8498 8524 9880
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8588 8906 8616 9862
rect 8680 9722 8708 10542
rect 9232 10418 9260 11750
rect 9312 11688 9364 11694
rect 9312 11630 9364 11636
rect 9140 10390 9260 10418
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 8944 10192 8996 10198
rect 8944 10134 8996 10140
rect 8852 10056 8904 10062
rect 8852 9998 8904 10004
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8772 9722 8800 9930
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8760 9716 8812 9722
rect 8760 9658 8812 9664
rect 8668 9580 8720 9586
rect 8864 9568 8892 9998
rect 8720 9540 8892 9568
rect 8668 9522 8720 9528
rect 8680 9042 8708 9522
rect 8956 9518 8984 10134
rect 8944 9512 8996 9518
rect 8772 9460 8944 9466
rect 8772 9454 8996 9460
rect 8772 9450 8984 9454
rect 8760 9444 8984 9450
rect 8812 9438 8984 9444
rect 8760 9386 8812 9392
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 9140 9160 9168 10390
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9048 9132 9168 9160
rect 8668 9036 8720 9042
rect 8668 8978 8720 8984
rect 8576 8900 8628 8906
rect 8576 8842 8628 8848
rect 8944 8832 8996 8838
rect 8944 8774 8996 8780
rect 8956 8634 8984 8774
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8392 8424 8444 8430
rect 9048 8401 9076 9132
rect 9128 8832 9180 8838
rect 9128 8774 9180 8780
rect 8392 8366 8444 8372
rect 8574 8392 8630 8401
rect 8404 7886 8432 8366
rect 8574 8327 8630 8336
rect 9034 8392 9090 8401
rect 9034 8327 9090 8336
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7002 8432 7686
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8392 6996 8444 7002
rect 8392 6938 8444 6944
rect 8300 6928 8352 6934
rect 8352 6876 8432 6882
rect 8300 6870 8432 6876
rect 8312 6854 8432 6870
rect 8300 6656 8352 6662
rect 8220 6616 8300 6644
rect 8300 6598 8352 6604
rect 8208 6452 8260 6458
rect 8208 6394 8260 6400
rect 8220 5778 8248 6394
rect 8208 5772 8260 5778
rect 8208 5714 8260 5720
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8116 5364 8168 5370
rect 8116 5306 8168 5312
rect 8024 5228 8076 5234
rect 8024 5170 8076 5176
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 7932 4616 7984 4622
rect 7984 4576 8064 4604
rect 7932 4558 7984 4564
rect 7932 4480 7984 4486
rect 7932 4422 7984 4428
rect 7944 3534 7972 4422
rect 8036 4146 8064 4576
rect 8220 4486 8248 5034
rect 8312 5030 8340 5646
rect 8404 5166 8432 6854
rect 8496 6225 8524 7482
rect 8588 6934 8616 8327
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8956 7274 8984 7822
rect 9140 7546 9168 8774
rect 9232 8566 9260 9862
rect 9324 9568 9352 11630
rect 9508 11150 9536 12038
rect 9496 11144 9548 11150
rect 9496 11086 9548 11092
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9416 10810 9444 11018
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9600 10656 9628 12242
rect 9692 11830 9720 13126
rect 9876 12986 9904 13874
rect 10336 13870 10364 14214
rect 11072 14090 11100 14350
rect 11256 14278 11284 16544
rect 11716 16454 11744 18226
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 15752 17808 15804 17814
rect 15752 17750 15804 17756
rect 12900 17672 12952 17678
rect 12530 17640 12586 17649
rect 12900 17614 12952 17620
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 12530 17575 12532 17584
rect 12584 17575 12586 17584
rect 12532 17546 12584 17552
rect 11796 17536 11848 17542
rect 11796 17478 11848 17484
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11808 17202 11836 17478
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11992 16590 12020 17478
rect 12912 16998 12940 17614
rect 12900 16992 12952 16998
rect 12900 16934 12952 16940
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11704 16448 11756 16454
rect 11704 16390 11756 16396
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 12912 16046 12940 16934
rect 13280 16794 13308 17614
rect 13544 17536 13596 17542
rect 13544 17478 13596 17484
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13556 16590 13584 17478
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 13544 16584 13596 16590
rect 13544 16526 13596 16532
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 12900 16040 12952 16046
rect 12900 15982 12952 15988
rect 11704 15700 11756 15706
rect 11704 15642 11756 15648
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11716 14482 11744 15642
rect 11796 15088 11848 15094
rect 11796 15030 11848 15036
rect 11704 14476 11756 14482
rect 11704 14418 11756 14424
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11072 14062 11284 14090
rect 10692 13932 10744 13938
rect 10692 13874 10744 13880
rect 10324 13864 10376 13870
rect 10324 13806 10376 13812
rect 9956 13796 10008 13802
rect 9956 13738 10008 13744
rect 9968 13530 9996 13738
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 10244 12918 10272 13398
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10416 12776 10468 12782
rect 10416 12718 10468 12724
rect 10428 12442 10456 12718
rect 10416 12436 10468 12442
rect 10416 12378 10468 12384
rect 10416 12232 10468 12238
rect 10416 12174 10468 12180
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9508 10628 9628 10656
rect 9680 10668 9732 10674
rect 9324 9540 9444 9568
rect 9312 9444 9364 9450
rect 9312 9386 9364 9392
rect 9324 9178 9352 9386
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9312 7812 9364 7818
rect 9312 7754 9364 7760
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9324 7410 9352 7754
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8944 7268 8996 7274
rect 8944 7210 8996 7216
rect 8747 7100 9055 7120
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 9416 6984 9444 9540
rect 9508 8634 9536 10628
rect 9680 10610 9732 10616
rect 9588 10532 9640 10538
rect 9588 10474 9640 10480
rect 9600 10198 9628 10474
rect 9588 10192 9640 10198
rect 9588 10134 9640 10140
rect 9692 9654 9720 10610
rect 10048 9988 10100 9994
rect 10048 9930 10100 9936
rect 9864 9920 9916 9926
rect 9864 9862 9916 9868
rect 9680 9648 9732 9654
rect 9680 9590 9732 9596
rect 9588 9580 9640 9586
rect 9588 9522 9640 9528
rect 9600 9042 9628 9522
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9496 8628 9548 8634
rect 9496 8570 9548 8576
rect 9496 8424 9548 8430
rect 9494 8392 9496 8401
rect 9548 8392 9550 8401
rect 9494 8327 9550 8336
rect 9586 7984 9642 7993
rect 9586 7919 9642 7928
rect 9496 7404 9548 7410
rect 9496 7346 9548 7352
rect 9232 6956 9444 6984
rect 8576 6928 8628 6934
rect 8576 6870 8628 6876
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8482 6216 8538 6225
rect 8482 6151 8538 6160
rect 8496 5234 8524 6151
rect 8680 6118 8708 6802
rect 9128 6316 9180 6322
rect 9128 6258 9180 6264
rect 8668 6112 8720 6118
rect 8668 6054 8720 6060
rect 8747 6012 9055 6032
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8484 5228 8536 5234
rect 8484 5170 8536 5176
rect 8392 5160 8444 5166
rect 8392 5102 8444 5108
rect 8576 5160 8628 5166
rect 8576 5102 8628 5108
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8588 4690 8616 5102
rect 8576 4684 8628 4690
rect 8576 4626 8628 4632
rect 8208 4480 8260 4486
rect 8208 4422 8260 4428
rect 8220 4282 8248 4422
rect 8208 4276 8260 4282
rect 8208 4218 8260 4224
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 8114 4040 8170 4049
rect 8114 3975 8170 3984
rect 8576 4004 8628 4010
rect 8024 3596 8076 3602
rect 8024 3538 8076 3544
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8036 3126 8064 3538
rect 8024 3120 8076 3126
rect 8024 3062 8076 3068
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 2650 8064 2790
rect 7564 2644 7616 2650
rect 7564 2586 7616 2592
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7484 2502 7696 2530
rect 7012 1896 7064 1902
rect 7012 1838 7064 1844
rect 7208 800 7236 2502
rect 7288 2304 7340 2310
rect 7288 2246 7340 2252
rect 7300 1766 7328 2246
rect 7288 1760 7340 1766
rect 7288 1702 7340 1708
rect 7668 800 7696 2502
rect 8128 800 8156 3975
rect 8576 3946 8628 3952
rect 8300 3936 8352 3942
rect 8300 3878 8352 3884
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8220 2038 8248 2518
rect 8312 2446 8340 3878
rect 8496 3602 8524 3878
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 8588 3482 8616 3946
rect 8404 3454 8616 3482
rect 8404 2530 8432 3454
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8404 2502 8524 2530
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8404 1630 8432 2382
rect 8496 1986 8524 2502
rect 8588 2106 8616 3334
rect 8680 2446 8708 5510
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9048 5137 9076 5170
rect 9034 5128 9090 5137
rect 9034 5063 9090 5072
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 9140 4690 9168 6258
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9232 4282 9260 6956
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 9220 3528 9272 3534
rect 9220 3470 9272 3476
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 9140 2564 9168 2994
rect 9048 2536 9168 2564
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8576 2100 8628 2106
rect 8576 2042 8628 2048
rect 8496 1958 8616 1986
rect 8392 1624 8444 1630
rect 8392 1566 8444 1572
rect 8588 800 8616 1958
rect 9048 800 9076 2536
rect 9232 1698 9260 3470
rect 9324 2514 9352 6802
rect 9404 6656 9456 6662
rect 9404 6598 9456 6604
rect 9416 5370 9444 6598
rect 9508 6254 9536 7346
rect 9496 6248 9548 6254
rect 9496 6190 9548 6196
rect 9508 5370 9536 6190
rect 9404 5364 9456 5370
rect 9404 5306 9456 5312
rect 9496 5364 9548 5370
rect 9496 5306 9548 5312
rect 9496 4480 9548 4486
rect 9496 4422 9548 4428
rect 9508 3058 9536 4422
rect 9496 3052 9548 3058
rect 9496 2994 9548 3000
rect 9600 2774 9628 7919
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9678 7032 9734 7041
rect 9678 6967 9734 6976
rect 9692 6610 9720 6967
rect 9784 6730 9812 7278
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9692 6582 9812 6610
rect 9680 6452 9732 6458
rect 9680 6394 9732 6400
rect 9692 5778 9720 6394
rect 9680 5772 9732 5778
rect 9680 5714 9732 5720
rect 9680 5568 9732 5574
rect 9680 5510 9732 5516
rect 9692 4865 9720 5510
rect 9678 4856 9734 4865
rect 9678 4791 9734 4800
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9692 3058 9720 4014
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9692 2825 9720 2994
rect 9416 2746 9628 2774
rect 9678 2816 9734 2825
rect 9678 2751 9734 2760
rect 9784 2774 9812 6582
rect 9876 4622 9904 9862
rect 10060 9518 10088 9930
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 9110 10088 9454
rect 10048 9104 10100 9110
rect 9968 9052 10048 9058
rect 9968 9046 10100 9052
rect 9968 9030 10088 9046
rect 9968 8430 9996 9030
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10138 8936 10194 8945
rect 9956 8424 10008 8430
rect 9956 8366 10008 8372
rect 9956 7268 10008 7274
rect 9956 7210 10008 7216
rect 9968 6798 9996 7210
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10060 6458 10088 8910
rect 10138 8871 10140 8880
rect 10192 8871 10194 8880
rect 10140 8842 10192 8848
rect 10244 8838 10272 12038
rect 10428 11150 10456 12174
rect 10600 11756 10652 11762
rect 10600 11698 10652 11704
rect 10612 11354 10640 11698
rect 10600 11348 10652 11354
rect 10600 11290 10652 11296
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10612 9110 10640 9454
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10232 8832 10284 8838
rect 10232 8774 10284 8780
rect 10324 8492 10376 8498
rect 10324 8434 10376 8440
rect 10336 7750 10364 8434
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10152 7274 10180 7686
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10140 6180 10192 6186
rect 10140 6122 10192 6128
rect 9956 5840 10008 5846
rect 9956 5782 10008 5788
rect 9968 5574 9996 5782
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9864 4616 9916 4622
rect 9864 4558 9916 4564
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 9864 4208 9916 4214
rect 9862 4176 9864 4185
rect 9916 4176 9918 4185
rect 9862 4111 9918 4120
rect 9864 4072 9916 4078
rect 9864 4014 9916 4020
rect 9876 3194 9904 4014
rect 9864 3188 9916 3194
rect 9864 3130 9916 3136
rect 9312 2508 9364 2514
rect 9312 2450 9364 2456
rect 9220 1692 9272 1698
rect 9220 1634 9272 1640
rect 9416 800 9444 2746
rect 9692 2582 9720 2751
rect 9784 2746 9904 2774
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9692 1834 9720 2382
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9680 1828 9732 1834
rect 9680 1770 9732 1776
rect 9784 1766 9812 2246
rect 9772 1760 9824 1766
rect 9772 1702 9824 1708
rect 9876 800 9904 2746
rect 9968 2446 9996 4490
rect 10060 3505 10088 5170
rect 10152 4826 10180 6122
rect 10230 5672 10286 5681
rect 10230 5607 10286 5616
rect 10140 4820 10192 4826
rect 10140 4762 10192 4768
rect 10140 4208 10192 4214
rect 10140 4150 10192 4156
rect 10046 3496 10102 3505
rect 10046 3431 10102 3440
rect 10060 3194 10088 3431
rect 10048 3188 10100 3194
rect 10048 3130 10100 3136
rect 10152 2650 10180 4150
rect 10244 3398 10272 5607
rect 10336 4690 10364 7686
rect 10324 4684 10376 4690
rect 10324 4626 10376 4632
rect 10324 4548 10376 4554
rect 10324 4490 10376 4496
rect 10336 4282 10364 4490
rect 10428 4486 10456 8842
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10612 6866 10640 7822
rect 10600 6860 10652 6866
rect 10600 6802 10652 6808
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10324 4276 10376 4282
rect 10324 4218 10376 4224
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10416 4208 10468 4214
rect 10414 4176 10416 4185
rect 10468 4176 10470 4185
rect 10324 4140 10376 4146
rect 10414 4111 10470 4120
rect 10324 4082 10376 4088
rect 10336 3398 10364 4082
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10232 3392 10284 3398
rect 10232 3334 10284 3340
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 9956 2440 10008 2446
rect 9956 2382 10008 2388
rect 10140 2304 10192 2310
rect 10140 2246 10192 2252
rect 10152 1698 10180 2246
rect 10140 1692 10192 1698
rect 10140 1634 10192 1640
rect 10336 800 10364 3334
rect 10428 2650 10456 3946
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10520 2446 10548 4218
rect 10612 3890 10640 5850
rect 10704 4010 10732 13874
rect 11256 13326 11284 14062
rect 11244 13320 11296 13326
rect 11244 13262 11296 13268
rect 11058 12472 11114 12481
rect 11256 12458 11284 13262
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11520 12640 11572 12646
rect 11518 12608 11520 12617
rect 11572 12608 11574 12617
rect 11518 12543 11574 12552
rect 11114 12430 11284 12458
rect 11808 12434 11836 15030
rect 11992 13870 12020 15982
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 12440 15360 12492 15366
rect 12440 15302 12492 15308
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 11980 13864 12032 13870
rect 11980 13806 12032 13812
rect 12268 13530 12296 14282
rect 12256 13524 12308 13530
rect 12256 13466 12308 13472
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 12084 12442 12112 13194
rect 12072 12436 12124 12442
rect 11058 12407 11114 12416
rect 11072 12238 11100 12407
rect 11808 12406 11928 12434
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 10784 11552 10836 11558
rect 10784 11494 10836 11500
rect 11060 11552 11112 11558
rect 11060 11494 11112 11500
rect 10796 11218 10824 11494
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10784 9512 10836 9518
rect 11072 9466 11100 11494
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11336 10464 11388 10470
rect 11336 10406 11388 10412
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9586 11192 9998
rect 11256 9654 11284 10202
rect 11348 9994 11376 10406
rect 11716 10010 11744 10542
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11808 10198 11836 10406
rect 11796 10192 11848 10198
rect 11796 10134 11848 10140
rect 11336 9988 11388 9994
rect 11716 9982 11836 10010
rect 11336 9930 11388 9936
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11808 9674 11836 9982
rect 11244 9648 11296 9654
rect 11244 9590 11296 9596
rect 11716 9646 11836 9674
rect 11152 9580 11204 9586
rect 11152 9522 11204 9528
rect 10784 9454 10836 9460
rect 10796 6662 10824 9454
rect 10888 9438 11100 9466
rect 10888 7721 10916 9438
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 11072 8838 11100 9318
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10968 8356 11020 8362
rect 10968 8298 11020 8304
rect 10874 7712 10930 7721
rect 10874 7647 10930 7656
rect 10784 6656 10836 6662
rect 10784 6598 10836 6604
rect 10980 5302 11008 8298
rect 11072 7954 11100 8434
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7410 11100 7686
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11060 7200 11112 7206
rect 11060 7142 11112 7148
rect 10968 5296 11020 5302
rect 10968 5238 11020 5244
rect 11072 4554 11100 7142
rect 11164 5234 11192 9522
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11244 8424 11296 8430
rect 11244 8366 11296 8372
rect 11256 7546 11284 8366
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 11244 7540 11296 7546
rect 11244 7482 11296 7488
rect 11428 7404 11480 7410
rect 11428 7346 11480 7352
rect 11334 7304 11390 7313
rect 11334 7239 11390 7248
rect 11348 6798 11376 7239
rect 11440 6934 11468 7346
rect 11428 6928 11480 6934
rect 11428 6870 11480 6876
rect 11336 6792 11388 6798
rect 11336 6734 11388 6740
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11152 5228 11204 5234
rect 11152 5170 11204 5176
rect 11164 4622 11192 5170
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11060 4548 11112 4554
rect 11060 4490 11112 4496
rect 10782 4176 10838 4185
rect 10782 4111 10838 4120
rect 10692 4004 10744 4010
rect 10692 3946 10744 3952
rect 10612 3862 10732 3890
rect 10600 3460 10652 3466
rect 10600 3402 10652 3408
rect 10508 2440 10560 2446
rect 10612 2417 10640 3402
rect 10508 2382 10560 2388
rect 10598 2408 10654 2417
rect 10598 2343 10654 2352
rect 10704 1766 10732 3862
rect 10692 1760 10744 1766
rect 10692 1702 10744 1708
rect 10796 800 10824 4111
rect 10874 4040 10930 4049
rect 10874 3975 10930 3984
rect 11058 4040 11114 4049
rect 11058 3975 11114 3984
rect 10888 3777 10916 3975
rect 10874 3768 10930 3777
rect 10874 3703 10930 3712
rect 11072 3670 11100 3975
rect 11164 3738 11192 4558
rect 11152 3732 11204 3738
rect 11152 3674 11204 3680
rect 11060 3664 11112 3670
rect 11060 3606 11112 3612
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 11060 3528 11112 3534
rect 11060 3470 11112 3476
rect 10888 2650 10916 3470
rect 11072 2854 11100 3470
rect 11164 2990 11192 3674
rect 11256 3602 11284 6598
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 11716 5642 11744 9646
rect 11900 9382 11928 12406
rect 12072 12378 12124 12384
rect 12164 12164 12216 12170
rect 12164 12106 12216 12112
rect 12176 11898 12204 12106
rect 12452 11898 12480 15302
rect 12714 14920 12770 14929
rect 12714 14855 12770 14864
rect 12622 12200 12678 12209
rect 12622 12135 12678 12144
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12636 11762 12664 12135
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12164 11144 12216 11150
rect 12164 11086 12216 11092
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 11978 10160 12034 10169
rect 11978 10095 12034 10104
rect 11992 9926 12020 10095
rect 11980 9920 12032 9926
rect 11980 9862 12032 9868
rect 11796 9376 11848 9382
rect 11796 9318 11848 9324
rect 11888 9376 11940 9382
rect 11888 9318 11940 9324
rect 11808 8838 11836 9318
rect 11796 8832 11848 8838
rect 11796 8774 11848 8780
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11808 6662 11836 8366
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11900 7410 11928 7822
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11888 7404 11940 7410
rect 11888 7346 11940 7352
rect 11888 7268 11940 7274
rect 11888 7210 11940 7216
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5636 11756 5642
rect 11704 5578 11756 5584
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 11716 5302 11744 5578
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11704 5024 11756 5030
rect 11704 4966 11756 4972
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 11716 4282 11744 4966
rect 11704 4276 11756 4282
rect 11704 4218 11756 4224
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 11702 3496 11758 3505
rect 11702 3431 11758 3440
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 11244 3120 11296 3126
rect 11244 3062 11296 3068
rect 11152 2984 11204 2990
rect 11152 2926 11204 2932
rect 11060 2848 11112 2854
rect 10966 2816 11022 2825
rect 11060 2790 11112 2796
rect 10966 2751 11022 2760
rect 10876 2644 10928 2650
rect 10876 2586 10928 2592
rect 10980 2514 11008 2751
rect 11150 2680 11206 2689
rect 11150 2615 11206 2624
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10966 2408 11022 2417
rect 10966 2343 11022 2352
rect 10980 2310 11008 2343
rect 10968 2304 11020 2310
rect 11164 2281 11192 2615
rect 10968 2246 11020 2252
rect 11150 2272 11206 2281
rect 11150 2207 11206 2216
rect 11256 800 11284 3062
rect 11716 3058 11744 3431
rect 11808 3346 11836 6054
rect 11900 5914 11928 7210
rect 11992 6798 12020 7482
rect 11980 6792 12032 6798
rect 11980 6734 12032 6740
rect 12084 6361 12112 11018
rect 12176 8566 12204 11086
rect 12268 9489 12296 11086
rect 12254 9480 12310 9489
rect 12254 9415 12310 9424
rect 12624 9376 12676 9382
rect 12624 9318 12676 9324
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12360 8650 12388 8842
rect 12636 8838 12664 9318
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12360 8622 12572 8650
rect 12728 8634 12756 14855
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 12992 12096 13044 12102
rect 12992 12038 13044 12044
rect 13452 12096 13504 12102
rect 13452 12038 13504 12044
rect 12808 10668 12860 10674
rect 12808 10610 12860 10616
rect 12820 9178 12848 10610
rect 12900 9580 12952 9586
rect 12900 9522 12952 9528
rect 12912 9382 12940 9522
rect 12900 9376 12952 9382
rect 12900 9318 12952 9324
rect 12808 9172 12860 9178
rect 12808 9114 12860 9120
rect 12912 9042 12940 9318
rect 12900 9036 12952 9042
rect 12900 8978 12952 8984
rect 12164 8560 12216 8566
rect 12164 8502 12216 8508
rect 12256 8288 12308 8294
rect 12256 8230 12308 8236
rect 12268 7206 12296 8230
rect 12440 7812 12492 7818
rect 12440 7754 12492 7760
rect 12256 7200 12308 7206
rect 12256 7142 12308 7148
rect 12452 6866 12480 7754
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12070 6352 12126 6361
rect 12070 6287 12126 6296
rect 12348 6248 12400 6254
rect 12348 6190 12400 6196
rect 12070 6080 12126 6089
rect 12070 6015 12126 6024
rect 11888 5908 11940 5914
rect 11888 5850 11940 5856
rect 11888 5704 11940 5710
rect 11888 5646 11940 5652
rect 11900 4826 11928 5646
rect 11978 5264 12034 5273
rect 11978 5199 12034 5208
rect 11992 5001 12020 5199
rect 11978 4992 12034 5001
rect 11978 4927 12034 4936
rect 11978 4856 12034 4865
rect 11888 4820 11940 4826
rect 11978 4791 12034 4800
rect 11888 4762 11940 4768
rect 11900 4010 11928 4762
rect 11992 4185 12020 4791
rect 11978 4176 12034 4185
rect 11978 4111 12034 4120
rect 11888 4004 11940 4010
rect 11888 3946 11940 3952
rect 11808 3318 11928 3346
rect 11796 3188 11848 3194
rect 11796 3130 11848 3136
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11808 2774 11836 3130
rect 11900 2854 11928 3318
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 11716 2746 11836 2774
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 11716 800 11744 2746
rect 11992 2417 12020 4111
rect 12084 3913 12112 6015
rect 12256 5568 12308 5574
rect 12256 5510 12308 5516
rect 12164 5296 12216 5302
rect 12164 5238 12216 5244
rect 12070 3904 12126 3913
rect 12070 3839 12126 3848
rect 12072 3664 12124 3670
rect 12072 3606 12124 3612
rect 12084 3058 12112 3606
rect 12176 3534 12204 5238
rect 12268 5166 12296 5510
rect 12360 5234 12388 6190
rect 12348 5228 12400 5234
rect 12348 5170 12400 5176
rect 12256 5160 12308 5166
rect 12256 5102 12308 5108
rect 12544 4622 12572 8622
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7410 12848 7822
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12716 6112 12768 6118
rect 13004 6089 13032 12038
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13280 11121 13308 11494
rect 13266 11112 13322 11121
rect 13266 11047 13322 11056
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13096 6866 13124 7346
rect 13084 6860 13136 6866
rect 13084 6802 13136 6808
rect 13096 6458 13124 6802
rect 13084 6452 13136 6458
rect 13084 6394 13136 6400
rect 13188 6338 13216 10406
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13280 6662 13308 8366
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 13372 7886 13400 8230
rect 13360 7880 13412 7886
rect 13360 7822 13412 7828
rect 13268 6656 13320 6662
rect 13268 6598 13320 6604
rect 13096 6322 13216 6338
rect 13084 6316 13216 6322
rect 13136 6310 13216 6316
rect 13084 6258 13136 6264
rect 12716 6054 12768 6060
rect 12990 6080 13046 6089
rect 12728 5642 12756 6054
rect 12990 6015 13046 6024
rect 13280 5953 13308 6598
rect 13266 5944 13322 5953
rect 13266 5879 13322 5888
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12622 4720 12678 4729
rect 12622 4655 12678 4664
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12636 4434 12664 4655
rect 12544 4406 12664 4434
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12544 3194 12572 4406
rect 12728 4146 12756 5578
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3534 12940 3878
rect 12900 3528 12952 3534
rect 12900 3470 12952 3476
rect 12532 3188 12584 3194
rect 12532 3130 12584 3136
rect 13096 3126 13124 5510
rect 13464 4865 13492 12038
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 14292 11121 14320 11494
rect 14830 11248 14886 11257
rect 14830 11183 14832 11192
rect 14884 11183 14886 11192
rect 14832 11154 14884 11160
rect 15304 11150 15332 13126
rect 15658 11656 15714 11665
rect 15658 11591 15714 11600
rect 15200 11144 15252 11150
rect 14278 11112 14334 11121
rect 13728 11076 13780 11082
rect 15200 11086 15252 11092
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 14278 11047 14334 11056
rect 14464 11076 14516 11082
rect 13728 11018 13780 11024
rect 14464 11018 14516 11024
rect 13740 10674 13768 11018
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13832 10146 13860 10746
rect 14370 10704 14426 10713
rect 14370 10639 14372 10648
rect 14424 10639 14426 10648
rect 14372 10610 14424 10616
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 13832 10118 13952 10146
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13648 8430 13676 9998
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 13832 9654 13860 9930
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13924 9364 13952 10118
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 13832 9336 13952 9364
rect 13636 8424 13688 8430
rect 13636 8366 13688 8372
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13556 6798 13584 8230
rect 13648 7342 13676 8366
rect 13636 7336 13688 7342
rect 13636 7278 13688 7284
rect 13648 6798 13676 7278
rect 13544 6792 13596 6798
rect 13544 6734 13596 6740
rect 13636 6792 13688 6798
rect 13636 6734 13688 6740
rect 13648 6254 13676 6734
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13740 6066 13768 6122
rect 13556 6038 13768 6066
rect 13556 5710 13584 6038
rect 13544 5704 13596 5710
rect 13544 5646 13596 5652
rect 13636 5704 13688 5710
rect 13636 5646 13688 5652
rect 13450 4856 13506 4865
rect 13450 4791 13506 4800
rect 13360 3936 13412 3942
rect 13360 3878 13412 3884
rect 13372 3398 13400 3878
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 13084 3120 13136 3126
rect 13556 3097 13584 5646
rect 13648 5030 13676 5646
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4758 13676 4966
rect 13636 4752 13688 4758
rect 13636 4694 13688 4700
rect 13832 4282 13860 9336
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 14292 9110 14320 9522
rect 14280 9104 14332 9110
rect 14280 9046 14332 9052
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 13912 7812 13964 7818
rect 13912 7754 13964 7760
rect 13924 7546 13952 7754
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14292 7206 14320 7958
rect 14476 7857 14504 11018
rect 14648 10532 14700 10538
rect 14648 10474 14700 10480
rect 14554 10024 14610 10033
rect 14554 9959 14556 9968
rect 14608 9959 14610 9968
rect 14556 9930 14608 9936
rect 14462 7848 14518 7857
rect 14462 7783 14518 7792
rect 14372 7268 14424 7274
rect 14372 7210 14424 7216
rect 14280 7200 14332 7206
rect 14280 7142 14332 7148
rect 13945 7100 14253 7120
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 14292 6730 14320 7142
rect 14384 6798 14412 7210
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14464 6656 14516 6662
rect 14464 6598 14516 6604
rect 14476 6458 14504 6598
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14108 4282 14136 4558
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13728 3936 13780 3942
rect 13726 3904 13728 3913
rect 13780 3904 13782 3913
rect 13726 3839 13782 3848
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13648 3194 13676 3538
rect 13832 3194 13860 4082
rect 14108 4026 14136 4218
rect 14384 4146 14412 5238
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 14108 3998 14320 4026
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 14292 3602 14320 3998
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14280 3596 14332 3602
rect 14280 3538 14332 3544
rect 14372 3392 14424 3398
rect 14372 3334 14424 3340
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 3120 13780 3126
rect 13084 3062 13136 3068
rect 13542 3088 13598 3097
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12360 2961 12388 3062
rect 13728 3062 13780 3068
rect 13542 3023 13598 3032
rect 12346 2952 12402 2961
rect 12164 2916 12216 2922
rect 12346 2887 12402 2896
rect 12164 2858 12216 2864
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12084 2689 12112 2790
rect 12070 2680 12126 2689
rect 12070 2615 12126 2624
rect 11978 2408 12034 2417
rect 11978 2343 12034 2352
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 2106 11928 2246
rect 11888 2100 11940 2106
rect 11888 2042 11940 2048
rect 12084 800 12112 2615
rect 12176 2514 12204 2858
rect 13740 2825 13768 3062
rect 14280 2984 14332 2990
rect 14280 2926 14332 2932
rect 13726 2816 13782 2825
rect 13726 2751 13782 2760
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 12532 2576 12584 2582
rect 12532 2518 12584 2524
rect 12164 2508 12216 2514
rect 12164 2450 12216 2456
rect 12544 800 12572 2518
rect 12992 2372 13044 2378
rect 12992 2314 13044 2320
rect 13004 800 13032 2314
rect 13176 2304 13228 2310
rect 13176 2246 13228 2252
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13188 1970 13216 2246
rect 13280 2038 13308 2246
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 13176 1964 13228 1970
rect 13176 1906 13228 1912
rect 13464 800 13492 2586
rect 13636 2576 13688 2582
rect 13636 2518 13688 2524
rect 13648 2446 13676 2518
rect 13636 2440 13688 2446
rect 13636 2382 13688 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 14096 2440 14148 2446
rect 14096 2382 14148 2388
rect 13832 1970 13860 2382
rect 13912 2032 13964 2038
rect 13912 1974 13964 1980
rect 13820 1964 13872 1970
rect 13820 1906 13872 1912
rect 13924 800 13952 1974
rect 14108 1902 14136 2382
rect 14096 1896 14148 1902
rect 14096 1838 14148 1844
rect 14292 800 14320 2926
rect 14384 1766 14412 3334
rect 14568 3058 14596 3878
rect 14660 3466 14688 10474
rect 15212 10266 15240 11086
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15200 10260 15252 10266
rect 15200 10202 15252 10208
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15108 9920 15160 9926
rect 15108 9862 15160 9868
rect 15120 9722 15148 9862
rect 15108 9716 15160 9722
rect 15108 9658 15160 9664
rect 14922 9616 14978 9625
rect 14922 9551 14978 9560
rect 14936 9518 14964 9551
rect 14924 9512 14976 9518
rect 14924 9454 14976 9460
rect 15016 8900 15068 8906
rect 15016 8842 15068 8848
rect 15028 8634 15056 8842
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14936 7886 14964 8366
rect 15028 7954 15056 8570
rect 15016 7948 15068 7954
rect 15016 7890 15068 7896
rect 15108 7948 15160 7954
rect 15108 7890 15160 7896
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 15120 7478 15148 7890
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 14740 6316 14792 6322
rect 14740 6258 14792 6264
rect 14752 5914 14780 6258
rect 15016 6112 15068 6118
rect 15016 6054 15068 6060
rect 14740 5908 14792 5914
rect 14740 5850 14792 5856
rect 15028 5710 15056 6054
rect 15016 5704 15068 5710
rect 15016 5646 15068 5652
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14752 4214 14780 4422
rect 14740 4208 14792 4214
rect 14740 4150 14792 4156
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 15212 3233 15240 9930
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 5914 15332 6122
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15396 4706 15424 10406
rect 15672 9382 15700 11591
rect 15764 11121 15792 17750
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 21284 17241 21312 17478
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19984 14476 20036 14482
rect 19984 14418 20036 14424
rect 18144 14272 18196 14278
rect 18144 14214 18196 14220
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15750 11112 15806 11121
rect 15750 11047 15806 11056
rect 15750 10568 15806 10577
rect 15750 10503 15752 10512
rect 15804 10503 15806 10512
rect 15752 10474 15804 10480
rect 15752 9580 15804 9586
rect 15752 9522 15804 9528
rect 15476 9376 15528 9382
rect 15660 9376 15712 9382
rect 15528 9324 15608 9330
rect 15476 9318 15608 9324
rect 15660 9318 15712 9324
rect 15488 9302 15608 9318
rect 15580 9110 15608 9302
rect 15568 9104 15620 9110
rect 15764 9081 15792 9522
rect 15568 9046 15620 9052
rect 15750 9072 15806 9081
rect 15750 9007 15806 9016
rect 15660 8492 15712 8498
rect 15660 8434 15712 8440
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 15568 8288 15620 8294
rect 15568 8230 15620 8236
rect 15580 8090 15608 8230
rect 15672 8090 15700 8434
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15764 7818 15792 8434
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15660 7472 15712 7478
rect 15660 7414 15712 7420
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15488 6254 15516 6598
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5710 15516 6190
rect 15672 5914 15700 7414
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 6458 15792 6598
rect 15752 6452 15804 6458
rect 15752 6394 15804 6400
rect 15660 5908 15712 5914
rect 15660 5850 15712 5856
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15856 5234 15884 11222
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 16120 10600 16172 10606
rect 16120 10542 16172 10548
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15948 5817 15976 8434
rect 16132 7750 16160 10542
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16212 8424 16264 8430
rect 16212 8366 16264 8372
rect 16028 7744 16080 7750
rect 16028 7686 16080 7692
rect 16120 7744 16172 7750
rect 16120 7686 16172 7692
rect 16040 7478 16068 7686
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 15934 5808 15990 5817
rect 16224 5778 16252 8366
rect 16316 7886 16344 8978
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16396 8084 16448 8090
rect 16396 8026 16448 8032
rect 16304 7880 16356 7886
rect 16304 7822 16356 7828
rect 16316 7342 16344 7822
rect 16408 7410 16436 8026
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 16960 7546 16988 8502
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 16304 7336 16356 7342
rect 16304 7278 16356 7284
rect 17040 7336 17092 7342
rect 17040 7278 17092 7284
rect 16316 6798 16344 7278
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 15934 5743 15990 5752
rect 16212 5772 16264 5778
rect 16212 5714 16264 5720
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 15844 5228 15896 5234
rect 15844 5170 15896 5176
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15568 5160 15620 5166
rect 15568 5102 15620 5108
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15304 4678 15424 4706
rect 15198 3224 15254 3233
rect 15198 3159 15254 3168
rect 14556 3052 14608 3058
rect 14556 2994 14608 3000
rect 14740 2916 14792 2922
rect 14740 2858 14792 2864
rect 14372 1760 14424 1766
rect 14372 1702 14424 1708
rect 14752 800 14780 2858
rect 15304 2854 15332 4678
rect 15382 4584 15438 4593
rect 15382 4519 15438 4528
rect 15396 3194 15424 4519
rect 15580 4486 15608 5102
rect 15764 4826 15792 5102
rect 15752 4820 15804 4826
rect 15752 4762 15804 4768
rect 15948 4554 15976 5170
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15936 4548 15988 4554
rect 15936 4490 15988 4496
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15476 3596 15528 3602
rect 15476 3538 15528 3544
rect 15488 3398 15516 3538
rect 15764 3534 15792 3878
rect 15752 3528 15804 3534
rect 15752 3470 15804 3476
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15292 2848 15344 2854
rect 15292 2790 15344 2796
rect 15382 2680 15438 2689
rect 15382 2615 15438 2624
rect 15292 2440 15344 2446
rect 15292 2382 15344 2388
rect 15200 2372 15252 2378
rect 15200 2314 15252 2320
rect 15212 800 15240 2314
rect 15304 2106 15332 2382
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15396 1737 15424 2615
rect 15382 1728 15438 1737
rect 15382 1663 15438 1672
rect 15672 800 15700 3130
rect 15856 1834 15884 3878
rect 15934 3768 15990 3777
rect 15934 3703 15990 3712
rect 15948 3398 15976 3703
rect 16040 3602 16068 4762
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 16132 3058 16160 5646
rect 16316 5302 16344 6734
rect 16948 6724 17000 6730
rect 16948 6666 17000 6672
rect 16396 6656 16448 6662
rect 16396 6598 16448 6604
rect 16408 6322 16436 6598
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16960 6338 16988 6666
rect 17052 6458 17080 7278
rect 17144 6458 17172 9386
rect 17972 8634 18000 10678
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17314 8528 17370 8537
rect 17314 8463 17316 8472
rect 17368 8463 17370 8472
rect 17316 8434 17368 8440
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17684 6656 17736 6662
rect 17684 6598 17736 6604
rect 17040 6452 17092 6458
rect 17040 6394 17092 6400
rect 17132 6452 17184 6458
rect 17132 6394 17184 6400
rect 16868 6322 16988 6338
rect 16396 6316 16448 6322
rect 16396 6258 16448 6264
rect 16856 6316 16988 6322
rect 16908 6310 16988 6316
rect 17316 6316 17368 6322
rect 16856 6258 16908 6264
rect 17316 6258 17368 6264
rect 16868 5914 16896 6258
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 17224 6248 17276 6254
rect 17224 6190 17276 6196
rect 16856 5908 16908 5914
rect 16856 5850 16908 5856
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16394 5400 16450 5409
rect 16544 5392 16852 5412
rect 16960 5370 16988 6190
rect 16394 5335 16450 5344
rect 16948 5364 17000 5370
rect 16304 5296 16356 5302
rect 16304 5238 16356 5244
rect 16316 4622 16344 5238
rect 16408 5001 16436 5335
rect 16948 5306 17000 5312
rect 17236 5166 17264 6190
rect 17132 5160 17184 5166
rect 17132 5102 17184 5108
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17040 5092 17092 5098
rect 17040 5034 17092 5040
rect 16394 4992 16450 5001
rect 16394 4927 16450 4936
rect 17052 4706 17080 5034
rect 17144 4808 17172 5102
rect 17144 4780 17264 4808
rect 17052 4678 17172 4706
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16396 4480 16448 4486
rect 16396 4422 16448 4428
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16408 4162 16436 4422
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 16960 4214 16988 4422
rect 16948 4208 17000 4214
rect 16212 4140 16264 4146
rect 16408 4134 16620 4162
rect 16212 4082 16264 4088
rect 16120 3052 16172 3058
rect 16120 2994 16172 3000
rect 16224 2689 16252 4082
rect 16592 3534 16620 4134
rect 16868 4156 16948 4162
rect 16868 4150 17000 4156
rect 16868 4134 16988 4150
rect 16868 4078 16896 4134
rect 16960 4085 16988 4134
rect 16856 4072 16908 4078
rect 16856 4014 16908 4020
rect 17052 3738 17080 4490
rect 17144 4078 17172 4678
rect 17236 4321 17264 4780
rect 17222 4312 17278 4321
rect 17222 4247 17278 4256
rect 17328 4162 17356 6258
rect 17696 6066 17724 6598
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17420 6038 17724 6066
rect 17420 5914 17448 6038
rect 17408 5908 17460 5914
rect 17684 5908 17736 5914
rect 17408 5850 17460 5856
rect 17604 5868 17684 5896
rect 17500 5568 17552 5574
rect 17500 5510 17552 5516
rect 17408 5228 17460 5234
rect 17408 5170 17460 5176
rect 17236 4134 17356 4162
rect 17132 4072 17184 4078
rect 17132 4014 17184 4020
rect 17236 3942 17264 4134
rect 17316 4004 17368 4010
rect 17316 3946 17368 3952
rect 17224 3936 17276 3942
rect 17224 3878 17276 3884
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16946 3496 17002 3505
rect 16946 3431 17002 3440
rect 16960 3398 16988 3431
rect 16948 3392 17000 3398
rect 16948 3334 17000 3340
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 17328 3058 17356 3946
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 16396 2916 16448 2922
rect 16396 2858 16448 2864
rect 16210 2680 16266 2689
rect 16120 2644 16172 2650
rect 16210 2615 16266 2624
rect 16120 2586 16172 2592
rect 15844 1828 15896 1834
rect 15844 1770 15896 1776
rect 16132 800 16160 2586
rect 16212 2576 16264 2582
rect 16212 2518 16264 2524
rect 16224 2038 16252 2518
rect 16212 2032 16264 2038
rect 16212 1974 16264 1980
rect 16408 1442 16436 2858
rect 17420 2774 17448 5170
rect 17512 3058 17540 5510
rect 17604 3942 17632 5868
rect 17684 5850 17736 5856
rect 17788 5370 17816 6326
rect 17868 6316 17920 6322
rect 17868 6258 17920 6264
rect 17880 5545 17908 6258
rect 17866 5536 17922 5545
rect 17866 5471 17922 5480
rect 17776 5364 17828 5370
rect 17776 5306 17828 5312
rect 17880 5216 17908 5471
rect 17972 5234 18000 8298
rect 18156 6458 18184 14214
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 18326 13424 18382 13433
rect 18326 13359 18382 13368
rect 18340 10674 18368 13359
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18248 8106 18276 8774
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18326 8392 18382 8401
rect 18326 8327 18328 8336
rect 18380 8327 18382 8336
rect 18328 8298 18380 8304
rect 18248 8078 18368 8106
rect 18234 7984 18290 7993
rect 18234 7919 18290 7928
rect 18248 7886 18276 7919
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18248 5930 18276 6394
rect 18156 5902 18276 5930
rect 18052 5772 18104 5778
rect 18052 5714 18104 5720
rect 17788 5188 17908 5216
rect 17960 5228 18012 5234
rect 17788 4593 17816 5188
rect 17960 5170 18012 5176
rect 17866 5128 17922 5137
rect 17866 5063 17922 5072
rect 17774 4584 17830 4593
rect 17684 4548 17736 4554
rect 17774 4519 17830 4528
rect 17684 4490 17736 4496
rect 17592 3936 17644 3942
rect 17592 3878 17644 3884
rect 17696 3534 17724 4490
rect 17880 4486 17908 5063
rect 17960 5024 18012 5030
rect 17960 4966 18012 4972
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17972 4214 18000 4966
rect 18064 4690 18092 5714
rect 18156 5710 18184 5902
rect 18236 5840 18288 5846
rect 18236 5782 18288 5788
rect 18144 5704 18196 5710
rect 18144 5646 18196 5652
rect 18144 5024 18196 5030
rect 18144 4966 18196 4972
rect 18052 4684 18104 4690
rect 18052 4626 18104 4632
rect 18052 4480 18104 4486
rect 18052 4422 18104 4428
rect 17868 4208 17920 4214
rect 17868 4150 17920 4156
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17776 4072 17828 4078
rect 17774 4040 17776 4049
rect 17828 4040 17830 4049
rect 17774 3975 17830 3984
rect 17776 3936 17828 3942
rect 17776 3878 17828 3884
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17328 2746 17448 2774
rect 16948 2372 17000 2378
rect 16948 2314 17000 2320
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 16408 1414 16528 1442
rect 16500 800 16528 1414
rect 16960 800 16988 2314
rect 17328 2009 17356 2746
rect 17500 2644 17552 2650
rect 17420 2604 17500 2632
rect 17314 2000 17370 2009
rect 17314 1935 17370 1944
rect 17420 800 17448 2604
rect 17500 2586 17552 2592
rect 17788 1970 17816 3878
rect 17880 3670 17908 4150
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 17868 3664 17920 3670
rect 17868 3606 17920 3612
rect 17868 3188 17920 3194
rect 17868 3130 17920 3136
rect 17776 1964 17828 1970
rect 17776 1906 17828 1912
rect 17880 800 17908 3130
rect 17972 2446 18000 3674
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18064 2106 18092 4422
rect 18156 2446 18184 4966
rect 18248 3738 18276 5782
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18340 2774 18368 8078
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18432 6866 18460 7754
rect 18510 7304 18566 7313
rect 18510 7239 18512 7248
rect 18564 7239 18566 7248
rect 18512 7210 18564 7216
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18420 6316 18472 6322
rect 18420 6258 18472 6264
rect 18432 3777 18460 6258
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18524 5681 18552 6190
rect 18616 5710 18644 8502
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18694 7440 18750 7449
rect 18694 7375 18696 7384
rect 18748 7375 18750 7384
rect 18696 7346 18748 7352
rect 18708 7002 18736 7346
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18696 6112 18748 6118
rect 18696 6054 18748 6060
rect 18708 5778 18736 6054
rect 18696 5772 18748 5778
rect 18696 5714 18748 5720
rect 18604 5704 18656 5710
rect 18510 5672 18566 5681
rect 18604 5646 18656 5652
rect 18510 5607 18566 5616
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18512 5568 18564 5574
rect 18510 5536 18512 5545
rect 18564 5536 18566 5545
rect 18510 5471 18566 5480
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18604 5228 18656 5234
rect 18524 4622 18552 5199
rect 18604 5170 18656 5176
rect 18616 4729 18644 5170
rect 18602 4720 18658 4729
rect 18602 4655 18658 4664
rect 18512 4616 18564 4622
rect 18512 4558 18564 4564
rect 18708 4146 18736 5578
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18694 4040 18750 4049
rect 18694 3975 18750 3984
rect 18418 3768 18474 3777
rect 18418 3703 18474 3712
rect 18602 3632 18658 3641
rect 18602 3567 18658 3576
rect 18616 3534 18644 3567
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18708 3466 18736 3975
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 18512 3392 18564 3398
rect 18512 3334 18564 3340
rect 18340 2746 18460 2774
rect 18328 2576 18380 2582
rect 18328 2518 18380 2524
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18052 2100 18104 2106
rect 18052 2042 18104 2048
rect 18340 800 18368 2518
rect 18432 1358 18460 2746
rect 18524 2689 18552 3334
rect 18708 2961 18736 3402
rect 18694 2952 18750 2961
rect 18694 2887 18750 2896
rect 18696 2848 18748 2854
rect 18696 2790 18748 2796
rect 18510 2680 18566 2689
rect 18510 2615 18566 2624
rect 18420 1352 18472 1358
rect 18420 1294 18472 1300
rect 18708 800 18736 2790
rect 18800 2774 18828 8298
rect 18892 7546 18920 12854
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18984 7410 19012 7686
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 18880 7200 18932 7206
rect 18880 7142 18932 7148
rect 18892 5710 18920 7142
rect 18984 7041 19012 7346
rect 18970 7032 19026 7041
rect 18970 6967 19026 6976
rect 18972 6112 19024 6118
rect 18972 6054 19024 6060
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18984 5302 19012 6054
rect 19076 5370 19104 13806
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19706 13288 19762 13297
rect 19706 13223 19762 13232
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19720 12238 19748 13223
rect 19708 12232 19760 12238
rect 19708 12174 19760 12180
rect 19246 11792 19302 11801
rect 19246 11727 19248 11736
rect 19300 11727 19302 11736
rect 19248 11698 19300 11704
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19616 11280 19668 11286
rect 19616 11222 19668 11228
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19524 7268 19576 7274
rect 19524 7210 19576 7216
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 19432 6792 19484 6798
rect 19430 6760 19432 6769
rect 19484 6760 19486 6769
rect 19430 6695 19486 6704
rect 19156 6452 19208 6458
rect 19156 6394 19208 6400
rect 19168 6254 19196 6394
rect 19156 6248 19208 6254
rect 19156 6190 19208 6196
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 19536 5896 19564 7210
rect 19168 5868 19564 5896
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18972 5296 19024 5302
rect 18972 5238 19024 5244
rect 19168 5234 19196 5868
rect 19156 5228 19208 5234
rect 19156 5170 19208 5176
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 18880 5092 18932 5098
rect 18880 5034 18932 5040
rect 18892 3058 18920 5034
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18984 3126 19012 4422
rect 19536 4282 19564 5102
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 19248 4072 19300 4078
rect 19246 4040 19248 4049
rect 19300 4040 19302 4049
rect 19246 3975 19302 3984
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 18972 3120 19024 3126
rect 18972 3062 19024 3068
rect 18880 3052 18932 3058
rect 18880 2994 18932 3000
rect 18800 2746 18920 2774
rect 18892 2553 18920 2746
rect 18878 2544 18934 2553
rect 18878 2479 18934 2488
rect 19076 1714 19104 3606
rect 19628 3058 19656 11222
rect 19892 9104 19944 9110
rect 19892 9046 19944 9052
rect 19904 7410 19932 9046
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19708 6656 19760 6662
rect 19708 6598 19760 6604
rect 19616 3052 19668 3058
rect 19616 2994 19668 3000
rect 19616 2848 19668 2854
rect 19616 2790 19668 2796
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19076 1686 19196 1714
rect 19168 800 19196 1686
rect 19628 800 19656 2790
rect 19720 2446 19748 6598
rect 19812 3126 19840 7142
rect 19892 6792 19944 6798
rect 19892 6734 19944 6740
rect 19904 5914 19932 6734
rect 19996 6458 20024 14418
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20168 11552 20220 11558
rect 20168 11494 20220 11500
rect 20076 10464 20128 10470
rect 20076 10406 20128 10412
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19984 6112 20036 6118
rect 19984 6054 20036 6060
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19892 5568 19944 5574
rect 19892 5510 19944 5516
rect 19904 5234 19932 5510
rect 19892 5228 19944 5234
rect 19892 5170 19944 5176
rect 19890 4040 19946 4049
rect 19890 3975 19892 3984
rect 19944 3975 19946 3984
rect 19892 3946 19944 3952
rect 19890 3904 19946 3913
rect 19890 3839 19946 3848
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 19904 2774 19932 3839
rect 19996 2990 20024 6054
rect 20088 3602 20116 10406
rect 20076 3596 20128 3602
rect 20076 3538 20128 3544
rect 20180 3534 20208 11494
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20272 6798 20300 8230
rect 20444 7200 20496 7206
rect 20444 7142 20496 7148
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20350 5400 20406 5409
rect 20350 5335 20352 5344
rect 20404 5335 20406 5344
rect 20352 5306 20404 5312
rect 20456 5234 20484 7142
rect 20444 5228 20496 5234
rect 20444 5170 20496 5176
rect 20456 5137 20484 5170
rect 20442 5128 20498 5137
rect 20442 5063 20498 5072
rect 20548 3534 20576 12038
rect 20720 8628 20772 8634
rect 20720 8570 20772 8576
rect 20628 5568 20680 5574
rect 20628 5510 20680 5516
rect 20168 3528 20220 3534
rect 20168 3470 20220 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 20076 3392 20128 3398
rect 20076 3334 20128 3340
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19904 2746 20024 2774
rect 19996 2582 20024 2746
rect 19984 2576 20036 2582
rect 19984 2518 20036 2524
rect 19708 2440 19760 2446
rect 19708 2382 19760 2388
rect 20088 800 20116 3334
rect 20548 800 20576 3334
rect 20640 2446 20668 5510
rect 20732 2990 20760 8570
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21272 7472 21324 7478
rect 21272 7414 21324 7420
rect 20996 7200 21048 7206
rect 20996 7142 21048 7148
rect 20904 6724 20956 6730
rect 20904 6666 20956 6672
rect 20812 6656 20864 6662
rect 20812 6598 20864 6604
rect 20824 6322 20852 6598
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 4146 20852 6054
rect 20916 5386 20944 6666
rect 21008 5710 21036 7142
rect 21088 6316 21140 6322
rect 21088 6258 21140 6264
rect 21100 5914 21128 6258
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 20916 5358 21036 5386
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20916 3890 20944 4966
rect 21008 4146 21036 5358
rect 21192 4554 21220 6054
rect 21284 5846 21312 7414
rect 21272 5840 21324 5846
rect 21272 5782 21324 5788
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 20996 4140 21048 4146
rect 20996 4082 21048 4088
rect 20824 3862 20944 3890
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20824 2514 20852 3862
rect 21008 2774 21036 3878
rect 21376 3058 21404 7686
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21468 6322 21496 7142
rect 21456 6316 21508 6322
rect 21456 6258 21508 6264
rect 21468 5817 21496 6258
rect 21454 5808 21510 5817
rect 21454 5743 21510 5752
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 21560 2774 21588 7754
rect 21824 5704 21876 5710
rect 21824 5646 21876 5652
rect 20916 2746 21036 2774
rect 21468 2746 21588 2774
rect 20812 2508 20864 2514
rect 20812 2450 20864 2456
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20916 800 20944 2746
rect 21468 2514 21496 2746
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21468 2394 21496 2450
rect 21376 2366 21496 2394
rect 21376 800 21404 2366
rect 21836 800 21864 5646
rect 22284 4004 22336 4010
rect 22284 3946 22336 3952
rect 22296 800 22324 3946
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22756 800 22784 2994
rect 5552 734 5856 762
rect 5906 0 5962 800
rect 6366 0 6422 800
rect 6826 0 6882 800
rect 7194 0 7250 800
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 9034 0 9090 800
rect 9402 0 9458 800
rect 9862 0 9918 800
rect 10322 0 10378 800
rect 10782 0 10838 800
rect 11242 0 11298 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12530 0 12586 800
rect 12990 0 13046 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14278 0 14334 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
rect 17406 0 17462 800
rect 17866 0 17922 800
rect 18326 0 18382 800
rect 18694 0 18750 800
rect 19154 0 19210 800
rect 19614 0 19670 800
rect 20074 0 20130 800
rect 20534 0 20590 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 1490 22616 1546 22672
rect 3146 22208 3202 22264
rect 2594 21664 2650 21720
rect 1950 21256 2006 21312
rect 1490 19352 1546 19408
rect 1490 18808 1546 18864
rect 1490 18400 1546 18456
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17484 1492 17504
rect 1492 17484 1544 17504
rect 1544 17484 1546 17504
rect 1490 17448 1546 17484
rect 1490 17060 1546 17096
rect 1490 17040 1492 17060
rect 1492 17040 1544 17060
rect 1544 17040 1546 17060
rect 1490 16088 1546 16144
rect 1490 15544 1546 15600
rect 2042 20324 2098 20360
rect 2042 20304 2044 20324
rect 2044 20304 2096 20324
rect 2096 20304 2098 20324
rect 2042 19760 2098 19816
rect 2778 20712 2834 20768
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 2042 16496 2098 16552
rect 1490 15136 1546 15192
rect 1490 14592 1546 14648
rect 1214 12280 1270 12336
rect 1490 13776 1546 13832
rect 1490 13232 1546 13288
rect 2042 14220 2044 14240
rect 2044 14220 2096 14240
rect 2096 14220 2098 14240
rect 2042 14184 2098 14220
rect 1582 9172 1638 9208
rect 1582 9152 1584 9172
rect 1584 9152 1636 9172
rect 1636 9152 1638 9172
rect 1674 8744 1730 8800
rect 1490 6316 1546 6352
rect 1490 6296 1492 6316
rect 1492 6296 1544 6316
rect 1544 6296 1546 6316
rect 1582 5616 1638 5672
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3790 12824 3846 12880
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3422 11348 3478 11384
rect 3422 11328 3424 11348
rect 3424 11328 3476 11348
rect 3476 11328 3478 11348
rect 2226 9868 2228 9888
rect 2228 9868 2280 9888
rect 2280 9868 2282 9888
rect 2226 9832 2282 9868
rect 3422 10376 3478 10432
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 2042 5752 2098 5808
rect 1490 3304 1546 3360
rect 1398 2488 1454 2544
rect 1030 1944 1086 2000
rect 2134 4120 2190 4176
rect 1950 2760 2006 2816
rect 1490 1672 1546 1728
rect 2226 4020 2228 4040
rect 2228 4020 2280 4040
rect 2280 4020 2282 4040
rect 2226 3984 2282 4020
rect 2778 8200 2834 8256
rect 2778 7656 2834 7712
rect 2778 5208 2834 5264
rect 3146 9696 3202 9752
rect 3422 9560 3478 9616
rect 3054 7928 3110 7984
rect 2962 4392 3018 4448
rect 2686 3188 2742 3224
rect 2686 3168 2688 3188
rect 2688 3168 2740 3188
rect 2740 3168 2742 3188
rect 2778 3032 2834 3088
rect 2134 2080 2190 2136
rect 2502 2352 2558 2408
rect 2870 584 2926 640
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3422 8608 3478 8664
rect 3422 8472 3478 8528
rect 3422 8200 3478 8256
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3422 8064 3478 8120
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 4066 11872 4122 11928
rect 4066 10920 4122 10976
rect 4342 10104 4398 10160
rect 4618 11092 4620 11112
rect 4620 11092 4672 11112
rect 4672 11092 4674 11112
rect 4618 11056 4674 11092
rect 4066 10004 4068 10024
rect 4068 10004 4120 10024
rect 4120 10004 4122 10024
rect 4066 9968 4122 10004
rect 4066 9016 4122 9072
rect 4158 8744 4214 8800
rect 3974 8608 4030 8664
rect 4066 7828 4068 7848
rect 4068 7828 4120 7848
rect 4120 7828 4122 7848
rect 4066 7792 4122 7828
rect 3054 3440 3110 3496
rect 3146 2488 3202 2544
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3422 3848 3478 3904
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 4066 5652 4068 5672
rect 4068 5652 4120 5672
rect 4120 5652 4122 5672
rect 4066 5616 4122 5652
rect 4802 9696 4858 9752
rect 4710 9152 4766 9208
rect 3974 4820 4030 4856
rect 3974 4800 3976 4820
rect 3976 4800 4028 4820
rect 4028 4800 4030 4820
rect 3974 4004 4030 4040
rect 3974 3984 3976 4004
rect 3976 3984 4028 4004
rect 4028 3984 4030 4004
rect 3422 3168 3478 3224
rect 3882 2896 3938 2952
rect 3422 2760 3478 2816
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3330 2508 3386 2544
rect 3330 2488 3332 2508
rect 3332 2488 3384 2508
rect 3384 2488 3386 2508
rect 4066 1536 4122 1592
rect 4802 5652 4804 5672
rect 4804 5652 4856 5672
rect 4856 5652 4858 5672
rect 4802 5616 4858 5652
rect 5354 11636 5356 11656
rect 5356 11636 5408 11656
rect 5408 11636 5410 11656
rect 5354 11600 5410 11636
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6550 14884 6606 14920
rect 6550 14864 6552 14884
rect 6552 14864 6604 14884
rect 6604 14864 6606 14884
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 5722 10648 5778 10704
rect 5446 10512 5502 10568
rect 5630 9016 5686 9072
rect 5722 8472 5778 8528
rect 5630 7248 5686 7304
rect 4526 992 4582 1048
rect 5446 4548 5502 4584
rect 5446 4528 5448 4548
rect 5448 4528 5500 4548
rect 5500 4528 5502 4548
rect 4986 2624 5042 2680
rect 5538 3304 5594 3360
rect 2962 176 3018 232
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6826 11092 6828 11112
rect 6828 11092 6880 11112
rect 6880 11092 6882 11112
rect 6826 11056 6882 11092
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6274 9288 6330 9344
rect 6182 9152 6238 9208
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6734 8608 6790 8664
rect 6826 8472 6882 8528
rect 6366 6316 6422 6352
rect 6366 6296 6368 6316
rect 6368 6296 6420 6316
rect 6420 6296 6422 6316
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 7286 12144 7342 12200
rect 7286 8336 7342 8392
rect 6826 6840 6882 6896
rect 7470 7792 7526 7848
rect 6918 6432 6974 6488
rect 6918 6160 6974 6216
rect 5998 3576 6054 3632
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6826 3168 6882 3224
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6366 1808 6422 1864
rect 8206 12824 8262 12880
rect 7838 12280 7894 12336
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8666 13232 8722 13288
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9218 12416 9274 12472
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 9678 13368 9734 13424
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8114 9288 8170 9344
rect 8022 8608 8078 8664
rect 7930 7248 7986 7304
rect 7654 5208 7710 5264
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8574 8336 8630 8392
rect 9034 8336 9090 8392
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 12530 17604 12586 17640
rect 12530 17584 12532 17604
rect 12532 17584 12584 17604
rect 12584 17584 12586 17604
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9494 8372 9496 8392
rect 9496 8372 9548 8392
rect 9548 8372 9550 8392
rect 9494 8336 9550 8372
rect 9586 7928 9642 7984
rect 8482 6160 8538 6216
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8114 3984 8170 4040
rect 9034 5072 9090 5128
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9678 6976 9734 7032
rect 9678 4800 9734 4856
rect 9678 2760 9734 2816
rect 10138 8900 10194 8936
rect 10138 8880 10140 8900
rect 10140 8880 10192 8900
rect 10192 8880 10194 8900
rect 9862 4156 9864 4176
rect 9864 4156 9916 4176
rect 9916 4156 9918 4176
rect 9862 4120 9918 4156
rect 10230 5616 10286 5672
rect 10046 3440 10102 3496
rect 10414 4156 10416 4176
rect 10416 4156 10468 4176
rect 10468 4156 10470 4176
rect 10414 4120 10470 4156
rect 11058 12416 11114 12472
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11518 12588 11520 12608
rect 11520 12588 11572 12608
rect 11572 12588 11574 12608
rect 11518 12552 11574 12588
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 10874 7656 10930 7712
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11334 7248 11390 7304
rect 10782 4120 10838 4176
rect 10598 2352 10654 2408
rect 10874 3984 10930 4040
rect 11058 3984 11114 4040
rect 10874 3712 10930 3768
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 12714 14864 12770 14920
rect 12622 12144 12678 12200
rect 11978 10104 12034 10160
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11702 3440 11758 3496
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 10966 2760 11022 2816
rect 11150 2624 11206 2680
rect 10966 2352 11022 2408
rect 11150 2216 11206 2272
rect 12254 9424 12310 9480
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 12070 6296 12126 6352
rect 12070 6024 12126 6080
rect 11978 5208 12034 5264
rect 11978 4936 12034 4992
rect 11978 4800 12034 4856
rect 11978 4120 12034 4176
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12070 3848 12126 3904
rect 13266 11056 13322 11112
rect 12990 6024 13046 6080
rect 13266 5888 13322 5944
rect 12622 4664 12678 4720
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14830 11212 14886 11248
rect 14830 11192 14832 11212
rect 14832 11192 14884 11212
rect 14884 11192 14886 11212
rect 15658 11600 15714 11656
rect 14278 11056 14334 11112
rect 14370 10668 14426 10704
rect 14370 10648 14372 10668
rect 14372 10648 14424 10668
rect 14424 10648 14426 10668
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13450 4800 13506 4856
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 14554 9988 14610 10024
rect 14554 9968 14556 9988
rect 14556 9968 14608 9988
rect 14608 9968 14610 9988
rect 14462 7792 14518 7848
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13726 3884 13728 3904
rect 13728 3884 13780 3904
rect 13780 3884 13782 3904
rect 13726 3848 13782 3884
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13542 3032 13598 3088
rect 12346 2896 12402 2952
rect 12070 2624 12126 2680
rect 11978 2352 12034 2408
rect 13726 2760 13782 2816
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14922 9560 14978 9616
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 21270 17176 21326 17232
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 15750 11056 15806 11112
rect 15750 10532 15806 10568
rect 15750 10512 15752 10532
rect 15752 10512 15804 10532
rect 15804 10512 15806 10532
rect 15750 9016 15806 9072
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 15934 5752 15990 5808
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 15198 3168 15254 3224
rect 15382 4528 15438 4584
rect 15382 2624 15438 2680
rect 15382 1672 15438 1728
rect 15934 3712 15990 3768
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 17314 8492 17370 8528
rect 17314 8472 17316 8492
rect 17316 8472 17368 8492
rect 17368 8472 17370 8492
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16394 5344 16450 5400
rect 16394 4936 16450 4992
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 17222 4256 17278 4312
rect 16946 3440 17002 3496
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16210 2624 16266 2680
rect 17866 5480 17922 5536
rect 18326 13368 18382 13424
rect 18326 8356 18382 8392
rect 18326 8336 18328 8356
rect 18328 8336 18380 8356
rect 18380 8336 18382 8356
rect 18234 7928 18290 7984
rect 17866 5072 17922 5128
rect 17774 4528 17830 4584
rect 17774 4020 17776 4040
rect 17776 4020 17828 4040
rect 17828 4020 17830 4040
rect 17774 3984 17830 4020
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17314 1944 17370 2000
rect 18510 7268 18566 7304
rect 18510 7248 18512 7268
rect 18512 7248 18564 7268
rect 18564 7248 18566 7268
rect 18694 7404 18750 7440
rect 18694 7384 18696 7404
rect 18696 7384 18748 7404
rect 18748 7384 18750 7404
rect 18510 5616 18566 5672
rect 18510 5516 18512 5536
rect 18512 5516 18564 5536
rect 18564 5516 18566 5536
rect 18510 5480 18566 5516
rect 18510 5208 18566 5264
rect 18602 4664 18658 4720
rect 18694 3984 18750 4040
rect 18418 3712 18474 3768
rect 18602 3576 18658 3632
rect 18694 2896 18750 2952
rect 18510 2624 18566 2680
rect 18970 6976 19026 7032
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19706 13232 19762 13288
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19246 11756 19302 11792
rect 19246 11736 19248 11756
rect 19248 11736 19300 11756
rect 19300 11736 19302 11756
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19430 6740 19432 6760
rect 19432 6740 19484 6760
rect 19484 6740 19486 6760
rect 19430 6704 19486 6740
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19246 4020 19248 4040
rect 19248 4020 19300 4040
rect 19300 4020 19302 4040
rect 19246 3984 19302 4020
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 18878 2488 18934 2544
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19890 4004 19946 4040
rect 19890 3984 19892 4004
rect 19892 3984 19944 4004
rect 19944 3984 19946 4004
rect 19890 3848 19946 3904
rect 20350 5364 20406 5400
rect 20350 5344 20352 5364
rect 20352 5344 20404 5364
rect 20404 5344 20406 5364
rect 20442 5072 20498 5128
rect 21454 5752 21510 5808
<< metal3 >>
rect 0 22674 800 22704
rect 1485 22674 1551 22677
rect 0 22672 1551 22674
rect 0 22616 1490 22672
rect 1546 22616 1551 22672
rect 0 22614 1551 22616
rect 0 22584 800 22614
rect 1485 22611 1551 22614
rect 0 22266 800 22296
rect 3141 22266 3207 22269
rect 0 22264 3207 22266
rect 0 22208 3146 22264
rect 3202 22208 3207 22264
rect 0 22206 3207 22208
rect 0 22176 800 22206
rect 3141 22203 3207 22206
rect 0 21722 800 21752
rect 2589 21722 2655 21725
rect 0 21720 2655 21722
rect 0 21664 2594 21720
rect 2650 21664 2655 21720
rect 0 21662 2655 21664
rect 0 21632 800 21662
rect 2589 21659 2655 21662
rect 0 21314 800 21344
rect 1945 21314 2011 21317
rect 0 21312 2011 21314
rect 0 21256 1950 21312
rect 2006 21256 2011 21312
rect 0 21254 2011 21256
rect 0 21224 800 21254
rect 1945 21251 2011 21254
rect 0 20770 800 20800
rect 2773 20770 2839 20773
rect 0 20768 2839 20770
rect 0 20712 2778 20768
rect 2834 20712 2839 20768
rect 0 20710 2839 20712
rect 0 20680 800 20710
rect 2773 20707 2839 20710
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 20639 16858 20640
rect 0 20362 800 20392
rect 2037 20362 2103 20365
rect 0 20360 2103 20362
rect 0 20304 2042 20360
rect 2098 20304 2103 20360
rect 0 20302 2103 20304
rect 0 20272 800 20302
rect 2037 20299 2103 20302
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 0 19818 800 19848
rect 2037 19818 2103 19821
rect 0 19816 2103 19818
rect 0 19760 2042 19816
rect 2098 19760 2103 19816
rect 0 19758 2103 19760
rect 0 19728 800 19758
rect 2037 19755 2103 19758
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 6142 18528 6462 18529
rect 0 18458 800 18488
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 18463 16858 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 17919 19457 17920
rect 12525 17642 12591 17645
rect 19926 17642 19932 17644
rect 12525 17640 19932 17642
rect 12525 17584 12530 17640
rect 12586 17584 19932 17640
rect 12525 17582 19932 17584
rect 12525 17579 12591 17582
rect 19926 17580 19932 17582
rect 19996 17580 20002 17644
rect 0 17506 800 17536
rect 1485 17506 1551 17509
rect 0 17504 1551 17506
rect 0 17448 1490 17504
rect 1546 17448 1551 17504
rect 0 17446 1551 17448
rect 0 17416 800 17446
rect 1485 17443 1551 17446
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 17375 16858 17376
rect 21265 17234 21331 17237
rect 22200 17234 23000 17264
rect 21265 17232 23000 17234
rect 21265 17176 21270 17232
rect 21326 17176 23000 17232
rect 21265 17174 23000 17176
rect 21265 17171 21331 17174
rect 22200 17144 23000 17174
rect 0 17098 800 17128
rect 1485 17098 1551 17101
rect 0 17096 1551 17098
rect 0 17040 1490 17096
rect 1546 17040 1551 17096
rect 0 17038 1551 17040
rect 0 17008 800 17038
rect 1485 17035 1551 17038
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 0 16554 800 16584
rect 2037 16554 2103 16557
rect 0 16552 2103 16554
rect 0 16496 2042 16552
rect 2098 16496 2103 16552
rect 0 16494 2103 16496
rect 0 16464 800 16494
rect 2037 16491 2103 16494
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 0 16146 800 16176
rect 1485 16146 1551 16149
rect 0 16144 1551 16146
rect 0 16088 1490 16144
rect 1546 16088 1551 16144
rect 0 16086 1551 16088
rect 0 16056 800 16086
rect 1485 16083 1551 16086
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 6142 15264 6462 15265
rect 0 15194 800 15224
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 15199 16858 15200
rect 1485 15194 1551 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 6545 14922 6611 14925
rect 12709 14922 12775 14925
rect 6545 14920 12775 14922
rect 6545 14864 6550 14920
rect 6606 14864 12714 14920
rect 12770 14864 12775 14920
rect 6545 14862 12775 14864
rect 6545 14859 6611 14862
rect 12709 14859 12775 14862
rect 3543 14720 3863 14721
rect 0 14650 800 14680
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 800 14590
rect 1485 14587 1551 14590
rect 0 14242 800 14272
rect 2037 14242 2103 14245
rect 0 14240 2103 14242
rect 0 14184 2042 14240
rect 2098 14184 2103 14240
rect 0 14182 2103 14184
rect 0 14152 800 14182
rect 2037 14179 2103 14182
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 14111 16858 14112
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 9673 13426 9739 13429
rect 18321 13426 18387 13429
rect 9673 13424 18387 13426
rect 9673 13368 9678 13424
rect 9734 13368 18326 13424
rect 18382 13368 18387 13424
rect 9673 13366 18387 13368
rect 9673 13363 9739 13366
rect 18321 13363 18387 13366
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 8661 13290 8727 13293
rect 19701 13290 19767 13293
rect 8661 13288 19767 13290
rect 8661 13232 8666 13288
rect 8722 13232 19706 13288
rect 19762 13232 19767 13288
rect 8661 13230 19767 13232
rect 8661 13227 8727 13230
rect 19701 13227 19767 13230
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 0 12882 800 12912
rect 3785 12882 3851 12885
rect 0 12880 3851 12882
rect 0 12824 3790 12880
rect 3846 12824 3851 12880
rect 0 12822 3851 12824
rect 0 12792 800 12822
rect 3785 12819 3851 12822
rect 3918 12820 3924 12884
rect 3988 12882 3994 12884
rect 8201 12882 8267 12885
rect 3988 12880 8267 12882
rect 3988 12824 8206 12880
rect 8262 12824 8267 12880
rect 3988 12822 8267 12824
rect 3988 12820 3994 12822
rect 8201 12819 8267 12822
rect 11094 12548 11100 12612
rect 11164 12610 11170 12612
rect 11513 12610 11579 12613
rect 11164 12608 11579 12610
rect 11164 12552 11518 12608
rect 11574 12552 11579 12608
rect 11164 12550 11579 12552
rect 11164 12548 11170 12550
rect 11513 12547 11579 12550
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 12479 19457 12480
rect 9213 12474 9279 12477
rect 11053 12474 11119 12477
rect 9213 12472 11119 12474
rect 9213 12416 9218 12472
rect 9274 12416 11058 12472
rect 11114 12416 11119 12472
rect 9213 12414 11119 12416
rect 9213 12411 9279 12414
rect 11053 12411 11119 12414
rect 0 12338 800 12368
rect 1209 12338 1275 12341
rect 7833 12338 7899 12341
rect 0 12336 7899 12338
rect 0 12280 1214 12336
rect 1270 12280 7838 12336
rect 7894 12280 7899 12336
rect 0 12278 7899 12280
rect 0 12248 800 12278
rect 1209 12275 1275 12278
rect 7833 12275 7899 12278
rect 7281 12202 7347 12205
rect 12617 12202 12683 12205
rect 7281 12200 12683 12202
rect 7281 12144 7286 12200
rect 7342 12144 12622 12200
rect 12678 12144 12683 12200
rect 7281 12142 12683 12144
rect 7281 12139 7347 12142
rect 12617 12139 12683 12142
rect 6142 12000 6462 12001
rect 0 11930 800 11960
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 11935 16858 11936
rect 4061 11930 4127 11933
rect 0 11928 4127 11930
rect 0 11872 4066 11928
rect 4122 11872 4127 11928
rect 0 11870 4127 11872
rect 0 11840 800 11870
rect 4061 11867 4127 11870
rect 1710 11732 1716 11796
rect 1780 11794 1786 11796
rect 19241 11794 19307 11797
rect 1780 11792 19307 11794
rect 1780 11736 19246 11792
rect 19302 11736 19307 11792
rect 1780 11734 19307 11736
rect 1780 11732 1786 11734
rect 19241 11731 19307 11734
rect 5349 11658 5415 11661
rect 15653 11658 15719 11661
rect 5349 11656 15719 11658
rect 5349 11600 5354 11656
rect 5410 11600 15658 11656
rect 15714 11600 15719 11656
rect 5349 11598 15719 11600
rect 5349 11595 5415 11598
rect 15653 11595 15719 11598
rect 3543 11456 3863 11457
rect 0 11386 800 11416
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 3417 11386 3483 11389
rect 0 11384 3483 11386
rect 0 11328 3422 11384
rect 3478 11328 3483 11384
rect 0 11326 3483 11328
rect 0 11296 800 11326
rect 3417 11323 3483 11326
rect 14825 11250 14891 11253
rect 2730 11248 14891 11250
rect 2730 11192 14830 11248
rect 14886 11192 14891 11248
rect 2730 11190 14891 11192
rect 2262 11052 2268 11116
rect 2332 11114 2338 11116
rect 2730 11114 2790 11190
rect 14825 11187 14891 11190
rect 2332 11054 2790 11114
rect 4613 11114 4679 11117
rect 6821 11114 6887 11117
rect 4613 11112 6887 11114
rect 4613 11056 4618 11112
rect 4674 11056 6826 11112
rect 6882 11056 6887 11112
rect 4613 11054 6887 11056
rect 2332 11052 2338 11054
rect 4613 11051 4679 11054
rect 6821 11051 6887 11054
rect 13261 11116 13327 11117
rect 13261 11112 13308 11116
rect 13372 11114 13378 11116
rect 14273 11114 14339 11117
rect 14406 11114 14412 11116
rect 13261 11056 13266 11112
rect 13261 11052 13308 11056
rect 13372 11054 13418 11114
rect 14273 11112 14412 11114
rect 14273 11056 14278 11112
rect 14334 11056 14412 11112
rect 14273 11054 14412 11056
rect 13372 11052 13378 11054
rect 13261 11051 13327 11052
rect 14273 11051 14339 11054
rect 14406 11052 14412 11054
rect 14476 11052 14482 11116
rect 15745 11114 15811 11117
rect 20294 11114 20300 11116
rect 15745 11112 20300 11114
rect 15745 11056 15750 11112
rect 15806 11056 20300 11112
rect 15745 11054 20300 11056
rect 15745 11051 15811 11054
rect 20294 11052 20300 11054
rect 20364 11052 20370 11116
rect 0 10978 800 11008
rect 4061 10978 4127 10981
rect 0 10976 4127 10978
rect 0 10920 4066 10976
rect 4122 10920 4127 10976
rect 0 10918 4127 10920
rect 0 10888 800 10918
rect 4061 10915 4127 10918
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 5717 10706 5783 10709
rect 14365 10706 14431 10709
rect 5717 10704 14431 10706
rect 5717 10648 5722 10704
rect 5778 10648 14370 10704
rect 14426 10648 14431 10704
rect 5717 10646 14431 10648
rect 5717 10643 5783 10646
rect 14365 10643 14431 10646
rect 5441 10570 5507 10573
rect 15745 10570 15811 10573
rect 5441 10568 15811 10570
rect 5441 10512 5446 10568
rect 5502 10512 15750 10568
rect 15806 10512 15811 10568
rect 5441 10510 15811 10512
rect 5441 10507 5507 10510
rect 15745 10507 15811 10510
rect 0 10434 800 10464
rect 3417 10434 3483 10437
rect 0 10432 3483 10434
rect 0 10376 3422 10432
rect 3478 10376 3483 10432
rect 0 10374 3483 10376
rect 0 10344 800 10374
rect 3417 10371 3483 10374
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 10303 19457 10304
rect 4337 10162 4403 10165
rect 11973 10162 12039 10165
rect 4337 10160 12039 10162
rect 4337 10104 4342 10160
rect 4398 10104 11978 10160
rect 12034 10104 12039 10160
rect 4337 10102 12039 10104
rect 4337 10099 4403 10102
rect 11973 10099 12039 10102
rect 0 10026 800 10056
rect 4061 10026 4127 10029
rect 14549 10026 14615 10029
rect 0 10024 4127 10026
rect 0 9968 4066 10024
rect 4122 9968 4127 10024
rect 0 9966 4127 9968
rect 0 9936 800 9966
rect 4061 9963 4127 9966
rect 5950 10024 14615 10026
rect 5950 9968 14554 10024
rect 14610 9968 14615 10024
rect 5950 9966 14615 9968
rect 2221 9890 2287 9893
rect 5950 9890 6010 9966
rect 14549 9963 14615 9966
rect 2221 9888 6010 9890
rect 2221 9832 2226 9888
rect 2282 9832 6010 9888
rect 2221 9830 6010 9832
rect 2221 9827 2287 9830
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 3141 9754 3207 9757
rect 4797 9754 4863 9757
rect 3141 9752 4863 9754
rect 3141 9696 3146 9752
rect 3202 9696 4802 9752
rect 4858 9696 4863 9752
rect 3141 9694 4863 9696
rect 3141 9691 3207 9694
rect 4797 9691 4863 9694
rect 3417 9618 3483 9621
rect 14917 9618 14983 9621
rect 3417 9616 14983 9618
rect 3417 9560 3422 9616
rect 3478 9560 14922 9616
rect 14978 9560 14983 9616
rect 3417 9558 14983 9560
rect 3417 9555 3483 9558
rect 14917 9555 14983 9558
rect 0 9482 800 9512
rect 12249 9482 12315 9485
rect 0 9480 12315 9482
rect 0 9424 12254 9480
rect 12310 9424 12315 9480
rect 0 9422 12315 9424
rect 0 9392 800 9422
rect 12249 9419 12315 9422
rect 6269 9346 6335 9349
rect 8109 9346 8175 9349
rect 6269 9344 8175 9346
rect 6269 9288 6274 9344
rect 6330 9288 8114 9344
rect 8170 9288 8175 9344
rect 6269 9286 8175 9288
rect 6269 9283 6335 9286
rect 8109 9283 8175 9286
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 9215 19457 9216
rect 1577 9210 1643 9213
rect 1710 9210 1716 9212
rect 1577 9208 1716 9210
rect 1577 9152 1582 9208
rect 1638 9152 1716 9208
rect 1577 9150 1716 9152
rect 1577 9147 1643 9150
rect 1710 9148 1716 9150
rect 1780 9148 1786 9212
rect 4705 9210 4771 9213
rect 6177 9210 6243 9213
rect 4705 9208 6243 9210
rect 4705 9152 4710 9208
rect 4766 9152 6182 9208
rect 6238 9152 6243 9208
rect 4705 9150 6243 9152
rect 4705 9147 4771 9150
rect 6177 9147 6243 9150
rect 0 9074 800 9104
rect 4061 9074 4127 9077
rect 0 9072 4127 9074
rect 0 9016 4066 9072
rect 4122 9016 4127 9072
rect 0 9014 4127 9016
rect 0 8984 800 9014
rect 4061 9011 4127 9014
rect 5625 9074 5691 9077
rect 15745 9074 15811 9077
rect 5625 9072 15811 9074
rect 5625 9016 5630 9072
rect 5686 9016 15750 9072
rect 15806 9016 15811 9072
rect 5625 9014 15811 9016
rect 5625 9011 5691 9014
rect 15745 9011 15811 9014
rect 2446 8876 2452 8940
rect 2516 8938 2522 8940
rect 10133 8938 10199 8941
rect 2516 8936 10199 8938
rect 2516 8880 10138 8936
rect 10194 8880 10199 8936
rect 2516 8878 10199 8880
rect 2516 8876 2522 8878
rect 10133 8875 10199 8878
rect 1669 8802 1735 8805
rect 4153 8802 4219 8805
rect 1669 8800 4219 8802
rect 1669 8744 1674 8800
rect 1730 8744 4158 8800
rect 4214 8744 4219 8800
rect 1669 8742 4219 8744
rect 1669 8739 1735 8742
rect 4153 8739 4219 8742
rect 6142 8736 6462 8737
rect 0 8666 800 8696
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 3417 8666 3483 8669
rect 3969 8666 4035 8669
rect 0 8664 4035 8666
rect 0 8608 3422 8664
rect 3478 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 800 8606
rect 3417 8603 3483 8606
rect 3969 8603 4035 8606
rect 6729 8666 6795 8669
rect 8017 8666 8083 8669
rect 6729 8664 8083 8666
rect 6729 8608 6734 8664
rect 6790 8608 8022 8664
rect 8078 8608 8083 8664
rect 6729 8606 8083 8608
rect 6729 8603 6795 8606
rect 8017 8603 8083 8606
rect 3417 8530 3483 8533
rect 5717 8530 5783 8533
rect 3417 8528 5783 8530
rect 3417 8472 3422 8528
rect 3478 8472 5722 8528
rect 5778 8472 5783 8528
rect 3417 8470 5783 8472
rect 3417 8467 3483 8470
rect 5717 8467 5783 8470
rect 6821 8530 6887 8533
rect 17309 8530 17375 8533
rect 6821 8528 17375 8530
rect 6821 8472 6826 8528
rect 6882 8472 17314 8528
rect 17370 8472 17375 8528
rect 6821 8470 17375 8472
rect 6821 8467 6887 8470
rect 17309 8467 17375 8470
rect 6678 8332 6684 8396
rect 6748 8394 6754 8396
rect 7281 8394 7347 8397
rect 6748 8392 7347 8394
rect 6748 8336 7286 8392
rect 7342 8336 7347 8392
rect 6748 8334 7347 8336
rect 6748 8332 6754 8334
rect 7281 8331 7347 8334
rect 8569 8394 8635 8397
rect 9029 8394 9095 8397
rect 9489 8394 9555 8397
rect 18321 8394 18387 8397
rect 8569 8392 18387 8394
rect 8569 8336 8574 8392
rect 8630 8336 9034 8392
rect 9090 8336 9494 8392
rect 9550 8336 18326 8392
rect 18382 8336 18387 8392
rect 8569 8334 18387 8336
rect 8569 8331 8635 8334
rect 9029 8331 9095 8334
rect 9489 8331 9555 8334
rect 18321 8331 18387 8334
rect 2773 8258 2839 8261
rect 3417 8258 3483 8261
rect 2773 8256 3483 8258
rect 2773 8200 2778 8256
rect 2834 8200 3422 8256
rect 3478 8200 3483 8256
rect 2773 8198 3483 8200
rect 2773 8195 2839 8198
rect 3417 8195 3483 8198
rect 3543 8192 3863 8193
rect 0 8122 800 8152
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 3417 8122 3483 8125
rect 0 8120 3483 8122
rect 0 8064 3422 8120
rect 3478 8064 3483 8120
rect 0 8062 3483 8064
rect 0 8032 800 8062
rect 3417 8059 3483 8062
rect 3049 7986 3115 7989
rect 9581 7986 9647 7989
rect 18229 7986 18295 7989
rect 3049 7984 7850 7986
rect 3049 7928 3054 7984
rect 3110 7928 7850 7984
rect 3049 7926 7850 7928
rect 3049 7923 3115 7926
rect 4061 7850 4127 7853
rect 4470 7850 4476 7852
rect 4061 7848 4476 7850
rect 4061 7792 4066 7848
rect 4122 7792 4476 7848
rect 4061 7790 4476 7792
rect 4061 7787 4127 7790
rect 4470 7788 4476 7790
rect 4540 7850 4546 7852
rect 7465 7850 7531 7853
rect 7598 7850 7604 7852
rect 4540 7790 6746 7850
rect 4540 7788 4546 7790
rect 0 7714 800 7744
rect 2773 7714 2839 7717
rect 0 7712 2839 7714
rect 0 7656 2778 7712
rect 2834 7656 2839 7712
rect 0 7654 2839 7656
rect 6686 7714 6746 7790
rect 7465 7848 7604 7850
rect 7465 7792 7470 7848
rect 7526 7792 7604 7848
rect 7465 7790 7604 7792
rect 7465 7787 7531 7790
rect 7598 7788 7604 7790
rect 7668 7788 7674 7852
rect 7790 7850 7850 7926
rect 9581 7984 18295 7986
rect 9581 7928 9586 7984
rect 9642 7928 18234 7984
rect 18290 7928 18295 7984
rect 9581 7926 18295 7928
rect 9581 7923 9647 7926
rect 18229 7923 18295 7926
rect 14457 7850 14523 7853
rect 7790 7848 14523 7850
rect 7790 7792 14462 7848
rect 14518 7792 14523 7848
rect 7790 7790 14523 7792
rect 14457 7787 14523 7790
rect 10869 7714 10935 7717
rect 6686 7712 10935 7714
rect 6686 7656 10874 7712
rect 10930 7656 10935 7712
rect 6686 7654 10935 7656
rect 0 7624 800 7654
rect 2773 7651 2839 7654
rect 10869 7651 10935 7654
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 18689 7442 18755 7445
rect 2730 7440 18755 7442
rect 2730 7384 18694 7440
rect 18750 7384 18755 7440
rect 2730 7382 18755 7384
rect 0 7170 800 7200
rect 2730 7170 2790 7382
rect 18689 7379 18755 7382
rect 5625 7306 5691 7309
rect 5942 7306 5948 7308
rect 5625 7304 5948 7306
rect 5625 7248 5630 7304
rect 5686 7248 5948 7304
rect 5625 7246 5948 7248
rect 5625 7243 5691 7246
rect 5942 7244 5948 7246
rect 6012 7244 6018 7308
rect 7925 7306 7991 7309
rect 9622 7306 9628 7308
rect 7925 7304 9628 7306
rect 7925 7248 7930 7304
rect 7986 7248 9628 7304
rect 7925 7246 9628 7248
rect 7925 7243 7991 7246
rect 9622 7244 9628 7246
rect 9692 7244 9698 7308
rect 11329 7306 11395 7309
rect 18505 7306 18571 7309
rect 11329 7304 18571 7306
rect 11329 7248 11334 7304
rect 11390 7248 18510 7304
rect 18566 7248 18571 7304
rect 11329 7246 18571 7248
rect 11329 7243 11395 7246
rect 18505 7243 18571 7246
rect 0 7110 2790 7170
rect 0 7080 800 7110
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 9673 7034 9739 7037
rect 18965 7034 19031 7037
rect 9673 7032 13738 7034
rect 9673 6976 9678 7032
rect 9734 6976 13738 7032
rect 9673 6974 13738 6976
rect 9673 6971 9739 6974
rect 6821 6898 6887 6901
rect 2730 6896 6887 6898
rect 2730 6840 6826 6896
rect 6882 6840 6887 6896
rect 2730 6838 6887 6840
rect 13678 6898 13738 6974
rect 14414 7032 19031 7034
rect 14414 6976 18970 7032
rect 19026 6976 19031 7032
rect 14414 6974 19031 6976
rect 14414 6898 14474 6974
rect 18965 6971 19031 6974
rect 13678 6838 14474 6898
rect 0 6762 800 6792
rect 2730 6762 2790 6838
rect 6821 6835 6887 6838
rect 19425 6762 19491 6765
rect 0 6702 2790 6762
rect 5950 6760 19491 6762
rect 5950 6704 19430 6760
rect 19486 6704 19491 6760
rect 5950 6702 19491 6704
rect 0 6672 800 6702
rect 5950 6490 6010 6702
rect 19425 6699 19491 6702
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 6495 16858 6496
rect 1350 6430 6010 6490
rect 6913 6490 6979 6493
rect 11094 6490 11100 6492
rect 6913 6488 11100 6490
rect 6913 6432 6918 6488
rect 6974 6432 11100 6488
rect 6913 6430 11100 6432
rect 0 6218 800 6248
rect 1350 6218 1410 6430
rect 6913 6427 6979 6430
rect 11094 6428 11100 6430
rect 11164 6428 11170 6492
rect 1485 6354 1551 6357
rect 6361 6354 6427 6357
rect 12065 6354 12131 6357
rect 1485 6352 2790 6354
rect 1485 6296 1490 6352
rect 1546 6296 2790 6352
rect 1485 6294 2790 6296
rect 1485 6291 1551 6294
rect 0 6158 1410 6218
rect 2730 6218 2790 6294
rect 6361 6352 12131 6354
rect 6361 6296 6366 6352
rect 6422 6296 12070 6352
rect 12126 6296 12131 6352
rect 6361 6294 12131 6296
rect 6361 6291 6427 6294
rect 12065 6291 12131 6294
rect 6913 6218 6979 6221
rect 2730 6216 6979 6218
rect 2730 6160 6918 6216
rect 6974 6160 6979 6216
rect 2730 6158 6979 6160
rect 0 6128 800 6158
rect 6913 6155 6979 6158
rect 8477 6218 8543 6221
rect 8477 6216 9276 6218
rect 8477 6160 8482 6216
rect 8538 6160 9276 6216
rect 8477 6158 9276 6160
rect 8477 6155 8543 6158
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 9216 5946 9276 6158
rect 12065 6082 12131 6085
rect 12985 6082 13051 6085
rect 12065 6080 13051 6082
rect 12065 6024 12070 6080
rect 12126 6024 12990 6080
rect 13046 6024 13051 6080
rect 12065 6022 13051 6024
rect 12065 6019 12131 6022
rect 12985 6019 13051 6022
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 5951 19457 5952
rect 13261 5946 13327 5949
rect 9216 5944 13327 5946
rect 9216 5888 13266 5944
rect 13322 5888 13327 5944
rect 9216 5886 13327 5888
rect 13261 5883 13327 5886
rect 0 5810 800 5840
rect 2037 5810 2103 5813
rect 15929 5810 15995 5813
rect 0 5750 1594 5810
rect 0 5720 800 5750
rect 1534 5677 1594 5750
rect 2037 5808 15995 5810
rect 2037 5752 2042 5808
rect 2098 5752 15934 5808
rect 15990 5752 15995 5808
rect 2037 5750 15995 5752
rect 2037 5747 2103 5750
rect 15929 5747 15995 5750
rect 21449 5810 21515 5813
rect 22200 5810 23000 5840
rect 21449 5808 23000 5810
rect 21449 5752 21454 5808
rect 21510 5752 23000 5808
rect 21449 5750 23000 5752
rect 21449 5747 21515 5750
rect 22200 5720 23000 5750
rect 1534 5674 1643 5677
rect 4061 5674 4127 5677
rect 1534 5672 4127 5674
rect 1534 5616 1582 5672
rect 1638 5616 4066 5672
rect 4122 5616 4127 5672
rect 1534 5614 4127 5616
rect 1577 5611 1643 5614
rect 4061 5611 4127 5614
rect 4797 5674 4863 5677
rect 6862 5674 6868 5676
rect 4797 5672 6868 5674
rect 4797 5616 4802 5672
rect 4858 5616 6868 5672
rect 4797 5614 6868 5616
rect 4797 5611 4863 5614
rect 6862 5612 6868 5614
rect 6932 5612 6938 5676
rect 10225 5674 10291 5677
rect 18505 5674 18571 5677
rect 10225 5672 18571 5674
rect 10225 5616 10230 5672
rect 10286 5616 18510 5672
rect 18566 5616 18571 5672
rect 10225 5614 18571 5616
rect 10225 5611 10291 5614
rect 18505 5611 18571 5614
rect 17861 5538 17927 5541
rect 18505 5538 18571 5541
rect 17861 5536 18571 5538
rect 17861 5480 17866 5536
rect 17922 5480 18510 5536
rect 18566 5480 18571 5536
rect 17861 5478 18571 5480
rect 17861 5475 17927 5478
rect 18505 5475 18571 5478
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 16389 5402 16455 5405
rect 20345 5404 20411 5405
rect 11838 5400 16455 5402
rect 11838 5344 16394 5400
rect 16450 5344 16455 5400
rect 11838 5342 16455 5344
rect 0 5266 800 5296
rect 2773 5266 2839 5269
rect 0 5264 2839 5266
rect 0 5208 2778 5264
rect 2834 5208 2839 5264
rect 0 5206 2839 5208
rect 0 5176 800 5206
rect 2773 5203 2839 5206
rect 7649 5266 7715 5269
rect 11838 5266 11898 5342
rect 16389 5339 16455 5342
rect 20294 5340 20300 5404
rect 20364 5402 20411 5404
rect 20364 5400 20456 5402
rect 20406 5344 20456 5400
rect 20364 5342 20456 5344
rect 20364 5340 20411 5342
rect 20345 5339 20411 5340
rect 7649 5264 11898 5266
rect 7649 5208 7654 5264
rect 7710 5208 11898 5264
rect 7649 5206 11898 5208
rect 11973 5266 12039 5269
rect 18505 5266 18571 5269
rect 11973 5264 18571 5266
rect 11973 5208 11978 5264
rect 12034 5208 18510 5264
rect 18566 5208 18571 5264
rect 11973 5206 18571 5208
rect 7649 5203 7715 5206
rect 11973 5203 12039 5206
rect 18505 5203 18571 5206
rect 9029 5130 9095 5133
rect 17861 5130 17927 5133
rect 20437 5130 20503 5133
rect 2730 5128 17927 5130
rect 2730 5072 9034 5128
rect 9090 5072 17866 5128
rect 17922 5072 17927 5128
rect 2730 5070 17927 5072
rect 0 4858 800 4888
rect 2730 4858 2790 5070
rect 9029 5067 9095 5070
rect 17861 5067 17927 5070
rect 19014 5128 20503 5130
rect 19014 5072 20442 5128
rect 20498 5072 20503 5128
rect 19014 5070 20503 5072
rect 9622 4932 9628 4996
rect 9692 4994 9698 4996
rect 11973 4994 12039 4997
rect 9692 4992 12039 4994
rect 9692 4936 11978 4992
rect 12034 4936 12039 4992
rect 9692 4934 12039 4936
rect 9692 4932 9698 4934
rect 11973 4931 12039 4934
rect 16389 4994 16455 4997
rect 19014 4994 19074 5070
rect 20437 5067 20503 5070
rect 16389 4992 19074 4994
rect 16389 4936 16394 4992
rect 16450 4936 19074 4992
rect 16389 4934 19074 4936
rect 16389 4931 16455 4934
rect 3543 4928 3863 4929
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 0 4798 2790 4858
rect 3969 4858 4035 4861
rect 7598 4858 7604 4860
rect 3969 4856 7604 4858
rect 3969 4800 3974 4856
rect 4030 4800 7604 4856
rect 3969 4798 7604 4800
rect 0 4768 800 4798
rect 3969 4795 4035 4798
rect 7598 4796 7604 4798
rect 7668 4796 7674 4860
rect 9673 4858 9739 4861
rect 11973 4858 12039 4861
rect 13445 4858 13511 4861
rect 9673 4856 12039 4858
rect 9673 4800 9678 4856
rect 9734 4800 11978 4856
rect 12034 4800 12039 4856
rect 9673 4798 12039 4800
rect 9673 4795 9739 4798
rect 11973 4795 12039 4798
rect 12390 4856 13511 4858
rect 12390 4800 13450 4856
rect 13506 4800 13511 4856
rect 12390 4798 13511 4800
rect 12390 4722 12450 4798
rect 13445 4795 13511 4798
rect 5214 4662 12450 4722
rect 12617 4722 12683 4725
rect 18597 4722 18663 4725
rect 12617 4720 18663 4722
rect 12617 4664 12622 4720
rect 12678 4664 18602 4720
rect 18658 4664 18663 4720
rect 12617 4662 18663 4664
rect 0 4450 800 4480
rect 2957 4450 3023 4453
rect 0 4448 3023 4450
rect 0 4392 2962 4448
rect 3018 4392 3023 4448
rect 0 4390 3023 4392
rect 0 4360 800 4390
rect 2957 4387 3023 4390
rect 2129 4178 2195 4181
rect 5214 4178 5274 4662
rect 12617 4659 12683 4662
rect 18597 4659 18663 4662
rect 5441 4586 5507 4589
rect 15377 4586 15443 4589
rect 17769 4586 17835 4589
rect 5441 4584 15443 4586
rect 5441 4528 5446 4584
rect 5502 4528 15382 4584
rect 15438 4528 15443 4584
rect 5441 4526 15443 4528
rect 5441 4523 5507 4526
rect 15377 4523 15443 4526
rect 16254 4584 17835 4586
rect 16254 4528 17774 4584
rect 17830 4528 17835 4584
rect 16254 4526 17835 4528
rect 16254 4450 16314 4526
rect 17769 4523 17835 4526
rect 12390 4390 16314 4450
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 12390 4314 12450 4390
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 4319 16858 4320
rect 17217 4314 17283 4317
rect 11838 4254 12450 4314
rect 17174 4312 17283 4314
rect 17174 4256 17222 4312
rect 17278 4256 17283 4312
rect 2129 4176 5274 4178
rect 2129 4120 2134 4176
rect 2190 4120 5274 4176
rect 2129 4118 5274 4120
rect 2129 4115 2195 4118
rect 7598 4116 7604 4180
rect 7668 4178 7674 4180
rect 9857 4178 9923 4181
rect 10409 4178 10475 4181
rect 7668 4118 9506 4178
rect 7668 4116 7674 4118
rect 2221 4044 2287 4045
rect 3969 4044 4035 4045
rect 2221 4040 2268 4044
rect 2332 4042 2338 4044
rect 2221 3984 2226 4040
rect 2221 3980 2268 3984
rect 2332 3982 2378 4042
rect 2332 3980 2338 3982
rect 3918 3980 3924 4044
rect 3988 4042 4035 4044
rect 3988 4040 4080 4042
rect 4030 3984 4080 4040
rect 3988 3982 4080 3984
rect 3988 3980 4035 3982
rect 6862 3980 6868 4044
rect 6932 4042 6938 4044
rect 8109 4042 8175 4045
rect 9446 4042 9506 4118
rect 9857 4176 10475 4178
rect 9857 4120 9862 4176
rect 9918 4120 10414 4176
rect 10470 4120 10475 4176
rect 9857 4118 10475 4120
rect 9857 4115 9923 4118
rect 10409 4115 10475 4118
rect 10777 4178 10843 4181
rect 11838 4178 11898 4254
rect 17174 4251 17283 4256
rect 10777 4176 11898 4178
rect 10777 4120 10782 4176
rect 10838 4120 11898 4176
rect 10777 4118 11898 4120
rect 11973 4178 12039 4181
rect 17174 4178 17234 4251
rect 11973 4176 19626 4178
rect 11973 4120 11978 4176
rect 12034 4120 19626 4176
rect 11973 4118 19626 4120
rect 10777 4115 10843 4118
rect 11973 4115 12039 4118
rect 10869 4042 10935 4045
rect 6932 4040 9276 4042
rect 6932 3984 8114 4040
rect 8170 3984 9276 4040
rect 6932 3982 9276 3984
rect 9446 4040 10935 4042
rect 9446 3984 10874 4040
rect 10930 3984 10935 4040
rect 9446 3982 10935 3984
rect 6932 3980 6938 3982
rect 2221 3979 2287 3980
rect 3969 3979 4035 3980
rect 8109 3979 8175 3982
rect 0 3906 800 3936
rect 3417 3906 3483 3909
rect 0 3904 3483 3906
rect 0 3848 3422 3904
rect 3478 3848 3483 3904
rect 0 3846 3483 3848
rect 9216 3906 9276 3982
rect 10869 3979 10935 3982
rect 11053 4042 11119 4045
rect 17769 4042 17835 4045
rect 11053 4040 17835 4042
rect 11053 3984 11058 4040
rect 11114 3984 17774 4040
rect 17830 3984 17835 4040
rect 11053 3982 17835 3984
rect 11053 3979 11119 3982
rect 17769 3979 17835 3982
rect 18689 4042 18755 4045
rect 19241 4042 19307 4045
rect 18689 4040 19307 4042
rect 18689 3984 18694 4040
rect 18750 3984 19246 4040
rect 19302 3984 19307 4040
rect 18689 3982 19307 3984
rect 18689 3979 18755 3982
rect 19241 3979 19307 3982
rect 12065 3906 12131 3909
rect 13721 3906 13787 3909
rect 9216 3904 12131 3906
rect 9216 3848 12070 3904
rect 12126 3848 12131 3904
rect 9216 3846 12131 3848
rect 0 3816 800 3846
rect 3417 3843 3483 3846
rect 12065 3843 12131 3846
rect 12390 3904 13787 3906
rect 12390 3848 13726 3904
rect 13782 3848 13787 3904
rect 12390 3846 13787 3848
rect 19566 3906 19626 4118
rect 19885 4044 19951 4045
rect 19885 4042 19932 4044
rect 19840 4040 19932 4042
rect 19840 3984 19890 4040
rect 19840 3982 19932 3984
rect 19885 3980 19932 3982
rect 19996 3980 20002 4044
rect 19885 3979 19951 3980
rect 19885 3906 19951 3909
rect 19566 3904 19951 3906
rect 19566 3848 19890 3904
rect 19946 3848 19951 3904
rect 19566 3846 19951 3848
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 10869 3770 10935 3773
rect 12390 3770 12450 3846
rect 13721 3843 13787 3846
rect 19885 3843 19951 3846
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 10869 3768 12450 3770
rect 10869 3712 10874 3768
rect 10930 3712 12450 3768
rect 10869 3710 12450 3712
rect 15929 3770 15995 3773
rect 18413 3770 18479 3773
rect 15929 3768 18479 3770
rect 15929 3712 15934 3768
rect 15990 3712 18418 3768
rect 18474 3712 18479 3768
rect 15929 3710 18479 3712
rect 10869 3707 10935 3710
rect 15929 3707 15995 3710
rect 18413 3707 18479 3710
rect 5993 3634 6059 3637
rect 18597 3634 18663 3637
rect 5993 3632 18663 3634
rect 5993 3576 5998 3632
rect 6054 3576 18602 3632
rect 18658 3576 18663 3632
rect 5993 3574 18663 3576
rect 5993 3571 6059 3574
rect 18597 3571 18663 3574
rect 0 3498 800 3528
rect 3049 3498 3115 3501
rect 4102 3498 4108 3500
rect 0 3496 4108 3498
rect 0 3440 3054 3496
rect 3110 3440 4108 3496
rect 0 3438 4108 3440
rect 0 3408 800 3438
rect 3049 3435 3115 3438
rect 4102 3436 4108 3438
rect 4172 3436 4178 3500
rect 10041 3498 10107 3501
rect 5950 3496 10107 3498
rect 5950 3440 10046 3496
rect 10102 3440 10107 3496
rect 5950 3438 10107 3440
rect 1485 3362 1551 3365
rect 5533 3362 5599 3365
rect 1485 3360 5599 3362
rect 1485 3304 1490 3360
rect 1546 3304 5538 3360
rect 5594 3304 5599 3360
rect 1485 3302 5599 3304
rect 1485 3299 1551 3302
rect 5533 3299 5599 3302
rect 2446 3164 2452 3228
rect 2516 3226 2522 3228
rect 2681 3226 2747 3229
rect 2516 3224 2747 3226
rect 2516 3168 2686 3224
rect 2742 3168 2747 3224
rect 2516 3166 2747 3168
rect 2516 3164 2522 3166
rect 2681 3163 2747 3166
rect 3417 3226 3483 3229
rect 5950 3226 6010 3438
rect 10041 3435 10107 3438
rect 11697 3498 11763 3501
rect 16941 3498 17007 3501
rect 11697 3496 17007 3498
rect 11697 3440 11702 3496
rect 11758 3440 16946 3496
rect 17002 3440 17007 3496
rect 11697 3438 17007 3440
rect 11697 3435 11763 3438
rect 16941 3435 17007 3438
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 3231 16858 3232
rect 3417 3224 6010 3226
rect 3417 3168 3422 3224
rect 3478 3168 6010 3224
rect 3417 3166 6010 3168
rect 3417 3163 3483 3166
rect 6678 3164 6684 3228
rect 6748 3226 6754 3228
rect 6821 3226 6887 3229
rect 15193 3226 15259 3229
rect 6748 3224 6887 3226
rect 6748 3168 6826 3224
rect 6882 3168 6887 3224
rect 6748 3166 6887 3168
rect 6748 3164 6754 3166
rect 6821 3163 6887 3166
rect 11838 3224 15259 3226
rect 11838 3168 15198 3224
rect 15254 3168 15259 3224
rect 11838 3166 15259 3168
rect 2773 3090 2839 3093
rect 11838 3090 11898 3166
rect 15193 3163 15259 3166
rect 13537 3090 13603 3093
rect 2638 3088 11898 3090
rect 2638 3032 2778 3088
rect 2834 3032 11898 3088
rect 2638 3030 11898 3032
rect 11976 3088 13603 3090
rect 11976 3032 13542 3088
rect 13598 3032 13603 3088
rect 11976 3030 13603 3032
rect 0 2954 800 2984
rect 2638 2954 2698 3030
rect 2773 3027 2839 3030
rect 0 2894 2698 2954
rect 3877 2954 3943 2957
rect 11976 2954 12036 3030
rect 13537 3027 13603 3030
rect 3877 2952 12036 2954
rect 3877 2896 3882 2952
rect 3938 2896 12036 2952
rect 3877 2894 12036 2896
rect 12341 2954 12407 2957
rect 18689 2954 18755 2957
rect 12341 2952 18755 2954
rect 12341 2896 12346 2952
rect 12402 2896 18694 2952
rect 18750 2896 18755 2952
rect 12341 2894 18755 2896
rect 0 2864 800 2894
rect 3877 2891 3943 2894
rect 12341 2891 12407 2894
rect 18689 2891 18755 2894
rect 1945 2818 2011 2821
rect 3417 2818 3483 2821
rect 1945 2816 3483 2818
rect 1945 2760 1950 2816
rect 2006 2760 3422 2816
rect 3478 2760 3483 2816
rect 1945 2758 3483 2760
rect 1945 2755 2011 2758
rect 3417 2755 3483 2758
rect 9673 2818 9739 2821
rect 10961 2818 11027 2821
rect 13721 2818 13787 2821
rect 9673 2816 13787 2818
rect 9673 2760 9678 2816
rect 9734 2760 10966 2816
rect 11022 2760 13726 2816
rect 13782 2760 13787 2816
rect 9673 2758 13787 2760
rect 9673 2755 9739 2758
rect 10961 2755 11027 2758
rect 13721 2755 13787 2758
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 4470 2620 4476 2684
rect 4540 2682 4546 2684
rect 4981 2682 5047 2685
rect 4540 2680 5047 2682
rect 4540 2624 4986 2680
rect 5042 2624 5047 2680
rect 4540 2622 5047 2624
rect 4540 2620 4546 2622
rect 4981 2619 5047 2622
rect 11145 2682 11211 2685
rect 12065 2682 12131 2685
rect 11145 2680 12131 2682
rect 11145 2624 11150 2680
rect 11206 2624 12070 2680
rect 12126 2624 12131 2680
rect 11145 2622 12131 2624
rect 11145 2619 11211 2622
rect 12065 2619 12131 2622
rect 15377 2682 15443 2685
rect 16205 2682 16271 2685
rect 18505 2682 18571 2685
rect 15377 2680 18571 2682
rect 15377 2624 15382 2680
rect 15438 2624 16210 2680
rect 16266 2624 18510 2680
rect 18566 2624 18571 2680
rect 15377 2622 18571 2624
rect 15377 2619 15443 2622
rect 16205 2619 16271 2622
rect 18505 2619 18571 2622
rect 0 2546 800 2576
rect 1393 2546 1459 2549
rect 3141 2546 3207 2549
rect 0 2544 3207 2546
rect 0 2488 1398 2544
rect 1454 2488 3146 2544
rect 3202 2488 3207 2544
rect 0 2486 3207 2488
rect 0 2456 800 2486
rect 1393 2483 1459 2486
rect 3141 2483 3207 2486
rect 3325 2546 3391 2549
rect 18873 2546 18939 2549
rect 3325 2544 18939 2546
rect 3325 2488 3330 2544
rect 3386 2488 18878 2544
rect 18934 2488 18939 2544
rect 3325 2486 18939 2488
rect 3325 2483 3391 2486
rect 18873 2483 18939 2486
rect 2497 2410 2563 2413
rect 10593 2410 10659 2413
rect 10961 2410 11027 2413
rect 11973 2410 12039 2413
rect 2497 2408 6930 2410
rect 2497 2352 2502 2408
rect 2558 2352 6930 2408
rect 2497 2350 6930 2352
rect 2497 2347 2563 2350
rect 6870 2274 6930 2350
rect 10593 2408 12039 2410
rect 10593 2352 10598 2408
rect 10654 2352 10966 2408
rect 11022 2352 11978 2408
rect 12034 2352 12039 2408
rect 10593 2350 12039 2352
rect 10593 2347 10659 2350
rect 10961 2347 11027 2350
rect 11973 2347 12039 2350
rect 11145 2274 11211 2277
rect 6870 2272 11211 2274
rect 6870 2216 11150 2272
rect 11206 2216 11211 2272
rect 6870 2214 11211 2216
rect 11145 2211 11211 2214
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 2129 2138 2195 2141
rect 798 2136 2195 2138
rect 798 2080 2134 2136
rect 2190 2080 2195 2136
rect 798 2078 2195 2080
rect 798 2032 858 2078
rect 2129 2075 2195 2078
rect 0 1942 858 2032
rect 1025 2002 1091 2005
rect 17309 2002 17375 2005
rect 1025 2000 17375 2002
rect 1025 1944 1030 2000
rect 1086 1944 17314 2000
rect 17370 1944 17375 2000
rect 1025 1942 17375 1944
rect 0 1912 800 1942
rect 1025 1939 1091 1942
rect 17309 1939 17375 1942
rect 5942 1804 5948 1868
rect 6012 1866 6018 1868
rect 6361 1866 6427 1869
rect 6012 1864 6427 1866
rect 6012 1808 6366 1864
rect 6422 1808 6427 1864
rect 6012 1806 6427 1808
rect 6012 1804 6018 1806
rect 6361 1803 6427 1806
rect 1485 1730 1551 1733
rect 15377 1730 15443 1733
rect 1485 1728 15443 1730
rect 1485 1672 1490 1728
rect 1546 1672 15382 1728
rect 15438 1672 15443 1728
rect 1485 1670 15443 1672
rect 1485 1667 1551 1670
rect 15377 1667 15443 1670
rect 0 1594 800 1624
rect 4061 1594 4127 1597
rect 0 1592 4127 1594
rect 0 1536 4066 1592
rect 4122 1536 4127 1592
rect 0 1534 4127 1536
rect 0 1504 800 1534
rect 4061 1531 4127 1534
rect 0 1050 800 1080
rect 4521 1050 4587 1053
rect 13302 1050 13308 1052
rect 0 1048 13308 1050
rect 0 992 4526 1048
rect 4582 992 13308 1048
rect 0 990 13308 992
rect 0 960 800 990
rect 4521 987 4587 990
rect 13302 988 13308 990
rect 13372 988 13378 1052
rect 0 642 800 672
rect 2865 642 2931 645
rect 0 640 2931 642
rect 0 584 2870 640
rect 2926 584 2931 640
rect 0 582 2931 584
rect 0 552 800 582
rect 2865 579 2931 582
rect 0 234 800 264
rect 2957 234 3023 237
rect 0 232 3023 234
rect 0 176 2962 232
rect 3018 176 3023 232
rect 0 174 3023 176
rect 0 144 800 174
rect 2957 171 3023 174
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 19932 17580 19996 17644
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 3924 12820 3988 12884
rect 11100 12548 11164 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 1716 11732 1780 11796
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 2268 11052 2332 11116
rect 13308 11112 13372 11116
rect 13308 11056 13322 11112
rect 13322 11056 13372 11112
rect 13308 11052 13372 11056
rect 14412 11052 14476 11116
rect 20300 11052 20364 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 1716 9148 1780 9212
rect 2452 8876 2516 8940
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 6684 8332 6748 8396
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 4476 7788 4540 7852
rect 7604 7788 7668 7852
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 5948 7244 6012 7308
rect 9628 7244 9692 7308
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 11100 6428 11164 6492
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 6868 5612 6932 5676
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 20300 5400 20364 5404
rect 20300 5344 20350 5400
rect 20350 5344 20364 5400
rect 20300 5340 20364 5344
rect 9628 4932 9692 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 7604 4796 7668 4860
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 7604 4116 7668 4180
rect 2268 4040 2332 4044
rect 2268 3984 2282 4040
rect 2282 3984 2332 4040
rect 2268 3980 2332 3984
rect 3924 4040 3988 4044
rect 3924 3984 3974 4040
rect 3974 3984 3988 4040
rect 3924 3980 3988 3984
rect 6868 3980 6932 4044
rect 19932 4040 19996 4044
rect 19932 3984 19946 4040
rect 19946 3984 19996 4040
rect 19932 3980 19996 3984
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 4108 3436 4172 3500
rect 2452 3164 2516 3228
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 6684 3164 6748 3228
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 4476 2620 4540 2684
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 5948 1804 6012 1868
rect 13308 988 13372 1052
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 3923 12884 3989 12885
rect 3923 12820 3924 12884
rect 3988 12820 3989 12884
rect 3923 12819 3989 12820
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 1715 11796 1781 11797
rect 1715 11732 1716 11796
rect 1780 11732 1781 11796
rect 1715 11731 1781 11732
rect 1718 9213 1778 11731
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 2267 11116 2333 11117
rect 2267 11052 2268 11116
rect 2332 11052 2333 11116
rect 2267 11051 2333 11052
rect 1715 9212 1781 9213
rect 1715 9148 1716 9212
rect 1780 9148 1781 9212
rect 1715 9147 1781 9148
rect 2270 4045 2330 11051
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 2451 8940 2517 8941
rect 2451 8876 2452 8940
rect 2516 8876 2517 8940
rect 2451 8875 2517 8876
rect 2267 4044 2333 4045
rect 2267 3980 2268 4044
rect 2332 3980 2333 4044
rect 2267 3979 2333 3980
rect 2454 3229 2514 8875
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3926 4045 3986 12819
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 4475 7852 4541 7853
rect 4475 7788 4476 7852
rect 4540 7788 4541 7852
rect 4475 7787 4541 7788
rect 3923 4044 3989 4045
rect 3923 3980 3924 4044
rect 3988 3980 3989 4044
rect 3923 3979 3989 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 2451 3228 2517 3229
rect 2451 3164 2452 3228
rect 2516 3164 2517 3228
rect 2451 3163 2517 3164
rect 3543 2752 3863 3776
rect 4110 3501 4170 3622
rect 4107 3500 4173 3501
rect 4107 3436 4108 3500
rect 4172 3436 4173 3500
rect 4107 3435 4173 3436
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 4478 2685 4538 7787
rect 6142 7648 6462 8672
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11099 12612 11165 12613
rect 11099 12548 11100 12612
rect 11164 12548 11165 12612
rect 11099 12547 11165 12548
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 6683 8396 6749 8397
rect 6683 8332 6684 8396
rect 6748 8332 6749 8396
rect 6683 8331 6749 8332
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 5947 7308 6013 7309
rect 5947 7244 5948 7308
rect 6012 7244 6013 7308
rect 5947 7243 6013 7244
rect 4475 2684 4541 2685
rect 4475 2620 4476 2684
rect 4540 2620 4541 2684
rect 4475 2619 4541 2620
rect 5950 1869 6010 7243
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6686 3229 6746 8331
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 7603 7852 7669 7853
rect 7603 7788 7604 7852
rect 7668 7788 7669 7852
rect 7603 7787 7669 7788
rect 6867 5676 6933 5677
rect 6867 5612 6868 5676
rect 6932 5612 6933 5676
rect 6867 5611 6933 5612
rect 6870 4045 6930 5611
rect 7606 4861 7666 7787
rect 8741 7104 9061 8128
rect 9627 7308 9693 7309
rect 9627 7244 9628 7308
rect 9692 7244 9693 7308
rect 9627 7243 9693 7244
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 9630 4997 9690 7243
rect 11102 6493 11162 12547
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13307 11116 13373 11117
rect 13307 11052 13308 11116
rect 13372 11052 13373 11116
rect 13307 11051 13373 11052
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11099 6492 11165 6493
rect 11099 6428 11100 6492
rect 11164 6428 11165 6492
rect 11099 6427 11165 6428
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 9627 4996 9693 4997
rect 9627 4932 9628 4996
rect 9692 4932 9693 4996
rect 9627 4931 9693 4932
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 7603 4860 7669 4861
rect 7603 4796 7604 4860
rect 7668 4796 7669 4860
rect 7603 4795 7669 4796
rect 7606 4181 7666 4795
rect 7603 4180 7669 4181
rect 7603 4116 7604 4180
rect 7668 4116 7669 4180
rect 7603 4115 7669 4116
rect 6867 4044 6933 4045
rect 6867 3980 6868 4044
rect 6932 3980 6933 4044
rect 6867 3979 6933 3980
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 6683 3228 6749 3229
rect 6683 3164 6684 3228
rect 6748 3164 6749 3228
rect 6683 3163 6749 3164
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 5947 1868 6013 1869
rect 5947 1804 5948 1868
rect 6012 1804 6013 1868
rect 5947 1803 6013 1804
rect 13310 1053 13370 11051
rect 13939 10368 14259 11392
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 14411 11116 14477 11117
rect 14411 11052 14412 11116
rect 14476 11052 14477 11116
rect 14411 11051 14477 11052
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 14414 3858 14474 11051
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19931 17644 19997 17645
rect 19931 17580 19932 17644
rect 19996 17580 19997 17644
rect 19931 17579 19997 17580
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19934 4045 19994 17579
rect 20299 11116 20365 11117
rect 20299 11052 20300 11116
rect 20364 11052 20365 11116
rect 20299 11051 20365 11052
rect 20302 5405 20362 11051
rect 20299 5404 20365 5405
rect 20299 5340 20300 5404
rect 20364 5340 20365 5404
rect 20299 5339 20365 5340
rect 19931 4044 19997 4045
rect 19931 3980 19932 4044
rect 19996 3980 19997 4044
rect 19931 3979 19997 3980
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 13307 1052 13373 1053
rect 13307 988 13308 1052
rect 13372 988 13373 1052
rect 13307 987 13373 988
<< via4 >>
rect 4022 3622 4258 3858
rect 14326 3622 14562 3858
<< metal5 >>
rect 3980 3858 14604 3900
rect 3980 3622 4022 3858
rect 4258 3622 14326 3858
rect 14562 3622 14604 3858
rect 3980 3580 14604 3622
use sky130_fd_sc_hd__diode_2  ANTENNA__108__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19872 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform 1 0 10580 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 16836 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 13708 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 6532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 6992 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform 1 0 4232 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 1564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 20792 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 9568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 18676 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 17848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 21160 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 14996 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 18032 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 16284 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 4876 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 3312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 4968 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5980 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6992 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8188 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 10488 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12604 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp 1649977179
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_149
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_155
timestamp 1649977179
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_161
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 1649977179
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_207
timestamp 1649977179
transform 1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_18
timestamp 1649977179
transform 1 0 2760 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1649977179
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_83
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_119
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 1649977179
transform 1 0 14628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_157
timestamp 1649977179
transform 1 0 15548 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_179
timestamp 1649977179
transform 1 0 17572 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_197
timestamp 1649977179
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_201
timestamp 1649977179
transform 1 0 19596 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1649977179
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_43
timestamp 1649977179
transform 1 0 5060 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_60
timestamp 1649977179
transform 1 0 6624 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_99
timestamp 1649977179
transform 1 0 10212 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_150
timestamp 1649977179
transform 1 0 14904 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_161
timestamp 1649977179
transform 1 0 15916 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_171
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_181
timestamp 1649977179
transform 1 0 17756 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_186
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_191
timestamp 1649977179
transform 1 0 18676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_199
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_205
timestamp 1649977179
transform 1 0 19964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_211
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_25
timestamp 1649977179
transform 1 0 3404 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_32
timestamp 1649977179
transform 1 0 4048 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_43
timestamp 1649977179
transform 1 0 5060 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_80
timestamp 1649977179
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_92
timestamp 1649977179
transform 1 0 9568 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_103
timestamp 1649977179
transform 1 0 10580 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_142
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_160
timestamp 1649977179
transform 1 0 15824 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_165
timestamp 1649977179
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_178
timestamp 1649977179
transform 1 0 17480 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_182
timestamp 1649977179
transform 1 0 17848 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_192
timestamp 1649977179
transform 1 0 18768 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_197
timestamp 1649977179
transform 1 0 19228 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_202
timestamp 1649977179
transform 1 0 19688 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_207
timestamp 1649977179
transform 1 0 20148 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_214
timestamp 1649977179
transform 1 0 20792 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 1649977179
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_25
timestamp 1649977179
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_45
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_70
timestamp 1649977179
transform 1 0 7544 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1649977179
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_88
timestamp 1649977179
transform 1 0 9200 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_99
timestamp 1649977179
transform 1 0 10212 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_118
timestamp 1649977179
transform 1 0 11960 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 1649977179
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1649977179
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 1649977179
transform 1 0 16468 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_185
timestamp 1649977179
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_190
timestamp 1649977179
transform 1 0 18584 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1649977179
transform 1 0 19504 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_204
timestamp 1649977179
transform 1 0 19872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_13
timestamp 1649977179
transform 1 0 2300 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_17
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_5_73
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_84
timestamp 1649977179
transform 1 0 8832 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_89
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_107
timestamp 1649977179
transform 1 0 10948 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_116
timestamp 1649977179
transform 1 0 11776 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 1649977179
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_183
timestamp 1649977179
transform 1 0 17940 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_188
timestamp 1649977179
transform 1 0 18400 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_198
timestamp 1649977179
transform 1 0 19320 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_203
timestamp 1649977179
transform 1 0 19780 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_208
timestamp 1649977179
transform 1 0 20240 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_213
timestamp 1649977179
transform 1 0 20700 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_38
timestamp 1649977179
transform 1 0 4600 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_43
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_70
timestamp 1649977179
transform 1 0 7544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1649977179
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_88
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_131
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_136
timestamp 1649977179
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_6_149
timestamp 1649977179
transform 1 0 14812 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 1649977179
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_164
timestamp 1649977179
transform 1 0 16192 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_168
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_185
timestamp 1649977179
transform 1 0 18124 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_190
timestamp 1649977179
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_200
timestamp 1649977179
transform 1 0 19504 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1649977179
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_210
timestamp 1649977179
transform 1 0 20424 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_215
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_220
timestamp 1649977179
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_18
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 1649977179
transform 1 0 4416 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_95
timestamp 1649977179
transform 1 0 9844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1649977179
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_119
timestamp 1649977179
transform 1 0 12052 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_141
timestamp 1649977179
transform 1 0 14076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_151
timestamp 1649977179
transform 1 0 14996 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_155
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_183
timestamp 1649977179
transform 1 0 17940 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_188
timestamp 1649977179
transform 1 0 18400 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_198
timestamp 1649977179
transform 1 0 19320 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_203
timestamp 1649977179
transform 1 0 19780 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_212
timestamp 1649977179
transform 1 0 20608 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_216
timestamp 1649977179
transform 1 0 20976 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_38
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_43
timestamp 1649977179
transform 1 0 5060 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_78
timestamp 1649977179
transform 1 0 8280 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_104
timestamp 1649977179
transform 1 0 10672 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_116
timestamp 1649977179
transform 1 0 11776 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_126
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_157
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_180
timestamp 1649977179
transform 1 0 17664 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 1649977179
transform 1 0 18584 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_200
timestamp 1649977179
transform 1 0 19504 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_205
timestamp 1649977179
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_210
timestamp 1649977179
transform 1 0 20424 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_214
timestamp 1649977179
transform 1 0 20792 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_218
timestamp 1649977179
transform 1 0 21160 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_5
timestamp 1649977179
transform 1 0 1564 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_23
timestamp 1649977179
transform 1 0 3220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_32
timestamp 1649977179
transform 1 0 4048 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_89
timestamp 1649977179
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_100
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_129
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_141
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_159
timestamp 1649977179
transform 1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_164
timestamp 1649977179
transform 1 0 16192 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_177
timestamp 1649977179
transform 1 0 17388 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_182
timestamp 1649977179
transform 1 0 17848 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_187
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_192
timestamp 1649977179
transform 1 0 18768 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_201
timestamp 1649977179
transform 1 0 19596 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_213
timestamp 1649977179
transform 1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp 1649977179
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_76
timestamp 1649977179
transform 1 0 8096 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 1649977179
transform 1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1649977179
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_136
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_152
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_162
timestamp 1649977179
transform 1 0 16008 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_182
timestamp 1649977179
transform 1 0 17848 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_191
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_199 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_217
timestamp 1649977179
transform 1 0 21068 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_29
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_34
timestamp 1649977179
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_52
timestamp 1649977179
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_95
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_108
timestamp 1649977179
transform 1 0 11040 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_122
timestamp 1649977179
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_134
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_152
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_157
timestamp 1649977179
transform 1 0 15548 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 1649977179
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 1649977179
transform 1 0 16928 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1649977179
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_18
timestamp 1649977179
transform 1 0 2760 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_22
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_52
timestamp 1649977179
transform 1 0 5888 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_63
timestamp 1649977179
transform 1 0 6900 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1649977179
transform 1 0 9200 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_102
timestamp 1649977179
transform 1 0 10488 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_117
timestamp 1649977179
transform 1 0 11868 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_129
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_167
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 1649977179
transform 1 0 16836 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_176
timestamp 1649977179
transform 1 0 17296 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_180
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_184
timestamp 1649977179
transform 1 0 18032 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_20
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_31
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_43
timestamp 1649977179
transform 1 0 5060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_64
timestamp 1649977179
transform 1 0 6992 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_75
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_88
timestamp 1649977179
transform 1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_99
timestamp 1649977179
transform 1 0 10212 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_139
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_150
timestamp 1649977179
transform 1 0 14904 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_160
timestamp 1649977179
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_183
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_195
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_207
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_14
timestamp 1649977179
transform 1 0 2392 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 1649977179
transform 1 0 3404 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_31
timestamp 1649977179
transform 1 0 3956 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_58
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_92
timestamp 1649977179
transform 1 0 9568 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_110
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_144
timestamp 1649977179
transform 1 0 14352 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_149
timestamp 1649977179
transform 1 0 14812 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_22
timestamp 1649977179
transform 1 0 3128 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_31
timestamp 1649977179
transform 1 0 3956 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_53
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1649977179
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_75
timestamp 1649977179
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_86
timestamp 1649977179
transform 1 0 9016 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_109
timestamp 1649977179
transform 1 0 11132 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1649977179
transform 1 0 13524 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_145
timestamp 1649977179
transform 1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_190
timestamp 1649977179
transform 1 0 18584 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_202
timestamp 1649977179
transform 1 0 19688 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_214 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_222
timestamp 1649977179
transform 1 0 21528 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_6
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_36
timestamp 1649977179
transform 1 0 4416 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_58
timestamp 1649977179
transform 1 0 6440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_62
timestamp 1649977179
transform 1 0 6808 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_87
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_98
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_108
timestamp 1649977179
transform 1 0 11040 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_118
timestamp 1649977179
transform 1 0 11960 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_137
timestamp 1649977179
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_147
timestamp 1649977179
transform 1 0 14628 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_151
timestamp 1649977179
transform 1 0 14996 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_163
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_175
timestamp 1649977179
transform 1 0 17204 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_187
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_200
timestamp 1649977179
transform 1 0 19504 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_212
timestamp 1649977179
transform 1 0 20608 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_220
timestamp 1649977179
transform 1 0 21344 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_18
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_36
timestamp 1649977179
transform 1 0 4416 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_41
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1649977179
transform 1 0 7544 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_121
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_126
timestamp 1649977179
transform 1 0 12696 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_130
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_134
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_138
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_142
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_154
timestamp 1649977179
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_204
timestamp 1649977179
transform 1 0 19872 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_222
timestamp 1649977179
transform 1 0 21528 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_9
timestamp 1649977179
transform 1 0 1932 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_20
timestamp 1649977179
transform 1 0 2944 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_38
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_56
timestamp 1649977179
transform 1 0 6256 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_76
timestamp 1649977179
transform 1 0 8096 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_87
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_92
timestamp 1649977179
transform 1 0 9568 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_110
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_124
timestamp 1649977179
transform 1 0 12512 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_128
timestamp 1649977179
transform 1 0 12880 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_132
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_201
timestamp 1649977179
transform 1 0 19596 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_205
timestamp 1649977179
transform 1 0 19964 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_217
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_11
timestamp 1649977179
transform 1 0 2116 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1649977179
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_30
timestamp 1649977179
transform 1 0 3864 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_48
timestamp 1649977179
transform 1 0 5520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 1649977179
transform 1 0 5980 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1649977179
transform 1 0 6532 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_70
timestamp 1649977179
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_104
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 1649977179
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_115
timestamp 1649977179
transform 1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_119
timestamp 1649977179
transform 1 0 12052 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_131
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_143
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_155
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_13
timestamp 1649977179
transform 1 0 2300 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_17
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_31
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_42
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1649977179
transform 1 0 7544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_94
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_112
timestamp 1649977179
transform 1 0 11408 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_122
timestamp 1649977179
transform 1 0 12328 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_134
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_17
timestamp 1649977179
transform 1 0 2668 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_28
timestamp 1649977179
transform 1 0 3680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_46
timestamp 1649977179
transform 1 0 5336 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_60
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_79
timestamp 1649977179
transform 1 0 8372 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_92
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_103
timestamp 1649977179
transform 1 0 10580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_108
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_17
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_33
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_51
timestamp 1649977179
transform 1 0 5796 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_61
timestamp 1649977179
transform 1 0 6716 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_89
timestamp 1649977179
transform 1 0 9292 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_117
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_137
timestamp 1649977179
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_11
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_16
timestamp 1649977179
transform 1 0 2576 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_26
timestamp 1649977179
transform 1 0 3496 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_64
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_75
timestamp 1649977179
transform 1 0 8004 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_79
timestamp 1649977179
transform 1 0 8372 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_92
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_16
timestamp 1649977179
transform 1 0 2576 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_26
timestamp 1649977179
transform 1 0 3496 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_32
timestamp 1649977179
transform 1 0 4048 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_43
timestamp 1649977179
transform 1 0 5060 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_55
timestamp 1649977179
transform 1 0 6164 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_75
timestamp 1649977179
transform 1 0 8004 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_79
timestamp 1649977179
transform 1 0 8372 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_111
timestamp 1649977179
transform 1 0 11316 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_123
timestamp 1649977179
transform 1 0 12420 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_135
timestamp 1649977179
transform 1 0 13524 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_17
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_47
timestamp 1649977179
transform 1 0 5428 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_70
timestamp 1649977179
transform 1 0 7544 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_99
timestamp 1649977179
transform 1 0 10212 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_122
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_134
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_146
timestamp 1649977179
transform 1 0 14536 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_158
timestamp 1649977179
transform 1 0 15640 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_18
timestamp 1649977179
transform 1 0 2760 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_23
timestamp 1649977179
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_43
timestamp 1649977179
transform 1 0 5060 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_61
timestamp 1649977179
transform 1 0 6716 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_71
timestamp 1649977179
transform 1 0 7636 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_94
timestamp 1649977179
transform 1 0 9752 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1649977179
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_102
timestamp 1649977179
transform 1 0 10488 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_17
timestamp 1649977179
transform 1 0 2668 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_23
timestamp 1649977179
transform 1 0 3220 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_33
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_91
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_129
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_141
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_153
timestamp 1649977179
transform 1 0 15180 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1649977179
transform 1 0 2668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_51
timestamp 1649977179
transform 1 0 5796 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_62
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_72
timestamp 1649977179
transform 1 0 7728 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_94
timestamp 1649977179
transform 1 0 9752 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_105
timestamp 1649977179
transform 1 0 10764 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_116
timestamp 1649977179
transform 1 0 11776 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_125
timestamp 1649977179
transform 1 0 12604 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1649977179
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_18
timestamp 1649977179
transform 1 0 2760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_23
timestamp 1649977179
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_28
timestamp 1649977179
transform 1 0 3680 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_38
timestamp 1649977179
transform 1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_42
timestamp 1649977179
transform 1 0 4968 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_66
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_76
timestamp 1649977179
transform 1 0 8096 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_29_82
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_88
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1649977179
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_102
timestamp 1649977179
transform 1 0 10488 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_106
timestamp 1649977179
transform 1 0 10856 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1649977179
transform 1 0 11224 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_116
timestamp 1649977179
transform 1 0 11776 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_128
timestamp 1649977179
transform 1 0 12880 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_140
timestamp 1649977179
transform 1 0 13984 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_152
timestamp 1649977179
transform 1 0 15088 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1649977179
transform 1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_32
timestamp 1649977179
transform 1 0 4048 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_37
timestamp 1649977179
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_42
timestamp 1649977179
transform 1 0 4968 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_50
timestamp 1649977179
transform 1 0 5704 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_61
timestamp 1649977179
transform 1 0 6716 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_64
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_76
timestamp 1649977179
transform 1 0 8096 0 1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_101
timestamp 1649977179
transform 1 0 10396 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_105
timestamp 1649977179
transform 1 0 10764 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_117
timestamp 1649977179
transform 1 0 11868 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_129
timestamp 1649977179
transform 1 0 12972 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_137
timestamp 1649977179
transform 1 0 13708 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_28
timestamp 1649977179
transform 1 0 3680 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_33
timestamp 1649977179
transform 1 0 4140 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_38
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_50
timestamp 1649977179
transform 1 0 5704 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_19
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_32
timestamp 1649977179
transform 1 0 4048 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_37
timestamp 1649977179
transform 1 0 4508 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_42
timestamp 1649977179
transform 1 0 4968 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_54
timestamp 1649977179
transform 1 0 6072 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_66
timestamp 1649977179
transform 1 0 7176 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_78
timestamp 1649977179
transform 1 0 8280 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_25
timestamp 1649977179
transform 1 0 3404 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1649977179
transform 1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1649977179
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_53
timestamp 1649977179
transform 1 0 5980 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _070_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform 1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform 1 0 4232 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform 1 0 3404 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 3864 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform 1 0 4232 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform 1 0 4692 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform 1 0 18308 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform 1 0 19044 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform 1 0 18308 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform 1 0 19044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform 1 0 19504 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform 1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform 1 0 19688 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 18584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 19504 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 20424 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13524 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 11224 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 7636 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform -1 0 6716 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 12512 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 10672 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 10304 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform -1 0 8832 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 12144 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform -1 0 7084 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 9016 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 9936 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform -1 0 17388 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform 1 0 12420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform 1 0 9476 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform 1 0 13340 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform 1 0 16100 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform -1 0 11316 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform -1 0 4416 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform 1 0 12880 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform 1 0 7360 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform -1 0 4600 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform 1 0 1564 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform -1 0 6072 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform 1 0 11040 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform 1 0 18032 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1649977179
transform 1 0 11408 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1649977179
transform -1 0 3864 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1649977179
transform -1 0 3496 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1649977179
transform -1 0 4140 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1649977179
transform 1 0 7912 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1649977179
transform 1 0 3864 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1649977179
transform -1 0 2944 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1649977179
transform -1 0 3496 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1649977179
transform 1 0 6992 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1649977179
transform -1 0 3496 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1649977179
transform -1 0 2116 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1649977179
transform -1 0 2208 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1649977179
transform 1 0 10396 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1649977179
transform 1 0 10304 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 1649977179
transform -1 0 3404 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 11776 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 6440 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 1649977179
transform -1 0 21436 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 8556 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 3496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 15364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 7544 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 5796 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 4876 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 9292 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 3496 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 7268 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 17112 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 5060 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 4048 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 18952 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 10948 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 19872 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 4784 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1649977179
transform -1 0 4692 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1649977179
transform -1 0 5796 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform -1 0 2300 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input57 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3036 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8740 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 2852 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 1932 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5152 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6716 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8372 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13708 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15732 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12696 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10948 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10488 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14352 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 16468 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16192 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17848 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13340 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6808 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8556 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6072 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4416 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3772 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 2944 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 1840 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4048 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4600 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6256 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3864 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6072 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2944 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5244 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4324 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5244 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6900 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8372 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6624 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6992 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7728 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10948 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9292 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8004 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11868 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10396 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10212 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8740 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_1__127 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 5888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10212 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8464 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_1__103
timestamp 1649977179
transform -1 0 6992 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8096 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8004 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7452 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_1__104
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2484 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6072 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8004 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_7.mux_l2_in_1__105
timestamp 1649977179
transform -1 0 4048 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7452 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8556 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_0__106
timestamp 1649977179
transform -1 0 12052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12788 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_11.mux_l2_in_0__128
timestamp 1649977179
transform 1 0 15732 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14996 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11776 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_13.mux_l2_in_0__129
timestamp 1649977179
transform -1 0 11040 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8280 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_15.mux_l2_in_0__130
timestamp 1649977179
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10304 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11132 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_0__131
timestamp 1649977179
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18400 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_19.mux_l2_in_0__132
timestamp 1649977179
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13432 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_21.mux_l2_in_0__133
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15916 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16284 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_23.mux_l2_in_0__134
timestamp 1649977179
transform 1 0 19504 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20148 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l1_in_1__135
timestamp 1649977179
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13432 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_27.mux_l2_in_0__136
timestamp 1649977179
transform 1 0 15272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15088 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_29.mux_l2_in_0__137
timestamp 1649977179
transform 1 0 13156 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_29.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17296 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8372 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_1__107
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6900 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5060 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_1__118
timestamp 1649977179
transform -1 0 4232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform -1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3864 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_1__124
timestamp 1649977179
transform 1 0 14536 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2392 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3128 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_7.mux_l2_in_1__125
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2576 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2760 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l1_in_1__126
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 4968 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_11.mux_l2_in_0__108
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5152 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_13.mux_l2_in_0__109
timestamp 1649977179
transform 1 0 5704 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2300 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_15.mux_l2_in_0__110
timestamp 1649977179
transform -1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2760 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5336 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_19.mux_l2_in_0__112
timestamp 1649977179
transform -1 0 3220 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 6808 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_21.mux_l2_in_0__113
timestamp 1649977179
transform -1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3220 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_23.mux_l2_in_0__114
timestamp 1649977179
transform -1 0 6072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_1__115
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7544 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_27.mux_l2_in_0__116
timestamp 1649977179
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_29.mux_l2_in_0__117
timestamp 1649977179
transform -1 0 9568 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_31.mux_l2_in_0__119
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3680 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9752 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_0__120
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4508 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_35.mux_l2_in_0__121
timestamp 1649977179
transform 1 0 8372 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9936 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_37.mux_l2_in_0__122
timestamp 1649977179
transform 1 0 10948 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_39.mux_l2_in_0__123
timestamp 1649977179
transform 1 0 11960 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11684 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output61 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20792 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 3404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 13800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 20148 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 19596 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 19688 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 20148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 20976 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 15364 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 17572 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 17572 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 18124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 -1 3264
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 0 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 3 nsew power input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 4 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 5 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 6 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 7 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 8 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 9 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 bottom_left_grid_pin_48_
port 10 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 bottom_left_grid_pin_49_
port 11 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 bottom_right_grid_pin_1_
port 12 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 ccff_head
port 13 nsew signal input
rlabel metal3 s 22200 17144 23000 17264 6 ccff_tail
port 14 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 15 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 16 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 17 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 18 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 19 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 20 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 21 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 22 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 23 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 24 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 25 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 26 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 27 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 28 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 29 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 30 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 31 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 32 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 33 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 34 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 35 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 36 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 37 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 38 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 39 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 40 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 41 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 42 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 43 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 44 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 45 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 46 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 47 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 48 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 49 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 50 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 51 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 52 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 53 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 54 nsew signal tristate
rlabel metal2 s 3698 0 3754 800 6 chany_bottom_in[0]
port 55 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[10]
port 56 nsew signal input
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[11]
port 57 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 chany_bottom_in[12]
port 58 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[13]
port 59 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 chany_bottom_in[14]
port 60 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 chany_bottom_in[15]
port 61 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 chany_bottom_in[16]
port 62 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 chany_bottom_in[17]
port 63 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_in[18]
port 64 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 chany_bottom_in[19]
port 65 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 chany_bottom_in[1]
port 66 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 chany_bottom_in[2]
port 67 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 chany_bottom_in[3]
port 68 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 chany_bottom_in[4]
port 69 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 chany_bottom_in[5]
port 70 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 chany_bottom_in[6]
port 71 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[7]
port 72 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 chany_bottom_in[8]
port 73 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[9]
port 74 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 chany_bottom_out[0]
port 75 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_out[10]
port 76 nsew signal tristate
rlabel metal2 s 17406 0 17462 800 6 chany_bottom_out[11]
port 77 nsew signal tristate
rlabel metal2 s 17866 0 17922 800 6 chany_bottom_out[12]
port 78 nsew signal tristate
rlabel metal2 s 18326 0 18382 800 6 chany_bottom_out[13]
port 79 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 chany_bottom_out[14]
port 80 nsew signal tristate
rlabel metal2 s 19154 0 19210 800 6 chany_bottom_out[15]
port 81 nsew signal tristate
rlabel metal2 s 19614 0 19670 800 6 chany_bottom_out[16]
port 82 nsew signal tristate
rlabel metal2 s 20074 0 20130 800 6 chany_bottom_out[17]
port 83 nsew signal tristate
rlabel metal2 s 20534 0 20590 800 6 chany_bottom_out[18]
port 84 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[19]
port 85 nsew signal tristate
rlabel metal2 s 12990 0 13046 800 6 chany_bottom_out[1]
port 86 nsew signal tristate
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_out[2]
port 87 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_out[3]
port 88 nsew signal tristate
rlabel metal2 s 14278 0 14334 800 6 chany_bottom_out[4]
port 89 nsew signal tristate
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_out[5]
port 90 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[6]
port 91 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[7]
port 92 nsew signal tristate
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_out[8]
port 93 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 94 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 95 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 96 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 97 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 98 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 99 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 100 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 101 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 102 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 103 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 104 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
