magic
tech sky130A
magscale 1 2
timestamp 1650626062
<< viali >>
rect 2789 14569 2823 14603
rect 3157 14569 3191 14603
rect 4261 14569 4295 14603
rect 4629 14569 4663 14603
rect 5733 14569 5767 14603
rect 6561 14569 6595 14603
rect 7113 14569 7147 14603
rect 7389 14569 7423 14603
rect 12173 14569 12207 14603
rect 12449 14569 12483 14603
rect 12633 14569 12667 14603
rect 12817 14569 12851 14603
rect 13001 14569 13035 14603
rect 13185 14569 13219 14603
rect 14105 14569 14139 14603
rect 14473 14569 14507 14603
rect 5089 14501 5123 14535
rect 5273 14501 5307 14535
rect 6009 14501 6043 14535
rect 6101 14501 6135 14535
rect 6745 14501 6779 14535
rect 6929 14501 6963 14535
rect 15117 14501 15151 14535
rect 1961 14433 1995 14467
rect 13737 14433 13771 14467
rect 17325 14433 17359 14467
rect 17601 14433 17635 14467
rect 18521 14433 18555 14467
rect 2237 14365 2271 14399
rect 2605 14365 2639 14399
rect 2973 14365 3007 14399
rect 3341 14365 3375 14399
rect 3617 14365 3651 14399
rect 3801 14365 3835 14399
rect 4077 14365 4111 14399
rect 4353 14365 4387 14399
rect 4789 14365 4823 14399
rect 4905 14365 4939 14399
rect 5549 14365 5583 14399
rect 6377 14365 6411 14399
rect 9965 14365 9999 14399
rect 14289 14365 14323 14399
rect 14565 14365 14599 14399
rect 15025 14365 15059 14399
rect 15301 14365 15335 14399
rect 15669 14365 15703 14399
rect 15853 14365 15887 14399
rect 16037 14365 16071 14399
rect 16405 14365 16439 14399
rect 18245 14365 18279 14399
rect 13461 14297 13495 14331
rect 13829 14297 13863 14331
rect 15485 14297 15519 14331
rect 2421 14229 2455 14263
rect 3433 14229 3467 14263
rect 3985 14229 4019 14263
rect 4537 14229 4571 14263
rect 5365 14229 5399 14263
rect 10149 14229 10183 14263
rect 11989 14229 12023 14263
rect 13369 14229 13403 14263
rect 14749 14229 14783 14263
rect 14841 14229 14875 14263
rect 16313 14229 16347 14263
rect 2789 14025 2823 14059
rect 3433 14025 3467 14059
rect 3617 14025 3651 14059
rect 4169 14025 4203 14059
rect 4445 14025 4479 14059
rect 4813 14025 4847 14059
rect 5365 14025 5399 14059
rect 6377 14025 6411 14059
rect 6653 14025 6687 14059
rect 7205 14025 7239 14059
rect 8125 14025 8159 14059
rect 9781 14025 9815 14059
rect 13737 14025 13771 14059
rect 14013 14025 14047 14059
rect 14841 14025 14875 14059
rect 15761 14025 15795 14059
rect 2605 13957 2639 13991
rect 5181 13957 5215 13991
rect 5917 13957 5951 13991
rect 6929 13957 6963 13991
rect 7113 13957 7147 13991
rect 7481 13957 7515 13991
rect 12081 13957 12115 13991
rect 12357 13957 12391 13991
rect 12541 13957 12575 13991
rect 12725 13957 12759 13991
rect 12909 13957 12943 13991
rect 16221 13957 16255 13991
rect 2237 13889 2271 13923
rect 2421 13889 2455 13923
rect 2973 13889 3007 13923
rect 3249 13889 3283 13923
rect 3801 13889 3835 13923
rect 3893 13889 3927 13923
rect 4353 13889 4387 13923
rect 4629 13889 4663 13923
rect 6009 13889 6043 13923
rect 6561 13889 6595 13923
rect 7941 13889 7975 13923
rect 9597 13873 9631 13907
rect 13093 13889 13127 13923
rect 13553 13889 13587 13923
rect 13829 13889 13863 13923
rect 14289 13889 14323 13923
rect 14565 13889 14599 13923
rect 15025 13889 15059 13923
rect 15301 13889 15335 13923
rect 15393 13889 15427 13923
rect 15853 13889 15887 13923
rect 16497 13889 16531 13923
rect 1961 13821 1995 13855
rect 3065 13821 3099 13855
rect 4905 13821 4939 13855
rect 7573 13821 7607 13855
rect 11529 13821 11563 13855
rect 13277 13821 13311 13855
rect 16773 13821 16807 13855
rect 17049 13821 17083 13855
rect 17693 13821 17727 13855
rect 17969 13821 18003 13855
rect 5641 13753 5675 13787
rect 13369 13753 13403 13787
rect 14105 13753 14139 13787
rect 14381 13753 14415 13787
rect 15577 13753 15611 13787
rect 4077 13685 4111 13719
rect 5549 13685 5583 13719
rect 7849 13685 7883 13719
rect 11713 13685 11747 13719
rect 11897 13685 11931 13719
rect 14657 13685 14691 13719
rect 15117 13685 15151 13719
rect 4629 13481 4663 13515
rect 6285 13481 6319 13515
rect 6653 13481 6687 13515
rect 8033 13481 8067 13515
rect 8309 13481 8343 13515
rect 8585 13481 8619 13515
rect 9045 13481 9079 13515
rect 11437 13481 11471 13515
rect 12817 13481 12851 13515
rect 16129 13481 16163 13515
rect 3157 13413 3191 13447
rect 3801 13413 3835 13447
rect 11805 13413 11839 13447
rect 12265 13413 12299 13447
rect 15025 13413 15059 13447
rect 2237 13345 2271 13379
rect 5733 13345 5767 13379
rect 7205 13345 7239 13379
rect 8769 13345 8803 13379
rect 11529 13345 11563 13379
rect 13001 13345 13035 13379
rect 15301 13345 15335 13379
rect 17693 13345 17727 13379
rect 1961 13277 1995 13311
rect 2605 13277 2639 13311
rect 2973 13277 3007 13311
rect 3341 13277 3375 13311
rect 3433 13277 3467 13311
rect 3985 13277 4019 13311
rect 4077 13277 4111 13311
rect 4353 13277 4387 13311
rect 4813 13277 4847 13311
rect 4905 13277 4939 13311
rect 5181 13277 5215 13311
rect 5365 13277 5399 13311
rect 11069 13277 11103 13311
rect 11897 13277 11931 13311
rect 12725 13277 12759 13311
rect 13177 13273 13211 13307
rect 13469 13273 13503 13307
rect 13737 13277 13771 13311
rect 14473 13277 14507 13311
rect 14565 13277 14599 13311
rect 14841 13277 14875 13311
rect 15393 13277 15427 13311
rect 17509 13277 17543 13311
rect 17969 13277 18003 13311
rect 6469 13209 6503 13243
rect 7021 13209 7055 13243
rect 10885 13209 10919 13243
rect 11161 13209 11195 13243
rect 12541 13209 12575 13243
rect 14105 13209 14139 13243
rect 17417 13209 17451 13243
rect 2421 13141 2455 13175
rect 2789 13141 2823 13175
rect 3617 13141 3651 13175
rect 4261 13141 4295 13175
rect 4537 13141 4571 13175
rect 5089 13141 5123 13175
rect 5917 13141 5951 13175
rect 6193 13141 6227 13175
rect 6929 13141 6963 13175
rect 7389 13141 7423 13175
rect 7573 13141 7607 13175
rect 7757 13141 7791 13175
rect 8125 13141 8159 13175
rect 10609 13141 10643 13175
rect 12081 13141 12115 13175
rect 13369 13141 13403 13175
rect 13645 13141 13679 13175
rect 13921 13141 13955 13175
rect 14289 13141 14323 13175
rect 14749 13141 14783 13175
rect 15577 13141 15611 13175
rect 4353 12937 4387 12971
rect 4813 12937 4847 12971
rect 5825 12937 5859 12971
rect 9137 12937 9171 12971
rect 9505 12937 9539 12971
rect 10057 12937 10091 12971
rect 10425 12937 10459 12971
rect 10609 12937 10643 12971
rect 11529 12937 11563 12971
rect 11989 12937 12023 12971
rect 13185 12937 13219 12971
rect 13829 12937 13863 12971
rect 15577 12937 15611 12971
rect 4077 12869 4111 12903
rect 7665 12869 7699 12903
rect 8125 12869 8159 12903
rect 8309 12869 8343 12903
rect 8769 12869 8803 12903
rect 9045 12869 9079 12903
rect 10793 12869 10827 12903
rect 16681 12869 16715 12903
rect 2881 12801 2915 12835
rect 3525 12801 3559 12835
rect 3801 12801 3835 12835
rect 4997 12801 5031 12835
rect 5365 12801 5399 12835
rect 5641 12801 5675 12835
rect 5917 12801 5951 12835
rect 7849 12801 7883 12835
rect 8585 12801 8619 12835
rect 9321 12801 9355 12835
rect 12265 12801 12299 12835
rect 12609 12801 12643 12835
rect 12725 12801 12759 12835
rect 13001 12801 13035 12835
rect 13461 12801 13495 12835
rect 13553 12801 13587 12835
rect 14013 12801 14047 12835
rect 14265 12801 14299 12835
rect 14381 12801 14415 12835
rect 14749 12801 14783 12835
rect 15301 12801 15335 12835
rect 15669 12801 15703 12835
rect 16037 12801 16071 12835
rect 16405 12801 16439 12835
rect 1961 12733 1995 12767
rect 2237 12733 2271 12767
rect 3157 12733 3191 12767
rect 5273 12733 5307 12767
rect 6653 12733 6687 12767
rect 7205 12733 7239 12767
rect 7573 12733 7607 12767
rect 11069 12733 11103 12767
rect 12173 12733 12207 12767
rect 3617 12665 3651 12699
rect 4721 12665 4755 12699
rect 5549 12665 5583 12699
rect 6561 12665 6595 12699
rect 6929 12665 6963 12699
rect 10149 12665 10183 12699
rect 10885 12665 10919 12699
rect 11345 12665 11379 12699
rect 12449 12665 12483 12699
rect 12909 12665 12943 12699
rect 14933 12665 14967 12699
rect 15853 12665 15887 12699
rect 16221 12665 16255 12699
rect 3341 12597 3375 12631
rect 3985 12597 4019 12631
rect 6101 12597 6135 12631
rect 7021 12597 7055 12631
rect 8493 12597 8527 12631
rect 11805 12597 11839 12631
rect 13277 12597 13311 12631
rect 13737 12597 13771 12631
rect 14105 12597 14139 12631
rect 14565 12597 14599 12631
rect 15209 12597 15243 12631
rect 17969 12597 18003 12631
rect 9137 12393 9171 12427
rect 9781 12393 9815 12427
rect 10149 12393 10183 12427
rect 11161 12393 11195 12427
rect 17141 12393 17175 12427
rect 8677 12325 8711 12359
rect 11529 12325 11563 12359
rect 11897 12325 11931 12359
rect 13461 12325 13495 12359
rect 16129 12325 16163 12359
rect 16865 12325 16899 12359
rect 2421 12257 2455 12291
rect 3433 12257 3467 12291
rect 4629 12257 4663 12291
rect 10793 12257 10827 12291
rect 14841 12257 14875 12291
rect 17693 12257 17727 12291
rect 17969 12257 18003 12291
rect 1961 12189 1995 12223
rect 2237 12189 2271 12223
rect 3249 12189 3283 12223
rect 4445 12189 4479 12223
rect 5365 12189 5399 12223
rect 5457 12189 5491 12223
rect 6201 12189 6235 12223
rect 6469 12189 6503 12223
rect 7205 12189 7239 12223
rect 7481 12189 7515 12223
rect 9321 12189 9355 12223
rect 11345 12189 11379 12223
rect 12541 12189 12575 12223
rect 12817 12189 12851 12223
rect 12909 12189 12943 12223
rect 13185 12189 13219 12223
rect 13645 12189 13679 12223
rect 14105 12189 14139 12223
rect 14473 12189 14507 12223
rect 15577 12189 15611 12223
rect 15945 12189 15979 12223
rect 16681 12189 16715 12223
rect 17417 12189 17451 12223
rect 3893 12121 3927 12155
rect 8125 12121 8159 12155
rect 10057 12121 10091 12155
rect 10885 12121 10919 12155
rect 16497 12121 16531 12155
rect 17233 12121 17267 12155
rect 2605 12053 2639 12087
rect 2697 12053 2731 12087
rect 3065 12053 3099 12087
rect 3525 12053 3559 12087
rect 3985 12053 4019 12087
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 6101 12053 6135 12087
rect 6377 12053 6411 12087
rect 7113 12053 7147 12087
rect 7389 12053 7423 12087
rect 8217 12053 8251 12087
rect 8493 12053 8527 12087
rect 9045 12053 9079 12087
rect 9505 12053 9539 12087
rect 10333 12053 10367 12087
rect 10517 12053 10551 12087
rect 11713 12053 11747 12087
rect 11989 12053 12023 12087
rect 12173 12053 12207 12087
rect 12357 12053 12391 12087
rect 12633 12053 12667 12087
rect 13093 12053 13127 12087
rect 13369 12053 13403 12087
rect 13829 12053 13863 12087
rect 14289 12053 14323 12087
rect 15761 12053 15795 12087
rect 16405 12053 16439 12087
rect 17601 12053 17635 12087
rect 3065 11849 3099 11883
rect 3893 11849 3927 11883
rect 4261 11849 4295 11883
rect 4721 11849 4755 11883
rect 11345 11849 11379 11883
rect 17417 11849 17451 11883
rect 4353 11781 4387 11815
rect 6101 11781 6135 11815
rect 7757 11781 7791 11815
rect 12449 11781 12483 11815
rect 14749 11781 14783 11815
rect 2237 11713 2271 11747
rect 2697 11713 2731 11747
rect 3525 11713 3559 11747
rect 5089 11713 5123 11747
rect 6009 11713 6043 11747
rect 6837 11713 6871 11747
rect 7665 11713 7699 11747
rect 8125 11713 8159 11747
rect 8769 11713 8803 11747
rect 10618 11713 10652 11747
rect 10885 11713 10919 11747
rect 11805 11713 11839 11747
rect 11989 11713 12023 11747
rect 12541 11713 12575 11747
rect 13001 11713 13035 11747
rect 13277 11713 13311 11747
rect 13737 11713 13771 11747
rect 14117 11713 14151 11747
rect 14203 11713 14237 11747
rect 14933 11713 14967 11747
rect 16313 11713 16347 11747
rect 16681 11713 16715 11747
rect 17601 11713 17635 11747
rect 1961 11645 1995 11679
rect 2421 11645 2455 11679
rect 2605 11645 2639 11679
rect 3249 11645 3283 11679
rect 3433 11645 3467 11679
rect 4077 11645 4111 11679
rect 5273 11645 5307 11679
rect 6929 11645 6963 11679
rect 7021 11645 7055 11679
rect 7849 11645 7883 11679
rect 8401 11645 8435 11679
rect 11529 11645 11563 11679
rect 17739 11645 17773 11679
rect 17969 11645 18003 11679
rect 11161 11577 11195 11611
rect 12817 11577 12851 11611
rect 13093 11577 13127 11611
rect 4905 11509 4939 11543
rect 5365 11509 5399 11543
rect 6469 11509 6503 11543
rect 7297 11509 7331 11543
rect 8309 11509 8343 11543
rect 9413 11509 9447 11543
rect 9505 11509 9539 11543
rect 12173 11509 12207 11543
rect 12725 11509 12759 11543
rect 13553 11509 13587 11543
rect 13921 11509 13955 11543
rect 14381 11509 14415 11543
rect 14657 11509 14691 11543
rect 15577 11509 15611 11543
rect 15669 11509 15703 11543
rect 16405 11509 16439 11543
rect 17325 11509 17359 11543
rect 2145 11305 2179 11339
rect 3801 11305 3835 11339
rect 10425 11305 10459 11339
rect 12449 11305 12483 11339
rect 15485 11305 15519 11339
rect 2237 11237 2271 11271
rect 11621 11237 11655 11271
rect 13737 11237 13771 11271
rect 1593 11169 1627 11203
rect 1685 11169 1719 11203
rect 4261 11169 4295 11203
rect 4445 11169 4479 11203
rect 8125 11169 8159 11203
rect 10333 11169 10367 11203
rect 11253 11169 11287 11203
rect 11345 11169 11379 11203
rect 12173 11169 12207 11203
rect 12817 11169 12851 11203
rect 1777 11101 1811 11135
rect 3617 11101 3651 11135
rect 4629 11101 4663 11135
rect 6101 11101 6135 11135
rect 7941 11101 7975 11135
rect 8769 11101 8803 11135
rect 10609 11077 10643 11111
rect 11161 11101 11195 11135
rect 12633 11101 12667 11135
rect 12909 11101 12943 11135
rect 13921 11101 13955 11135
rect 14105 11101 14139 11135
rect 15577 11101 15611 11135
rect 17049 11101 17083 11135
rect 3372 11033 3406 11067
rect 4896 11033 4930 11067
rect 6346 11033 6380 11067
rect 8033 11033 8067 11067
rect 10088 11033 10122 11067
rect 11989 11033 12023 11067
rect 12081 11033 12115 11067
rect 13553 11033 13587 11067
rect 14350 11033 14384 11067
rect 15822 11033 15856 11067
rect 17316 11033 17350 11067
rect 4169 10965 4203 10999
rect 6009 10965 6043 10999
rect 7481 10965 7515 10999
rect 7573 10965 7607 10999
rect 8401 10965 8435 10999
rect 8585 10965 8619 10999
rect 8953 10965 8987 10999
rect 10793 10965 10827 10999
rect 16957 10965 16991 10999
rect 18429 10965 18463 10999
rect 1409 10761 1443 10795
rect 3525 10761 3559 10795
rect 3617 10761 3651 10795
rect 3985 10761 4019 10795
rect 6193 10761 6227 10795
rect 7297 10761 7331 10795
rect 8217 10761 8251 10795
rect 8585 10761 8619 10795
rect 9045 10761 9079 10795
rect 9413 10761 9447 10795
rect 9781 10761 9815 10795
rect 10241 10761 10275 10795
rect 10609 10761 10643 10795
rect 13461 10761 13495 10795
rect 17417 10761 17451 10795
rect 17785 10761 17819 10795
rect 2522 10693 2556 10727
rect 2973 10693 3007 10727
rect 5190 10693 5224 10727
rect 7205 10693 7239 10727
rect 8125 10693 8159 10727
rect 10701 10693 10735 10727
rect 11253 10693 11287 10727
rect 14749 10693 14783 10727
rect 5549 10625 5583 10659
rect 6377 10625 6411 10659
rect 8953 10625 8987 10659
rect 11529 10625 11563 10659
rect 12541 10625 12575 10659
rect 12909 10625 12943 10659
rect 15965 10625 15999 10659
rect 17325 10625 17359 10659
rect 18153 10625 18187 10659
rect 18245 10625 18279 10659
rect 2789 10557 2823 10591
rect 3433 10557 3467 10591
rect 5457 10557 5491 10591
rect 7389 10557 7423 10591
rect 8401 10557 8435 10591
rect 9229 10557 9263 10591
rect 9873 10557 9907 10591
rect 9965 10557 9999 10591
rect 10793 10557 10827 10591
rect 16221 10557 16255 10591
rect 16313 10557 16347 10591
rect 16865 10557 16899 10591
rect 17601 10557 17635 10591
rect 18337 10557 18371 10591
rect 12173 10489 12207 10523
rect 3065 10421 3099 10455
rect 4077 10421 4111 10455
rect 6561 10421 6595 10455
rect 6837 10421 6871 10455
rect 7757 10421 7791 10455
rect 11161 10421 11195 10455
rect 12357 10421 12391 10455
rect 12725 10421 12759 10455
rect 14841 10421 14875 10455
rect 16957 10421 16991 10455
rect 6101 10217 6135 10251
rect 7021 10217 7055 10251
rect 8769 10217 8803 10251
rect 8953 10217 8987 10251
rect 9505 10217 9539 10251
rect 11713 10217 11747 10251
rect 16589 10217 16623 10251
rect 6193 10149 6227 10183
rect 7849 10149 7883 10183
rect 2237 10081 2271 10115
rect 4997 10081 5031 10115
rect 5457 10081 5491 10115
rect 6653 10081 6687 10115
rect 6745 10081 6779 10115
rect 7573 10081 7607 10115
rect 8217 10081 8251 10115
rect 10149 10081 10183 10115
rect 12357 10081 12391 10115
rect 14289 10081 14323 10115
rect 15485 10081 15519 10115
rect 15853 10081 15887 10115
rect 16037 10081 16071 10115
rect 17141 10081 17175 10115
rect 17969 10081 18003 10115
rect 1961 10013 1995 10047
rect 2329 10013 2363 10047
rect 2605 10013 2639 10047
rect 3617 10013 3651 10047
rect 4077 10013 4111 10047
rect 4353 10013 4387 10047
rect 4813 10013 4847 10047
rect 6561 10013 6595 10047
rect 8401 10013 8435 10047
rect 9129 10013 9163 10047
rect 9229 10013 9263 10047
rect 9873 10013 9907 10047
rect 10333 10013 10367 10047
rect 11805 10013 11839 10047
rect 12265 10013 12299 10047
rect 14381 10013 14415 10047
rect 14473 10013 14507 10047
rect 16957 10013 16991 10047
rect 18245 10013 18279 10047
rect 5641 9945 5675 9979
rect 7481 9945 7515 9979
rect 8309 9945 8343 9979
rect 10578 9945 10612 9979
rect 12624 9945 12658 9979
rect 13921 9945 13955 9979
rect 15301 9945 15335 9979
rect 15393 9945 15427 9979
rect 16129 9945 16163 9979
rect 17877 9945 17911 9979
rect 3433 9877 3467 9911
rect 3893 9877 3927 9911
rect 4169 9877 4203 9911
rect 4445 9877 4479 9911
rect 4905 9877 4939 9911
rect 5733 9877 5767 9911
rect 7389 9877 7423 9911
rect 9413 9877 9447 9911
rect 9965 9877 9999 9911
rect 12081 9877 12115 9911
rect 13737 9877 13771 9911
rect 14841 9877 14875 9911
rect 14933 9877 14967 9911
rect 16497 9877 16531 9911
rect 17049 9877 17083 9911
rect 17417 9877 17451 9911
rect 17785 9877 17819 9911
rect 18429 9877 18463 9911
rect 4905 9673 4939 9707
rect 6377 9673 6411 9707
rect 8033 9673 8067 9707
rect 10333 9673 10367 9707
rect 14565 9673 14599 9707
rect 17417 9673 17451 9707
rect 17693 9673 17727 9707
rect 5917 9605 5951 9639
rect 7490 9605 7524 9639
rect 13032 9605 13066 9639
rect 15384 9605 15418 9639
rect 16957 9605 16991 9639
rect 17049 9605 17083 9639
rect 18061 9605 18095 9639
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 2421 9537 2455 9571
rect 3902 9537 3936 9571
rect 4169 9537 4203 9571
rect 4813 9537 4847 9571
rect 5825 9537 5859 9571
rect 7849 9537 7883 9571
rect 8381 9537 8415 9571
rect 9597 9537 9631 9571
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 11345 9537 11379 9571
rect 11805 9537 11839 9571
rect 13277 9537 13311 9571
rect 13737 9537 13771 9571
rect 14657 9537 14691 9571
rect 15117 9537 15151 9571
rect 17509 9537 17543 9571
rect 18153 9537 18187 9571
rect 4997 9469 5031 9503
rect 6101 9469 6135 9503
rect 7757 9469 7791 9503
rect 8125 9469 8159 9503
rect 10977 9469 11011 9503
rect 13829 9469 13863 9503
rect 13921 9469 13955 9503
rect 14749 9469 14783 9503
rect 16865 9469 16899 9503
rect 18245 9469 18279 9503
rect 4353 9401 4387 9435
rect 5457 9401 5491 9435
rect 9505 9401 9539 9435
rect 11161 9401 11195 9435
rect 11897 9401 11931 9435
rect 14197 9401 14231 9435
rect 16497 9401 16531 9435
rect 2513 9333 2547 9367
rect 2789 9333 2823 9367
rect 4445 9333 4479 9367
rect 5365 9333 5399 9367
rect 10241 9333 10275 9367
rect 11621 9333 11655 9367
rect 13369 9333 13403 9367
rect 3985 9129 4019 9163
rect 6469 9129 6503 9163
rect 7205 9129 7239 9163
rect 10793 9129 10827 9163
rect 13185 9129 13219 9163
rect 13921 9129 13955 9163
rect 14105 9129 14139 9163
rect 10701 9061 10735 9095
rect 1685 8993 1719 9027
rect 4537 8993 4571 9027
rect 5089 8993 5123 9027
rect 11345 8993 11379 9027
rect 12173 8993 12207 9027
rect 12633 8993 12667 9027
rect 15761 8993 15795 9027
rect 1501 8925 1535 8959
rect 2890 8925 2924 8959
rect 3157 8925 3191 8959
rect 3801 8925 3835 8959
rect 4997 8901 5031 8935
rect 5356 8925 5390 8959
rect 6561 8925 6595 8959
rect 7297 8925 7331 8959
rect 8953 8925 8987 8959
rect 9321 8925 9355 8959
rect 9577 8925 9611 8959
rect 11253 8925 11287 8959
rect 11989 8925 12023 8959
rect 12817 8925 12851 8959
rect 13277 8925 13311 8959
rect 15485 8925 15519 8959
rect 16497 8925 16531 8959
rect 16764 8925 16798 8959
rect 18245 8925 18279 8959
rect 18521 8925 18555 8959
rect 3341 8857 3375 8891
rect 4445 8857 4479 8891
rect 7564 8857 7598 8891
rect 15218 8857 15252 8891
rect 16037 8857 16071 8891
rect 1777 8789 1811 8823
rect 3433 8789 3467 8823
rect 4353 8789 4387 8823
rect 4813 8789 4847 8823
rect 8677 8789 8711 8823
rect 9137 8789 9171 8823
rect 11161 8789 11195 8823
rect 11621 8789 11655 8823
rect 12081 8789 12115 8823
rect 12725 8789 12759 8823
rect 15945 8789 15979 8823
rect 16405 8789 16439 8823
rect 17877 8789 17911 8823
rect 18061 8789 18095 8823
rect 18337 8789 18371 8823
rect 6193 8585 6227 8619
rect 12449 8585 12483 8619
rect 12633 8585 12667 8619
rect 13461 8585 13495 8619
rect 13829 8585 13863 8619
rect 14289 8585 14323 8619
rect 16313 8585 16347 8619
rect 17141 8585 17175 8619
rect 17509 8585 17543 8619
rect 18337 8585 18371 8619
rect 4241 8517 4275 8551
rect 9157 8517 9191 8551
rect 13001 8517 13035 8551
rect 15608 8517 15642 8551
rect 17877 8517 17911 8551
rect 17969 8517 18003 8551
rect 1501 8449 1535 8483
rect 1768 8449 1802 8483
rect 3525 8449 3559 8483
rect 3985 8449 4019 8483
rect 5825 8449 5859 8483
rect 7582 8449 7616 8483
rect 7849 8449 7883 8483
rect 9413 8449 9447 8483
rect 9505 8449 9539 8483
rect 11078 8449 11112 8483
rect 11805 8449 11839 8483
rect 15853 8449 15887 8483
rect 15945 8449 15979 8483
rect 16497 8449 16531 8483
rect 17049 8449 17083 8483
rect 18521 8449 18555 8483
rect 3801 8381 3835 8415
rect 5641 8381 5675 8415
rect 5733 8381 5767 8415
rect 11345 8381 11379 8415
rect 11529 8381 11563 8415
rect 13093 8381 13127 8415
rect 13277 8381 13311 8415
rect 13921 8381 13955 8415
rect 14105 8381 14139 8415
rect 17233 8381 17267 8415
rect 18061 8381 18095 8415
rect 2881 8313 2915 8347
rect 5365 8313 5399 8347
rect 6469 8313 6503 8347
rect 9689 8313 9723 8347
rect 16129 8313 16163 8347
rect 16681 8313 16715 8347
rect 8033 8245 8067 8279
rect 9965 8245 9999 8279
rect 14473 8245 14507 8279
rect 4353 8041 4387 8075
rect 5733 8041 5767 8075
rect 15853 8041 15887 8075
rect 3525 7973 3559 8007
rect 4445 7973 4479 8007
rect 10885 7973 10919 8007
rect 2237 7905 2271 7939
rect 4997 7905 5031 7939
rect 7757 7905 7791 7939
rect 8953 7905 8987 7939
rect 12357 7905 12391 7939
rect 16037 7905 16071 7939
rect 16221 7905 16255 7939
rect 17325 7905 17359 7939
rect 18153 7905 18187 7939
rect 1961 7837 1995 7871
rect 3157 7837 3191 7871
rect 4169 7837 4203 7871
rect 4813 7837 4847 7871
rect 7021 7837 7055 7871
rect 7481 7837 7515 7871
rect 7941 7837 7975 7871
rect 8263 7837 8297 7871
rect 9229 7837 9263 7871
rect 10333 7837 10367 7871
rect 12624 7837 12658 7871
rect 14105 7837 14139 7871
rect 14473 7837 14507 7871
rect 14740 7837 14774 7871
rect 18061 7837 18095 7871
rect 3341 7769 3375 7803
rect 3893 7769 3927 7803
rect 4077 7769 4111 7803
rect 12173 7769 12207 7803
rect 16313 7769 16347 7803
rect 17233 7769 17267 7803
rect 2927 7701 2961 7735
rect 4905 7701 4939 7735
rect 7113 7701 7147 7735
rect 7573 7701 7607 7735
rect 9873 7701 9907 7735
rect 10149 7701 10183 7735
rect 13737 7701 13771 7735
rect 13829 7701 13863 7735
rect 14289 7701 14323 7735
rect 16681 7701 16715 7735
rect 16773 7701 16807 7735
rect 17141 7701 17175 7735
rect 17601 7701 17635 7735
rect 17969 7701 18003 7735
rect 18521 7701 18555 7735
rect 2513 7497 2547 7531
rect 4905 7497 4939 7531
rect 6377 7497 6411 7531
rect 8033 7497 8067 7531
rect 8217 7497 8251 7531
rect 8861 7497 8895 7531
rect 9597 7497 9631 7531
rect 12909 7497 12943 7531
rect 14841 7497 14875 7531
rect 15669 7497 15703 7531
rect 17049 7497 17083 7531
rect 17509 7497 17543 7531
rect 17969 7497 18003 7531
rect 5641 7429 5675 7463
rect 11069 7429 11103 7463
rect 16037 7429 16071 7463
rect 16129 7429 16163 7463
rect 17141 7429 17175 7463
rect 1685 7361 1719 7395
rect 2145 7361 2179 7395
rect 2605 7361 2639 7395
rect 4353 7361 4387 7395
rect 4813 7361 4847 7395
rect 7501 7361 7535 7395
rect 7757 7361 7791 7395
rect 7849 7361 7883 7395
rect 8401 7361 8435 7395
rect 8953 7361 8987 7395
rect 11161 7361 11195 7395
rect 11796 7361 11830 7395
rect 13001 7361 13035 7395
rect 15209 7361 15243 7395
rect 17877 7361 17911 7395
rect 18521 7361 18555 7395
rect 1869 7293 1903 7327
rect 2053 7293 2087 7327
rect 5089 7293 5123 7327
rect 5733 7293 5767 7327
rect 5917 7293 5951 7327
rect 9137 7293 9171 7327
rect 11529 7293 11563 7327
rect 15301 7293 15335 7327
rect 15393 7293 15427 7327
rect 16221 7293 16255 7327
rect 17325 7293 17359 7327
rect 18061 7293 18095 7327
rect 6101 7225 6135 7259
rect 16681 7225 16715 7259
rect 1501 7157 1535 7191
rect 4445 7157 4479 7191
rect 5273 7157 5307 7191
rect 8493 7157 8527 7191
rect 11345 7157 11379 7191
rect 14289 7157 14323 7191
rect 18337 7157 18371 7191
rect 7205 6953 7239 6987
rect 10425 6953 10459 6987
rect 18245 6953 18279 6987
rect 2881 6885 2915 6919
rect 4721 6885 4755 6919
rect 4813 6885 4847 6919
rect 6377 6885 6411 6919
rect 3801 6817 3835 6851
rect 4169 6817 4203 6851
rect 4261 6817 4295 6851
rect 6193 6817 6227 6851
rect 6929 6817 6963 6851
rect 7665 6817 7699 6851
rect 7849 6817 7883 6851
rect 8125 6817 8159 6851
rect 8309 6817 8343 6851
rect 10977 6817 11011 6851
rect 13737 6817 13771 6851
rect 17601 6817 17635 6851
rect 17785 6817 17819 6851
rect 1501 6749 1535 6783
rect 3617 6749 3651 6783
rect 4353 6749 4387 6783
rect 6745 6749 6779 6783
rect 7573 6749 7607 6783
rect 10333 6749 10367 6783
rect 11529 6749 11563 6783
rect 13001 6749 13035 6783
rect 13553 6749 13587 6783
rect 15485 6749 15519 6783
rect 15669 6749 15703 6783
rect 17141 6749 17175 6783
rect 1746 6681 1780 6715
rect 5948 6681 5982 6715
rect 10066 6681 10100 6715
rect 10793 6681 10827 6715
rect 12756 6681 12790 6715
rect 15218 6681 15252 6715
rect 15936 6681 15970 6715
rect 17877 6681 17911 6715
rect 18337 6681 18371 6715
rect 2973 6613 3007 6647
rect 6837 6613 6871 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 8953 6613 8987 6647
rect 10885 6613 10919 6647
rect 11345 6613 11379 6647
rect 11621 6613 11655 6647
rect 13185 6613 13219 6647
rect 13645 6613 13679 6647
rect 14105 6613 14139 6647
rect 17049 6613 17083 6647
rect 17325 6613 17359 6647
rect 1593 6409 1627 6443
rect 4537 6409 4571 6443
rect 4813 6409 4847 6443
rect 6377 6409 6411 6443
rect 6745 6409 6779 6443
rect 7205 6409 7239 6443
rect 7665 6409 7699 6443
rect 9505 6409 9539 6443
rect 9873 6409 9907 6443
rect 9965 6409 9999 6443
rect 10333 6409 10367 6443
rect 10701 6409 10735 6443
rect 11345 6409 11379 6443
rect 11805 6409 11839 6443
rect 13185 6409 13219 6443
rect 15117 6409 15151 6443
rect 18337 6409 18371 6443
rect 2513 6341 2547 6375
rect 6837 6341 6871 6375
rect 8278 6341 8312 6375
rect 14381 6341 14415 6375
rect 14473 6341 14507 6375
rect 15209 6341 15243 6375
rect 16948 6341 16982 6375
rect 1961 6273 1995 6307
rect 2421 6273 2455 6307
rect 3148 6273 3182 6307
rect 4353 6273 4387 6307
rect 5926 6273 5960 6307
rect 7573 6273 7607 6307
rect 11897 6273 11931 6307
rect 12725 6273 12759 6307
rect 12817 6273 12851 6307
rect 13553 6273 13587 6307
rect 16037 6273 16071 6307
rect 18153 6273 18187 6307
rect 2605 6205 2639 6239
rect 2881 6205 2915 6239
rect 6193 6205 6227 6239
rect 6929 6205 6963 6239
rect 7849 6205 7883 6239
rect 8033 6205 8067 6239
rect 10057 6205 10091 6239
rect 10793 6205 10827 6239
rect 10977 6205 11011 6239
rect 11713 6205 11747 6239
rect 12909 6205 12943 6239
rect 13645 6205 13679 6239
rect 13829 6205 13863 6239
rect 14565 6205 14599 6239
rect 14933 6205 14967 6239
rect 16129 6205 16163 6239
rect 16221 6205 16255 6239
rect 16681 6205 16715 6239
rect 9413 6137 9447 6171
rect 12357 6137 12391 6171
rect 14013 6137 14047 6171
rect 15669 6137 15703 6171
rect 1777 6069 1811 6103
rect 2053 6069 2087 6103
rect 4261 6069 4295 6103
rect 12265 6069 12299 6103
rect 15577 6069 15611 6103
rect 18061 6069 18095 6103
rect 1961 5865 1995 5899
rect 3617 5865 3651 5899
rect 5457 5865 5491 5899
rect 16589 5865 16623 5899
rect 1685 5797 1719 5831
rect 2789 5797 2823 5831
rect 8769 5797 8803 5831
rect 13737 5797 13771 5831
rect 14105 5797 14139 5831
rect 17417 5797 17451 5831
rect 2237 5729 2271 5763
rect 2973 5729 3007 5763
rect 8125 5729 8159 5763
rect 14565 5729 14599 5763
rect 14657 5729 14691 5763
rect 15393 5729 15427 5763
rect 15485 5729 15519 5763
rect 16313 5729 16347 5763
rect 17141 5729 17175 5763
rect 17969 5729 18003 5763
rect 1777 5661 1811 5695
rect 2421 5661 2455 5695
rect 3249 5661 3283 5695
rect 4077 5661 4111 5695
rect 5549 5661 5583 5695
rect 5825 5661 5859 5695
rect 7941 5661 7975 5695
rect 8953 5661 8987 5695
rect 9220 5661 9254 5695
rect 12265 5661 12299 5695
rect 12521 5661 12555 5695
rect 13921 5661 13955 5695
rect 16221 5661 16255 5695
rect 17877 5661 17911 5695
rect 18245 5661 18279 5695
rect 1501 5593 1535 5627
rect 3157 5593 3191 5627
rect 4344 5593 4378 5627
rect 7696 5593 7730 5627
rect 10425 5593 10459 5627
rect 14473 5593 14507 5627
rect 16957 5593 16991 5627
rect 17785 5593 17819 5627
rect 2329 5525 2363 5559
rect 3985 5525 4019 5559
rect 6561 5525 6595 5559
rect 8309 5525 8343 5559
rect 8401 5525 8435 5559
rect 10333 5525 10367 5559
rect 11713 5525 11747 5559
rect 13645 5525 13679 5559
rect 14933 5525 14967 5559
rect 15301 5525 15335 5559
rect 15761 5525 15795 5559
rect 16129 5525 16163 5559
rect 17049 5525 17083 5559
rect 18429 5525 18463 5559
rect 2053 5321 2087 5355
rect 6101 5321 6135 5355
rect 6837 5321 6871 5355
rect 8585 5321 8619 5355
rect 9045 5321 9079 5355
rect 9413 5321 9447 5355
rect 9505 5321 9539 5355
rect 18429 5321 18463 5355
rect 1961 5253 1995 5287
rect 4896 5253 4930 5287
rect 8677 5253 8711 5287
rect 13001 5253 13035 5287
rect 14933 5253 14967 5287
rect 15292 5253 15326 5287
rect 1409 5185 1443 5219
rect 3626 5185 3660 5219
rect 3985 5185 4019 5219
rect 4261 5185 4295 5219
rect 6929 5185 6963 5219
rect 7757 5185 7791 5219
rect 10986 5185 11020 5219
rect 12653 5185 12687 5219
rect 16773 5185 16807 5219
rect 17509 5185 17543 5219
rect 17969 5185 18003 5219
rect 18245 5185 18279 5219
rect 1869 5117 1903 5151
rect 3893 5117 3927 5151
rect 4629 5117 4663 5151
rect 6469 5117 6503 5151
rect 6745 5117 6779 5151
rect 7849 5117 7883 5151
rect 8033 5117 8067 5151
rect 8861 5117 8895 5151
rect 9689 5117 9723 5151
rect 11253 5117 11287 5151
rect 12909 5117 12943 5151
rect 15025 5117 15059 5151
rect 17601 5117 17635 5151
rect 17693 5117 17727 5151
rect 2421 5049 2455 5083
rect 4169 5049 4203 5083
rect 7297 5049 7331 5083
rect 14289 5049 14323 5083
rect 1593 4981 1627 5015
rect 2513 4981 2547 5015
rect 4445 4981 4479 5015
rect 6009 4981 6043 5015
rect 7389 4981 7423 5015
rect 8217 4981 8251 5015
rect 9873 4981 9907 5015
rect 11529 4981 11563 5015
rect 16405 4981 16439 5015
rect 16957 4981 16991 5015
rect 17141 4981 17175 5015
rect 18153 4981 18187 5015
rect 1869 4777 1903 4811
rect 2881 4777 2915 4811
rect 3801 4777 3835 4811
rect 10425 4777 10459 4811
rect 12081 4777 12115 4811
rect 18429 4777 18463 4811
rect 6193 4709 6227 4743
rect 10333 4709 10367 4743
rect 14105 4709 14139 4743
rect 2145 4641 2179 4675
rect 2329 4641 2363 4675
rect 3433 4641 3467 4675
rect 4997 4641 5031 4675
rect 5273 4641 5307 4675
rect 8309 4641 8343 4675
rect 9321 4641 9355 4675
rect 9781 4641 9815 4675
rect 10885 4641 10919 4675
rect 10977 4641 11011 4675
rect 11805 4641 11839 4675
rect 12633 4641 12667 4675
rect 13553 4641 13587 4675
rect 16221 4641 16255 4675
rect 17141 4641 17175 4675
rect 17969 4641 18003 4675
rect 1409 4573 1443 4607
rect 1685 4573 1719 4607
rect 2421 4573 2455 4607
rect 3985 4573 4019 4607
rect 4353 4573 4387 4607
rect 5549 4573 5583 4607
rect 6837 4573 6871 4607
rect 8677 4573 8711 4607
rect 8953 4573 8987 4607
rect 9965 4573 9999 4607
rect 11621 4573 11655 4607
rect 13461 4573 13495 4607
rect 15485 4573 15519 4607
rect 15945 4573 15979 4607
rect 16957 4573 16991 4607
rect 18245 4573 18279 4607
rect 4813 4505 4847 4539
rect 8064 4505 8098 4539
rect 9873 4505 9907 4539
rect 12449 4505 12483 4539
rect 15218 4505 15252 4539
rect 16037 4505 16071 4539
rect 17049 4505 17083 4539
rect 17785 4505 17819 4539
rect 1593 4437 1627 4471
rect 2789 4437 2823 4471
rect 3249 4437 3283 4471
rect 3341 4437 3375 4471
rect 4169 4437 4203 4471
rect 4445 4437 4479 4471
rect 4905 4437 4939 4471
rect 6929 4437 6963 4471
rect 8493 4437 8527 4471
rect 9137 4437 9171 4471
rect 10793 4437 10827 4471
rect 11253 4437 11287 4471
rect 11713 4437 11747 4471
rect 12541 4437 12575 4471
rect 13001 4437 13035 4471
rect 13369 4437 13403 4471
rect 13921 4437 13955 4471
rect 15577 4437 15611 4471
rect 16405 4437 16439 4471
rect 16589 4437 16623 4471
rect 17417 4437 17451 4471
rect 17877 4437 17911 4471
rect 5089 4233 5123 4267
rect 5457 4233 5491 4267
rect 10057 4233 10091 4267
rect 10977 4233 11011 4267
rect 12633 4233 12667 4267
rect 13829 4233 13863 4267
rect 14197 4233 14231 4267
rect 17417 4233 17451 4267
rect 4997 4165 5031 4199
rect 11897 4165 11931 4199
rect 13001 4165 13035 4199
rect 17785 4165 17819 4199
rect 2533 4097 2567 4131
rect 4097 4097 4131 4131
rect 4353 4097 4387 4131
rect 4537 4097 4571 4131
rect 5825 4097 5859 4131
rect 7501 4097 7535 4131
rect 8125 4097 8159 4131
rect 8484 4097 8518 4131
rect 10885 4097 10919 4131
rect 12541 4097 12575 4131
rect 13461 4097 13495 4131
rect 14657 4097 14691 4131
rect 16149 4097 16183 4131
rect 16405 4097 16439 4131
rect 17325 4097 17359 4131
rect 17877 4097 17911 4131
rect 18245 4097 18279 4131
rect 2789 4029 2823 4063
rect 5273 4029 5307 4063
rect 5917 4029 5951 4063
rect 6101 4029 6135 4063
rect 7757 4029 7791 4063
rect 8217 4029 8251 4063
rect 9781 4029 9815 4063
rect 9965 4029 9999 4063
rect 11161 4029 11195 4063
rect 11989 4029 12023 4063
rect 12081 4029 12115 4063
rect 13093 4029 13127 4063
rect 13277 4029 13311 4063
rect 14289 4029 14323 4063
rect 14473 4029 14507 4063
rect 17969 4029 18003 4063
rect 10425 3961 10459 3995
rect 13645 3961 13679 3995
rect 14841 3961 14875 3995
rect 16681 3961 16715 3995
rect 18429 3961 18463 3995
rect 1409 3893 1443 3927
rect 2973 3893 3007 3927
rect 4629 3893 4663 3927
rect 6377 3893 6411 3927
rect 7941 3893 7975 3927
rect 9597 3893 9631 3927
rect 10517 3893 10551 3927
rect 11529 3893 11563 3927
rect 12357 3893 12391 3927
rect 15025 3893 15059 3927
rect 11069 3689 11103 3723
rect 13737 3689 13771 3723
rect 17601 3689 17635 3723
rect 18521 3689 18555 3723
rect 1501 3621 1535 3655
rect 6561 3621 6595 3655
rect 12541 3621 12575 3655
rect 14105 3621 14139 3655
rect 2513 3553 2547 3587
rect 3341 3553 3375 3587
rect 3985 3553 4019 3587
rect 4629 3553 4663 3587
rect 7113 3553 7147 3587
rect 7849 3553 7883 3587
rect 8033 3553 8067 3587
rect 8953 3553 8987 3587
rect 13185 3553 13219 3587
rect 14749 3553 14783 3587
rect 15485 3553 15519 3587
rect 16129 3553 16163 3587
rect 16865 3553 16899 3587
rect 17003 3553 17037 3587
rect 18153 3553 18187 3587
rect 1869 3485 1903 3519
rect 4169 3485 4203 3519
rect 4885 3485 4919 3519
rect 6469 3485 6503 3519
rect 6929 3485 6963 3519
rect 8493 3485 8527 3519
rect 10425 3485 10459 3519
rect 11161 3485 11195 3519
rect 12633 3485 12667 3519
rect 13829 3485 13863 3519
rect 14473 3485 14507 3519
rect 15761 3485 15795 3519
rect 16773 3485 16807 3519
rect 17233 3485 17267 3519
rect 18061 3485 18095 3519
rect 2421 3417 2455 3451
rect 9220 3417 9254 3451
rect 11428 3417 11462 3451
rect 17969 3417 18003 3451
rect 1685 3349 1719 3383
rect 1961 3349 1995 3383
rect 2329 3349 2363 3383
rect 2789 3349 2823 3383
rect 3157 3349 3191 3383
rect 3249 3349 3283 3383
rect 4077 3349 4111 3383
rect 4537 3349 4571 3383
rect 6009 3349 6043 3383
rect 6285 3349 6319 3383
rect 7021 3349 7055 3383
rect 7389 3349 7423 3383
rect 7757 3349 7791 3383
rect 8401 3349 8435 3383
rect 8677 3349 8711 3383
rect 10333 3349 10367 3383
rect 12817 3349 12851 3383
rect 13277 3349 13311 3383
rect 13369 3349 13403 3383
rect 14565 3349 14599 3383
rect 14933 3349 14967 3383
rect 15301 3349 15335 3383
rect 15393 3349 15427 3383
rect 15945 3349 15979 3383
rect 16405 3349 16439 3383
rect 17417 3349 17451 3383
rect 1593 3145 1627 3179
rect 1961 3145 1995 3179
rect 2053 3145 2087 3179
rect 6745 3145 6779 3179
rect 8309 3145 8343 3179
rect 10149 3145 10183 3179
rect 10885 3145 10919 3179
rect 11529 3145 11563 3179
rect 14105 3145 14139 3179
rect 14565 3145 14599 3179
rect 15117 3145 15151 3179
rect 15393 3145 15427 3179
rect 15761 3145 15795 3179
rect 15853 3145 15887 3179
rect 17509 3145 17543 3179
rect 17969 3145 18003 3179
rect 2789 3077 2823 3111
rect 4353 3077 4387 3111
rect 4997 3077 5031 3111
rect 7113 3077 7147 3111
rect 9597 3077 9631 3111
rect 10057 3077 10091 3111
rect 11897 3077 11931 3111
rect 11989 3077 12023 3111
rect 12900 3077 12934 3111
rect 17049 3077 17083 3111
rect 18429 3077 18463 3111
rect 1409 3009 1443 3043
rect 4905 3009 4939 3043
rect 5733 3009 5767 3043
rect 6653 3009 6687 3043
rect 7565 3013 7599 3047
rect 12541 3009 12575 3043
rect 14473 3009 14507 3043
rect 14933 3009 14967 3043
rect 16221 3009 16255 3043
rect 16681 3009 16715 3043
rect 17601 3009 17635 3043
rect 18061 3009 18095 3043
rect 1869 2941 1903 2975
rect 5181 2941 5215 2975
rect 5825 2941 5859 2975
rect 6009 2941 6043 2975
rect 7205 2941 7239 2975
rect 7389 2941 7423 2975
rect 10241 2941 10275 2975
rect 10977 2941 11011 2975
rect 11069 2941 11103 2975
rect 12081 2941 12115 2975
rect 12633 2941 12667 2975
rect 14657 2941 14691 2975
rect 15945 2941 15979 2975
rect 17417 2941 17451 2975
rect 2421 2873 2455 2907
rect 6469 2873 6503 2907
rect 7757 2873 7791 2907
rect 10517 2873 10551 2907
rect 12357 2873 12391 2907
rect 16405 2873 16439 2907
rect 16865 2873 16899 2907
rect 4537 2805 4571 2839
rect 5365 2805 5399 2839
rect 9689 2805 9723 2839
rect 14013 2805 14047 2839
rect 18245 2805 18279 2839
rect 3617 2601 3651 2635
rect 4629 2601 4663 2635
rect 7573 2601 7607 2635
rect 10701 2601 10735 2635
rect 14105 2601 14139 2635
rect 15577 2601 15611 2635
rect 3433 2533 3467 2567
rect 6193 2533 6227 2567
rect 16313 2533 16347 2567
rect 18061 2533 18095 2567
rect 2053 2465 2087 2499
rect 2145 2465 2179 2499
rect 2789 2465 2823 2499
rect 2973 2465 3007 2499
rect 3893 2465 3927 2499
rect 5273 2465 5307 2499
rect 5641 2465 5675 2499
rect 6929 2465 6963 2499
rect 8125 2465 8159 2499
rect 8953 2465 8987 2499
rect 9229 2465 9263 2499
rect 9413 2465 9447 2499
rect 10149 2465 10183 2499
rect 12081 2465 12115 2499
rect 12541 2465 12575 2499
rect 13277 2465 13311 2499
rect 14657 2465 14691 2499
rect 1777 2397 1811 2431
rect 3065 2397 3099 2431
rect 4169 2397 4203 2431
rect 4997 2397 5031 2431
rect 5825 2397 5859 2431
rect 6653 2397 6687 2431
rect 8493 2397 8527 2431
rect 9505 2397 9539 2431
rect 10333 2397 10367 2431
rect 10793 2397 10827 2431
rect 11345 2397 11379 2431
rect 11897 2397 11931 2431
rect 13461 2397 13495 2431
rect 14565 2397 14599 2431
rect 14933 2397 14967 2431
rect 15669 2397 15703 2431
rect 16681 2397 16715 2431
rect 17417 2397 17451 2431
rect 18153 2397 18187 2431
rect 4077 2329 4111 2363
rect 5733 2329 5767 2363
rect 8033 2329 8067 2363
rect 10241 2329 10275 2363
rect 13553 2329 13587 2363
rect 14473 2329 14507 2363
rect 1593 2261 1627 2295
rect 2237 2261 2271 2295
rect 2605 2261 2639 2295
rect 4537 2261 4571 2295
rect 5089 2261 5123 2295
rect 6469 2261 6503 2295
rect 7021 2261 7055 2295
rect 7113 2261 7147 2295
rect 7481 2261 7515 2295
rect 7941 2261 7975 2295
rect 8677 2261 8711 2295
rect 9873 2261 9907 2295
rect 10977 2261 11011 2295
rect 11161 2261 11195 2295
rect 11529 2261 11563 2295
rect 11989 2261 12023 2295
rect 12633 2261 12667 2295
rect 12725 2261 12759 2295
rect 13093 2261 13127 2295
rect 13921 2261 13955 2295
rect 16405 2261 16439 2295
rect 17325 2261 17359 2295
rect 18337 2261 18371 2295
<< metal1 >>
rect 6546 15784 6552 15836
rect 6604 15824 6610 15836
rect 14826 15824 14832 15836
rect 6604 15796 14832 15824
rect 6604 15784 6610 15796
rect 14826 15784 14832 15796
rect 14884 15784 14890 15836
rect 4246 15648 4252 15700
rect 4304 15688 4310 15700
rect 14550 15688 14556 15700
rect 4304 15660 14556 15688
rect 4304 15648 4310 15660
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 2682 15580 2688 15632
rect 2740 15620 2746 15632
rect 14642 15620 14648 15632
rect 2740 15592 14648 15620
rect 2740 15580 2746 15592
rect 14642 15580 14648 15592
rect 14700 15580 14706 15632
rect 5258 15512 5264 15564
rect 5316 15552 5322 15564
rect 17954 15552 17960 15564
rect 5316 15524 17960 15552
rect 5316 15512 5322 15524
rect 17954 15512 17960 15524
rect 18012 15512 18018 15564
rect 750 15444 756 15496
rect 808 15484 814 15496
rect 8110 15484 8116 15496
rect 808 15456 8116 15484
rect 808 15444 814 15456
rect 8110 15444 8116 15456
rect 8168 15444 8174 15496
rect 13354 15444 13360 15496
rect 13412 15484 13418 15496
rect 13906 15484 13912 15496
rect 13412 15456 13912 15484
rect 13412 15444 13418 15456
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14 15376 20 15428
rect 72 15416 78 15428
rect 8478 15416 8484 15428
rect 72 15388 8484 15416
rect 72 15376 78 15388
rect 8478 15376 8484 15388
rect 8536 15376 8542 15428
rect 10318 15376 10324 15428
rect 10376 15416 10382 15428
rect 19886 15416 19892 15428
rect 10376 15388 19892 15416
rect 10376 15376 10382 15388
rect 19886 15376 19892 15388
rect 19944 15376 19950 15428
rect 2314 15308 2320 15360
rect 2372 15348 2378 15360
rect 6454 15348 6460 15360
rect 2372 15320 6460 15348
rect 2372 15308 2378 15320
rect 6454 15308 6460 15320
rect 6512 15308 6518 15360
rect 11974 15308 11980 15360
rect 12032 15348 12038 15360
rect 18506 15348 18512 15360
rect 12032 15320 18512 15348
rect 12032 15308 12038 15320
rect 18506 15308 18512 15320
rect 18564 15308 18570 15360
rect 2038 15240 2044 15292
rect 2096 15280 2102 15292
rect 5810 15280 5816 15292
rect 2096 15252 5816 15280
rect 2096 15240 2102 15252
rect 5810 15240 5816 15252
rect 5868 15240 5874 15292
rect 12434 15240 12440 15292
rect 12492 15280 12498 15292
rect 15470 15280 15476 15292
rect 12492 15252 15476 15280
rect 12492 15240 12498 15252
rect 15470 15240 15476 15252
rect 15528 15240 15534 15292
rect 2130 15172 2136 15224
rect 2188 15212 2194 15224
rect 6638 15212 6644 15224
rect 2188 15184 6644 15212
rect 2188 15172 2194 15184
rect 6638 15172 6644 15184
rect 6696 15172 6702 15224
rect 12618 15172 12624 15224
rect 12676 15212 12682 15224
rect 12676 15184 15240 15212
rect 12676 15172 12682 15184
rect 7190 15144 7196 15156
rect 2746 15116 7196 15144
rect 2498 15036 2504 15088
rect 2556 15076 2562 15088
rect 2746 15076 2774 15116
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 10502 15104 10508 15156
rect 10560 15144 10566 15156
rect 15212 15144 15240 15184
rect 17586 15144 17592 15156
rect 10560 15116 15148 15144
rect 15212 15116 17592 15144
rect 10560 15104 10566 15116
rect 2556 15048 2774 15076
rect 2556 15036 2562 15048
rect 3786 15036 3792 15088
rect 3844 15076 3850 15088
rect 6914 15076 6920 15088
rect 3844 15048 6920 15076
rect 3844 15036 3850 15048
rect 6914 15036 6920 15048
rect 6972 15036 6978 15088
rect 11606 15036 11612 15088
rect 11664 15076 11670 15088
rect 15010 15076 15016 15088
rect 11664 15048 15016 15076
rect 11664 15036 11670 15048
rect 15010 15036 15016 15048
rect 15068 15036 15074 15088
rect 15120 15076 15148 15116
rect 17586 15104 17592 15116
rect 17644 15104 17650 15156
rect 15286 15076 15292 15088
rect 15120 15048 15292 15076
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 15470 15036 15476 15088
rect 15528 15076 15534 15088
rect 17678 15076 17684 15088
rect 15528 15048 17684 15076
rect 15528 15036 15534 15048
rect 17678 15036 17684 15048
rect 17736 15036 17742 15088
rect 4062 14968 4068 15020
rect 4120 15008 4126 15020
rect 6730 15008 6736 15020
rect 4120 14980 6736 15008
rect 4120 14968 4126 14980
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 12802 14968 12808 15020
rect 12860 15008 12866 15020
rect 16298 15008 16304 15020
rect 12860 14980 16304 15008
rect 12860 14968 12866 14980
rect 16298 14968 16304 14980
rect 16356 14968 16362 15020
rect 4338 14900 4344 14952
rect 4396 14940 4402 14952
rect 6086 14940 6092 14952
rect 4396 14912 6092 14940
rect 4396 14900 4402 14912
rect 6086 14900 6092 14912
rect 6144 14900 6150 14952
rect 7098 14900 7104 14952
rect 7156 14940 7162 14952
rect 10594 14940 10600 14952
rect 7156 14912 10600 14940
rect 7156 14900 7162 14912
rect 10594 14900 10600 14912
rect 10652 14940 10658 14952
rect 12894 14940 12900 14952
rect 10652 14912 12900 14940
rect 10652 14900 10658 14912
rect 12894 14900 12900 14912
rect 12952 14900 12958 14952
rect 13170 14900 13176 14952
rect 13228 14940 13234 14952
rect 15654 14940 15660 14952
rect 13228 14912 15660 14940
rect 13228 14900 13234 14912
rect 15654 14900 15660 14912
rect 15712 14900 15718 14952
rect 3878 14832 3884 14884
rect 3936 14872 3942 14884
rect 5994 14872 6000 14884
rect 3936 14844 6000 14872
rect 3936 14832 3942 14844
rect 5994 14832 6000 14844
rect 6052 14832 6058 14884
rect 6178 14832 6184 14884
rect 6236 14872 6242 14884
rect 11422 14872 11428 14884
rect 6236 14844 11428 14872
rect 6236 14832 6242 14844
rect 11422 14832 11428 14844
rect 11480 14832 11486 14884
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 16390 14872 16396 14884
rect 12584 14844 16396 14872
rect 12584 14832 12590 14844
rect 16390 14832 16396 14844
rect 16448 14832 16454 14884
rect 2866 14764 2872 14816
rect 2924 14804 2930 14816
rect 4430 14804 4436 14816
rect 2924 14776 4436 14804
rect 2924 14764 2930 14776
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 12986 14764 12992 14816
rect 13044 14804 13050 14816
rect 16022 14804 16028 14816
rect 13044 14776 16028 14804
rect 13044 14764 13050 14776
rect 16022 14764 16028 14776
rect 16080 14764 16086 14816
rect 1104 14714 18860 14736
rect 1104 14662 3174 14714
rect 3226 14662 3238 14714
rect 3290 14662 3302 14714
rect 3354 14662 3366 14714
rect 3418 14662 3430 14714
rect 3482 14662 7622 14714
rect 7674 14662 7686 14714
rect 7738 14662 7750 14714
rect 7802 14662 7814 14714
rect 7866 14662 7878 14714
rect 7930 14662 12070 14714
rect 12122 14662 12134 14714
rect 12186 14662 12198 14714
rect 12250 14662 12262 14714
rect 12314 14662 12326 14714
rect 12378 14662 16518 14714
rect 16570 14662 16582 14714
rect 16634 14662 16646 14714
rect 16698 14662 16710 14714
rect 16762 14662 16774 14714
rect 16826 14662 18860 14714
rect 1104 14640 18860 14662
rect 2774 14560 2780 14612
rect 2832 14600 2838 14612
rect 2832 14572 2877 14600
rect 2832 14560 2838 14572
rect 2958 14560 2964 14612
rect 3016 14600 3022 14612
rect 3145 14603 3203 14609
rect 3145 14600 3157 14603
rect 3016 14572 3157 14600
rect 3016 14560 3022 14572
rect 3145 14569 3157 14572
rect 3191 14569 3203 14603
rect 3145 14563 3203 14569
rect 3988 14572 4200 14600
rect 2222 14492 2228 14544
rect 2280 14532 2286 14544
rect 3988 14532 4016 14572
rect 2280 14504 4016 14532
rect 4172 14532 4200 14572
rect 4246 14560 4252 14612
rect 4304 14600 4310 14612
rect 4522 14600 4528 14612
rect 4304 14572 4528 14600
rect 4304 14560 4310 14572
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 4617 14603 4675 14609
rect 4617 14569 4629 14603
rect 4663 14600 4675 14603
rect 4706 14600 4712 14612
rect 4663 14572 4712 14600
rect 4663 14569 4675 14572
rect 4617 14563 4675 14569
rect 4706 14560 4712 14572
rect 4764 14560 4770 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5721 14603 5779 14609
rect 5721 14600 5733 14603
rect 4856 14572 5733 14600
rect 4856 14560 4862 14572
rect 5721 14569 5733 14572
rect 5767 14569 5779 14603
rect 5721 14563 5779 14569
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 6549 14603 6607 14609
rect 6549 14600 6561 14603
rect 5960 14572 6561 14600
rect 5960 14560 5966 14572
rect 6549 14569 6561 14572
rect 6595 14569 6607 14603
rect 6549 14563 6607 14569
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 7101 14603 7159 14609
rect 7101 14600 7113 14603
rect 6696 14572 7113 14600
rect 6696 14560 6702 14572
rect 7101 14569 7113 14572
rect 7147 14569 7159 14603
rect 7374 14600 7380 14612
rect 7287 14572 7380 14600
rect 7101 14563 7159 14569
rect 7374 14560 7380 14572
rect 7432 14600 7438 14612
rect 11882 14600 11888 14612
rect 7432 14572 11888 14600
rect 7432 14560 7438 14572
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 11974 14560 11980 14612
rect 12032 14600 12038 14612
rect 12161 14603 12219 14609
rect 12161 14600 12173 14603
rect 12032 14572 12173 14600
rect 12032 14560 12038 14572
rect 12161 14569 12173 14572
rect 12207 14569 12219 14603
rect 12161 14563 12219 14569
rect 12434 14560 12440 14612
rect 12492 14600 12498 14612
rect 12618 14600 12624 14612
rect 12492 14572 12537 14600
rect 12579 14572 12624 14600
rect 12492 14560 12498 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 12802 14600 12808 14612
rect 12763 14572 12808 14600
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 12986 14600 12992 14612
rect 12947 14572 12992 14600
rect 12986 14560 12992 14572
rect 13044 14560 13050 14612
rect 13170 14600 13176 14612
rect 13131 14572 13176 14600
rect 13170 14560 13176 14572
rect 13228 14560 13234 14612
rect 13998 14600 14004 14612
rect 13280 14572 14004 14600
rect 5077 14535 5135 14541
rect 4172 14504 4936 14532
rect 2280 14492 2286 14504
rect 1946 14464 1952 14476
rect 1907 14436 1952 14464
rect 1946 14424 1952 14436
rect 2004 14424 2010 14476
rect 2866 14464 2872 14476
rect 2608 14436 2872 14464
rect 2130 14356 2136 14408
rect 2188 14396 2194 14408
rect 2608 14405 2636 14436
rect 2866 14424 2872 14436
rect 2924 14424 2930 14476
rect 3970 14464 3976 14476
rect 3344 14436 3976 14464
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 2188 14368 2237 14396
rect 2188 14356 2194 14368
rect 2225 14365 2237 14368
rect 2271 14365 2283 14399
rect 2225 14359 2283 14365
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14365 2651 14399
rect 2593 14359 2651 14365
rect 2961 14399 3019 14405
rect 2961 14365 2973 14399
rect 3007 14396 3019 14399
rect 3234 14396 3240 14408
rect 3007 14368 3240 14396
rect 3007 14365 3019 14368
rect 2961 14359 3019 14365
rect 3234 14356 3240 14368
rect 3292 14356 3298 14408
rect 3344 14405 3372 14436
rect 3970 14424 3976 14436
rect 4028 14424 4034 14476
rect 3329 14399 3387 14405
rect 3329 14365 3341 14399
rect 3375 14365 3387 14399
rect 3329 14359 3387 14365
rect 3418 14356 3424 14408
rect 3476 14396 3482 14408
rect 3605 14399 3663 14405
rect 3605 14396 3617 14399
rect 3476 14368 3617 14396
rect 3476 14356 3482 14368
rect 3605 14365 3617 14368
rect 3651 14365 3663 14399
rect 3786 14396 3792 14408
rect 3747 14368 3792 14396
rect 3605 14359 3663 14365
rect 3786 14356 3792 14368
rect 3844 14356 3850 14408
rect 4062 14396 4068 14408
rect 4023 14368 4068 14396
rect 4062 14356 4068 14368
rect 4120 14356 4126 14408
rect 4338 14396 4344 14408
rect 4299 14368 4344 14396
rect 4338 14356 4344 14368
rect 4396 14356 4402 14408
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4908 14405 4936 14504
rect 5077 14501 5089 14535
rect 5123 14501 5135 14535
rect 5077 14495 5135 14501
rect 5261 14535 5319 14541
rect 5261 14501 5273 14535
rect 5307 14532 5319 14535
rect 5350 14532 5356 14544
rect 5307 14504 5356 14532
rect 5307 14501 5319 14504
rect 5261 14495 5319 14501
rect 5092 14464 5120 14495
rect 5350 14492 5356 14504
rect 5408 14492 5414 14544
rect 5994 14532 6000 14544
rect 5955 14504 6000 14532
rect 5994 14492 6000 14504
rect 6052 14492 6058 14544
rect 6086 14492 6092 14544
rect 6144 14532 6150 14544
rect 6730 14532 6736 14544
rect 6144 14504 6189 14532
rect 6691 14504 6736 14532
rect 6144 14492 6150 14504
rect 6730 14492 6736 14504
rect 6788 14492 6794 14544
rect 6914 14532 6920 14544
rect 6875 14504 6920 14532
rect 6914 14492 6920 14504
rect 6972 14492 6978 14544
rect 7006 14492 7012 14544
rect 7064 14532 7070 14544
rect 11606 14532 11612 14544
rect 7064 14504 11612 14532
rect 7064 14492 7070 14504
rect 11606 14492 11612 14504
rect 11664 14492 11670 14544
rect 11790 14492 11796 14544
rect 11848 14532 11854 14544
rect 13280 14532 13308 14572
rect 13998 14560 14004 14572
rect 14056 14600 14062 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 14056 14572 14105 14600
rect 14056 14560 14062 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 14461 14603 14519 14609
rect 14461 14569 14473 14603
rect 14507 14600 14519 14603
rect 17862 14600 17868 14612
rect 14507 14572 17868 14600
rect 14507 14569 14519 14572
rect 14461 14563 14519 14569
rect 17862 14560 17868 14572
rect 17920 14560 17926 14612
rect 15010 14532 15016 14544
rect 11848 14504 13308 14532
rect 13464 14504 15016 14532
rect 11848 14492 11854 14504
rect 13170 14464 13176 14476
rect 5092 14436 6960 14464
rect 4777 14399 4835 14405
rect 4777 14396 4789 14399
rect 4672 14368 4789 14396
rect 4672 14356 4678 14368
rect 4777 14365 4789 14368
rect 4823 14365 4835 14399
rect 4777 14359 4835 14365
rect 4893 14399 4951 14405
rect 4893 14365 4905 14399
rect 4939 14396 4951 14399
rect 5537 14399 5595 14405
rect 5537 14396 5549 14399
rect 4939 14368 5549 14396
rect 4939 14365 4951 14368
rect 4893 14359 4951 14365
rect 5537 14365 5549 14368
rect 5583 14365 5595 14399
rect 6362 14396 6368 14408
rect 6323 14368 6368 14396
rect 5537 14359 5595 14365
rect 6362 14356 6368 14368
rect 6420 14356 6426 14408
rect 6932 14396 6960 14436
rect 9324 14436 13176 14464
rect 9324 14396 9352 14436
rect 13170 14424 13176 14436
rect 13228 14424 13234 14476
rect 6932 14368 9352 14396
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 9953 14399 10011 14405
rect 9953 14396 9965 14399
rect 9824 14368 9965 14396
rect 9824 14356 9830 14368
rect 9953 14365 9965 14368
rect 9999 14365 10011 14399
rect 9953 14359 10011 14365
rect 9674 14328 9680 14340
rect 2746 14300 3464 14328
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 2590 14220 2596 14272
rect 2648 14260 2654 14272
rect 2746 14260 2774 14300
rect 3436 14269 3464 14300
rect 3988 14300 9680 14328
rect 3988 14269 4016 14300
rect 9674 14288 9680 14300
rect 9732 14288 9738 14340
rect 13464 14337 13492 14504
rect 15010 14492 15016 14504
rect 15068 14492 15074 14544
rect 15102 14492 15108 14544
rect 15160 14532 15166 14544
rect 15160 14504 15205 14532
rect 15160 14492 15166 14504
rect 13725 14467 13783 14473
rect 13725 14433 13737 14467
rect 13771 14464 13783 14467
rect 13906 14464 13912 14476
rect 13771 14436 13912 14464
rect 13771 14433 13783 14436
rect 13725 14427 13783 14433
rect 13906 14424 13912 14436
rect 13964 14424 13970 14476
rect 16942 14464 16948 14476
rect 14200 14436 16948 14464
rect 13449 14331 13507 14337
rect 13449 14328 13461 14331
rect 10060 14300 13461 14328
rect 2648 14232 2774 14260
rect 3421 14263 3479 14269
rect 2648 14220 2654 14232
rect 3421 14229 3433 14263
rect 3467 14229 3479 14263
rect 3421 14223 3479 14229
rect 3973 14263 4031 14269
rect 3973 14229 3985 14263
rect 4019 14229 4031 14263
rect 3973 14223 4031 14229
rect 4525 14263 4583 14269
rect 4525 14229 4537 14263
rect 4571 14260 4583 14263
rect 4614 14260 4620 14272
rect 4571 14232 4620 14260
rect 4571 14229 4583 14232
rect 4525 14223 4583 14229
rect 4614 14220 4620 14232
rect 4672 14220 4678 14272
rect 4890 14220 4896 14272
rect 4948 14260 4954 14272
rect 5353 14263 5411 14269
rect 5353 14260 5365 14263
rect 4948 14232 5365 14260
rect 4948 14220 4954 14232
rect 5353 14229 5365 14232
rect 5399 14260 5411 14263
rect 8570 14260 8576 14272
rect 5399 14232 8576 14260
rect 5399 14229 5411 14232
rect 5353 14223 5411 14229
rect 8570 14220 8576 14232
rect 8628 14220 8634 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 10060 14260 10088 14300
rect 13449 14297 13461 14300
rect 13495 14297 13507 14331
rect 13814 14328 13820 14340
rect 13775 14300 13820 14328
rect 13449 14291 13507 14297
rect 13814 14288 13820 14300
rect 13872 14328 13878 14340
rect 14090 14328 14096 14340
rect 13872 14300 14096 14328
rect 13872 14288 13878 14300
rect 14090 14288 14096 14300
rect 14148 14288 14154 14340
rect 9088 14232 10088 14260
rect 10137 14263 10195 14269
rect 9088 14220 9094 14232
rect 10137 14229 10149 14263
rect 10183 14260 10195 14263
rect 10410 14260 10416 14272
rect 10183 14232 10416 14260
rect 10183 14229 10195 14232
rect 10137 14223 10195 14229
rect 10410 14220 10416 14232
rect 10468 14220 10474 14272
rect 11974 14260 11980 14272
rect 11935 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 13357 14263 13415 14269
rect 13357 14229 13369 14263
rect 13403 14260 13415 14263
rect 14200 14260 14228 14436
rect 14277 14399 14335 14405
rect 14277 14365 14289 14399
rect 14323 14365 14335 14399
rect 14550 14396 14556 14408
rect 14511 14368 14556 14396
rect 14277 14359 14335 14365
rect 14292 14328 14320 14359
rect 14550 14356 14556 14368
rect 14608 14356 14614 14408
rect 15010 14356 15016 14408
rect 15068 14396 15074 14408
rect 15304 14405 15332 14436
rect 16942 14424 16948 14436
rect 17000 14424 17006 14476
rect 17310 14464 17316 14476
rect 17271 14436 17316 14464
rect 17310 14424 17316 14436
rect 17368 14424 17374 14476
rect 17586 14464 17592 14476
rect 17547 14436 17592 14464
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 18506 14464 18512 14476
rect 18467 14436 18512 14464
rect 18506 14424 18512 14436
rect 18564 14424 18570 14476
rect 15289 14399 15347 14405
rect 15068 14368 15113 14396
rect 15068 14356 15074 14368
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15654 14396 15660 14408
rect 15615 14368 15660 14396
rect 15289 14359 15347 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15838 14396 15844 14408
rect 15799 14368 15844 14396
rect 15838 14356 15844 14368
rect 15896 14356 15902 14408
rect 16022 14396 16028 14408
rect 15983 14368 16028 14396
rect 16022 14356 16028 14368
rect 16080 14356 16086 14408
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16393 14399 16451 14405
rect 16393 14396 16405 14399
rect 16356 14368 16405 14396
rect 16356 14356 16362 14368
rect 16393 14365 16405 14368
rect 16439 14365 16451 14399
rect 18230 14396 18236 14408
rect 18143 14368 18236 14396
rect 16393 14359 16451 14365
rect 18230 14356 18236 14368
rect 18288 14396 18294 14408
rect 19610 14396 19616 14408
rect 18288 14368 19616 14396
rect 18288 14356 18294 14368
rect 19610 14356 19616 14368
rect 19668 14356 19674 14408
rect 15102 14328 15108 14340
rect 14292 14300 15108 14328
rect 15102 14288 15108 14300
rect 15160 14288 15166 14340
rect 15194 14288 15200 14340
rect 15252 14328 15258 14340
rect 15473 14331 15531 14337
rect 15473 14328 15485 14331
rect 15252 14300 15485 14328
rect 15252 14288 15258 14300
rect 15473 14297 15485 14300
rect 15519 14328 15531 14331
rect 17402 14328 17408 14340
rect 15519 14300 17408 14328
rect 15519 14297 15531 14300
rect 15473 14291 15531 14297
rect 17402 14288 17408 14300
rect 17460 14288 17466 14340
rect 14734 14260 14740 14272
rect 13403 14232 14228 14260
rect 14695 14232 14740 14260
rect 13403 14229 13415 14232
rect 13357 14223 13415 14229
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 14829 14263 14887 14269
rect 14829 14229 14841 14263
rect 14875 14260 14887 14263
rect 15010 14260 15016 14272
rect 14875 14232 15016 14260
rect 14875 14229 14887 14232
rect 14829 14223 14887 14229
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 15286 14220 15292 14272
rect 15344 14260 15350 14272
rect 16301 14263 16359 14269
rect 16301 14260 16313 14263
rect 15344 14232 16313 14260
rect 15344 14220 15350 14232
rect 16301 14229 16313 14232
rect 16347 14260 16359 14263
rect 17586 14260 17592 14272
rect 16347 14232 17592 14260
rect 16347 14229 16359 14232
rect 16301 14223 16359 14229
rect 17586 14220 17592 14232
rect 17644 14220 17650 14272
rect 1104 14170 18860 14192
rect 1104 14118 5398 14170
rect 5450 14118 5462 14170
rect 5514 14118 5526 14170
rect 5578 14118 5590 14170
rect 5642 14118 5654 14170
rect 5706 14118 9846 14170
rect 9898 14118 9910 14170
rect 9962 14118 9974 14170
rect 10026 14118 10038 14170
rect 10090 14118 10102 14170
rect 10154 14118 14294 14170
rect 14346 14118 14358 14170
rect 14410 14118 14422 14170
rect 14474 14118 14486 14170
rect 14538 14118 14550 14170
rect 14602 14118 18860 14170
rect 1104 14096 18860 14118
rect 2774 14056 2780 14068
rect 2735 14028 2780 14056
rect 2774 14016 2780 14028
rect 2832 14016 2838 14068
rect 3418 14056 3424 14068
rect 3379 14028 3424 14056
rect 3418 14016 3424 14028
rect 3476 14016 3482 14068
rect 3605 14059 3663 14065
rect 3605 14025 3617 14059
rect 3651 14025 3663 14059
rect 4157 14059 4215 14065
rect 4157 14056 4169 14059
rect 3605 14019 3663 14025
rect 3712 14028 4169 14056
rect 1578 13948 1584 14000
rect 1636 13988 1642 14000
rect 2593 13991 2651 13997
rect 1636 13960 2553 13988
rect 1636 13948 1642 13960
rect 1118 13880 1124 13932
rect 1176 13920 1182 13932
rect 2222 13920 2228 13932
rect 1176 13892 2228 13920
rect 1176 13880 1182 13892
rect 2222 13880 2228 13892
rect 2280 13880 2286 13932
rect 2409 13923 2467 13929
rect 2409 13889 2421 13923
rect 2455 13889 2467 13923
rect 2525 13920 2553 13960
rect 2593 13957 2605 13991
rect 2639 13988 2651 13991
rect 2682 13988 2688 14000
rect 2639 13960 2688 13988
rect 2639 13957 2651 13960
rect 2593 13951 2651 13957
rect 2682 13948 2688 13960
rect 2740 13948 2746 14000
rect 3620 13988 3648 14019
rect 2976 13960 3648 13988
rect 2976 13929 3004 13960
rect 2961 13923 3019 13929
rect 2525 13892 2921 13920
rect 2409 13883 2467 13889
rect 1949 13855 2007 13861
rect 1949 13821 1961 13855
rect 1995 13852 2007 13855
rect 2038 13852 2044 13864
rect 1995 13824 2044 13852
rect 1995 13821 2007 13824
rect 1949 13815 2007 13821
rect 2038 13812 2044 13824
rect 2096 13812 2102 13864
rect 2424 13852 2452 13883
rect 2893 13852 2921 13892
rect 2961 13889 2973 13923
rect 3007 13889 3019 13923
rect 3234 13920 3240 13932
rect 3195 13892 3240 13920
rect 2961 13883 3019 13889
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 3326 13880 3332 13932
rect 3384 13920 3390 13932
rect 3712 13920 3740 14028
rect 4157 14025 4169 14028
rect 4203 14025 4215 14059
rect 4430 14056 4436 14068
rect 4391 14028 4436 14056
rect 4157 14019 4215 14025
rect 4430 14016 4436 14028
rect 4488 14016 4494 14068
rect 4706 14016 4712 14068
rect 4764 14016 4770 14068
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 4982 14056 4988 14068
rect 4847 14028 4988 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 4982 14016 4988 14028
rect 5040 14016 5046 14068
rect 5353 14059 5411 14065
rect 5353 14025 5365 14059
rect 5399 14056 5411 14059
rect 5810 14056 5816 14068
rect 5399 14028 5816 14056
rect 5399 14025 5411 14028
rect 5353 14019 5411 14025
rect 5810 14016 5816 14028
rect 5868 14016 5874 14068
rect 6362 14056 6368 14068
rect 6323 14028 6368 14056
rect 6362 14016 6368 14028
rect 6420 14016 6426 14068
rect 6454 14016 6460 14068
rect 6512 14056 6518 14068
rect 6641 14059 6699 14065
rect 6641 14056 6653 14059
rect 6512 14028 6653 14056
rect 6512 14016 6518 14028
rect 6641 14025 6653 14028
rect 6687 14025 6699 14059
rect 7006 14056 7012 14068
rect 6641 14019 6699 14025
rect 6748 14028 7012 14056
rect 4724 13988 4752 14016
rect 5166 13988 5172 14000
rect 3804 13960 4752 13988
rect 5079 13960 5172 13988
rect 3804 13929 3832 13960
rect 5166 13948 5172 13960
rect 5224 13988 5230 14000
rect 5626 13988 5632 14000
rect 5224 13960 5632 13988
rect 5224 13948 5230 13960
rect 5626 13948 5632 13960
rect 5684 13948 5690 14000
rect 5718 13948 5724 14000
rect 5776 13988 5782 14000
rect 5905 13991 5963 13997
rect 5905 13988 5917 13991
rect 5776 13960 5917 13988
rect 5776 13948 5782 13960
rect 5905 13957 5917 13960
rect 5951 13988 5963 13991
rect 6748 13988 6776 14028
rect 7006 14016 7012 14028
rect 7064 14016 7070 14068
rect 7190 14056 7196 14068
rect 7151 14028 7196 14056
rect 7190 14016 7196 14028
rect 7248 14016 7254 14068
rect 8110 14056 8116 14068
rect 8071 14028 8116 14056
rect 8110 14016 8116 14028
rect 8168 14016 8174 14068
rect 9306 14016 9312 14068
rect 9364 14056 9370 14068
rect 9766 14056 9772 14068
rect 9364 14028 9674 14056
rect 9727 14028 9772 14056
rect 9364 14016 9370 14028
rect 6914 13988 6920 14000
rect 5951 13960 6776 13988
rect 6875 13960 6920 13988
rect 5951 13957 5963 13960
rect 5905 13951 5963 13957
rect 6914 13948 6920 13960
rect 6972 13948 6978 14000
rect 7098 13988 7104 14000
rect 7059 13960 7104 13988
rect 7098 13948 7104 13960
rect 7156 13948 7162 14000
rect 7469 13991 7527 13997
rect 7469 13957 7481 13991
rect 7515 13988 7527 13991
rect 9398 13988 9404 14000
rect 7515 13960 9404 13988
rect 7515 13957 7527 13960
rect 7469 13951 7527 13957
rect 9398 13948 9404 13960
rect 9456 13948 9462 14000
rect 9646 13988 9674 14028
rect 9766 14016 9772 14028
rect 9824 14016 9830 14068
rect 13630 14056 13636 14068
rect 10581 14028 13636 14056
rect 10226 13988 10232 14000
rect 9646 13960 10232 13988
rect 10226 13948 10232 13960
rect 10284 13948 10290 14000
rect 3384 13892 3740 13920
rect 3789 13923 3847 13929
rect 3384 13880 3390 13892
rect 3789 13889 3801 13923
rect 3835 13889 3847 13923
rect 3789 13883 3847 13889
rect 3053 13855 3111 13861
rect 3053 13852 3065 13855
rect 2424 13824 2544 13852
rect 2893 13824 3065 13852
rect 2516 13716 2544 13824
rect 3053 13821 3065 13824
rect 3099 13821 3111 13855
rect 3053 13815 3111 13821
rect 3804 13716 3832 13883
rect 3878 13880 3884 13932
rect 3936 13920 3942 13932
rect 4341 13923 4399 13929
rect 3936 13892 3981 13920
rect 3936 13880 3942 13892
rect 4341 13889 4353 13923
rect 4387 13920 4399 13923
rect 4522 13920 4528 13932
rect 4387 13892 4528 13920
rect 4387 13889 4399 13892
rect 4341 13883 4399 13889
rect 4522 13880 4528 13892
rect 4580 13880 4586 13932
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4706 13920 4712 13932
rect 4663 13892 4712 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 5074 13880 5080 13932
rect 5132 13920 5138 13932
rect 5994 13920 6000 13932
rect 5132 13892 5764 13920
rect 5955 13892 6000 13920
rect 5132 13880 5138 13892
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 4212 13824 4905 13852
rect 4212 13812 4218 13824
rect 4893 13821 4905 13824
rect 4939 13821 4951 13855
rect 5736 13852 5764 13892
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 6546 13920 6552 13932
rect 6507 13892 6552 13920
rect 6546 13880 6552 13892
rect 6604 13880 6610 13932
rect 6822 13880 6828 13932
rect 6880 13920 6886 13932
rect 7929 13923 7987 13929
rect 7929 13920 7941 13923
rect 6880 13892 7941 13920
rect 6880 13880 6886 13892
rect 7929 13889 7941 13892
rect 7975 13920 7987 13923
rect 9306 13920 9312 13932
rect 7975 13892 9312 13920
rect 7975 13889 7987 13892
rect 7929 13883 7987 13889
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 9585 13907 9643 13913
rect 9585 13873 9597 13907
rect 9631 13904 9643 13907
rect 9766 13904 9772 13932
rect 9631 13880 9772 13904
rect 9824 13920 9830 13932
rect 10581 13920 10609 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 13722 14016 13728 14068
rect 13780 14056 13786 14068
rect 13780 14028 13825 14056
rect 13780 14016 13786 14028
rect 13906 14016 13912 14068
rect 13964 14056 13970 14068
rect 14001 14059 14059 14065
rect 14001 14056 14013 14059
rect 13964 14028 14013 14056
rect 13964 14016 13970 14028
rect 14001 14025 14013 14028
rect 14047 14025 14059 14059
rect 14826 14056 14832 14068
rect 14787 14028 14832 14056
rect 14001 14019 14059 14025
rect 14826 14016 14832 14028
rect 14884 14016 14890 14068
rect 14918 14016 14924 14068
rect 14976 14056 14982 14068
rect 15654 14056 15660 14068
rect 14976 14028 15660 14056
rect 14976 14016 14982 14028
rect 12069 13991 12127 13997
rect 12069 13988 12081 13991
rect 9824 13892 10609 13920
rect 10704 13960 12081 13988
rect 9824 13880 9830 13892
rect 9631 13876 9812 13880
rect 9631 13873 9643 13876
rect 9585 13867 9643 13873
rect 7561 13855 7619 13861
rect 7561 13852 7573 13855
rect 5736 13824 7573 13852
rect 4893 13815 4951 13821
rect 7561 13821 7573 13824
rect 7607 13821 7619 13855
rect 7561 13815 7619 13821
rect 8018 13812 8024 13864
rect 8076 13852 8082 13864
rect 9398 13852 9404 13864
rect 8076 13824 9404 13852
rect 8076 13812 8082 13824
rect 9398 13812 9404 13824
rect 9456 13812 9462 13864
rect 4522 13744 4528 13796
rect 4580 13784 4586 13796
rect 5629 13787 5687 13793
rect 5629 13784 5641 13787
rect 4580 13756 5641 13784
rect 4580 13744 4586 13756
rect 5629 13753 5641 13756
rect 5675 13753 5687 13787
rect 5629 13747 5687 13753
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 10704 13784 10732 13960
rect 12069 13957 12081 13960
rect 12115 13957 12127 13991
rect 12342 13988 12348 14000
rect 12303 13960 12348 13988
rect 12069 13951 12127 13957
rect 12342 13948 12348 13960
rect 12400 13948 12406 14000
rect 12526 13988 12532 14000
rect 12487 13960 12532 13988
rect 12526 13948 12532 13960
rect 12584 13948 12590 14000
rect 12710 13988 12716 14000
rect 12671 13960 12716 13988
rect 12710 13948 12716 13960
rect 12768 13948 12774 14000
rect 12897 13991 12955 13997
rect 12897 13957 12909 13991
rect 12943 13988 12955 13991
rect 12943 13960 14964 13988
rect 12943 13957 12955 13960
rect 12897 13951 12955 13957
rect 12158 13880 12164 13932
rect 12216 13920 12222 13932
rect 13078 13920 13084 13932
rect 12216 13892 13084 13920
rect 12216 13880 12222 13892
rect 13078 13880 13084 13892
rect 13136 13880 13142 13932
rect 13170 13880 13176 13932
rect 13228 13920 13234 13932
rect 13541 13923 13599 13929
rect 13541 13920 13553 13923
rect 13228 13892 13553 13920
rect 13228 13880 13234 13892
rect 13541 13889 13553 13892
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 13630 13880 13636 13932
rect 13688 13920 13694 13932
rect 13817 13923 13875 13929
rect 13817 13920 13829 13923
rect 13688 13892 13829 13920
rect 13688 13880 13694 13892
rect 13817 13889 13829 13892
rect 13863 13889 13875 13923
rect 14277 13923 14335 13929
rect 14277 13920 14289 13923
rect 13817 13883 13875 13889
rect 13924 13892 14289 13920
rect 10778 13812 10784 13864
rect 10836 13852 10842 13864
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 10836 13824 11529 13852
rect 10836 13812 10842 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 11808 13824 12020 13852
rect 8628 13756 10732 13784
rect 8628 13744 8634 13756
rect 11146 13744 11152 13796
rect 11204 13784 11210 13796
rect 11808 13784 11836 13824
rect 11204 13756 11836 13784
rect 11992 13784 12020 13824
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 13265 13855 13323 13861
rect 13265 13852 13277 13855
rect 12124 13824 13277 13852
rect 12124 13812 12130 13824
rect 13265 13821 13277 13824
rect 13311 13852 13323 13855
rect 13924 13852 13952 13892
rect 14277 13889 14289 13892
rect 14323 13889 14335 13923
rect 14277 13883 14335 13889
rect 14553 13923 14611 13929
rect 14553 13889 14565 13923
rect 14599 13920 14611 13923
rect 14599 13892 14872 13920
rect 14599 13889 14611 13892
rect 14553 13883 14611 13889
rect 14642 13852 14648 13864
rect 13311 13824 13952 13852
rect 14108 13824 14648 13852
rect 13311 13821 13323 13824
rect 13265 13815 13323 13821
rect 13357 13787 13415 13793
rect 13357 13784 13369 13787
rect 11992 13756 13369 13784
rect 11204 13744 11210 13756
rect 13357 13753 13369 13756
rect 13403 13784 13415 13787
rect 13630 13784 13636 13796
rect 13403 13756 13636 13784
rect 13403 13753 13415 13756
rect 13357 13747 13415 13753
rect 13630 13744 13636 13756
rect 13688 13744 13694 13796
rect 14108 13793 14136 13824
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 14093 13787 14151 13793
rect 14093 13753 14105 13787
rect 14139 13753 14151 13787
rect 14366 13784 14372 13796
rect 14327 13756 14372 13784
rect 14093 13747 14151 13753
rect 14366 13744 14372 13756
rect 14424 13744 14430 13796
rect 14844 13784 14872 13892
rect 14936 13852 14964 13960
rect 15028 13929 15056 14028
rect 15654 14016 15660 14028
rect 15712 14016 15718 14068
rect 15749 14059 15807 14065
rect 15749 14025 15761 14059
rect 15795 14056 15807 14059
rect 19426 14056 19432 14068
rect 15795 14028 19432 14056
rect 15795 14025 15807 14028
rect 15749 14019 15807 14025
rect 19426 14016 19432 14028
rect 19484 14016 19490 14068
rect 15102 13948 15108 14000
rect 15160 13988 15166 14000
rect 16209 13991 16267 13997
rect 16209 13988 16221 13991
rect 15160 13960 16221 13988
rect 15160 13948 15166 13960
rect 16209 13957 16221 13960
rect 16255 13957 16267 13991
rect 16209 13951 16267 13957
rect 15013 13923 15071 13929
rect 15013 13889 15025 13923
rect 15059 13889 15071 13923
rect 15286 13920 15292 13932
rect 15247 13892 15292 13920
rect 15013 13883 15071 13889
rect 15286 13880 15292 13892
rect 15344 13880 15350 13932
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 15838 13920 15844 13932
rect 15436 13892 15481 13920
rect 15799 13892 15844 13920
rect 15436 13880 15442 13892
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 16114 13880 16120 13932
rect 16172 13920 16178 13932
rect 16485 13923 16543 13929
rect 16485 13920 16497 13923
rect 16172 13892 16497 13920
rect 16172 13880 16178 13892
rect 16485 13889 16497 13892
rect 16531 13889 16543 13923
rect 19058 13920 19064 13932
rect 16485 13883 16543 13889
rect 16868 13892 19064 13920
rect 15856 13852 15884 13880
rect 14936 13824 15884 13852
rect 16390 13812 16396 13864
rect 16448 13852 16454 13864
rect 16761 13855 16819 13861
rect 16761 13852 16773 13855
rect 16448 13824 16773 13852
rect 16448 13812 16454 13824
rect 16761 13821 16773 13824
rect 16807 13821 16819 13855
rect 16761 13815 16819 13821
rect 15565 13787 15623 13793
rect 14476 13756 14780 13784
rect 14844 13756 15516 13784
rect 4062 13716 4068 13728
rect 2516 13688 3832 13716
rect 4023 13688 4068 13716
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 5074 13676 5080 13728
rect 5132 13716 5138 13728
rect 5350 13716 5356 13728
rect 5132 13688 5356 13716
rect 5132 13676 5138 13688
rect 5350 13676 5356 13688
rect 5408 13676 5414 13728
rect 5534 13716 5540 13728
rect 5495 13688 5540 13716
rect 5534 13676 5540 13688
rect 5592 13676 5598 13728
rect 5902 13676 5908 13728
rect 5960 13716 5966 13728
rect 6638 13716 6644 13728
rect 5960 13688 6644 13716
rect 5960 13676 5966 13688
rect 6638 13676 6644 13688
rect 6696 13676 6702 13728
rect 6822 13676 6828 13728
rect 6880 13716 6886 13728
rect 7837 13719 7895 13725
rect 7837 13716 7849 13719
rect 6880 13688 7849 13716
rect 6880 13676 6886 13688
rect 7837 13685 7849 13688
rect 7883 13716 7895 13719
rect 11330 13716 11336 13728
rect 7883 13688 11336 13716
rect 7883 13685 7895 13688
rect 7837 13679 7895 13685
rect 11330 13676 11336 13688
rect 11388 13676 11394 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 11701 13719 11759 13725
rect 11701 13716 11713 13719
rect 11664 13688 11713 13716
rect 11664 13676 11670 13688
rect 11701 13685 11713 13688
rect 11747 13685 11759 13719
rect 11882 13716 11888 13728
rect 11843 13688 11888 13716
rect 11701 13679 11759 13685
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 13170 13676 13176 13728
rect 13228 13716 13234 13728
rect 14476 13716 14504 13756
rect 13228 13688 14504 13716
rect 13228 13676 13234 13688
rect 14550 13676 14556 13728
rect 14608 13716 14614 13728
rect 14645 13719 14703 13725
rect 14645 13716 14657 13719
rect 14608 13688 14657 13716
rect 14608 13676 14614 13688
rect 14645 13685 14657 13688
rect 14691 13685 14703 13719
rect 14752 13716 14780 13756
rect 14918 13716 14924 13728
rect 14752 13688 14924 13716
rect 14645 13679 14703 13685
rect 14918 13676 14924 13688
rect 14976 13676 14982 13728
rect 15102 13716 15108 13728
rect 15063 13688 15108 13716
rect 15102 13676 15108 13688
rect 15160 13676 15166 13728
rect 15488 13716 15516 13756
rect 15565 13753 15577 13787
rect 15611 13784 15623 13787
rect 16868 13784 16896 13892
rect 19058 13880 19064 13892
rect 19116 13880 19122 13932
rect 17037 13855 17095 13861
rect 17037 13821 17049 13855
rect 17083 13852 17095 13855
rect 17126 13852 17132 13864
rect 17083 13824 17132 13852
rect 17083 13821 17095 13824
rect 17037 13815 17095 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17678 13852 17684 13864
rect 17639 13824 17684 13852
rect 17678 13812 17684 13824
rect 17736 13812 17742 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13852 18015 13855
rect 18598 13852 18604 13864
rect 18003 13824 18604 13852
rect 18003 13821 18015 13824
rect 17957 13815 18015 13821
rect 18598 13812 18604 13824
rect 18656 13812 18662 13864
rect 15611 13756 16896 13784
rect 15611 13753 15623 13756
rect 15565 13747 15623 13753
rect 17034 13716 17040 13728
rect 15488 13688 17040 13716
rect 17034 13676 17040 13688
rect 17092 13676 17098 13728
rect 1104 13626 18860 13648
rect 1104 13574 3174 13626
rect 3226 13574 3238 13626
rect 3290 13574 3302 13626
rect 3354 13574 3366 13626
rect 3418 13574 3430 13626
rect 3482 13574 7622 13626
rect 7674 13574 7686 13626
rect 7738 13574 7750 13626
rect 7802 13574 7814 13626
rect 7866 13574 7878 13626
rect 7930 13574 12070 13626
rect 12122 13574 12134 13626
rect 12186 13574 12198 13626
rect 12250 13574 12262 13626
rect 12314 13574 12326 13626
rect 12378 13574 16518 13626
rect 16570 13574 16582 13626
rect 16634 13574 16646 13626
rect 16698 13574 16710 13626
rect 16762 13574 16774 13626
rect 16826 13574 18860 13626
rect 1104 13552 18860 13574
rect 842 13472 848 13524
rect 900 13512 906 13524
rect 900 13484 4200 13512
rect 900 13472 906 13484
rect 1210 13404 1216 13456
rect 1268 13444 1274 13456
rect 3145 13447 3203 13453
rect 3145 13444 3157 13447
rect 1268 13416 3157 13444
rect 1268 13404 1274 13416
rect 3145 13413 3157 13416
rect 3191 13413 3203 13447
rect 3145 13407 3203 13413
rect 3789 13447 3847 13453
rect 3789 13413 3801 13447
rect 3835 13413 3847 13447
rect 3789 13407 3847 13413
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13376 2283 13379
rect 2498 13376 2504 13388
rect 2271 13348 2504 13376
rect 2271 13345 2283 13348
rect 2225 13339 2283 13345
rect 2498 13336 2504 13348
rect 2556 13336 2562 13388
rect 3804 13376 3832 13407
rect 2976 13348 3832 13376
rect 4172 13376 4200 13484
rect 4246 13472 4252 13524
rect 4304 13512 4310 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4304 13484 4629 13512
rect 4304 13472 4310 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 4617 13475 4675 13481
rect 5350 13472 5356 13524
rect 5408 13512 5414 13524
rect 6273 13515 6331 13521
rect 6273 13512 6285 13515
rect 5408 13484 6285 13512
rect 5408 13472 5414 13484
rect 6273 13481 6285 13484
rect 6319 13481 6331 13515
rect 6638 13512 6644 13524
rect 6599 13484 6644 13512
rect 6273 13475 6331 13481
rect 6638 13472 6644 13484
rect 6696 13512 6702 13524
rect 7282 13512 7288 13524
rect 6696 13484 7288 13512
rect 6696 13472 6702 13484
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 8018 13512 8024 13524
rect 7979 13484 8024 13512
rect 8018 13472 8024 13484
rect 8076 13472 8082 13524
rect 8294 13512 8300 13524
rect 8255 13484 8300 13512
rect 8294 13472 8300 13484
rect 8352 13472 8358 13524
rect 8570 13512 8576 13524
rect 8531 13484 8576 13512
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 9030 13512 9036 13524
rect 8991 13484 9036 13512
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10870 13512 10876 13524
rect 10468 13484 10876 13512
rect 10468 13472 10474 13484
rect 10870 13472 10876 13484
rect 10928 13472 10934 13524
rect 11422 13512 11428 13524
rect 11383 13484 11428 13512
rect 11422 13472 11428 13484
rect 11480 13472 11486 13524
rect 11606 13472 11612 13524
rect 11664 13512 11670 13524
rect 12802 13512 12808 13524
rect 11664 13484 11836 13512
rect 12763 13484 12808 13512
rect 11664 13472 11670 13484
rect 4798 13404 4804 13456
rect 4856 13444 4862 13456
rect 11808 13453 11836 13484
rect 12802 13472 12808 13484
rect 12860 13472 12866 13524
rect 13538 13472 13544 13524
rect 13596 13512 13602 13524
rect 15654 13512 15660 13524
rect 13596 13484 15660 13512
rect 13596 13472 13602 13484
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 16114 13512 16120 13524
rect 16075 13484 16120 13512
rect 16114 13472 16120 13484
rect 16172 13472 16178 13524
rect 16206 13472 16212 13524
rect 16264 13512 16270 13524
rect 16264 13484 17724 13512
rect 16264 13472 16270 13484
rect 11793 13447 11851 13453
rect 4856 13416 11652 13444
rect 4856 13404 4862 13416
rect 5534 13376 5540 13388
rect 4172 13348 5540 13376
rect 1949 13311 2007 13317
rect 1949 13277 1961 13311
rect 1995 13308 2007 13311
rect 2130 13308 2136 13320
rect 1995 13280 2136 13308
rect 1995 13277 2007 13280
rect 1949 13271 2007 13277
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2590 13308 2596 13320
rect 2551 13280 2596 13308
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 2976 13317 3004 13348
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 3326 13308 3332 13320
rect 3287 13280 3332 13308
rect 2961 13271 3019 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 3418 13268 3424 13320
rect 3476 13308 3482 13320
rect 3476 13280 3521 13308
rect 3476 13268 3482 13280
rect 3878 13268 3884 13320
rect 3936 13308 3942 13320
rect 3973 13311 4031 13317
rect 3973 13308 3985 13311
rect 3936 13280 3985 13308
rect 3936 13268 3942 13280
rect 3973 13277 3985 13280
rect 4019 13277 4031 13311
rect 3973 13271 4031 13277
rect 4062 13268 4068 13320
rect 4120 13308 4126 13320
rect 4356 13317 4384 13348
rect 5534 13336 5540 13348
rect 5592 13336 5598 13388
rect 5626 13336 5632 13388
rect 5684 13376 5690 13388
rect 5721 13379 5779 13385
rect 5721 13376 5733 13379
rect 5684 13348 5733 13376
rect 5684 13336 5690 13348
rect 5721 13345 5733 13348
rect 5767 13376 5779 13379
rect 6730 13376 6736 13388
rect 5767 13348 6736 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 7190 13376 7196 13388
rect 7151 13348 7196 13376
rect 7190 13336 7196 13348
rect 7248 13336 7254 13388
rect 8294 13336 8300 13388
rect 8352 13376 8358 13388
rect 8757 13379 8815 13385
rect 8757 13376 8769 13379
rect 8352 13348 8769 13376
rect 8352 13336 8358 13348
rect 8757 13345 8769 13348
rect 8803 13376 8815 13379
rect 11514 13376 11520 13388
rect 8803 13348 11520 13376
rect 8803 13345 8815 13348
rect 8757 13339 8815 13345
rect 11514 13336 11520 13348
rect 11572 13336 11578 13388
rect 11624 13376 11652 13416
rect 11793 13413 11805 13447
rect 11839 13444 11851 13447
rect 12066 13444 12072 13456
rect 11839 13416 12072 13444
rect 11839 13413 11851 13416
rect 11793 13407 11851 13413
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 12253 13447 12311 13453
rect 12253 13413 12265 13447
rect 12299 13444 12311 13447
rect 13078 13444 13084 13456
rect 12299 13416 13084 13444
rect 12299 13413 12311 13416
rect 12253 13407 12311 13413
rect 13078 13404 13084 13416
rect 13136 13404 13142 13456
rect 13814 13404 13820 13456
rect 13872 13444 13878 13456
rect 14918 13444 14924 13456
rect 13872 13416 14924 13444
rect 13872 13404 13878 13416
rect 14918 13404 14924 13416
rect 14976 13404 14982 13456
rect 15013 13447 15071 13453
rect 15013 13413 15025 13447
rect 15059 13444 15071 13447
rect 15562 13444 15568 13456
rect 15059 13416 15568 13444
rect 15059 13413 15071 13416
rect 15013 13407 15071 13413
rect 15562 13404 15568 13416
rect 15620 13404 15626 13456
rect 12342 13376 12348 13388
rect 11624 13348 12348 13376
rect 12342 13336 12348 13348
rect 12400 13336 12406 13388
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 12986 13376 12992 13388
rect 12584 13348 12992 13376
rect 12584 13336 12590 13348
rect 12986 13336 12992 13348
rect 13044 13336 13050 13388
rect 14274 13336 14280 13388
rect 14332 13376 14338 13388
rect 15194 13376 15200 13388
rect 14332 13348 15200 13376
rect 14332 13336 14338 13348
rect 4341 13311 4399 13317
rect 4120 13280 4165 13308
rect 4120 13268 4126 13280
rect 4341 13277 4353 13311
rect 4387 13277 4399 13311
rect 4341 13271 4399 13277
rect 4614 13268 4620 13320
rect 4672 13308 4678 13320
rect 4798 13308 4804 13320
rect 4672 13280 4804 13308
rect 4672 13268 4678 13280
rect 4798 13268 4804 13280
rect 4856 13268 4862 13320
rect 4890 13268 4896 13320
rect 4948 13308 4954 13320
rect 4948 13280 4993 13308
rect 4948 13268 4954 13280
rect 5074 13268 5080 13320
rect 5132 13308 5138 13320
rect 5169 13311 5227 13317
rect 5169 13308 5181 13311
rect 5132 13280 5181 13308
rect 5132 13268 5138 13280
rect 5169 13277 5181 13280
rect 5215 13277 5227 13311
rect 5169 13271 5227 13277
rect 5258 13268 5264 13320
rect 5316 13308 5322 13320
rect 5353 13311 5411 13317
rect 5353 13308 5365 13311
rect 5316 13280 5365 13308
rect 5316 13268 5322 13280
rect 5353 13277 5365 13280
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 10226 13308 10232 13320
rect 5868 13280 10232 13308
rect 5868 13268 5874 13280
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 11054 13268 11060 13320
rect 11112 13308 11118 13320
rect 11885 13311 11943 13317
rect 11885 13308 11897 13311
rect 11112 13280 11897 13308
rect 11112 13268 11118 13280
rect 11885 13277 11897 13280
rect 11931 13277 11943 13311
rect 11885 13271 11943 13277
rect 12066 13268 12072 13320
rect 12124 13308 12130 13320
rect 12434 13308 12440 13320
rect 12124 13280 12440 13308
rect 12124 13268 12130 13280
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12713 13311 12771 13317
rect 12713 13277 12725 13311
rect 12759 13308 12771 13311
rect 12894 13308 12900 13320
rect 12759 13280 12900 13308
rect 12759 13277 12771 13280
rect 12713 13271 12771 13277
rect 12894 13268 12900 13280
rect 12952 13308 12958 13320
rect 12952 13304 13124 13308
rect 13165 13307 13223 13313
rect 13165 13304 13177 13307
rect 12952 13280 13177 13304
rect 12952 13268 12958 13280
rect 13096 13276 13177 13280
rect 13165 13273 13177 13276
rect 13211 13273 13223 13307
rect 13165 13267 13223 13273
rect 13280 13304 13400 13308
rect 13457 13307 13515 13313
rect 13457 13304 13469 13307
rect 13280 13280 13469 13304
rect 1302 13200 1308 13252
rect 1360 13240 1366 13252
rect 1360 13212 3648 13240
rect 1360 13200 1366 13212
rect 2406 13172 2412 13184
rect 2367 13144 2412 13172
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3620 13181 3648 13212
rect 3786 13200 3792 13252
rect 3844 13240 3850 13252
rect 6457 13243 6515 13249
rect 6457 13240 6469 13243
rect 3844 13212 6469 13240
rect 3844 13200 3850 13212
rect 6457 13209 6469 13212
rect 6503 13209 6515 13243
rect 6457 13203 6515 13209
rect 6546 13200 6552 13252
rect 6604 13240 6610 13252
rect 7009 13243 7067 13249
rect 7009 13240 7021 13243
rect 6604 13212 7021 13240
rect 6604 13200 6610 13212
rect 7009 13209 7021 13212
rect 7055 13209 7067 13243
rect 7009 13203 7067 13209
rect 7282 13200 7288 13252
rect 7340 13240 7346 13252
rect 10686 13240 10692 13252
rect 7340 13212 10692 13240
rect 7340 13200 7346 13212
rect 10686 13200 10692 13212
rect 10744 13200 10750 13252
rect 10873 13243 10931 13249
rect 10873 13209 10885 13243
rect 10919 13240 10931 13243
rect 10962 13240 10968 13252
rect 10919 13212 10968 13240
rect 10919 13209 10931 13212
rect 10873 13203 10931 13209
rect 10962 13200 10968 13212
rect 11020 13200 11026 13252
rect 11146 13240 11152 13252
rect 11107 13212 11152 13240
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 12526 13240 12532 13252
rect 11296 13212 12204 13240
rect 12487 13212 12532 13240
rect 11296 13200 11302 13212
rect 3605 13175 3663 13181
rect 2832 13144 2877 13172
rect 2832 13132 2838 13144
rect 3605 13141 3617 13175
rect 3651 13141 3663 13175
rect 3605 13135 3663 13141
rect 3694 13132 3700 13184
rect 3752 13172 3758 13184
rect 4062 13172 4068 13184
rect 3752 13144 4068 13172
rect 3752 13132 3758 13144
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 4246 13172 4252 13184
rect 4207 13144 4252 13172
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 4430 13132 4436 13184
rect 4488 13172 4494 13184
rect 4525 13175 4583 13181
rect 4525 13172 4537 13175
rect 4488 13144 4537 13172
rect 4488 13132 4494 13144
rect 4525 13141 4537 13144
rect 4571 13141 4583 13175
rect 4525 13135 4583 13141
rect 5077 13175 5135 13181
rect 5077 13141 5089 13175
rect 5123 13172 5135 13175
rect 5258 13172 5264 13184
rect 5123 13144 5264 13172
rect 5123 13141 5135 13144
rect 5077 13135 5135 13141
rect 5258 13132 5264 13144
rect 5316 13132 5322 13184
rect 5902 13172 5908 13184
rect 5863 13144 5908 13172
rect 5902 13132 5908 13144
rect 5960 13132 5966 13184
rect 6178 13172 6184 13184
rect 6139 13144 6184 13172
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 6914 13172 6920 13184
rect 6875 13144 6920 13172
rect 6914 13132 6920 13144
rect 6972 13132 6978 13184
rect 7374 13172 7380 13184
rect 7335 13144 7380 13172
rect 7374 13132 7380 13144
rect 7432 13132 7438 13184
rect 7466 13132 7472 13184
rect 7524 13172 7530 13184
rect 7561 13175 7619 13181
rect 7561 13172 7573 13175
rect 7524 13144 7573 13172
rect 7524 13132 7530 13144
rect 7561 13141 7573 13144
rect 7607 13141 7619 13175
rect 7742 13172 7748 13184
rect 7703 13144 7748 13172
rect 7561 13135 7619 13141
rect 7742 13132 7748 13144
rect 7800 13132 7806 13184
rect 8018 13132 8024 13184
rect 8076 13172 8082 13184
rect 8113 13175 8171 13181
rect 8113 13172 8125 13175
rect 8076 13144 8125 13172
rect 8076 13132 8082 13144
rect 8113 13141 8125 13144
rect 8159 13141 8171 13175
rect 10594 13172 10600 13184
rect 10555 13144 10600 13172
rect 8113 13135 8171 13141
rect 10594 13132 10600 13144
rect 10652 13132 10658 13184
rect 12066 13172 12072 13184
rect 12027 13144 12072 13172
rect 12066 13132 12072 13144
rect 12124 13132 12130 13184
rect 12176 13172 12204 13212
rect 12526 13200 12532 13212
rect 12584 13200 12590 13252
rect 13280 13172 13308 13280
rect 13372 13276 13469 13280
rect 13457 13273 13469 13276
rect 13503 13304 13515 13307
rect 13503 13276 13584 13304
rect 13503 13273 13515 13276
rect 13457 13267 13515 13273
rect 13556 13240 13584 13276
rect 13630 13268 13636 13320
rect 13688 13308 13694 13320
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 13688 13280 13737 13308
rect 13688 13268 13694 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 14182 13268 14188 13320
rect 14240 13308 14246 13320
rect 14568 13317 14596 13348
rect 15194 13336 15200 13348
rect 15252 13336 15258 13388
rect 15289 13379 15347 13385
rect 15289 13345 15301 13379
rect 15335 13376 15347 13379
rect 16850 13376 16856 13388
rect 15335 13348 16856 13376
rect 15335 13345 15347 13348
rect 15289 13339 15347 13345
rect 16850 13336 16856 13348
rect 16908 13336 16914 13388
rect 17696 13385 17724 13484
rect 17681 13379 17739 13385
rect 17681 13345 17693 13379
rect 17727 13376 17739 13379
rect 17862 13376 17868 13388
rect 17727 13348 17868 13376
rect 17727 13345 17739 13348
rect 17681 13339 17739 13345
rect 17862 13336 17868 13348
rect 17920 13336 17926 13388
rect 14461 13311 14519 13317
rect 14461 13308 14473 13311
rect 14240 13280 14473 13308
rect 14240 13268 14246 13280
rect 14461 13277 14473 13280
rect 14507 13277 14519 13311
rect 14461 13271 14519 13277
rect 14553 13311 14611 13317
rect 14553 13277 14565 13311
rect 14599 13277 14611 13311
rect 14553 13271 14611 13277
rect 14829 13311 14887 13317
rect 14829 13277 14841 13311
rect 14875 13308 14887 13311
rect 15378 13308 15384 13320
rect 14875 13280 15384 13308
rect 14875 13277 14887 13280
rect 14829 13271 14887 13277
rect 15378 13268 15384 13280
rect 15436 13268 15442 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 15528 13280 17509 13308
rect 15528 13268 15534 13280
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18046 13308 18052 13320
rect 18003 13280 18052 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 14093 13243 14151 13249
rect 14093 13240 14105 13243
rect 13556 13212 14105 13240
rect 14093 13209 14105 13212
rect 14139 13240 14151 13243
rect 14918 13240 14924 13252
rect 14139 13212 14924 13240
rect 14139 13209 14151 13212
rect 14093 13203 14151 13209
rect 14918 13200 14924 13212
rect 14976 13200 14982 13252
rect 16390 13200 16396 13252
rect 16448 13240 16454 13252
rect 17405 13243 17463 13249
rect 17405 13240 17417 13243
rect 16448 13212 17417 13240
rect 16448 13200 16454 13212
rect 17405 13209 17417 13212
rect 17451 13209 17463 13243
rect 17512 13240 17540 13271
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 17770 13240 17776 13252
rect 17512 13212 17776 13240
rect 17405 13203 17463 13209
rect 17770 13200 17776 13212
rect 17828 13200 17834 13252
rect 12176 13144 13308 13172
rect 13357 13175 13415 13181
rect 13357 13141 13369 13175
rect 13403 13172 13415 13175
rect 13446 13172 13452 13184
rect 13403 13144 13452 13172
rect 13403 13141 13415 13144
rect 13357 13135 13415 13141
rect 13446 13132 13452 13144
rect 13504 13132 13510 13184
rect 13630 13172 13636 13184
rect 13591 13144 13636 13172
rect 13630 13132 13636 13144
rect 13688 13132 13694 13184
rect 13909 13175 13967 13181
rect 13909 13141 13921 13175
rect 13955 13172 13967 13175
rect 13998 13172 14004 13184
rect 13955 13144 14004 13172
rect 13955 13141 13967 13144
rect 13909 13135 13967 13141
rect 13998 13132 14004 13144
rect 14056 13132 14062 13184
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14277 13175 14335 13181
rect 14277 13172 14289 13175
rect 14240 13144 14289 13172
rect 14240 13132 14246 13144
rect 14277 13141 14289 13144
rect 14323 13141 14335 13175
rect 14277 13135 14335 13141
rect 14737 13175 14795 13181
rect 14737 13141 14749 13175
rect 14783 13172 14795 13175
rect 15378 13172 15384 13184
rect 14783 13144 15384 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 15378 13132 15384 13144
rect 15436 13132 15442 13184
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 15746 13132 15752 13184
rect 15804 13172 15810 13184
rect 19150 13172 19156 13184
rect 15804 13144 19156 13172
rect 15804 13132 15810 13144
rect 19150 13132 19156 13144
rect 19208 13132 19214 13184
rect 1104 13082 18860 13104
rect 1104 13030 5398 13082
rect 5450 13030 5462 13082
rect 5514 13030 5526 13082
rect 5578 13030 5590 13082
rect 5642 13030 5654 13082
rect 5706 13030 9846 13082
rect 9898 13030 9910 13082
rect 9962 13030 9974 13082
rect 10026 13030 10038 13082
rect 10090 13030 10102 13082
rect 10154 13030 14294 13082
rect 14346 13030 14358 13082
rect 14410 13030 14422 13082
rect 14474 13030 14486 13082
rect 14538 13030 14550 13082
rect 14602 13030 18860 13082
rect 1104 13008 18860 13030
rect 2314 12928 2320 12980
rect 2372 12968 2378 12980
rect 4338 12968 4344 12980
rect 2372 12940 4200 12968
rect 4299 12940 4344 12968
rect 2372 12928 2378 12940
rect 1762 12860 1768 12912
rect 1820 12900 1826 12912
rect 4065 12903 4123 12909
rect 4065 12900 4077 12903
rect 1820 12872 4077 12900
rect 1820 12860 1826 12872
rect 4065 12869 4077 12872
rect 4111 12869 4123 12903
rect 4172 12900 4200 12940
rect 4338 12928 4344 12940
rect 4396 12928 4402 12980
rect 4801 12971 4859 12977
rect 4801 12937 4813 12971
rect 4847 12937 4859 12971
rect 5810 12968 5816 12980
rect 5771 12940 5816 12968
rect 4801 12931 4859 12937
rect 4816 12900 4844 12931
rect 5810 12928 5816 12940
rect 5868 12928 5874 12980
rect 6546 12928 6552 12980
rect 6604 12968 6610 12980
rect 6914 12968 6920 12980
rect 6604 12940 6920 12968
rect 6604 12928 6610 12940
rect 6914 12928 6920 12940
rect 6972 12968 6978 12980
rect 9125 12971 9183 12977
rect 9125 12968 9137 12971
rect 6972 12940 9137 12968
rect 6972 12928 6978 12940
rect 9125 12937 9137 12940
rect 9171 12937 9183 12971
rect 9490 12968 9496 12980
rect 9451 12940 9496 12968
rect 9125 12931 9183 12937
rect 9490 12928 9496 12940
rect 9548 12928 9554 12980
rect 10045 12971 10103 12977
rect 10045 12937 10057 12971
rect 10091 12968 10103 12971
rect 10318 12968 10324 12980
rect 10091 12940 10324 12968
rect 10091 12937 10103 12940
rect 10045 12931 10103 12937
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10410 12928 10416 12980
rect 10468 12968 10474 12980
rect 10597 12971 10655 12977
rect 10468 12940 10513 12968
rect 10468 12928 10474 12940
rect 10597 12937 10609 12971
rect 10643 12968 10655 12971
rect 10686 12968 10692 12980
rect 10643 12940 10692 12968
rect 10643 12937 10655 12940
rect 10597 12931 10655 12937
rect 10686 12928 10692 12940
rect 10744 12928 10750 12980
rect 11422 12928 11428 12980
rect 11480 12968 11486 12980
rect 11517 12971 11575 12977
rect 11517 12968 11529 12971
rect 11480 12940 11529 12968
rect 11480 12928 11486 12940
rect 11517 12937 11529 12940
rect 11563 12937 11575 12971
rect 11517 12931 11575 12937
rect 11977 12971 12035 12977
rect 11977 12937 11989 12971
rect 12023 12968 12035 12971
rect 12710 12968 12716 12980
rect 12023 12940 12388 12968
rect 12023 12937 12035 12940
rect 11977 12931 12035 12937
rect 6086 12900 6092 12912
rect 4172 12872 4844 12900
rect 4899 12872 6092 12900
rect 4065 12863 4123 12869
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3050 12832 3056 12844
rect 2915 12804 3056 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3050 12792 3056 12804
rect 3108 12792 3114 12844
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 3694 12832 3700 12844
rect 3559 12804 3700 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 3694 12792 3700 12804
rect 3752 12792 3758 12844
rect 3789 12835 3847 12841
rect 3789 12801 3801 12835
rect 3835 12832 3847 12835
rect 3835 12816 4016 12832
rect 3835 12804 4108 12816
rect 3835 12801 3847 12804
rect 3789 12795 3847 12801
rect 3988 12788 4108 12804
rect 4246 12792 4252 12844
rect 4304 12832 4310 12844
rect 4899 12832 4927 12872
rect 6086 12860 6092 12872
rect 6144 12860 6150 12912
rect 7282 12860 7288 12912
rect 7340 12900 7346 12912
rect 7653 12903 7711 12909
rect 7653 12900 7665 12903
rect 7340 12872 7665 12900
rect 7340 12860 7346 12872
rect 7653 12869 7665 12872
rect 7699 12869 7711 12903
rect 8110 12900 8116 12912
rect 8071 12872 8116 12900
rect 7653 12863 7711 12869
rect 8110 12860 8116 12872
rect 8168 12860 8174 12912
rect 8294 12860 8300 12912
rect 8352 12900 8358 12912
rect 8352 12872 8397 12900
rect 8352 12860 8358 12872
rect 8754 12860 8760 12912
rect 8812 12900 8818 12912
rect 9030 12900 9036 12912
rect 8812 12872 8857 12900
rect 8991 12872 9036 12900
rect 8812 12860 8818 12872
rect 9030 12860 9036 12872
rect 9088 12860 9094 12912
rect 9582 12860 9588 12912
rect 9640 12900 9646 12912
rect 10781 12903 10839 12909
rect 10781 12900 10793 12903
rect 9640 12872 10793 12900
rect 9640 12860 9646 12872
rect 10781 12869 10793 12872
rect 10827 12900 10839 12903
rect 12158 12900 12164 12912
rect 10827 12872 12164 12900
rect 10827 12869 10839 12872
rect 10781 12863 10839 12869
rect 12158 12860 12164 12872
rect 12216 12860 12222 12912
rect 12360 12900 12388 12940
rect 12544 12940 12716 12968
rect 12544 12900 12572 12940
rect 12710 12928 12716 12940
rect 12768 12928 12774 12980
rect 13170 12968 13176 12980
rect 13131 12940 13176 12968
rect 13170 12928 13176 12940
rect 13228 12928 13234 12980
rect 13814 12928 13820 12980
rect 13872 12968 13878 12980
rect 13872 12940 13917 12968
rect 13872 12928 13878 12940
rect 14090 12928 14096 12980
rect 14148 12968 14154 12980
rect 15565 12971 15623 12977
rect 14148 12940 14320 12968
rect 14148 12928 14154 12940
rect 12360 12872 12572 12900
rect 4304 12804 4927 12832
rect 4304 12792 4310 12804
rect 4982 12792 4988 12844
rect 5040 12832 5046 12844
rect 5040 12804 5085 12832
rect 5040 12792 5046 12804
rect 5166 12792 5172 12844
rect 5224 12832 5230 12844
rect 5350 12832 5356 12844
rect 5224 12804 5356 12832
rect 5224 12792 5230 12804
rect 5350 12792 5356 12804
rect 5408 12792 5414 12844
rect 5629 12835 5687 12841
rect 5629 12801 5641 12835
rect 5675 12801 5687 12835
rect 5629 12795 5687 12801
rect 5905 12835 5963 12841
rect 5905 12801 5917 12835
rect 5951 12832 5963 12835
rect 6270 12832 6276 12844
rect 5951 12804 6276 12832
rect 5951 12801 5963 12804
rect 5905 12795 5963 12801
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 1949 12767 2007 12773
rect 1949 12764 1961 12767
rect 1544 12736 1961 12764
rect 1544 12724 1550 12736
rect 1949 12733 1961 12736
rect 1995 12733 2007 12767
rect 1949 12727 2007 12733
rect 2225 12767 2283 12773
rect 2225 12733 2237 12767
rect 2271 12764 2283 12767
rect 2774 12764 2780 12776
rect 2271 12736 2780 12764
rect 2271 12733 2283 12736
rect 2225 12727 2283 12733
rect 2774 12724 2780 12736
rect 2832 12724 2838 12776
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3145 12767 3203 12773
rect 3145 12764 3157 12767
rect 3016 12736 3157 12764
rect 3016 12724 3022 12736
rect 3145 12733 3157 12736
rect 3191 12764 3203 12767
rect 3234 12764 3240 12776
rect 3191 12736 3240 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3234 12724 3240 12736
rect 3292 12724 3298 12776
rect 3602 12696 3608 12708
rect 3563 12668 3608 12696
rect 3602 12656 3608 12668
rect 3660 12656 3666 12708
rect 4080 12696 4108 12788
rect 4080 12668 4292 12696
rect 2958 12588 2964 12640
rect 3016 12628 3022 12640
rect 3329 12631 3387 12637
rect 3329 12628 3341 12631
rect 3016 12600 3341 12628
rect 3016 12588 3022 12600
rect 3329 12597 3341 12600
rect 3375 12597 3387 12631
rect 3329 12591 3387 12597
rect 3973 12631 4031 12637
rect 3973 12597 3985 12631
rect 4019 12628 4031 12631
rect 4062 12628 4068 12640
rect 4019 12600 4068 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4062 12588 4068 12600
rect 4120 12588 4126 12640
rect 4264 12628 4292 12668
rect 4338 12656 4344 12708
rect 4396 12696 4402 12708
rect 4709 12699 4767 12705
rect 4709 12696 4721 12699
rect 4396 12668 4721 12696
rect 4396 12656 4402 12668
rect 4709 12665 4721 12668
rect 4755 12696 4767 12699
rect 5000 12696 5028 12792
rect 5261 12767 5319 12773
rect 5261 12764 5273 12767
rect 5184 12736 5273 12764
rect 5184 12708 5212 12736
rect 5261 12733 5273 12736
rect 5307 12733 5319 12767
rect 5644 12764 5672 12795
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 6730 12792 6736 12844
rect 6788 12832 6794 12844
rect 7837 12835 7895 12841
rect 7837 12832 7849 12835
rect 6788 12804 7849 12832
rect 6788 12792 6794 12804
rect 7837 12801 7849 12804
rect 7883 12801 7895 12835
rect 7837 12795 7895 12801
rect 8386 12792 8392 12844
rect 8444 12832 8450 12844
rect 8573 12835 8631 12841
rect 8573 12832 8585 12835
rect 8444 12804 8585 12832
rect 8444 12792 8450 12804
rect 8573 12801 8585 12804
rect 8619 12801 8631 12835
rect 8573 12795 8631 12801
rect 6454 12764 6460 12776
rect 5644 12736 6460 12764
rect 5261 12727 5319 12733
rect 6454 12724 6460 12736
rect 6512 12764 6518 12776
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6512 12736 6653 12764
rect 6512 12724 6518 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 7190 12764 7196 12776
rect 7151 12736 7196 12764
rect 6641 12727 6699 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 7561 12767 7619 12773
rect 7561 12733 7573 12767
rect 7607 12764 7619 12767
rect 8110 12764 8116 12776
rect 7607 12736 8116 12764
rect 7607 12733 7619 12736
rect 7561 12727 7619 12733
rect 8110 12724 8116 12736
rect 8168 12724 8174 12776
rect 8588 12764 8616 12795
rect 8846 12792 8852 12844
rect 8904 12832 8910 12844
rect 9309 12835 9367 12841
rect 9309 12832 9321 12835
rect 8904 12804 9321 12832
rect 8904 12792 8910 12804
rect 9309 12801 9321 12804
rect 9355 12832 9367 12835
rect 9398 12832 9404 12844
rect 9355 12804 9404 12832
rect 9355 12801 9367 12804
rect 9309 12795 9367 12801
rect 9398 12792 9404 12804
rect 9456 12792 9462 12844
rect 10686 12832 10692 12844
rect 9646 12804 10692 12832
rect 9646 12764 9674 12804
rect 10686 12792 10692 12804
rect 10744 12792 10750 12844
rect 11974 12832 11980 12844
rect 11256 12804 11980 12832
rect 8588 12736 9674 12764
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10594 12764 10600 12776
rect 10008 12736 10600 12764
rect 10008 12724 10014 12736
rect 10594 12724 10600 12736
rect 10652 12764 10658 12776
rect 11057 12767 11115 12773
rect 11057 12764 11069 12767
rect 10652 12736 11069 12764
rect 10652 12724 10658 12736
rect 11057 12733 11069 12736
rect 11103 12733 11115 12767
rect 11057 12727 11115 12733
rect 4755 12668 5028 12696
rect 4755 12665 4767 12668
rect 4709 12659 4767 12665
rect 5166 12656 5172 12708
rect 5224 12656 5230 12708
rect 5537 12699 5595 12705
rect 5537 12665 5549 12699
rect 5583 12696 5595 12699
rect 6270 12696 6276 12708
rect 5583 12668 6276 12696
rect 5583 12665 5595 12668
rect 5537 12659 5595 12665
rect 6270 12656 6276 12668
rect 6328 12656 6334 12708
rect 6549 12699 6607 12705
rect 6549 12665 6561 12699
rect 6595 12696 6607 12699
rect 6822 12696 6828 12708
rect 6595 12668 6828 12696
rect 6595 12665 6607 12668
rect 6549 12659 6607 12665
rect 6822 12656 6828 12668
rect 6880 12656 6886 12708
rect 6914 12656 6920 12708
rect 6972 12696 6978 12708
rect 10137 12699 10195 12705
rect 10137 12696 10149 12699
rect 6972 12668 7236 12696
rect 6972 12656 6978 12668
rect 5902 12628 5908 12640
rect 4264 12600 5908 12628
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 6086 12628 6092 12640
rect 6047 12600 6092 12628
rect 6086 12588 6092 12600
rect 6144 12588 6150 12640
rect 7006 12628 7012 12640
rect 6967 12600 7012 12628
rect 7006 12588 7012 12600
rect 7064 12588 7070 12640
rect 7208 12628 7236 12668
rect 8312 12668 10149 12696
rect 8312 12628 8340 12668
rect 10137 12665 10149 12668
rect 10183 12665 10195 12699
rect 10870 12696 10876 12708
rect 10831 12668 10876 12696
rect 10137 12659 10195 12665
rect 8478 12628 8484 12640
rect 7208 12600 8340 12628
rect 8439 12600 8484 12628
rect 8478 12588 8484 12600
rect 8536 12588 8542 12640
rect 10152 12628 10180 12659
rect 10870 12656 10876 12668
rect 10928 12696 10934 12708
rect 11256 12696 11284 12804
rect 11974 12792 11980 12804
rect 12032 12832 12038 12844
rect 12253 12835 12311 12841
rect 12253 12832 12265 12835
rect 12032 12804 12265 12832
rect 12032 12792 12038 12804
rect 12253 12801 12265 12804
rect 12299 12801 12311 12835
rect 12253 12795 12311 12801
rect 11514 12724 11520 12776
rect 11572 12764 11578 12776
rect 12158 12764 12164 12776
rect 11572 12736 11744 12764
rect 12119 12736 12164 12764
rect 11572 12724 11578 12736
rect 10928 12668 11284 12696
rect 11333 12699 11391 12705
rect 10928 12656 10934 12668
rect 11333 12665 11345 12699
rect 11379 12696 11391 12699
rect 11606 12696 11612 12708
rect 11379 12668 11612 12696
rect 11379 12665 11391 12668
rect 11333 12659 11391 12665
rect 11606 12656 11612 12668
rect 11664 12656 11670 12708
rect 11716 12696 11744 12736
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 12268 12764 12296 12795
rect 12342 12792 12348 12844
rect 12400 12832 12406 12844
rect 12597 12835 12655 12841
rect 12597 12832 12609 12835
rect 12400 12804 12609 12832
rect 12400 12792 12406 12804
rect 12597 12801 12609 12804
rect 12643 12801 12655 12835
rect 12597 12795 12655 12801
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12801 12771 12835
rect 12713 12795 12771 12801
rect 12728 12764 12756 12795
rect 12802 12792 12808 12844
rect 12860 12832 12866 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12860 12804 13001 12832
rect 12860 12792 12866 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 12989 12795 13047 12801
rect 13078 12792 13084 12844
rect 13136 12832 13142 12844
rect 13449 12835 13507 12841
rect 13449 12832 13461 12835
rect 13136 12804 13461 12832
rect 13136 12792 13142 12804
rect 13449 12801 13461 12804
rect 13495 12801 13507 12835
rect 13449 12795 13507 12801
rect 13538 12792 13544 12844
rect 13596 12832 13602 12844
rect 14001 12835 14059 12841
rect 13596 12804 13641 12832
rect 13596 12792 13602 12804
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14090 12832 14096 12844
rect 14047 12804 14096 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 14090 12792 14096 12804
rect 14148 12792 14154 12844
rect 14292 12841 14320 12940
rect 15565 12937 15577 12971
rect 15611 12968 15623 12971
rect 15838 12968 15844 12980
rect 15611 12940 15844 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 15838 12928 15844 12940
rect 15896 12928 15902 12980
rect 16669 12903 16727 12909
rect 16669 12900 16681 12903
rect 14660 12872 16681 12900
rect 14253 12835 14320 12841
rect 14253 12801 14265 12835
rect 14299 12804 14320 12835
rect 14369 12835 14427 12841
rect 14299 12801 14311 12804
rect 14253 12795 14311 12801
rect 14369 12801 14381 12835
rect 14415 12832 14427 12835
rect 14550 12832 14556 12844
rect 14415 12804 14556 12832
rect 14415 12801 14427 12804
rect 14369 12795 14427 12801
rect 14550 12792 14556 12804
rect 14608 12792 14614 12844
rect 13354 12764 13360 12776
rect 12268 12736 12756 12764
rect 12820 12736 13360 12764
rect 12437 12699 12495 12705
rect 12437 12696 12449 12699
rect 11716 12668 12449 12696
rect 12437 12665 12449 12668
rect 12483 12665 12495 12699
rect 12437 12659 12495 12665
rect 12526 12656 12532 12708
rect 12584 12696 12590 12708
rect 12820 12696 12848 12736
rect 13354 12724 13360 12736
rect 13412 12764 13418 12776
rect 14660 12764 14688 12872
rect 16669 12869 16681 12872
rect 16715 12869 16727 12903
rect 16669 12863 16727 12869
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 15289 12835 15347 12841
rect 14792 12804 14837 12832
rect 14792 12792 14798 12804
rect 15289 12801 15301 12835
rect 15335 12832 15347 12835
rect 15470 12832 15476 12844
rect 15335 12804 15476 12832
rect 15335 12801 15347 12804
rect 15289 12795 15347 12801
rect 15470 12792 15476 12804
rect 15528 12792 15534 12844
rect 15654 12832 15660 12844
rect 15615 12804 15660 12832
rect 15654 12792 15660 12804
rect 15712 12792 15718 12844
rect 16022 12832 16028 12844
rect 15983 12804 16028 12832
rect 16022 12792 16028 12804
rect 16080 12792 16086 12844
rect 16393 12835 16451 12841
rect 16393 12801 16405 12835
rect 16439 12832 16451 12835
rect 16482 12832 16488 12844
rect 16439 12804 16488 12832
rect 16439 12801 16451 12804
rect 16393 12795 16451 12801
rect 16482 12792 16488 12804
rect 16540 12792 16546 12844
rect 18230 12764 18236 12776
rect 13412 12736 14688 12764
rect 15120 12736 18236 12764
rect 13412 12724 13418 12736
rect 12584 12668 12848 12696
rect 12897 12699 12955 12705
rect 12584 12656 12590 12668
rect 12897 12665 12909 12699
rect 12943 12696 12955 12699
rect 12986 12696 12992 12708
rect 12943 12668 12992 12696
rect 12943 12665 12955 12668
rect 12897 12659 12955 12665
rect 12986 12656 12992 12668
rect 13044 12656 13050 12708
rect 14182 12696 14188 12708
rect 13188 12668 14188 12696
rect 11514 12628 11520 12640
rect 10152 12600 11520 12628
rect 11514 12588 11520 12600
rect 11572 12588 11578 12640
rect 11793 12631 11851 12637
rect 11793 12597 11805 12631
rect 11839 12628 11851 12631
rect 13188 12628 13216 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 14274 12656 14280 12708
rect 14332 12696 14338 12708
rect 14921 12699 14979 12705
rect 14921 12696 14933 12699
rect 14332 12668 14933 12696
rect 14332 12656 14338 12668
rect 14921 12665 14933 12668
rect 14967 12665 14979 12699
rect 14921 12659 14979 12665
rect 11839 12600 13216 12628
rect 11839 12597 11851 12600
rect 11793 12591 11851 12597
rect 13262 12588 13268 12640
rect 13320 12628 13326 12640
rect 13320 12600 13365 12628
rect 13320 12588 13326 12600
rect 13630 12588 13636 12640
rect 13688 12628 13694 12640
rect 13725 12631 13783 12637
rect 13725 12628 13737 12631
rect 13688 12600 13737 12628
rect 13688 12588 13694 12600
rect 13725 12597 13737 12600
rect 13771 12597 13783 12631
rect 14090 12628 14096 12640
rect 14051 12600 14096 12628
rect 13725 12591 13783 12597
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14553 12631 14611 12637
rect 14553 12597 14565 12631
rect 14599 12628 14611 12631
rect 15120 12628 15148 12736
rect 18230 12724 18236 12736
rect 18288 12724 18294 12776
rect 15378 12656 15384 12708
rect 15436 12696 15442 12708
rect 15841 12699 15899 12705
rect 15841 12696 15853 12699
rect 15436 12668 15853 12696
rect 15436 12656 15442 12668
rect 15841 12665 15853 12668
rect 15887 12665 15899 12699
rect 16206 12696 16212 12708
rect 16119 12668 16212 12696
rect 15841 12659 15899 12665
rect 16206 12656 16212 12668
rect 16264 12696 16270 12708
rect 18138 12696 18144 12708
rect 16264 12668 18144 12696
rect 16264 12656 16270 12668
rect 18138 12656 18144 12668
rect 18196 12656 18202 12708
rect 14599 12600 15148 12628
rect 14599 12597 14611 12600
rect 14553 12591 14611 12597
rect 15194 12588 15200 12640
rect 15252 12628 15258 12640
rect 15252 12600 15297 12628
rect 15252 12588 15258 12600
rect 16390 12588 16396 12640
rect 16448 12628 16454 12640
rect 17957 12631 18015 12637
rect 17957 12628 17969 12631
rect 16448 12600 17969 12628
rect 16448 12588 16454 12600
rect 17957 12597 17969 12600
rect 18003 12597 18015 12631
rect 17957 12591 18015 12597
rect 1104 12538 18860 12560
rect 1104 12486 3174 12538
rect 3226 12486 3238 12538
rect 3290 12486 3302 12538
rect 3354 12486 3366 12538
rect 3418 12486 3430 12538
rect 3482 12486 7622 12538
rect 7674 12486 7686 12538
rect 7738 12486 7750 12538
rect 7802 12486 7814 12538
rect 7866 12486 7878 12538
rect 7930 12486 12070 12538
rect 12122 12486 12134 12538
rect 12186 12486 12198 12538
rect 12250 12486 12262 12538
rect 12314 12486 12326 12538
rect 12378 12486 16518 12538
rect 16570 12486 16582 12538
rect 16634 12486 16646 12538
rect 16698 12486 16710 12538
rect 16762 12486 16774 12538
rect 16826 12486 18860 12538
rect 1104 12464 18860 12486
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 7466 12424 7472 12436
rect 2832 12396 7472 12424
rect 2832 12384 2838 12396
rect 7466 12384 7472 12396
rect 7524 12384 7530 12436
rect 8570 12384 8576 12436
rect 8628 12424 8634 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8628 12396 9137 12424
rect 8628 12384 8634 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 9582 12424 9588 12436
rect 9125 12387 9183 12393
rect 9232 12396 9588 12424
rect 2866 12356 2872 12368
rect 2746 12328 2872 12356
rect 2406 12288 2412 12300
rect 2367 12260 2412 12288
rect 2406 12248 2412 12260
rect 2464 12248 2470 12300
rect 1946 12220 1952 12232
rect 1907 12192 1952 12220
rect 1946 12180 1952 12192
rect 2004 12180 2010 12232
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12220 2283 12223
rect 2746 12220 2774 12328
rect 2866 12316 2872 12328
rect 2924 12356 2930 12368
rect 6730 12356 6736 12368
rect 2924 12328 6736 12356
rect 2924 12316 2930 12328
rect 6730 12316 6736 12328
rect 6788 12316 6794 12368
rect 6914 12316 6920 12368
rect 6972 12356 6978 12368
rect 7190 12356 7196 12368
rect 6972 12328 7196 12356
rect 6972 12316 6978 12328
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 8665 12359 8723 12365
rect 8665 12356 8677 12359
rect 7300 12328 8677 12356
rect 3418 12288 3424 12300
rect 3379 12260 3424 12288
rect 3418 12248 3424 12260
rect 3476 12248 3482 12300
rect 4522 12288 4528 12300
rect 3528 12260 4528 12288
rect 2271 12192 2774 12220
rect 2271 12189 2283 12192
rect 2225 12183 2283 12189
rect 2958 12180 2964 12232
rect 3016 12220 3022 12232
rect 3237 12223 3295 12229
rect 3237 12220 3249 12223
rect 3016 12192 3249 12220
rect 3016 12180 3022 12192
rect 3237 12189 3249 12192
rect 3283 12220 3295 12223
rect 3528 12220 3556 12260
rect 4522 12248 4528 12260
rect 4580 12248 4586 12300
rect 4614 12248 4620 12300
rect 4672 12288 4678 12300
rect 5810 12288 5816 12300
rect 4672 12260 5816 12288
rect 4672 12248 4678 12260
rect 5810 12248 5816 12260
rect 5868 12248 5874 12300
rect 5902 12248 5908 12300
rect 5960 12288 5966 12300
rect 6638 12288 6644 12300
rect 5960 12260 6644 12288
rect 5960 12248 5966 12260
rect 6638 12248 6644 12260
rect 6696 12288 6702 12300
rect 7300 12288 7328 12328
rect 8665 12325 8677 12328
rect 8711 12356 8723 12359
rect 9232 12356 9260 12396
rect 9582 12384 9588 12396
rect 9640 12384 9646 12436
rect 9674 12384 9680 12436
rect 9732 12424 9738 12436
rect 9769 12427 9827 12433
rect 9769 12424 9781 12427
rect 9732 12396 9781 12424
rect 9732 12384 9738 12396
rect 9769 12393 9781 12396
rect 9815 12393 9827 12427
rect 10134 12424 10140 12436
rect 10095 12396 10140 12424
rect 9769 12387 9827 12393
rect 10134 12384 10140 12396
rect 10192 12384 10198 12436
rect 10226 12384 10232 12436
rect 10284 12424 10290 12436
rect 11149 12427 11207 12433
rect 10284 12396 10732 12424
rect 10284 12384 10290 12396
rect 8711 12328 9260 12356
rect 8711 12325 8723 12328
rect 8665 12319 8723 12325
rect 9398 12316 9404 12368
rect 9456 12356 9462 12368
rect 10042 12356 10048 12368
rect 9456 12328 10048 12356
rect 9456 12316 9462 12328
rect 10042 12316 10048 12328
rect 10100 12316 10106 12368
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 10594 12356 10600 12368
rect 10468 12328 10600 12356
rect 10468 12316 10474 12328
rect 10594 12316 10600 12328
rect 10652 12316 10658 12368
rect 10704 12356 10732 12396
rect 11149 12393 11161 12427
rect 11195 12424 11207 12427
rect 11238 12424 11244 12436
rect 11195 12396 11244 12424
rect 11195 12393 11207 12396
rect 11149 12387 11207 12393
rect 11238 12384 11244 12396
rect 11296 12384 11302 12436
rect 11330 12384 11336 12436
rect 11388 12424 11394 12436
rect 11790 12424 11796 12436
rect 11388 12396 11796 12424
rect 11388 12384 11394 12396
rect 11790 12384 11796 12396
rect 11848 12384 11854 12436
rect 14458 12424 14464 12436
rect 12360 12396 14464 12424
rect 11517 12359 11575 12365
rect 10704 12328 11284 12356
rect 11256 12300 11284 12328
rect 11517 12325 11529 12359
rect 11563 12356 11575 12359
rect 11698 12356 11704 12368
rect 11563 12328 11704 12356
rect 11563 12325 11575 12328
rect 11517 12319 11575 12325
rect 11698 12316 11704 12328
rect 11756 12316 11762 12368
rect 11882 12356 11888 12368
rect 11843 12328 11888 12356
rect 11882 12316 11888 12328
rect 11940 12316 11946 12368
rect 12360 12356 12388 12396
rect 14458 12384 14464 12396
rect 14516 12384 14522 12436
rect 14918 12384 14924 12436
rect 14976 12424 14982 12436
rect 14976 12396 16712 12424
rect 14976 12384 14982 12396
rect 12084 12328 12388 12356
rect 6696 12260 7328 12288
rect 6696 12248 6702 12260
rect 7650 12248 7656 12300
rect 7708 12288 7714 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 7708 12260 10793 12288
rect 7708 12248 7714 12260
rect 10781 12257 10793 12260
rect 10827 12288 10839 12291
rect 11054 12288 11060 12300
rect 10827 12260 11060 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11054 12248 11060 12260
rect 11112 12248 11118 12300
rect 11238 12248 11244 12300
rect 11296 12248 11302 12300
rect 12084 12288 12112 12328
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 13449 12359 13507 12365
rect 13449 12356 13461 12359
rect 12492 12328 13461 12356
rect 12492 12316 12498 12328
rect 13449 12325 13461 12328
rect 13495 12325 13507 12359
rect 13449 12319 13507 12325
rect 13722 12316 13728 12368
rect 13780 12356 13786 12368
rect 16117 12359 16175 12365
rect 13780 12328 15976 12356
rect 13780 12316 13786 12328
rect 11348 12260 12112 12288
rect 3283 12192 3556 12220
rect 4433 12223 4491 12229
rect 3283 12189 3295 12192
rect 3237 12183 3295 12189
rect 4433 12189 4445 12223
rect 4479 12189 4491 12223
rect 4433 12183 4491 12189
rect 2498 12112 2504 12164
rect 2556 12152 2562 12164
rect 2556 12124 3280 12152
rect 2556 12112 2562 12124
rect 2590 12084 2596 12096
rect 2551 12056 2596 12084
rect 2590 12044 2596 12056
rect 2648 12044 2654 12096
rect 2682 12044 2688 12096
rect 2740 12084 2746 12096
rect 3053 12087 3111 12093
rect 2740 12056 2785 12084
rect 2740 12044 2746 12056
rect 3053 12053 3065 12087
rect 3099 12084 3111 12087
rect 3142 12084 3148 12096
rect 3099 12056 3148 12084
rect 3099 12053 3111 12056
rect 3053 12047 3111 12053
rect 3142 12044 3148 12056
rect 3200 12044 3206 12096
rect 3252 12084 3280 12124
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 3881 12155 3939 12161
rect 3881 12152 3893 12155
rect 3384 12124 3893 12152
rect 3384 12112 3390 12124
rect 3881 12121 3893 12124
rect 3927 12152 3939 12155
rect 4062 12152 4068 12164
rect 3927 12124 4068 12152
rect 3927 12121 3939 12124
rect 3881 12115 3939 12121
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 4448 12152 4476 12183
rect 4798 12180 4804 12232
rect 4856 12220 4862 12232
rect 5353 12223 5411 12229
rect 5353 12220 5365 12223
rect 4856 12192 5365 12220
rect 4856 12180 4862 12192
rect 5353 12189 5365 12192
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 5442 12180 5448 12232
rect 5500 12220 5506 12232
rect 6189 12223 6247 12229
rect 5500 12192 5545 12220
rect 5500 12180 5506 12192
rect 6189 12189 6201 12223
rect 6235 12220 6247 12223
rect 6235 12192 6316 12220
rect 6235 12189 6247 12192
rect 6189 12183 6247 12189
rect 5994 12152 6000 12164
rect 4448 12124 6000 12152
rect 5994 12112 6000 12124
rect 6052 12112 6058 12164
rect 6288 12152 6316 12192
rect 6362 12180 6368 12232
rect 6420 12216 6426 12232
rect 6457 12223 6515 12229
rect 6457 12216 6469 12223
rect 6420 12189 6469 12216
rect 6503 12189 6515 12223
rect 6420 12188 6515 12189
rect 6420 12180 6426 12188
rect 6457 12183 6515 12188
rect 7193 12223 7251 12229
rect 7193 12189 7205 12223
rect 7239 12220 7251 12223
rect 7282 12220 7288 12232
rect 7239 12192 7288 12220
rect 7239 12189 7251 12192
rect 7193 12183 7251 12189
rect 7282 12180 7288 12192
rect 7340 12180 7346 12232
rect 7466 12220 7472 12232
rect 7427 12192 7472 12220
rect 7466 12180 7472 12192
rect 7524 12180 7530 12232
rect 8294 12180 8300 12232
rect 8352 12220 8358 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8352 12192 9321 12220
rect 8352 12180 8358 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 10962 12220 10968 12232
rect 9309 12183 9367 12189
rect 9600 12192 10968 12220
rect 8110 12152 8116 12164
rect 6196 12124 6316 12152
rect 8071 12124 8116 12152
rect 6196 12096 6224 12124
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 9600 12152 9628 12192
rect 10962 12180 10968 12192
rect 11020 12220 11026 12232
rect 11348 12229 11376 12260
rect 12986 12248 12992 12300
rect 13044 12288 13050 12300
rect 14826 12288 14832 12300
rect 13044 12260 14596 12288
rect 14787 12260 14832 12288
rect 13044 12248 13050 12260
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11020 12192 11345 12220
rect 11020 12180 11026 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 11790 12180 11796 12232
rect 11848 12220 11854 12232
rect 12360 12229 12572 12236
rect 12360 12223 12587 12229
rect 12360 12220 12541 12223
rect 11848 12208 12541 12220
rect 11848 12192 12388 12208
rect 11848 12180 11854 12192
rect 12529 12189 12541 12208
rect 12575 12189 12587 12223
rect 12802 12220 12808 12232
rect 12763 12192 12808 12220
rect 12529 12183 12587 12189
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 12894 12180 12900 12232
rect 12952 12220 12958 12232
rect 13170 12220 13176 12232
rect 12952 12192 12997 12220
rect 13131 12192 13176 12220
rect 12952 12180 12958 12192
rect 13170 12180 13176 12192
rect 13228 12180 13234 12232
rect 13633 12223 13691 12229
rect 13633 12189 13645 12223
rect 13679 12189 13691 12223
rect 13633 12183 13691 12189
rect 8220 12124 9628 12152
rect 10045 12155 10103 12161
rect 3513 12087 3571 12093
rect 3513 12084 3525 12087
rect 3252 12056 3525 12084
rect 3513 12053 3525 12056
rect 3559 12053 3571 12087
rect 3970 12084 3976 12096
rect 3931 12056 3976 12084
rect 3513 12047 3571 12053
rect 3970 12044 3976 12056
rect 4028 12044 4034 12096
rect 4246 12084 4252 12096
rect 4207 12056 4252 12084
rect 4246 12044 4252 12056
rect 4304 12044 4310 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 5810 12084 5816 12096
rect 4755 12056 5816 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6086 12084 6092 12096
rect 6047 12056 6092 12084
rect 6086 12044 6092 12056
rect 6144 12044 6150 12096
rect 6178 12044 6184 12096
rect 6236 12044 6242 12096
rect 6365 12087 6423 12093
rect 6365 12053 6377 12087
rect 6411 12084 6423 12087
rect 6546 12084 6552 12096
rect 6411 12056 6552 12084
rect 6411 12053 6423 12056
rect 6365 12047 6423 12053
rect 6546 12044 6552 12056
rect 6604 12044 6610 12096
rect 7098 12084 7104 12096
rect 7059 12056 7104 12084
rect 7098 12044 7104 12056
rect 7156 12044 7162 12096
rect 7377 12087 7435 12093
rect 7377 12053 7389 12087
rect 7423 12084 7435 12087
rect 7558 12084 7564 12096
rect 7423 12056 7564 12084
rect 7423 12053 7435 12056
rect 7377 12047 7435 12053
rect 7558 12044 7564 12056
rect 7616 12044 7622 12096
rect 7742 12044 7748 12096
rect 7800 12084 7806 12096
rect 8220 12093 8248 12124
rect 10045 12121 10057 12155
rect 10091 12152 10103 12155
rect 10134 12152 10140 12164
rect 10091 12124 10140 12152
rect 10091 12121 10103 12124
rect 10045 12115 10103 12121
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 10686 12112 10692 12164
rect 10744 12152 10750 12164
rect 10873 12155 10931 12161
rect 10873 12152 10885 12155
rect 10744 12124 10885 12152
rect 10744 12112 10750 12124
rect 10873 12121 10885 12124
rect 10919 12121 10931 12155
rect 10873 12115 10931 12121
rect 11238 12112 11244 12164
rect 11296 12152 11302 12164
rect 13648 12152 13676 12183
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13780 12192 14105 12220
rect 13780 12180 13786 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 14182 12180 14188 12232
rect 14240 12220 14246 12232
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 14240 12192 14473 12220
rect 14240 12180 14246 12192
rect 14461 12189 14473 12192
rect 14507 12189 14519 12223
rect 14568 12220 14596 12260
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 15948 12229 15976 12328
rect 16117 12325 16129 12359
rect 16163 12356 16175 12359
rect 16163 12328 16620 12356
rect 16163 12325 16175 12328
rect 16117 12319 16175 12325
rect 15565 12223 15623 12229
rect 15565 12220 15577 12223
rect 14568 12192 15577 12220
rect 14461 12183 14519 12189
rect 15565 12189 15577 12192
rect 15611 12189 15623 12223
rect 15565 12183 15623 12189
rect 15933 12223 15991 12229
rect 15933 12189 15945 12223
rect 15979 12189 15991 12223
rect 15933 12183 15991 12189
rect 11296 12124 13676 12152
rect 13740 12124 15976 12152
rect 11296 12112 11302 12124
rect 8205 12087 8263 12093
rect 8205 12084 8217 12087
rect 7800 12056 8217 12084
rect 7800 12044 7806 12056
rect 8205 12053 8217 12056
rect 8251 12053 8263 12087
rect 8478 12084 8484 12096
rect 8439 12056 8484 12084
rect 8205 12047 8263 12053
rect 8478 12044 8484 12056
rect 8536 12044 8542 12096
rect 9033 12087 9091 12093
rect 9033 12053 9045 12087
rect 9079 12084 9091 12087
rect 9214 12084 9220 12096
rect 9079 12056 9220 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 9214 12044 9220 12056
rect 9272 12044 9278 12096
rect 9490 12084 9496 12096
rect 9451 12056 9496 12084
rect 9490 12044 9496 12056
rect 9548 12044 9554 12096
rect 9582 12044 9588 12096
rect 9640 12084 9646 12096
rect 10318 12084 10324 12096
rect 9640 12056 10324 12084
rect 9640 12044 9646 12056
rect 10318 12044 10324 12056
rect 10376 12044 10382 12096
rect 10410 12044 10416 12096
rect 10468 12084 10474 12096
rect 10505 12087 10563 12093
rect 10505 12084 10517 12087
rect 10468 12056 10517 12084
rect 10468 12044 10474 12056
rect 10505 12053 10517 12056
rect 10551 12084 10563 12087
rect 11146 12084 11152 12096
rect 10551 12056 11152 12084
rect 10551 12053 10563 12056
rect 10505 12047 10563 12053
rect 11146 12044 11152 12056
rect 11204 12044 11210 12096
rect 11698 12084 11704 12096
rect 11659 12056 11704 12084
rect 11698 12044 11704 12056
rect 11756 12044 11762 12096
rect 11974 12084 11980 12096
rect 11935 12056 11980 12084
rect 11974 12044 11980 12056
rect 12032 12044 12038 12096
rect 12158 12084 12164 12096
rect 12119 12056 12164 12084
rect 12158 12044 12164 12056
rect 12216 12044 12222 12096
rect 12342 12084 12348 12096
rect 12303 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 12526 12044 12532 12096
rect 12584 12084 12590 12096
rect 12621 12087 12679 12093
rect 12621 12084 12633 12087
rect 12584 12056 12633 12084
rect 12584 12044 12590 12056
rect 12621 12053 12633 12056
rect 12667 12053 12679 12087
rect 13078 12084 13084 12096
rect 13039 12056 13084 12084
rect 12621 12047 12679 12053
rect 13078 12044 13084 12056
rect 13136 12044 13142 12096
rect 13357 12087 13415 12093
rect 13357 12053 13369 12087
rect 13403 12084 13415 12087
rect 13740 12084 13768 12124
rect 15948 12096 15976 12124
rect 16206 12112 16212 12164
rect 16264 12152 16270 12164
rect 16485 12155 16543 12161
rect 16485 12152 16497 12155
rect 16264 12124 16497 12152
rect 16264 12112 16270 12124
rect 16485 12121 16497 12124
rect 16531 12121 16543 12155
rect 16592 12152 16620 12328
rect 16684 12229 16712 12396
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17129 12427 17187 12433
rect 17129 12424 17141 12427
rect 17000 12396 17141 12424
rect 17000 12384 17006 12396
rect 17129 12393 17141 12396
rect 17175 12424 17187 12427
rect 18966 12424 18972 12436
rect 17175 12396 18972 12424
rect 17175 12393 17187 12396
rect 17129 12387 17187 12393
rect 18966 12384 18972 12396
rect 19024 12384 19030 12436
rect 16853 12359 16911 12365
rect 16853 12325 16865 12359
rect 16899 12356 16911 12359
rect 18874 12356 18880 12368
rect 16899 12328 18880 12356
rect 16899 12325 16911 12328
rect 16853 12319 16911 12325
rect 18874 12316 18880 12328
rect 18932 12316 18938 12368
rect 17678 12288 17684 12300
rect 17639 12260 17684 12288
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 17954 12288 17960 12300
rect 17915 12260 17960 12288
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18046 12248 18052 12300
rect 18104 12288 18110 12300
rect 18414 12288 18420 12300
rect 18104 12260 18420 12288
rect 18104 12248 18110 12260
rect 18414 12248 18420 12260
rect 18472 12248 18478 12300
rect 16669 12223 16727 12229
rect 16669 12189 16681 12223
rect 16715 12189 16727 12223
rect 17405 12223 17463 12229
rect 16669 12183 16727 12189
rect 17052 12192 17356 12220
rect 17052 12152 17080 12192
rect 17218 12152 17224 12164
rect 16592 12124 17080 12152
rect 17179 12124 17224 12152
rect 16485 12115 16543 12121
rect 17218 12112 17224 12124
rect 17276 12112 17282 12164
rect 17328 12152 17356 12192
rect 17405 12189 17417 12223
rect 17451 12220 17463 12223
rect 17494 12220 17500 12232
rect 17451 12192 17500 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 17494 12180 17500 12192
rect 17552 12180 17558 12232
rect 18046 12152 18052 12164
rect 17328 12124 18052 12152
rect 18046 12112 18052 12124
rect 18104 12112 18110 12164
rect 13403 12056 13768 12084
rect 13403 12053 13415 12056
rect 13357 12047 13415 12053
rect 13814 12044 13820 12096
rect 13872 12084 13878 12096
rect 14277 12087 14335 12093
rect 13872 12056 13917 12084
rect 13872 12044 13878 12056
rect 14277 12053 14289 12087
rect 14323 12084 14335 12087
rect 14918 12084 14924 12096
rect 14323 12056 14924 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 14918 12044 14924 12056
rect 14976 12044 14982 12096
rect 15010 12044 15016 12096
rect 15068 12084 15074 12096
rect 15286 12084 15292 12096
rect 15068 12056 15292 12084
rect 15068 12044 15074 12056
rect 15286 12044 15292 12056
rect 15344 12044 15350 12096
rect 15746 12044 15752 12096
rect 15804 12084 15810 12096
rect 15804 12056 15849 12084
rect 15804 12044 15810 12056
rect 15930 12044 15936 12096
rect 15988 12044 15994 12096
rect 16114 12044 16120 12096
rect 16172 12084 16178 12096
rect 16393 12087 16451 12093
rect 16393 12084 16405 12087
rect 16172 12056 16405 12084
rect 16172 12044 16178 12056
rect 16393 12053 16405 12056
rect 16439 12053 16451 12087
rect 16393 12047 16451 12053
rect 17589 12087 17647 12093
rect 17589 12053 17601 12087
rect 17635 12084 17647 12087
rect 18322 12084 18328 12096
rect 17635 12056 18328 12084
rect 17635 12053 17647 12056
rect 17589 12047 17647 12053
rect 18322 12044 18328 12056
rect 18380 12044 18386 12096
rect 1104 11994 18860 12016
rect 1104 11942 5398 11994
rect 5450 11942 5462 11994
rect 5514 11942 5526 11994
rect 5578 11942 5590 11994
rect 5642 11942 5654 11994
rect 5706 11942 9846 11994
rect 9898 11942 9910 11994
rect 9962 11942 9974 11994
rect 10026 11942 10038 11994
rect 10090 11942 10102 11994
rect 10154 11942 14294 11994
rect 14346 11942 14358 11994
rect 14410 11942 14422 11994
rect 14474 11942 14486 11994
rect 14538 11942 14550 11994
rect 14602 11942 18860 11994
rect 1104 11920 18860 11942
rect 2590 11840 2596 11892
rect 2648 11880 2654 11892
rect 3053 11883 3111 11889
rect 3053 11880 3065 11883
rect 2648 11852 3065 11880
rect 2648 11840 2654 11852
rect 3053 11849 3065 11852
rect 3099 11849 3111 11883
rect 3053 11843 3111 11849
rect 3881 11883 3939 11889
rect 3881 11849 3893 11883
rect 3927 11880 3939 11883
rect 4249 11883 4307 11889
rect 4249 11880 4261 11883
rect 3927 11852 4261 11880
rect 3927 11849 3939 11852
rect 3881 11843 3939 11849
rect 4249 11849 4261 11852
rect 4295 11849 4307 11883
rect 4249 11843 4307 11849
rect 4709 11883 4767 11889
rect 4709 11849 4721 11883
rect 4755 11880 4767 11883
rect 11333 11883 11391 11889
rect 4755 11852 11008 11880
rect 4755 11849 4767 11852
rect 4709 11843 4767 11849
rect 2038 11772 2044 11824
rect 2096 11812 2102 11824
rect 2096 11784 2636 11812
rect 2096 11772 2102 11784
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2608 11744 2636 11784
rect 3142 11772 3148 11824
rect 3200 11812 3206 11824
rect 4341 11815 4399 11821
rect 4341 11812 4353 11815
rect 3200 11784 4353 11812
rect 3200 11772 3206 11784
rect 4341 11781 4353 11784
rect 4387 11781 4399 11815
rect 4341 11775 4399 11781
rect 5902 11772 5908 11824
rect 5960 11812 5966 11824
rect 6089 11815 6147 11821
rect 6089 11812 6101 11815
rect 5960 11784 6101 11812
rect 5960 11772 5966 11784
rect 6089 11781 6101 11784
rect 6135 11781 6147 11815
rect 6089 11775 6147 11781
rect 2685 11747 2743 11753
rect 2685 11744 2697 11747
rect 2608 11716 2697 11744
rect 2685 11713 2697 11716
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 3513 11747 3571 11753
rect 3513 11713 3525 11747
rect 3559 11744 3571 11747
rect 3786 11744 3792 11756
rect 3559 11716 3792 11744
rect 3559 11713 3571 11716
rect 3513 11707 3571 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 5077 11747 5135 11753
rect 5077 11713 5089 11747
rect 5123 11744 5135 11747
rect 5718 11744 5724 11756
rect 5123 11716 5724 11744
rect 5123 11713 5135 11716
rect 5077 11707 5135 11713
rect 5718 11704 5724 11716
rect 5776 11704 5782 11756
rect 5994 11744 6000 11756
rect 5955 11716 6000 11744
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 1118 11636 1124 11688
rect 1176 11676 1182 11688
rect 1949 11679 2007 11685
rect 1949 11676 1961 11679
rect 1176 11648 1961 11676
rect 1176 11636 1182 11648
rect 1949 11645 1961 11648
rect 1995 11645 2007 11679
rect 1949 11639 2007 11645
rect 2130 11636 2136 11688
rect 2188 11676 2194 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 2188 11648 2421 11676
rect 2188 11636 2194 11648
rect 2409 11645 2421 11648
rect 2455 11645 2467 11679
rect 2409 11639 2467 11645
rect 2593 11679 2651 11685
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3050 11676 3056 11688
rect 2639 11648 3056 11676
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3050 11636 3056 11648
rect 3108 11636 3114 11688
rect 3237 11679 3295 11685
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3970 11676 3976 11688
rect 3467 11648 3976 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 2038 11568 2044 11620
rect 2096 11608 2102 11620
rect 3252 11608 3280 11639
rect 3970 11636 3976 11648
rect 4028 11636 4034 11688
rect 4065 11679 4123 11685
rect 4065 11645 4077 11679
rect 4111 11645 4123 11679
rect 4065 11639 4123 11645
rect 2096 11580 3280 11608
rect 2096 11568 2102 11580
rect 1394 11500 1400 11552
rect 1452 11540 1458 11552
rect 2590 11540 2596 11552
rect 1452 11512 2596 11540
rect 1452 11500 1458 11512
rect 2590 11500 2596 11512
rect 2648 11540 2654 11552
rect 4080 11540 4108 11639
rect 4338 11636 4344 11688
rect 4396 11676 4402 11688
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 4396 11648 5273 11676
rect 4396 11636 4402 11648
rect 5261 11645 5273 11648
rect 5307 11676 5319 11679
rect 5350 11676 5356 11688
rect 5307 11648 5356 11676
rect 5307 11645 5319 11648
rect 5261 11639 5319 11645
rect 5350 11636 5356 11648
rect 5408 11636 5414 11688
rect 6104 11608 6132 11775
rect 6270 11772 6276 11824
rect 6328 11812 6334 11824
rect 7006 11812 7012 11824
rect 6328 11784 7012 11812
rect 6328 11772 6334 11784
rect 7006 11772 7012 11784
rect 7064 11772 7070 11824
rect 7742 11812 7748 11824
rect 7703 11784 7748 11812
rect 7742 11772 7748 11784
rect 7800 11772 7806 11824
rect 8018 11772 8024 11824
rect 8076 11812 8082 11824
rect 8076 11784 8156 11812
rect 8076 11772 8082 11784
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6454 11744 6460 11756
rect 6236 11716 6460 11744
rect 6236 11704 6242 11716
rect 6454 11704 6460 11716
rect 6512 11704 6518 11756
rect 6730 11704 6736 11756
rect 6788 11744 6794 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6788 11716 6837 11744
rect 6788 11704 6794 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 7650 11744 7656 11756
rect 6825 11707 6883 11713
rect 7116 11716 7656 11744
rect 6270 11636 6276 11688
rect 6328 11676 6334 11688
rect 6917 11679 6975 11685
rect 6917 11676 6929 11679
rect 6328 11648 6929 11676
rect 6328 11636 6334 11648
rect 6917 11645 6929 11648
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 7009 11679 7067 11685
rect 7009 11645 7021 11679
rect 7055 11645 7067 11679
rect 7009 11639 7067 11645
rect 6104 11580 6776 11608
rect 2648 11512 4108 11540
rect 2648 11500 2654 11512
rect 4154 11500 4160 11552
rect 4212 11540 4218 11552
rect 4614 11540 4620 11552
rect 4212 11512 4620 11540
rect 4212 11500 4218 11512
rect 4614 11500 4620 11512
rect 4672 11500 4678 11552
rect 4890 11540 4896 11552
rect 4851 11512 4896 11540
rect 4890 11500 4896 11512
rect 4948 11500 4954 11552
rect 5258 11500 5264 11552
rect 5316 11540 5322 11552
rect 5353 11543 5411 11549
rect 5353 11540 5365 11543
rect 5316 11512 5365 11540
rect 5316 11500 5322 11512
rect 5353 11509 5365 11512
rect 5399 11509 5411 11543
rect 5353 11503 5411 11509
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6178 11540 6184 11552
rect 5960 11512 6184 11540
rect 5960 11500 5966 11512
rect 6178 11500 6184 11512
rect 6236 11500 6242 11552
rect 6454 11540 6460 11552
rect 6415 11512 6460 11540
rect 6454 11500 6460 11512
rect 6512 11500 6518 11552
rect 6748 11540 6776 11580
rect 6822 11568 6828 11620
rect 6880 11608 6886 11620
rect 7024 11608 7052 11639
rect 6880 11580 7052 11608
rect 6880 11568 6886 11580
rect 7116 11540 7144 11716
rect 7650 11704 7656 11716
rect 7708 11704 7714 11756
rect 8128 11753 8156 11784
rect 9122 11772 9128 11824
rect 9180 11812 9186 11824
rect 9180 11784 10364 11812
rect 9180 11772 9186 11784
rect 8113 11747 8171 11753
rect 8113 11713 8125 11747
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 8757 11747 8815 11753
rect 8757 11713 8769 11747
rect 8803 11744 8815 11747
rect 8846 11744 8852 11756
rect 8803 11716 8852 11744
rect 8803 11713 8815 11716
rect 8757 11707 8815 11713
rect 8846 11704 8852 11716
rect 8904 11704 8910 11756
rect 10226 11744 10232 11756
rect 9646 11716 10232 11744
rect 7282 11636 7288 11688
rect 7340 11636 7346 11688
rect 7837 11679 7895 11685
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8018 11676 8024 11688
rect 7883 11648 8024 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8018 11636 8024 11648
rect 8076 11636 8082 11688
rect 8386 11676 8392 11688
rect 8347 11648 8392 11676
rect 8386 11636 8392 11648
rect 8444 11636 8450 11688
rect 7300 11608 7328 11636
rect 7926 11608 7932 11620
rect 7300 11580 7932 11608
rect 7926 11568 7932 11580
rect 7984 11608 7990 11620
rect 9646 11608 9674 11716
rect 10226 11704 10232 11716
rect 10284 11704 10290 11756
rect 10336 11744 10364 11784
rect 10410 11772 10416 11824
rect 10468 11812 10474 11824
rect 10980 11812 11008 11852
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11514 11880 11520 11892
rect 11379 11852 11520 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11514 11840 11520 11852
rect 11572 11880 11578 11892
rect 11974 11880 11980 11892
rect 11572 11852 11980 11880
rect 11572 11840 11578 11852
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 14918 11880 14924 11892
rect 12084 11852 13032 11880
rect 12084 11812 12112 11852
rect 10468 11784 10916 11812
rect 10980 11784 12112 11812
rect 12437 11815 12495 11821
rect 10468 11772 10474 11784
rect 10888 11753 10916 11784
rect 12437 11781 12449 11815
rect 12483 11812 12495 11815
rect 12894 11812 12900 11824
rect 12483 11784 12900 11812
rect 12483 11781 12495 11784
rect 12437 11775 12495 11781
rect 12894 11772 12900 11784
rect 12952 11772 12958 11824
rect 10606 11747 10664 11753
rect 10606 11744 10618 11747
rect 10336 11716 10618 11744
rect 10606 11713 10618 11716
rect 10652 11744 10664 11747
rect 10873 11747 10931 11753
rect 10652 11716 10824 11744
rect 10652 11713 10664 11716
rect 10606 11707 10664 11713
rect 10796 11676 10824 11716
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 11054 11704 11060 11756
rect 11112 11744 11118 11756
rect 11793 11747 11851 11753
rect 11793 11744 11805 11747
rect 11112 11716 11805 11744
rect 11112 11704 11118 11716
rect 11793 11713 11805 11716
rect 11839 11713 11851 11747
rect 11974 11744 11980 11756
rect 11935 11716 11980 11744
rect 11793 11707 11851 11713
rect 11974 11704 11980 11716
rect 12032 11704 12038 11756
rect 12526 11744 12532 11756
rect 12487 11716 12532 11744
rect 12526 11704 12532 11716
rect 12584 11704 12590 11756
rect 13004 11753 13032 11852
rect 13740 11852 14320 11880
rect 12989 11747 13047 11753
rect 12989 11713 13001 11747
rect 13035 11713 13047 11747
rect 12989 11707 13047 11713
rect 13265 11747 13323 11753
rect 13265 11713 13277 11747
rect 13311 11744 13323 11747
rect 13630 11744 13636 11756
rect 13311 11716 13636 11744
rect 13311 11713 13323 11716
rect 13265 11707 13323 11713
rect 13630 11704 13636 11716
rect 13688 11704 13694 11756
rect 13740 11753 13768 11852
rect 13998 11772 14004 11824
rect 14056 11812 14062 11824
rect 14056 11784 14228 11812
rect 14056 11772 14062 11784
rect 14200 11753 14228 11784
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 14105 11747 14163 11753
rect 14105 11740 14117 11747
rect 13725 11707 13783 11713
rect 14090 11688 14096 11740
rect 14151 11713 14163 11747
rect 14148 11707 14163 11713
rect 14191 11747 14249 11753
rect 14191 11713 14203 11747
rect 14237 11713 14249 11747
rect 14292 11744 14320 11852
rect 14568 11852 14924 11880
rect 14568 11824 14596 11852
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 16114 11880 16120 11892
rect 15344 11852 16120 11880
rect 15344 11840 15350 11852
rect 16114 11840 16120 11852
rect 16172 11840 16178 11892
rect 16206 11840 16212 11892
rect 16264 11880 16270 11892
rect 17405 11883 17463 11889
rect 17405 11880 17417 11883
rect 16264 11852 17417 11880
rect 16264 11840 16270 11852
rect 17405 11849 17417 11852
rect 17451 11849 17463 11883
rect 17405 11843 17463 11849
rect 14550 11772 14556 11824
rect 14608 11772 14614 11824
rect 14737 11815 14795 11821
rect 14737 11781 14749 11815
rect 14783 11812 14795 11815
rect 15102 11812 15108 11824
rect 14783 11784 15108 11812
rect 14783 11781 14795 11784
rect 14737 11775 14795 11781
rect 15102 11772 15108 11784
rect 15160 11772 15166 11824
rect 15746 11772 15752 11824
rect 15804 11812 15810 11824
rect 19242 11812 19248 11824
rect 15804 11784 19248 11812
rect 15804 11772 15810 11784
rect 19242 11772 19248 11784
rect 19300 11772 19306 11824
rect 14642 11744 14648 11756
rect 14292 11716 14648 11744
rect 14191 11707 14249 11713
rect 14148 11688 14154 11707
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 14918 11744 14924 11756
rect 14879 11716 14924 11744
rect 14918 11704 14924 11716
rect 14976 11704 14982 11756
rect 16298 11744 16304 11756
rect 16259 11716 16304 11744
rect 16298 11704 16304 11716
rect 16356 11704 16362 11756
rect 16669 11747 16727 11753
rect 16669 11713 16681 11747
rect 16715 11713 16727 11747
rect 16669 11707 16727 11713
rect 17589 11747 17647 11753
rect 17589 11713 17601 11747
rect 17635 11744 17647 11747
rect 18322 11744 18328 11756
rect 17635 11716 18328 11744
rect 17635 11713 17647 11716
rect 17589 11707 17647 11713
rect 11330 11676 11336 11688
rect 10796 11648 11336 11676
rect 11330 11636 11336 11648
rect 11388 11636 11394 11688
rect 11514 11676 11520 11688
rect 11475 11648 11520 11676
rect 11514 11636 11520 11648
rect 11572 11636 11578 11688
rect 12644 11648 14044 11676
rect 7984 11580 9674 11608
rect 11149 11611 11207 11617
rect 7984 11568 7990 11580
rect 11149 11577 11161 11611
rect 11195 11608 11207 11611
rect 12644 11608 12672 11648
rect 12802 11608 12808 11620
rect 11195 11580 12672 11608
rect 12763 11580 12808 11608
rect 11195 11577 11207 11580
rect 11149 11571 11207 11577
rect 12802 11568 12808 11580
rect 12860 11568 12866 11620
rect 13078 11608 13084 11620
rect 13039 11580 13084 11608
rect 13078 11568 13084 11580
rect 13136 11568 13142 11620
rect 14016 11608 14044 11648
rect 16114 11636 16120 11688
rect 16172 11676 16178 11688
rect 16684 11676 16712 11707
rect 18322 11704 18328 11716
rect 18380 11704 18386 11756
rect 17678 11676 17684 11688
rect 16172 11648 16712 11676
rect 16767 11648 17684 11676
rect 16172 11636 16178 11648
rect 16767 11608 16795 11648
rect 17678 11636 17684 11648
rect 17736 11685 17742 11688
rect 17736 11679 17785 11685
rect 17736 11645 17739 11679
rect 17773 11645 17785 11679
rect 17954 11676 17960 11688
rect 17915 11648 17960 11676
rect 17736 11639 17785 11645
rect 17736 11636 17742 11639
rect 17954 11636 17960 11648
rect 18012 11636 18018 11688
rect 14016 11580 16795 11608
rect 7282 11540 7288 11552
rect 6748 11512 7144 11540
rect 7243 11512 7288 11540
rect 7282 11500 7288 11512
rect 7340 11500 7346 11552
rect 8297 11543 8355 11549
rect 8297 11509 8309 11543
rect 8343 11540 8355 11543
rect 9030 11540 9036 11552
rect 8343 11512 9036 11540
rect 8343 11509 8355 11512
rect 8297 11503 8355 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 9398 11540 9404 11552
rect 9359 11512 9404 11540
rect 9398 11500 9404 11512
rect 9456 11500 9462 11552
rect 9493 11543 9551 11549
rect 9493 11509 9505 11543
rect 9539 11540 9551 11543
rect 10226 11540 10232 11552
rect 9539 11512 10232 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 10226 11500 10232 11512
rect 10284 11500 10290 11552
rect 11882 11500 11888 11552
rect 11940 11540 11946 11552
rect 12161 11543 12219 11549
rect 12161 11540 12173 11543
rect 11940 11512 12173 11540
rect 11940 11500 11946 11512
rect 12161 11509 12173 11512
rect 12207 11509 12219 11543
rect 12710 11540 12716 11552
rect 12671 11512 12716 11540
rect 12161 11503 12219 11509
rect 12710 11500 12716 11512
rect 12768 11500 12774 11552
rect 13541 11543 13599 11549
rect 13541 11509 13553 11543
rect 13587 11540 13599 11543
rect 13630 11540 13636 11552
rect 13587 11512 13636 11540
rect 13587 11509 13599 11512
rect 13541 11503 13599 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13814 11500 13820 11552
rect 13872 11540 13878 11552
rect 13909 11543 13967 11549
rect 13909 11540 13921 11543
rect 13872 11512 13921 11540
rect 13872 11500 13878 11512
rect 13909 11509 13921 11512
rect 13955 11509 13967 11543
rect 14366 11540 14372 11552
rect 14327 11512 14372 11540
rect 13909 11503 13967 11509
rect 14366 11500 14372 11512
rect 14424 11500 14430 11552
rect 14642 11540 14648 11552
rect 14603 11512 14648 11540
rect 14642 11500 14648 11512
rect 14700 11500 14706 11552
rect 15562 11540 15568 11552
rect 15523 11512 15568 11540
rect 15562 11500 15568 11512
rect 15620 11500 15626 11552
rect 15654 11500 15660 11552
rect 15712 11540 15718 11552
rect 15712 11512 15757 11540
rect 15712 11500 15718 11512
rect 16022 11500 16028 11552
rect 16080 11540 16086 11552
rect 16393 11543 16451 11549
rect 16393 11540 16405 11543
rect 16080 11512 16405 11540
rect 16080 11500 16086 11512
rect 16393 11509 16405 11512
rect 16439 11509 16451 11543
rect 16393 11503 16451 11509
rect 17126 11500 17132 11552
rect 17184 11540 17190 11552
rect 17313 11543 17371 11549
rect 17313 11540 17325 11543
rect 17184 11512 17325 11540
rect 17184 11500 17190 11512
rect 17313 11509 17325 11512
rect 17359 11509 17371 11543
rect 17313 11503 17371 11509
rect 1104 11450 18860 11472
rect 1104 11398 3174 11450
rect 3226 11398 3238 11450
rect 3290 11398 3302 11450
rect 3354 11398 3366 11450
rect 3418 11398 3430 11450
rect 3482 11398 7622 11450
rect 7674 11398 7686 11450
rect 7738 11398 7750 11450
rect 7802 11398 7814 11450
rect 7866 11398 7878 11450
rect 7930 11398 12070 11450
rect 12122 11398 12134 11450
rect 12186 11398 12198 11450
rect 12250 11398 12262 11450
rect 12314 11398 12326 11450
rect 12378 11398 16518 11450
rect 16570 11398 16582 11450
rect 16634 11398 16646 11450
rect 16698 11398 16710 11450
rect 16762 11398 16774 11450
rect 16826 11398 18860 11450
rect 1104 11376 18860 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2682 11336 2688 11348
rect 2179 11308 2688 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 5644 11308 7052 11336
rect 2038 11228 2044 11280
rect 2096 11268 2102 11280
rect 2225 11271 2283 11277
rect 2225 11268 2237 11271
rect 2096 11240 2237 11268
rect 2096 11228 2102 11240
rect 2225 11237 2237 11240
rect 2271 11268 2283 11271
rect 2406 11268 2412 11280
rect 2271 11240 2412 11268
rect 2271 11237 2283 11240
rect 2225 11231 2283 11237
rect 2406 11228 2412 11240
rect 2464 11228 2470 11280
rect 4264 11240 4568 11268
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11169 1639 11203
rect 1581 11163 1639 11169
rect 1596 11064 1624 11163
rect 1670 11160 1676 11212
rect 1728 11200 1734 11212
rect 1728 11172 1773 11200
rect 1728 11160 1734 11172
rect 3786 11160 3792 11212
rect 3844 11200 3850 11212
rect 4154 11200 4160 11212
rect 3844 11172 4160 11200
rect 3844 11160 3850 11172
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 4264 11209 4292 11240
rect 4540 11212 4568 11240
rect 4249 11203 4307 11209
rect 4249 11169 4261 11203
rect 4295 11169 4307 11203
rect 4430 11200 4436 11212
rect 4391 11172 4436 11200
rect 4249 11163 4307 11169
rect 4430 11160 4436 11172
rect 4488 11160 4494 11212
rect 4522 11160 4528 11212
rect 4580 11160 4586 11212
rect 1762 11132 1768 11144
rect 1723 11104 1768 11132
rect 1762 11092 1768 11104
rect 1820 11092 1826 11144
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 2924 11104 3617 11132
rect 2924 11092 2930 11104
rect 3605 11101 3617 11104
rect 3651 11132 3663 11135
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 3651 11104 4629 11132
rect 3651 11101 3663 11104
rect 3605 11095 3663 11101
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 2130 11064 2136 11076
rect 1596 11036 2136 11064
rect 2130 11024 2136 11036
rect 2188 11064 2194 11076
rect 3360 11067 3418 11073
rect 3360 11064 3372 11067
rect 2188 11036 3372 11064
rect 2188 11024 2194 11036
rect 3360 11033 3372 11036
rect 3406 11064 3418 11067
rect 4430 11064 4436 11076
rect 3406 11036 4436 11064
rect 3406 11033 3418 11036
rect 3360 11027 3418 11033
rect 4430 11024 4436 11036
rect 4488 11024 4494 11076
rect 4884 11067 4942 11073
rect 4884 11033 4896 11067
rect 4930 11064 4942 11067
rect 5074 11064 5080 11076
rect 4930 11036 5080 11064
rect 4930 11033 4942 11036
rect 4884 11027 4942 11033
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 2498 10956 2504 11008
rect 2556 10996 2562 11008
rect 3142 10996 3148 11008
rect 2556 10968 3148 10996
rect 2556 10956 2562 10968
rect 3142 10956 3148 10968
rect 3200 10996 3206 11008
rect 4157 10999 4215 11005
rect 4157 10996 4169 10999
rect 3200 10968 4169 10996
rect 3200 10956 3206 10968
rect 4157 10965 4169 10968
rect 4203 10996 4215 10999
rect 5644 10996 5672 11308
rect 7024 11268 7052 11308
rect 9306 11296 9312 11348
rect 9364 11336 9370 11348
rect 10413 11339 10471 11345
rect 10413 11336 10425 11339
rect 9364 11308 10425 11336
rect 9364 11296 9370 11308
rect 10413 11305 10425 11308
rect 10459 11305 10471 11339
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 10413 11299 10471 11305
rect 10520 11308 12449 11336
rect 8938 11268 8944 11280
rect 7024 11240 8944 11268
rect 8938 11228 8944 11240
rect 8996 11228 9002 11280
rect 8018 11160 8024 11212
rect 8076 11200 8082 11212
rect 8113 11203 8171 11209
rect 8113 11200 8125 11203
rect 8076 11172 8125 11200
rect 8076 11160 8082 11172
rect 8113 11169 8125 11172
rect 8159 11169 8171 11203
rect 8113 11163 8171 11169
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 10410 11200 10416 11212
rect 10367 11172 10416 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 10410 11160 10416 11172
rect 10468 11160 10474 11212
rect 6086 11132 6092 11144
rect 6047 11104 6092 11132
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 7929 11135 7987 11141
rect 7929 11101 7941 11135
rect 7975 11132 7987 11135
rect 8386 11132 8392 11144
rect 7975 11104 8392 11132
rect 7975 11101 7987 11104
rect 7929 11095 7987 11101
rect 8386 11092 8392 11104
rect 8444 11092 8450 11144
rect 8478 11092 8484 11144
rect 8536 11132 8542 11144
rect 8757 11135 8815 11141
rect 8757 11132 8769 11135
rect 8536 11104 8769 11132
rect 8536 11092 8542 11104
rect 8757 11101 8769 11104
rect 8803 11101 8815 11135
rect 8757 11095 8815 11101
rect 8938 11092 8944 11144
rect 8996 11132 9002 11144
rect 10520 11132 10548 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 12437 11299 12495 11305
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 13630 11336 13636 11348
rect 12860 11308 13636 11336
rect 12860 11296 12866 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 13998 11336 14004 11348
rect 13832 11308 14004 11336
rect 10686 11228 10692 11280
rect 10744 11268 10750 11280
rect 11609 11271 11667 11277
rect 11609 11268 11621 11271
rect 10744 11240 11621 11268
rect 10744 11228 10750 11240
rect 11609 11237 11621 11240
rect 11655 11237 11667 11271
rect 11609 11231 11667 11237
rect 13170 11228 13176 11280
rect 13228 11268 13234 11280
rect 13725 11271 13783 11277
rect 13725 11268 13737 11271
rect 13228 11240 13737 11268
rect 13228 11228 13234 11240
rect 13725 11237 13737 11240
rect 13771 11237 13783 11271
rect 13725 11231 13783 11237
rect 10962 11160 10968 11212
rect 11020 11200 11026 11212
rect 11241 11203 11299 11209
rect 11241 11200 11253 11203
rect 11020 11172 11253 11200
rect 11020 11160 11026 11172
rect 11241 11169 11253 11172
rect 11287 11169 11299 11203
rect 11241 11163 11299 11169
rect 11330 11160 11336 11212
rect 11388 11200 11394 11212
rect 12161 11203 12219 11209
rect 12161 11200 12173 11203
rect 11388 11172 12173 11200
rect 11388 11160 11394 11172
rect 12161 11169 12173 11172
rect 12207 11169 12219 11203
rect 12161 11163 12219 11169
rect 12250 11160 12256 11212
rect 12308 11200 12314 11212
rect 12805 11203 12863 11209
rect 12805 11200 12817 11203
rect 12308 11172 12817 11200
rect 12308 11160 12314 11172
rect 12805 11169 12817 11172
rect 12851 11200 12863 11203
rect 13832 11200 13860 11308
rect 13998 11296 14004 11308
rect 14056 11296 14062 11348
rect 15010 11336 15016 11348
rect 14108 11308 15016 11336
rect 14108 11200 14136 11308
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15473 11339 15531 11345
rect 15473 11305 15485 11339
rect 15519 11336 15531 11339
rect 15838 11336 15844 11348
rect 15519 11308 15844 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 15838 11296 15844 11308
rect 15896 11336 15902 11348
rect 16298 11336 16304 11348
rect 15896 11308 16304 11336
rect 15896 11296 15902 11308
rect 16298 11296 16304 11308
rect 16356 11296 16362 11348
rect 12851 11172 13860 11200
rect 13924 11172 14136 11200
rect 12851 11169 12863 11172
rect 12805 11163 12863 11169
rect 8996 11104 10548 11132
rect 11149 11135 11207 11141
rect 10597 11111 10655 11117
rect 8996 11092 9002 11104
rect 10597 11077 10609 11111
rect 10643 11077 10655 11111
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11514 11132 11520 11144
rect 11195 11128 11376 11132
rect 11440 11128 11520 11132
rect 11195 11104 11520 11128
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11348 11100 11468 11104
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12621 11135 12679 11141
rect 12621 11132 12633 11135
rect 12492 11104 12633 11132
rect 12492 11092 12498 11104
rect 12621 11101 12633 11104
rect 12667 11101 12679 11135
rect 12894 11132 12900 11144
rect 12855 11104 12900 11132
rect 12621 11095 12679 11101
rect 6178 11024 6184 11076
rect 6236 11064 6242 11076
rect 6334 11067 6392 11073
rect 6334 11064 6346 11067
rect 6236 11036 6346 11064
rect 6236 11024 6242 11036
rect 6334 11033 6346 11036
rect 6380 11033 6392 11067
rect 6334 11027 6392 11033
rect 6638 11024 6644 11076
rect 6696 11064 6702 11076
rect 8021 11067 8079 11073
rect 8021 11064 8033 11067
rect 6696 11036 8033 11064
rect 6696 11024 6702 11036
rect 8021 11033 8033 11036
rect 8067 11033 8079 11067
rect 8021 11027 8079 11033
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 9674 11064 9680 11076
rect 8168 11036 9680 11064
rect 8168 11024 8174 11036
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 10076 11067 10134 11073
rect 10076 11033 10088 11067
rect 10122 11064 10134 11067
rect 10226 11064 10232 11076
rect 10122 11036 10232 11064
rect 10122 11033 10134 11036
rect 10076 11027 10134 11033
rect 10226 11024 10232 11036
rect 10284 11024 10290 11076
rect 10597 11071 10655 11077
rect 10612 11008 10640 11071
rect 11054 11024 11060 11076
rect 11112 11064 11118 11076
rect 11977 11067 12035 11073
rect 11977 11064 11989 11067
rect 11112 11036 11192 11064
rect 11112 11024 11118 11036
rect 4203 10968 5672 10996
rect 5997 10999 6055 11005
rect 4203 10965 4215 10968
rect 4157 10959 4215 10965
rect 5997 10965 6009 10999
rect 6043 10996 6055 10999
rect 6822 10996 6828 11008
rect 6043 10968 6828 10996
rect 6043 10965 6055 10968
rect 5997 10959 6055 10965
rect 6822 10956 6828 10968
rect 6880 10956 6886 11008
rect 7466 10996 7472 11008
rect 7427 10968 7472 10996
rect 7466 10956 7472 10968
rect 7524 10956 7530 11008
rect 7558 10956 7564 11008
rect 7616 10996 7622 11008
rect 8386 10996 8392 11008
rect 7616 10968 7661 10996
rect 8347 10968 8392 10996
rect 7616 10956 7622 10968
rect 8386 10956 8392 10968
rect 8444 10956 8450 11008
rect 8570 10996 8576 11008
rect 8531 10968 8576 10996
rect 8570 10956 8576 10968
rect 8628 10956 8634 11008
rect 8846 10956 8852 11008
rect 8904 10996 8910 11008
rect 8941 10999 8999 11005
rect 8941 10996 8953 10999
rect 8904 10968 8953 10996
rect 8904 10956 8910 10968
rect 8941 10965 8953 10968
rect 8987 10965 8999 10999
rect 8941 10959 8999 10965
rect 10594 10956 10600 11008
rect 10652 10956 10658 11008
rect 10778 10996 10784 11008
rect 10739 10968 10784 10996
rect 10778 10956 10784 10968
rect 10836 10956 10842 11008
rect 11164 10996 11192 11036
rect 11900 11036 11989 11064
rect 11900 10996 11928 11036
rect 11977 11033 11989 11036
rect 12023 11033 12035 11067
rect 11977 11027 12035 11033
rect 12069 11067 12127 11073
rect 12069 11033 12081 11067
rect 12115 11064 12127 11067
rect 12636 11064 12664 11095
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13078 11092 13084 11144
rect 13136 11132 13142 11144
rect 13446 11132 13452 11144
rect 13136 11104 13452 11132
rect 13136 11092 13142 11104
rect 13446 11092 13452 11104
rect 13504 11092 13510 11144
rect 13924 11141 13952 11172
rect 13909 11135 13967 11141
rect 13909 11101 13921 11135
rect 13955 11101 13967 11135
rect 13909 11095 13967 11101
rect 14093 11135 14151 11141
rect 14093 11101 14105 11135
rect 14139 11132 14151 11135
rect 15565 11135 15623 11141
rect 15565 11132 15577 11135
rect 14139 11104 15577 11132
rect 14139 11101 14151 11104
rect 14093 11095 14151 11101
rect 15565 11101 15577 11104
rect 15611 11132 15623 11135
rect 16206 11132 16212 11144
rect 15611 11104 16212 11132
rect 15611 11101 15623 11104
rect 15565 11095 15623 11101
rect 16206 11092 16212 11104
rect 16264 11132 16270 11144
rect 17037 11135 17095 11141
rect 17037 11132 17049 11135
rect 16264 11104 17049 11132
rect 16264 11092 16270 11104
rect 17037 11101 17049 11104
rect 17083 11101 17095 11135
rect 17037 11095 17095 11101
rect 12986 11064 12992 11076
rect 12115 11036 12572 11064
rect 12636 11036 12992 11064
rect 12115 11033 12127 11036
rect 12069 11027 12127 11033
rect 12158 10996 12164 11008
rect 11164 10968 12164 10996
rect 12158 10956 12164 10968
rect 12216 10956 12222 11008
rect 12544 10996 12572 11036
rect 12986 11024 12992 11036
rect 13044 11024 13050 11076
rect 13538 11064 13544 11076
rect 13499 11036 13544 11064
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 13998 11024 14004 11076
rect 14056 11064 14062 11076
rect 14338 11067 14396 11073
rect 14338 11064 14350 11067
rect 14056 11036 14350 11064
rect 14056 11024 14062 11036
rect 14338 11033 14350 11036
rect 14384 11033 14396 11067
rect 14338 11027 14396 11033
rect 14550 11024 14556 11076
rect 14608 11064 14614 11076
rect 15010 11064 15016 11076
rect 14608 11036 15016 11064
rect 14608 11024 14614 11036
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 15654 11024 15660 11076
rect 15712 11064 15718 11076
rect 15810 11067 15868 11073
rect 15810 11064 15822 11067
rect 15712 11036 15822 11064
rect 15712 11024 15718 11036
rect 15810 11033 15822 11036
rect 15856 11033 15868 11067
rect 15810 11027 15868 11033
rect 17304 11067 17362 11073
rect 17304 11033 17316 11067
rect 17350 11033 17362 11067
rect 17304 11027 17362 11033
rect 12618 10996 12624 11008
rect 12544 10968 12624 10996
rect 12618 10956 12624 10968
rect 12676 10996 12682 11008
rect 15378 10996 15384 11008
rect 12676 10968 15384 10996
rect 12676 10956 12682 10968
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 16945 10999 17003 11005
rect 16945 10965 16957 10999
rect 16991 10996 17003 10999
rect 17328 10996 17356 11027
rect 17678 10996 17684 11008
rect 16991 10968 17684 10996
rect 16991 10965 17003 10968
rect 16945 10959 17003 10965
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 17954 10956 17960 11008
rect 18012 10996 18018 11008
rect 18417 10999 18475 11005
rect 18417 10996 18429 10999
rect 18012 10968 18429 10996
rect 18012 10956 18018 10968
rect 18417 10965 18429 10968
rect 18463 10965 18475 10999
rect 18417 10959 18475 10965
rect 1104 10906 18860 10928
rect 1104 10854 5398 10906
rect 5450 10854 5462 10906
rect 5514 10854 5526 10906
rect 5578 10854 5590 10906
rect 5642 10854 5654 10906
rect 5706 10854 9846 10906
rect 9898 10854 9910 10906
rect 9962 10854 9974 10906
rect 10026 10854 10038 10906
rect 10090 10854 10102 10906
rect 10154 10854 14294 10906
rect 14346 10854 14358 10906
rect 14410 10854 14422 10906
rect 14474 10854 14486 10906
rect 14538 10854 14550 10906
rect 14602 10854 18860 10906
rect 1104 10832 18860 10854
rect 1394 10792 1400 10804
rect 1355 10764 1400 10792
rect 1394 10752 1400 10764
rect 1452 10752 1458 10804
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 2038 10792 2044 10804
rect 1636 10764 2044 10792
rect 1636 10752 1642 10764
rect 2038 10752 2044 10764
rect 2096 10792 2102 10804
rect 3513 10795 3571 10801
rect 3513 10792 3525 10795
rect 2096 10764 3525 10792
rect 2096 10752 2102 10764
rect 3513 10761 3525 10764
rect 3559 10761 3571 10795
rect 3513 10755 3571 10761
rect 3605 10795 3663 10801
rect 3605 10761 3617 10795
rect 3651 10792 3663 10795
rect 3786 10792 3792 10804
rect 3651 10764 3792 10792
rect 3651 10761 3663 10764
rect 3605 10755 3663 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 3973 10795 4031 10801
rect 3973 10761 3985 10795
rect 4019 10792 4031 10795
rect 4522 10792 4528 10804
rect 4019 10764 4528 10792
rect 4019 10761 4031 10764
rect 3973 10755 4031 10761
rect 4522 10752 4528 10764
rect 4580 10752 4586 10804
rect 6178 10792 6184 10804
rect 6139 10764 6184 10792
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 7282 10792 7288 10804
rect 7243 10764 7288 10792
rect 7282 10752 7288 10764
rect 7340 10752 7346 10804
rect 8205 10795 8263 10801
rect 8205 10761 8217 10795
rect 8251 10792 8263 10795
rect 8573 10795 8631 10801
rect 8573 10792 8585 10795
rect 8251 10764 8585 10792
rect 8251 10761 8263 10764
rect 8205 10755 8263 10761
rect 8573 10761 8585 10764
rect 8619 10761 8631 10795
rect 8573 10755 8631 10761
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9401 10795 9459 10801
rect 9401 10792 9413 10795
rect 9079 10764 9413 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9401 10761 9413 10764
rect 9447 10761 9459 10795
rect 9401 10755 9459 10761
rect 9490 10752 9496 10804
rect 9548 10792 9554 10804
rect 9769 10795 9827 10801
rect 9769 10792 9781 10795
rect 9548 10764 9781 10792
rect 9548 10752 9554 10764
rect 9769 10761 9781 10764
rect 9815 10761 9827 10795
rect 9769 10755 9827 10761
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10761 10287 10795
rect 10229 10755 10287 10761
rect 10597 10795 10655 10801
rect 10597 10761 10609 10795
rect 10643 10792 10655 10795
rect 10778 10792 10784 10804
rect 10643 10764 10784 10792
rect 10643 10761 10655 10764
rect 10597 10755 10655 10761
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 2510 10727 2568 10733
rect 2510 10724 2522 10727
rect 2464 10696 2522 10724
rect 2464 10684 2470 10696
rect 2510 10693 2522 10696
rect 2556 10693 2568 10727
rect 2958 10724 2964 10736
rect 2919 10696 2964 10724
rect 2510 10687 2568 10693
rect 2958 10684 2964 10696
rect 3016 10684 3022 10736
rect 4982 10724 4988 10736
rect 3436 10696 4988 10724
rect 2777 10591 2835 10597
rect 2777 10557 2789 10591
rect 2823 10588 2835 10591
rect 2866 10588 2872 10600
rect 2823 10560 2872 10588
rect 2823 10557 2835 10560
rect 2777 10551 2835 10557
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 3436 10597 3464 10696
rect 4982 10684 4988 10696
rect 5040 10724 5046 10736
rect 5178 10727 5236 10733
rect 5178 10724 5190 10727
rect 5040 10696 5190 10724
rect 5040 10684 5046 10696
rect 5178 10693 5190 10696
rect 5224 10693 5236 10727
rect 5178 10687 5236 10693
rect 5902 10684 5908 10736
rect 5960 10724 5966 10736
rect 7193 10727 7251 10733
rect 5960 10696 6408 10724
rect 5960 10684 5966 10696
rect 6380 10665 6408 10696
rect 7193 10693 7205 10727
rect 7239 10724 7251 10727
rect 7558 10724 7564 10736
rect 7239 10696 7564 10724
rect 7239 10693 7251 10696
rect 7193 10687 7251 10693
rect 7558 10684 7564 10696
rect 7616 10684 7622 10736
rect 8113 10727 8171 10733
rect 8113 10693 8125 10727
rect 8159 10724 8171 10727
rect 10244 10724 10272 10755
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 12710 10752 12716 10804
rect 12768 10792 12774 10804
rect 12986 10792 12992 10804
rect 12768 10764 12992 10792
rect 12768 10752 12774 10764
rect 12986 10752 12992 10764
rect 13044 10752 13050 10804
rect 13449 10795 13507 10801
rect 13449 10761 13461 10795
rect 13495 10792 13507 10795
rect 14182 10792 14188 10804
rect 13495 10764 14188 10792
rect 13495 10761 13507 10764
rect 13449 10755 13507 10761
rect 14182 10752 14188 10764
rect 14240 10752 14246 10804
rect 17405 10795 17463 10801
rect 17405 10761 17417 10795
rect 17451 10792 17463 10795
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17451 10764 17785 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 18138 10752 18144 10804
rect 18196 10792 18202 10804
rect 18196 10764 18276 10792
rect 18196 10752 18202 10764
rect 10686 10724 10692 10736
rect 8159 10696 10272 10724
rect 10647 10696 10692 10724
rect 8159 10693 8171 10696
rect 8113 10687 8171 10693
rect 10686 10684 10692 10696
rect 10744 10684 10750 10736
rect 11241 10727 11299 10733
rect 11241 10693 11253 10727
rect 11287 10724 11299 10727
rect 14642 10724 14648 10736
rect 11287 10696 14648 10724
rect 11287 10693 11299 10696
rect 11241 10687 11299 10693
rect 5537 10659 5595 10665
rect 5537 10625 5549 10659
rect 5583 10656 5595 10659
rect 6365 10659 6423 10665
rect 5583 10628 6316 10656
rect 5583 10625 5595 10628
rect 5537 10619 5595 10625
rect 3421 10591 3479 10597
rect 3421 10557 3433 10591
rect 3467 10557 3479 10591
rect 3421 10551 3479 10557
rect 5445 10591 5503 10597
rect 5445 10557 5457 10591
rect 5491 10588 5503 10591
rect 5718 10588 5724 10600
rect 5491 10560 5724 10588
rect 5491 10557 5503 10560
rect 5445 10551 5503 10557
rect 5718 10548 5724 10560
rect 5776 10588 5782 10600
rect 6086 10588 6092 10600
rect 5776 10560 6092 10588
rect 5776 10548 5782 10560
rect 6086 10548 6092 10560
rect 6144 10548 6150 10600
rect 6288 10588 6316 10628
rect 6365 10625 6377 10659
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6546 10616 6552 10668
rect 6604 10656 6610 10668
rect 6914 10656 6920 10668
rect 6604 10628 6920 10656
rect 6604 10616 6610 10628
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 8754 10616 8760 10668
rect 8812 10656 8818 10668
rect 8941 10659 8999 10665
rect 8941 10656 8953 10659
rect 8812 10628 8953 10656
rect 8812 10616 8818 10628
rect 8941 10625 8953 10628
rect 8987 10625 8999 10659
rect 8941 10619 8999 10625
rect 9122 10616 9128 10668
rect 9180 10656 9186 10668
rect 9180 10628 9996 10656
rect 9180 10616 9186 10628
rect 6822 10588 6828 10600
rect 6288 10560 6828 10588
rect 6822 10548 6828 10560
rect 6880 10588 6886 10600
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 6880 10560 7389 10588
rect 6880 10548 6886 10560
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 8389 10591 8447 10597
rect 8389 10557 8401 10591
rect 8435 10588 8447 10591
rect 8846 10588 8852 10600
rect 8435 10560 8852 10588
rect 8435 10557 8447 10560
rect 8389 10551 8447 10557
rect 8846 10548 8852 10560
rect 8904 10548 8910 10600
rect 7190 10520 7196 10532
rect 2792 10492 4568 10520
rect 2792 10464 2820 10492
rect 2774 10412 2780 10464
rect 2832 10412 2838 10464
rect 3050 10452 3056 10464
rect 3011 10424 3056 10452
rect 3050 10412 3056 10424
rect 3108 10412 3114 10464
rect 4065 10455 4123 10461
rect 4065 10421 4077 10455
rect 4111 10452 4123 10455
rect 4430 10452 4436 10464
rect 4111 10424 4436 10452
rect 4111 10421 4123 10424
rect 4065 10415 4123 10421
rect 4430 10412 4436 10424
rect 4488 10412 4494 10464
rect 4540 10452 4568 10492
rect 5460 10492 7196 10520
rect 5460 10452 5488 10492
rect 7190 10480 7196 10492
rect 7248 10480 7254 10532
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 9140 10520 9168 10616
rect 9217 10591 9275 10597
rect 9217 10557 9229 10591
rect 9263 10557 9275 10591
rect 9217 10551 9275 10557
rect 8536 10492 9168 10520
rect 9232 10520 9260 10551
rect 9490 10548 9496 10600
rect 9548 10588 9554 10600
rect 9968 10597 9996 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 11256 10656 11284 10687
rect 14642 10684 14648 10696
rect 14700 10684 14706 10736
rect 14737 10727 14795 10733
rect 14737 10693 14749 10727
rect 14783 10724 14795 10727
rect 16390 10724 16396 10736
rect 14783 10696 16396 10724
rect 14783 10693 14795 10696
rect 14737 10687 14795 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 16850 10684 16856 10736
rect 16908 10724 16914 10736
rect 17586 10724 17592 10736
rect 16908 10696 17592 10724
rect 16908 10684 16914 10696
rect 17586 10684 17592 10696
rect 17644 10684 17650 10736
rect 11514 10656 11520 10668
rect 10192 10628 11284 10656
rect 11475 10628 11520 10656
rect 10192 10616 10198 10628
rect 11514 10616 11520 10628
rect 11572 10616 11578 10668
rect 12529 10659 12587 10665
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12897 10659 12955 10665
rect 12575 10628 12848 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 9861 10591 9919 10597
rect 9861 10588 9873 10591
rect 9548 10560 9873 10588
rect 9548 10548 9554 10560
rect 9861 10557 9873 10560
rect 9907 10557 9919 10591
rect 9861 10551 9919 10557
rect 9953 10591 10011 10597
rect 9953 10557 9965 10591
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10781 10591 10839 10597
rect 10781 10588 10793 10591
rect 10284 10560 10793 10588
rect 10284 10548 10290 10560
rect 10781 10557 10793 10560
rect 10827 10557 10839 10591
rect 10781 10551 10839 10557
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 11146 10588 11152 10600
rect 11020 10560 11152 10588
rect 11020 10548 11026 10560
rect 11146 10548 11152 10560
rect 11204 10548 11210 10600
rect 11698 10548 11704 10600
rect 11756 10588 11762 10600
rect 12820 10588 12848 10628
rect 12897 10625 12909 10659
rect 12943 10656 12955 10659
rect 13262 10656 13268 10668
rect 12943 10628 13268 10656
rect 12943 10625 12955 10628
rect 12897 10619 12955 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 15953 10659 16011 10665
rect 15953 10625 15965 10659
rect 15999 10656 16011 10659
rect 17310 10656 17316 10668
rect 15999 10628 17172 10656
rect 17271 10628 17316 10656
rect 15999 10625 16011 10628
rect 15953 10619 16011 10625
rect 13354 10588 13360 10600
rect 11756 10560 12756 10588
rect 12820 10560 13360 10588
rect 11756 10548 11762 10560
rect 10244 10520 10272 10548
rect 9232 10492 10272 10520
rect 8536 10480 8542 10492
rect 10502 10480 10508 10532
rect 10560 10520 10566 10532
rect 12158 10520 12164 10532
rect 10560 10492 11744 10520
rect 12119 10492 12164 10520
rect 10560 10480 10566 10492
rect 11716 10464 11744 10492
rect 12158 10480 12164 10492
rect 12216 10480 12222 10532
rect 12250 10480 12256 10532
rect 12308 10480 12314 10532
rect 12728 10520 12756 10560
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 14090 10548 14096 10600
rect 14148 10588 14154 10600
rect 15102 10588 15108 10600
rect 14148 10560 15108 10588
rect 14148 10548 14154 10560
rect 15102 10548 15108 10560
rect 15160 10548 15166 10600
rect 16206 10588 16212 10600
rect 16167 10560 16212 10588
rect 16206 10548 16212 10560
rect 16264 10548 16270 10600
rect 16298 10548 16304 10600
rect 16356 10588 16362 10600
rect 16850 10588 16856 10600
rect 16356 10560 16401 10588
rect 16811 10560 16856 10588
rect 16356 10548 16362 10560
rect 16850 10548 16856 10560
rect 16908 10548 16914 10600
rect 17144 10588 17172 10628
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 18138 10656 18144 10668
rect 18099 10628 18144 10656
rect 18138 10616 18144 10628
rect 18196 10616 18202 10668
rect 18248 10665 18276 10764
rect 18233 10659 18291 10665
rect 18233 10625 18245 10659
rect 18279 10656 18291 10659
rect 18782 10656 18788 10668
rect 18279 10628 18788 10656
rect 18279 10625 18291 10628
rect 18233 10619 18291 10625
rect 18782 10616 18788 10628
rect 18840 10616 18846 10668
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 17144 10560 17601 10588
rect 17589 10557 17601 10560
rect 17635 10588 17647 10591
rect 17954 10588 17960 10600
rect 17635 10560 17960 10588
rect 17635 10557 17647 10560
rect 17589 10551 17647 10557
rect 17954 10548 17960 10560
rect 18012 10548 18018 10600
rect 18325 10591 18383 10597
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 18325 10551 18383 10557
rect 17494 10520 17500 10532
rect 12728 10492 14964 10520
rect 4540 10424 5488 10452
rect 5534 10412 5540 10464
rect 5592 10452 5598 10464
rect 6549 10455 6607 10461
rect 6549 10452 6561 10455
rect 5592 10424 6561 10452
rect 5592 10412 5598 10424
rect 6549 10421 6561 10424
rect 6595 10421 6607 10455
rect 6822 10452 6828 10464
rect 6783 10424 6828 10452
rect 6549 10415 6607 10421
rect 6822 10412 6828 10424
rect 6880 10412 6886 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7745 10455 7803 10461
rect 7745 10452 7757 10455
rect 6972 10424 7757 10452
rect 6972 10412 6978 10424
rect 7745 10421 7757 10424
rect 7791 10421 7803 10455
rect 7745 10415 7803 10421
rect 8110 10412 8116 10464
rect 8168 10452 8174 10464
rect 10042 10452 10048 10464
rect 8168 10424 10048 10452
rect 8168 10412 8174 10424
rect 10042 10412 10048 10424
rect 10100 10412 10106 10464
rect 10686 10412 10692 10464
rect 10744 10452 10750 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 10744 10424 11161 10452
rect 10744 10412 10750 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 11698 10412 11704 10464
rect 11756 10452 11762 10464
rect 12268 10452 12296 10480
rect 11756 10424 12296 10452
rect 12345 10455 12403 10461
rect 11756 10412 11762 10424
rect 12345 10421 12357 10455
rect 12391 10452 12403 10455
rect 12618 10452 12624 10464
rect 12391 10424 12624 10452
rect 12391 10421 12403 10424
rect 12345 10415 12403 10421
rect 12618 10412 12624 10424
rect 12676 10412 12682 10464
rect 12713 10455 12771 10461
rect 12713 10421 12725 10455
rect 12759 10452 12771 10455
rect 13170 10452 13176 10464
rect 12759 10424 13176 10452
rect 12759 10421 12771 10424
rect 12713 10415 12771 10421
rect 13170 10412 13176 10424
rect 13228 10412 13234 10464
rect 14826 10452 14832 10464
rect 14787 10424 14832 10452
rect 14826 10412 14832 10424
rect 14884 10412 14890 10464
rect 14936 10452 14964 10492
rect 16224 10492 17500 10520
rect 16224 10452 16252 10492
rect 17494 10480 17500 10492
rect 17552 10480 17558 10532
rect 17678 10480 17684 10532
rect 17736 10520 17742 10532
rect 18340 10520 18368 10551
rect 17736 10492 18368 10520
rect 17736 10480 17742 10492
rect 18506 10480 18512 10532
rect 18564 10520 18570 10532
rect 19702 10520 19708 10532
rect 18564 10492 19708 10520
rect 18564 10480 18570 10492
rect 19702 10480 19708 10492
rect 19760 10480 19766 10532
rect 16942 10452 16948 10464
rect 14936 10424 16252 10452
rect 16903 10424 16948 10452
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 1104 10362 18860 10384
rect 1104 10310 3174 10362
rect 3226 10310 3238 10362
rect 3290 10310 3302 10362
rect 3354 10310 3366 10362
rect 3418 10310 3430 10362
rect 3482 10310 7622 10362
rect 7674 10310 7686 10362
rect 7738 10310 7750 10362
rect 7802 10310 7814 10362
rect 7866 10310 7878 10362
rect 7930 10310 12070 10362
rect 12122 10310 12134 10362
rect 12186 10310 12198 10362
rect 12250 10310 12262 10362
rect 12314 10310 12326 10362
rect 12378 10310 16518 10362
rect 16570 10310 16582 10362
rect 16634 10310 16646 10362
rect 16698 10310 16710 10362
rect 16762 10310 16774 10362
rect 16826 10310 18860 10362
rect 1104 10288 18860 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 3786 10248 3792 10260
rect 2004 10220 3792 10248
rect 2004 10208 2010 10220
rect 3786 10208 3792 10220
rect 3844 10208 3850 10260
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 6270 10248 6276 10260
rect 6135 10220 6276 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 6270 10208 6276 10220
rect 6328 10208 6334 10260
rect 6730 10208 6736 10260
rect 6788 10248 6794 10260
rect 7009 10251 7067 10257
rect 7009 10248 7021 10251
rect 6788 10220 7021 10248
rect 6788 10208 6794 10220
rect 7009 10217 7021 10220
rect 7055 10217 7067 10251
rect 8110 10248 8116 10260
rect 7009 10211 7067 10217
rect 7852 10220 8116 10248
rect 2498 10140 2504 10192
rect 2556 10180 2562 10192
rect 3602 10180 3608 10192
rect 2556 10152 3608 10180
rect 2556 10140 2562 10152
rect 3602 10140 3608 10152
rect 3660 10140 3666 10192
rect 3878 10140 3884 10192
rect 3936 10180 3942 10192
rect 6181 10183 6239 10189
rect 6181 10180 6193 10183
rect 3936 10152 6193 10180
rect 3936 10140 3942 10152
rect 6181 10149 6193 10152
rect 6227 10149 6239 10183
rect 6181 10143 6239 10149
rect 6546 10140 6552 10192
rect 6604 10180 6610 10192
rect 7852 10189 7880 10220
rect 8110 10208 8116 10220
rect 8168 10208 8174 10260
rect 8754 10248 8760 10260
rect 8715 10220 8760 10248
rect 8754 10208 8760 10220
rect 8812 10208 8818 10260
rect 8846 10208 8852 10260
rect 8904 10248 8910 10260
rect 8941 10251 8999 10257
rect 8941 10248 8953 10251
rect 8904 10220 8953 10248
rect 8904 10208 8910 10220
rect 8941 10217 8953 10220
rect 8987 10217 8999 10251
rect 9490 10248 9496 10260
rect 9451 10220 9496 10248
rect 8941 10211 8999 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 9582 10208 9588 10260
rect 9640 10248 9646 10260
rect 10502 10248 10508 10260
rect 9640 10220 10508 10248
rect 9640 10208 9646 10220
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11388 10220 11713 10248
rect 11388 10208 11394 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 14734 10248 14740 10260
rect 11701 10211 11759 10217
rect 13372 10220 14740 10248
rect 7837 10183 7895 10189
rect 7837 10180 7849 10183
rect 6604 10152 7849 10180
rect 6604 10140 6610 10152
rect 7837 10149 7849 10152
rect 7883 10149 7895 10183
rect 10226 10180 10232 10192
rect 7837 10143 7895 10149
rect 8128 10152 10232 10180
rect 2225 10115 2283 10121
rect 2225 10081 2237 10115
rect 2271 10112 2283 10115
rect 2774 10112 2780 10124
rect 2271 10084 2780 10112
rect 2271 10081 2283 10084
rect 2225 10075 2283 10081
rect 2774 10072 2780 10084
rect 2832 10072 2838 10124
rect 3050 10072 3056 10124
rect 3108 10112 3114 10124
rect 3510 10112 3516 10124
rect 3108 10084 3516 10112
rect 3108 10072 3114 10084
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 4982 10112 4988 10124
rect 4943 10084 4988 10112
rect 4982 10072 4988 10084
rect 5040 10072 5046 10124
rect 5074 10072 5080 10124
rect 5132 10112 5138 10124
rect 5445 10115 5503 10121
rect 5445 10112 5457 10115
rect 5132 10084 5457 10112
rect 5132 10072 5138 10084
rect 5445 10081 5457 10084
rect 5491 10081 5503 10115
rect 5445 10075 5503 10081
rect 5810 10072 5816 10124
rect 5868 10112 5874 10124
rect 6086 10112 6092 10124
rect 5868 10084 6092 10112
rect 5868 10072 5874 10084
rect 6086 10072 6092 10084
rect 6144 10072 6150 10124
rect 6454 10072 6460 10124
rect 6512 10112 6518 10124
rect 6641 10115 6699 10121
rect 6641 10112 6653 10115
rect 6512 10084 6653 10112
rect 6512 10072 6518 10084
rect 6641 10081 6653 10084
rect 6687 10081 6699 10115
rect 6641 10075 6699 10081
rect 6733 10115 6791 10121
rect 6733 10081 6745 10115
rect 6779 10112 6791 10115
rect 7466 10112 7472 10124
rect 6779 10084 7472 10112
rect 6779 10081 6791 10084
rect 6733 10075 6791 10081
rect 7466 10072 7472 10084
rect 7524 10072 7530 10124
rect 7558 10072 7564 10124
rect 7616 10112 7622 10124
rect 8018 10112 8024 10124
rect 7616 10084 8024 10112
rect 7616 10072 7622 10084
rect 8018 10072 8024 10084
rect 8076 10072 8082 10124
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10044 2007 10047
rect 2130 10044 2136 10056
rect 1995 10016 2136 10044
rect 1995 10013 2007 10016
rect 1949 10007 2007 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10013 2375 10047
rect 2317 10007 2375 10013
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 2682 10044 2688 10056
rect 2639 10016 2688 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 1854 9936 1860 9988
rect 1912 9976 1918 9988
rect 2332 9976 2360 10007
rect 2682 10004 2688 10016
rect 2740 10004 2746 10056
rect 3602 10044 3608 10056
rect 3563 10016 3608 10044
rect 3602 10004 3608 10016
rect 3660 10004 3666 10056
rect 4062 10044 4068 10056
rect 4023 10016 4068 10044
rect 4062 10004 4068 10016
rect 4120 10004 4126 10056
rect 4338 10044 4344 10056
rect 4299 10016 4344 10044
rect 4338 10004 4344 10016
rect 4396 10004 4402 10056
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10044 4859 10047
rect 6549 10047 6607 10053
rect 4847 10016 6500 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 1912 9948 2360 9976
rect 1912 9936 1918 9948
rect 4246 9936 4252 9988
rect 4304 9976 4310 9988
rect 5534 9976 5540 9988
rect 4304 9948 5540 9976
rect 4304 9936 4310 9948
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 5629 9979 5687 9985
rect 5629 9945 5641 9979
rect 5675 9976 5687 9979
rect 5810 9976 5816 9988
rect 5675 9948 5816 9976
rect 5675 9945 5687 9948
rect 5629 9939 5687 9945
rect 5810 9936 5816 9948
rect 5868 9936 5874 9988
rect 6472 9976 6500 10016
rect 6549 10013 6561 10047
rect 6595 10044 6607 10047
rect 6822 10044 6828 10056
rect 6595 10016 6828 10044
rect 6595 10013 6607 10016
rect 6549 10007 6607 10013
rect 6822 10004 6828 10016
rect 6880 10004 6886 10056
rect 8128 10044 8156 10152
rect 10226 10140 10232 10152
rect 10284 10140 10290 10192
rect 8205 10115 8263 10121
rect 8205 10081 8217 10115
rect 8251 10112 8263 10115
rect 8478 10112 8484 10124
rect 8251 10084 8484 10112
rect 8251 10081 8263 10084
rect 8205 10075 8263 10081
rect 8478 10072 8484 10084
rect 8536 10072 8542 10124
rect 9582 10112 9588 10124
rect 9160 10084 9588 10112
rect 8386 10044 8392 10056
rect 7484 10016 8156 10044
rect 8347 10016 8392 10044
rect 7484 9985 7512 10016
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 9160 10053 9188 10084
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 10137 10115 10195 10121
rect 10137 10081 10149 10115
rect 10183 10081 10195 10115
rect 12345 10115 12403 10121
rect 12345 10112 12357 10115
rect 10137 10075 10195 10081
rect 11348 10084 12357 10112
rect 9117 10047 9188 10053
rect 9117 10013 9129 10047
rect 9163 10013 9188 10047
rect 9117 10007 9188 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 9306 10044 9312 10056
rect 9263 10016 9312 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 7469 9979 7527 9985
rect 7469 9976 7481 9979
rect 6472 9948 7481 9976
rect 7469 9945 7481 9948
rect 7515 9945 7527 9979
rect 7469 9939 7527 9945
rect 8297 9979 8355 9985
rect 8297 9945 8309 9979
rect 8343 9976 8355 9979
rect 8662 9976 8668 9988
rect 8343 9948 8668 9976
rect 8343 9945 8355 9948
rect 8297 9939 8355 9945
rect 8662 9936 8668 9948
rect 8720 9936 8726 9988
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 3694 9908 3700 9920
rect 3467 9880 3700 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 3694 9868 3700 9880
rect 3752 9868 3758 9920
rect 3878 9908 3884 9920
rect 3839 9880 3884 9908
rect 3878 9868 3884 9880
rect 3936 9868 3942 9920
rect 4154 9908 4160 9920
rect 4115 9880 4160 9908
rect 4154 9868 4160 9880
rect 4212 9868 4218 9920
rect 4338 9868 4344 9920
rect 4396 9908 4402 9920
rect 4433 9911 4491 9917
rect 4433 9908 4445 9911
rect 4396 9880 4445 9908
rect 4396 9868 4402 9880
rect 4433 9877 4445 9880
rect 4479 9877 4491 9911
rect 4433 9871 4491 9877
rect 4893 9911 4951 9917
rect 4893 9877 4905 9911
rect 4939 9908 4951 9911
rect 5721 9911 5779 9917
rect 5721 9908 5733 9911
rect 4939 9880 5733 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 5721 9877 5733 9880
rect 5767 9908 5779 9911
rect 6454 9908 6460 9920
rect 5767 9880 6460 9908
rect 5767 9877 5779 9880
rect 5721 9871 5779 9877
rect 6454 9868 6460 9880
rect 6512 9868 6518 9920
rect 6914 9868 6920 9920
rect 6972 9908 6978 9920
rect 7377 9911 7435 9917
rect 7377 9908 7389 9911
rect 6972 9880 7389 9908
rect 6972 9868 6978 9880
rect 7377 9877 7389 9880
rect 7423 9877 7435 9911
rect 7377 9871 7435 9877
rect 7742 9868 7748 9920
rect 7800 9908 7806 9920
rect 9160 9908 9188 10007
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 9858 10044 9864 10056
rect 9819 10016 9864 10044
rect 9858 10004 9864 10016
rect 9916 10004 9922 10056
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 10152 9976 10180 10075
rect 11348 10056 11376 10084
rect 12345 10081 12357 10084
rect 12391 10081 12403 10115
rect 12345 10075 12403 10081
rect 10321 10047 10379 10053
rect 10321 10013 10333 10047
rect 10367 10044 10379 10047
rect 11330 10044 11336 10056
rect 10367 10016 11336 10044
rect 10367 10013 10379 10016
rect 10321 10007 10379 10013
rect 11330 10004 11336 10016
rect 11388 10004 11394 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11793 10047 11851 10053
rect 11793 10044 11805 10047
rect 11756 10016 11805 10044
rect 11756 10004 11762 10016
rect 11793 10013 11805 10016
rect 11839 10013 11851 10047
rect 11793 10007 11851 10013
rect 12253 10047 12311 10053
rect 12253 10013 12265 10047
rect 12299 10044 12311 10047
rect 13372 10044 13400 10220
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 16022 10248 16028 10260
rect 14844 10220 16028 10248
rect 14844 10180 14872 10220
rect 16022 10208 16028 10220
rect 16080 10208 16086 10260
rect 16577 10251 16635 10257
rect 16577 10217 16589 10251
rect 16623 10248 16635 10251
rect 17034 10248 17040 10260
rect 16623 10220 17040 10248
rect 16623 10217 16635 10220
rect 16577 10211 16635 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 12299 10016 13400 10044
rect 13464 10152 14872 10180
rect 12299 10013 12311 10016
rect 12253 10007 12311 10013
rect 12618 9985 12624 9988
rect 10566 9979 10624 9985
rect 10566 9976 10578 9979
rect 9548 9948 10578 9976
rect 9548 9936 9554 9948
rect 10566 9945 10578 9948
rect 10612 9945 10624 9979
rect 12612 9976 12624 9985
rect 10566 9939 10624 9945
rect 10704 9948 12480 9976
rect 12579 9948 12624 9976
rect 7800 9880 9188 9908
rect 9401 9911 9459 9917
rect 7800 9868 7806 9880
rect 9401 9877 9413 9911
rect 9447 9908 9459 9911
rect 9582 9908 9588 9920
rect 9447 9880 9588 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9953 9911 10011 9917
rect 9953 9877 9965 9911
rect 9999 9908 10011 9911
rect 10226 9908 10232 9920
rect 9999 9880 10232 9908
rect 9999 9877 10011 9880
rect 9953 9871 10011 9877
rect 10226 9868 10232 9880
rect 10284 9908 10290 9920
rect 10704 9908 10732 9948
rect 10284 9880 10732 9908
rect 12069 9911 12127 9917
rect 10284 9868 10290 9880
rect 12069 9877 12081 9911
rect 12115 9908 12127 9911
rect 12342 9908 12348 9920
rect 12115 9880 12348 9908
rect 12115 9877 12127 9880
rect 12069 9871 12127 9877
rect 12342 9868 12348 9880
rect 12400 9868 12406 9920
rect 12452 9908 12480 9948
rect 12612 9939 12624 9948
rect 12618 9936 12624 9939
rect 12676 9936 12682 9988
rect 13464 9908 13492 10152
rect 14918 10140 14924 10192
rect 14976 10180 14982 10192
rect 14976 10152 17172 10180
rect 14976 10140 14982 10152
rect 14090 10072 14096 10124
rect 14148 10112 14154 10124
rect 14277 10115 14335 10121
rect 14277 10112 14289 10115
rect 14148 10084 14289 10112
rect 14148 10072 14154 10084
rect 14277 10081 14289 10084
rect 14323 10112 14335 10115
rect 15473 10115 15531 10121
rect 15473 10112 15485 10115
rect 14323 10084 15485 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 15473 10081 15485 10084
rect 15519 10081 15531 10115
rect 15838 10112 15844 10124
rect 15799 10084 15844 10112
rect 15473 10075 15531 10081
rect 15838 10072 15844 10084
rect 15896 10072 15902 10124
rect 16022 10112 16028 10124
rect 15983 10084 16028 10112
rect 16022 10072 16028 10084
rect 16080 10072 16086 10124
rect 17144 10121 17172 10152
rect 17218 10140 17224 10192
rect 17276 10180 17282 10192
rect 18414 10180 18420 10192
rect 17276 10152 18420 10180
rect 17276 10140 17282 10152
rect 18414 10140 18420 10152
rect 18472 10140 18478 10192
rect 17129 10115 17187 10121
rect 17129 10081 17141 10115
rect 17175 10081 17187 10115
rect 17954 10112 17960 10124
rect 17915 10084 17960 10112
rect 17129 10075 17187 10081
rect 17954 10072 17960 10084
rect 18012 10072 18018 10124
rect 14366 10044 14372 10056
rect 14327 10016 14372 10044
rect 14366 10004 14372 10016
rect 14424 10004 14430 10056
rect 14461 10047 14519 10053
rect 14461 10013 14473 10047
rect 14507 10044 14519 10047
rect 16298 10044 16304 10056
rect 14507 10016 16304 10044
rect 14507 10013 14519 10016
rect 14461 10007 14519 10013
rect 16298 10004 16304 10016
rect 16356 10004 16362 10056
rect 16942 10044 16948 10056
rect 16903 10016 16948 10044
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 18230 10044 18236 10056
rect 17328 10016 18000 10044
rect 18191 10016 18236 10044
rect 13909 9979 13967 9985
rect 13909 9945 13921 9979
rect 13955 9976 13967 9979
rect 15194 9976 15200 9988
rect 13955 9948 15200 9976
rect 13955 9945 13967 9948
rect 13909 9939 13967 9945
rect 15194 9936 15200 9948
rect 15252 9976 15258 9988
rect 15289 9979 15347 9985
rect 15289 9976 15301 9979
rect 15252 9948 15301 9976
rect 15252 9936 15258 9948
rect 15289 9945 15301 9948
rect 15335 9945 15347 9979
rect 15289 9939 15347 9945
rect 15378 9936 15384 9988
rect 15436 9976 15442 9988
rect 15654 9976 15660 9988
rect 15436 9948 15660 9976
rect 15436 9936 15442 9948
rect 15654 9936 15660 9948
rect 15712 9936 15718 9988
rect 16117 9979 16175 9985
rect 16117 9945 16129 9979
rect 16163 9976 16175 9979
rect 17328 9976 17356 10016
rect 16163 9948 17356 9976
rect 16163 9945 16175 9948
rect 16117 9939 16175 9945
rect 17494 9936 17500 9988
rect 17552 9976 17558 9988
rect 17865 9979 17923 9985
rect 17865 9976 17877 9979
rect 17552 9948 17877 9976
rect 17552 9936 17558 9948
rect 17865 9945 17877 9948
rect 17911 9945 17923 9979
rect 17972 9976 18000 10016
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 18322 9976 18328 9988
rect 17972 9948 18328 9976
rect 17865 9939 17923 9945
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 13722 9908 13728 9920
rect 12452 9880 13492 9908
rect 13683 9880 13728 9908
rect 13722 9868 13728 9880
rect 13780 9868 13786 9920
rect 14826 9908 14832 9920
rect 14787 9880 14832 9908
rect 14826 9868 14832 9880
rect 14884 9868 14890 9920
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 16482 9908 16488 9920
rect 14976 9880 15021 9908
rect 16443 9880 16488 9908
rect 14976 9868 14982 9880
rect 16482 9868 16488 9880
rect 16540 9868 16546 9920
rect 17037 9911 17095 9917
rect 17037 9877 17049 9911
rect 17083 9908 17095 9911
rect 17405 9911 17463 9917
rect 17405 9908 17417 9911
rect 17083 9880 17417 9908
rect 17083 9877 17095 9880
rect 17037 9871 17095 9877
rect 17405 9877 17417 9880
rect 17451 9877 17463 9911
rect 17770 9908 17776 9920
rect 17731 9880 17776 9908
rect 17405 9871 17463 9877
rect 17770 9868 17776 9880
rect 17828 9868 17834 9920
rect 18414 9908 18420 9920
rect 18375 9880 18420 9908
rect 18414 9868 18420 9880
rect 18472 9868 18478 9920
rect 1104 9818 18860 9840
rect 1104 9766 5398 9818
rect 5450 9766 5462 9818
rect 5514 9766 5526 9818
rect 5578 9766 5590 9818
rect 5642 9766 5654 9818
rect 5706 9766 9846 9818
rect 9898 9766 9910 9818
rect 9962 9766 9974 9818
rect 10026 9766 10038 9818
rect 10090 9766 10102 9818
rect 10154 9766 14294 9818
rect 14346 9766 14358 9818
rect 14410 9766 14422 9818
rect 14474 9766 14486 9818
rect 14538 9766 14550 9818
rect 14602 9766 18860 9818
rect 1104 9744 18860 9766
rect 3786 9664 3792 9716
rect 3844 9704 3850 9716
rect 4893 9707 4951 9713
rect 4893 9704 4905 9707
rect 3844 9676 4905 9704
rect 3844 9664 3850 9676
rect 4893 9673 4905 9676
rect 4939 9673 4951 9707
rect 4893 9667 4951 9673
rect 2130 9596 2136 9648
rect 2188 9636 2194 9648
rect 4908 9636 4936 9667
rect 5074 9664 5080 9716
rect 5132 9704 5138 9716
rect 6365 9707 6423 9713
rect 6365 9704 6377 9707
rect 5132 9676 6377 9704
rect 5132 9664 5138 9676
rect 6365 9673 6377 9676
rect 6411 9704 6423 9707
rect 7558 9704 7564 9716
rect 6411 9676 7564 9704
rect 6411 9673 6423 9676
rect 6365 9667 6423 9673
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 8021 9707 8079 9713
rect 8021 9673 8033 9707
rect 8067 9704 8079 9707
rect 8110 9704 8116 9716
rect 8067 9676 8116 9704
rect 8067 9673 8079 9676
rect 8021 9667 8079 9673
rect 8110 9664 8116 9676
rect 8168 9664 8174 9716
rect 8662 9664 8668 9716
rect 8720 9704 8726 9716
rect 9674 9704 9680 9716
rect 8720 9676 9680 9704
rect 8720 9664 8726 9676
rect 9674 9664 9680 9676
rect 9732 9664 9738 9716
rect 9766 9664 9772 9716
rect 9824 9704 9830 9716
rect 10321 9707 10379 9713
rect 10321 9704 10333 9707
rect 9824 9676 10333 9704
rect 9824 9664 9830 9676
rect 10321 9673 10333 9676
rect 10367 9673 10379 9707
rect 10321 9667 10379 9673
rect 10410 9664 10416 9716
rect 10468 9704 10474 9716
rect 11606 9704 11612 9716
rect 10468 9676 11612 9704
rect 10468 9664 10474 9676
rect 11606 9664 11612 9676
rect 11664 9664 11670 9716
rect 14090 9704 14096 9716
rect 13188 9676 14096 9704
rect 5905 9639 5963 9645
rect 5905 9636 5917 9639
rect 2188 9608 4752 9636
rect 4908 9608 5917 9636
rect 2188 9596 2194 9608
rect 1946 9568 1952 9580
rect 1907 9540 1952 9568
rect 1946 9528 1952 9540
rect 2004 9528 2010 9580
rect 2222 9568 2228 9580
rect 2183 9540 2228 9568
rect 2222 9528 2228 9540
rect 2280 9528 2286 9580
rect 2409 9571 2467 9577
rect 2409 9537 2421 9571
rect 2455 9568 2467 9571
rect 2498 9568 2504 9580
rect 2455 9540 2504 9568
rect 2455 9537 2467 9540
rect 2409 9531 2467 9537
rect 1394 9460 1400 9512
rect 1452 9500 1458 9512
rect 2424 9500 2452 9531
rect 2498 9528 2504 9540
rect 2556 9528 2562 9580
rect 3878 9568 3884 9580
rect 3936 9577 3942 9580
rect 3848 9540 3884 9568
rect 3878 9528 3884 9540
rect 3936 9531 3948 9577
rect 3936 9528 3942 9531
rect 4062 9528 4068 9580
rect 4120 9568 4126 9580
rect 4157 9571 4215 9577
rect 4157 9568 4169 9571
rect 4120 9540 4169 9568
rect 4120 9528 4126 9540
rect 4157 9537 4169 9540
rect 4203 9537 4215 9571
rect 4157 9531 4215 9537
rect 1452 9472 2452 9500
rect 1452 9460 1458 9472
rect 1946 9392 1952 9444
rect 2004 9432 2010 9444
rect 4341 9435 4399 9441
rect 2004 9404 2912 9432
rect 2004 9392 2010 9404
rect 2222 9324 2228 9376
rect 2280 9364 2286 9376
rect 2501 9367 2559 9373
rect 2501 9364 2513 9367
rect 2280 9336 2513 9364
rect 2280 9324 2286 9336
rect 2501 9333 2513 9336
rect 2547 9333 2559 9367
rect 2774 9364 2780 9376
rect 2735 9336 2780 9364
rect 2501 9327 2559 9333
rect 2774 9324 2780 9336
rect 2832 9324 2838 9376
rect 2884 9364 2912 9404
rect 4341 9401 4353 9435
rect 4387 9432 4399 9435
rect 4724 9432 4752 9608
rect 5905 9605 5917 9608
rect 5951 9636 5963 9639
rect 6546 9636 6552 9648
rect 5951 9608 6552 9636
rect 5951 9605 5963 9608
rect 5905 9599 5963 9605
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 7098 9596 7104 9648
rect 7156 9636 7162 9648
rect 7478 9639 7536 9645
rect 7478 9636 7490 9639
rect 7156 9608 7490 9636
rect 7156 9596 7162 9608
rect 7478 9605 7490 9608
rect 7524 9605 7536 9639
rect 7478 9599 7536 9605
rect 8478 9596 8484 9648
rect 8536 9636 8542 9648
rect 12434 9636 12440 9648
rect 8536 9608 11376 9636
rect 8536 9596 8542 9608
rect 4801 9571 4859 9577
rect 4801 9537 4813 9571
rect 4847 9568 4859 9571
rect 5813 9571 5871 9577
rect 5813 9568 5825 9571
rect 4847 9540 5825 9568
rect 4847 9537 4859 9540
rect 4801 9531 4859 9537
rect 5813 9537 5825 9540
rect 5859 9568 5871 9571
rect 7650 9568 7656 9580
rect 5859 9540 7656 9568
rect 5859 9537 5871 9540
rect 5813 9531 5871 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7834 9568 7840 9580
rect 7795 9540 7840 9568
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8018 9528 8024 9580
rect 8076 9568 8082 9580
rect 8369 9571 8427 9577
rect 8369 9568 8381 9571
rect 8076 9540 8381 9568
rect 8076 9528 8082 9540
rect 8369 9537 8381 9540
rect 8415 9537 8427 9571
rect 8369 9531 8427 9537
rect 8662 9528 8668 9580
rect 8720 9568 8726 9580
rect 9585 9571 9643 9577
rect 9585 9568 9597 9571
rect 8720 9540 9597 9568
rect 8720 9528 8726 9540
rect 9585 9537 9597 9540
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 10226 9528 10232 9580
rect 10284 9568 10290 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10284 9540 10701 9568
rect 10284 9528 10290 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11348 9577 11376 9608
rect 11808 9608 12440 9636
rect 11808 9577 11836 9608
rect 12434 9596 12440 9608
rect 12492 9596 12498 9648
rect 13020 9639 13078 9645
rect 13020 9605 13032 9639
rect 13066 9636 13078 9639
rect 13188 9636 13216 9676
rect 14090 9664 14096 9676
rect 14148 9664 14154 9716
rect 14553 9707 14611 9713
rect 14553 9673 14565 9707
rect 14599 9704 14611 9707
rect 14826 9704 14832 9716
rect 14599 9676 14832 9704
rect 14599 9673 14611 9676
rect 14553 9667 14611 9673
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 17218 9704 17224 9716
rect 15344 9676 17224 9704
rect 15344 9664 15350 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17405 9707 17463 9713
rect 17405 9673 17417 9707
rect 17451 9704 17463 9707
rect 17494 9704 17500 9716
rect 17451 9676 17500 9704
rect 17451 9673 17463 9676
rect 17405 9667 17463 9673
rect 17494 9664 17500 9676
rect 17552 9664 17558 9716
rect 17681 9707 17739 9713
rect 17681 9673 17693 9707
rect 17727 9704 17739 9707
rect 17770 9704 17776 9716
rect 17727 9676 17776 9704
rect 17727 9673 17739 9676
rect 17681 9667 17739 9673
rect 17770 9664 17776 9676
rect 17828 9664 17834 9716
rect 14182 9636 14188 9648
rect 13066 9608 13216 9636
rect 13280 9608 14188 9636
rect 13066 9605 13078 9608
rect 13020 9599 13078 9605
rect 11333 9571 11391 9577
rect 10836 9540 10881 9568
rect 10836 9528 10842 9540
rect 11333 9537 11345 9571
rect 11379 9537 11391 9571
rect 11333 9531 11391 9537
rect 11793 9571 11851 9577
rect 11793 9537 11805 9571
rect 11839 9537 11851 9571
rect 12618 9568 12624 9580
rect 11793 9531 11851 9537
rect 11900 9540 12624 9568
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 6089 9503 6147 9509
rect 5040 9472 5085 9500
rect 5040 9460 5046 9472
rect 6089 9469 6101 9503
rect 6135 9500 6147 9503
rect 6362 9500 6368 9512
rect 6135 9472 6368 9500
rect 6135 9469 6147 9472
rect 6089 9463 6147 9469
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 7745 9503 7803 9509
rect 7745 9469 7757 9503
rect 7791 9500 7803 9503
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7791 9472 8125 9500
rect 7791 9469 7803 9472
rect 7745 9463 7803 9469
rect 8113 9469 8125 9472
rect 8159 9469 8171 9503
rect 10962 9500 10968 9512
rect 10923 9472 10968 9500
rect 8113 9463 8171 9469
rect 5445 9435 5503 9441
rect 4387 9404 4660 9432
rect 4724 9404 5396 9432
rect 4387 9401 4399 9404
rect 4341 9395 4399 9401
rect 4154 9364 4160 9376
rect 2884 9336 4160 9364
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4430 9364 4436 9376
rect 4391 9336 4436 9364
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4632 9364 4660 9404
rect 5074 9364 5080 9376
rect 4632 9336 5080 9364
rect 5074 9324 5080 9336
rect 5132 9324 5138 9376
rect 5368 9373 5396 9404
rect 5445 9401 5457 9435
rect 5491 9432 5503 9435
rect 5810 9432 5816 9444
rect 5491 9404 5816 9432
rect 5491 9401 5503 9404
rect 5445 9395 5503 9401
rect 5810 9392 5816 9404
rect 5868 9392 5874 9444
rect 5353 9367 5411 9373
rect 5353 9333 5365 9367
rect 5399 9364 5411 9367
rect 6178 9364 6184 9376
rect 5399 9336 6184 9364
rect 5399 9333 5411 9336
rect 5353 9327 5411 9333
rect 6178 9324 6184 9336
rect 6236 9324 6242 9376
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 7760 9364 7788 9463
rect 10962 9460 10968 9472
rect 11020 9460 11026 9512
rect 7926 9392 7932 9444
rect 7984 9392 7990 9444
rect 9490 9432 9496 9444
rect 9403 9404 9496 9432
rect 9490 9392 9496 9404
rect 9548 9432 9554 9444
rect 10980 9432 11008 9460
rect 9548 9404 11008 9432
rect 11149 9435 11207 9441
rect 9548 9392 9554 9404
rect 11149 9401 11161 9435
rect 11195 9432 11207 9435
rect 11698 9432 11704 9444
rect 11195 9404 11704 9432
rect 11195 9401 11207 9404
rect 11149 9395 11207 9401
rect 11698 9392 11704 9404
rect 11756 9392 11762 9444
rect 11900 9441 11928 9540
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13280 9577 13308 9608
rect 14182 9596 14188 9608
rect 14240 9636 14246 9648
rect 15372 9639 15430 9645
rect 14240 9608 15148 9636
rect 14240 9596 14246 9608
rect 13265 9571 13323 9577
rect 13265 9537 13277 9571
rect 13311 9537 13323 9571
rect 13265 9531 13323 9537
rect 13725 9571 13783 9577
rect 13725 9537 13737 9571
rect 13771 9568 13783 9571
rect 14645 9571 14703 9577
rect 13771 9540 14228 9568
rect 13771 9537 13783 9540
rect 13725 9531 13783 9537
rect 13354 9460 13360 9512
rect 13412 9500 13418 9512
rect 13817 9503 13875 9509
rect 13817 9500 13829 9503
rect 13412 9472 13829 9500
rect 13412 9460 13418 9472
rect 13817 9469 13829 9472
rect 13863 9469 13875 9503
rect 13817 9463 13875 9469
rect 13909 9503 13967 9509
rect 13909 9469 13921 9503
rect 13955 9469 13967 9503
rect 13909 9463 13967 9469
rect 11885 9435 11943 9441
rect 11885 9401 11897 9435
rect 11931 9401 11943 9435
rect 11885 9395 11943 9401
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 13924 9432 13952 9463
rect 14200 9441 14228 9540
rect 14645 9537 14657 9571
rect 14691 9568 14703 9571
rect 14918 9568 14924 9580
rect 14691 9540 14924 9568
rect 14691 9537 14703 9540
rect 14645 9531 14703 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 15120 9577 15148 9608
rect 15372 9605 15384 9639
rect 15418 9636 15430 9639
rect 15562 9636 15568 9648
rect 15418 9608 15568 9636
rect 15418 9605 15430 9608
rect 15372 9599 15430 9605
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 16482 9596 16488 9648
rect 16540 9636 16546 9648
rect 16945 9639 17003 9645
rect 16945 9636 16957 9639
rect 16540 9608 16957 9636
rect 16540 9596 16546 9608
rect 16945 9605 16957 9608
rect 16991 9605 17003 9639
rect 16945 9599 17003 9605
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 18049 9639 18107 9645
rect 17092 9608 17137 9636
rect 17092 9596 17098 9608
rect 18049 9605 18061 9639
rect 18095 9636 18107 9639
rect 18230 9636 18236 9648
rect 18095 9608 18236 9636
rect 18095 9605 18107 9608
rect 18049 9599 18107 9605
rect 18230 9596 18236 9608
rect 18288 9636 18294 9648
rect 19518 9636 19524 9648
rect 18288 9608 19524 9636
rect 18288 9596 18294 9608
rect 19518 9596 19524 9608
rect 19576 9596 19582 9648
rect 15105 9571 15163 9577
rect 15105 9537 15117 9571
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 16758 9528 16764 9580
rect 16816 9568 16822 9580
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 16816 9540 17509 9568
rect 16816 9528 16822 9540
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18966 9568 18972 9580
rect 18187 9540 18972 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 14734 9500 14740 9512
rect 14695 9472 14740 9500
rect 14734 9460 14740 9472
rect 14792 9460 14798 9512
rect 16853 9503 16911 9509
rect 16853 9469 16865 9503
rect 16899 9469 16911 9503
rect 16853 9463 16911 9469
rect 18233 9503 18291 9509
rect 18233 9469 18245 9503
rect 18279 9469 18291 9503
rect 18233 9463 18291 9469
rect 13780 9404 13952 9432
rect 14185 9435 14243 9441
rect 13780 9392 13786 9404
rect 14185 9401 14197 9435
rect 14231 9401 14243 9435
rect 14185 9395 14243 9401
rect 16114 9392 16120 9444
rect 16172 9432 16178 9444
rect 16485 9435 16543 9441
rect 16485 9432 16497 9435
rect 16172 9404 16497 9432
rect 16172 9392 16178 9404
rect 16485 9401 16497 9404
rect 16531 9401 16543 9435
rect 16868 9432 16896 9463
rect 17678 9432 17684 9444
rect 16868 9404 17684 9432
rect 16485 9395 16543 9401
rect 17678 9392 17684 9404
rect 17736 9432 17742 9444
rect 17862 9432 17868 9444
rect 17736 9404 17868 9432
rect 17736 9392 17742 9404
rect 17862 9392 17868 9404
rect 17920 9432 17926 9444
rect 18248 9432 18276 9463
rect 17920 9404 18276 9432
rect 17920 9392 17926 9404
rect 6880 9336 7788 9364
rect 7944 9364 7972 9392
rect 9766 9364 9772 9376
rect 7944 9336 9772 9364
rect 6880 9324 6886 9336
rect 9766 9324 9772 9336
rect 9824 9324 9830 9376
rect 10226 9364 10232 9376
rect 10187 9336 10232 9364
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 11606 9364 11612 9376
rect 11567 9336 11612 9364
rect 11606 9324 11612 9336
rect 11664 9324 11670 9376
rect 12526 9324 12532 9376
rect 12584 9364 12590 9376
rect 13357 9367 13415 9373
rect 13357 9364 13369 9367
rect 12584 9336 13369 9364
rect 12584 9324 12590 9336
rect 13357 9333 13369 9336
rect 13403 9333 13415 9367
rect 13357 9327 13415 9333
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 14734 9364 14740 9376
rect 13504 9336 14740 9364
rect 13504 9324 13510 9336
rect 14734 9324 14740 9336
rect 14792 9324 14798 9376
rect 1104 9274 18860 9296
rect 1104 9222 3174 9274
rect 3226 9222 3238 9274
rect 3290 9222 3302 9274
rect 3354 9222 3366 9274
rect 3418 9222 3430 9274
rect 3482 9222 7622 9274
rect 7674 9222 7686 9274
rect 7738 9222 7750 9274
rect 7802 9222 7814 9274
rect 7866 9222 7878 9274
rect 7930 9222 12070 9274
rect 12122 9222 12134 9274
rect 12186 9222 12198 9274
rect 12250 9222 12262 9274
rect 12314 9222 12326 9274
rect 12378 9222 16518 9274
rect 16570 9222 16582 9274
rect 16634 9222 16646 9274
rect 16698 9222 16710 9274
rect 16762 9222 16774 9274
rect 16826 9222 18860 9274
rect 1104 9200 18860 9222
rect 2866 9160 2872 9172
rect 1780 9132 2872 9160
rect 1780 9104 1808 9132
rect 2866 9120 2872 9132
rect 2924 9160 2930 9172
rect 3970 9160 3976 9172
rect 2924 9132 3188 9160
rect 3931 9132 3976 9160
rect 2924 9120 2930 9132
rect 1762 9052 1768 9104
rect 1820 9052 1826 9104
rect 3160 9092 3188 9132
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 4154 9120 4160 9172
rect 4212 9160 4218 9172
rect 4212 9132 6316 9160
rect 4212 9120 4218 9132
rect 4062 9092 4068 9104
rect 3160 9064 4068 9092
rect 1670 9024 1676 9036
rect 1631 8996 1676 9024
rect 1670 8984 1676 8996
rect 1728 8984 1734 9036
rect 1486 8956 1492 8968
rect 1447 8928 1492 8956
rect 1486 8916 1492 8928
rect 1544 8916 1550 8968
rect 2590 8916 2596 8968
rect 2648 8956 2654 8968
rect 3160 8965 3188 9064
rect 4062 9052 4068 9064
rect 4120 9092 4126 9104
rect 6288 9092 6316 9132
rect 6362 9120 6368 9172
rect 6420 9160 6426 9172
rect 6457 9163 6515 9169
rect 6457 9160 6469 9163
rect 6420 9132 6469 9160
rect 6420 9120 6426 9132
rect 6457 9129 6469 9132
rect 6503 9129 6515 9163
rect 6457 9123 6515 9129
rect 7193 9163 7251 9169
rect 7193 9129 7205 9163
rect 7239 9160 7251 9163
rect 8018 9160 8024 9172
rect 7239 9132 8024 9160
rect 7239 9129 7251 9132
rect 7193 9123 7251 9129
rect 8018 9120 8024 9132
rect 8076 9120 8082 9172
rect 9490 9160 9496 9172
rect 8496 9132 9496 9160
rect 6638 9092 6644 9104
rect 4120 9064 5120 9092
rect 6288 9064 6644 9092
rect 4120 9052 4126 9064
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 5092 9033 5120 9064
rect 6638 9052 6644 9064
rect 6696 9052 6702 9104
rect 5077 9027 5135 9033
rect 4580 8996 4625 9024
rect 4580 8984 4586 8996
rect 5077 8993 5089 9027
rect 5123 8993 5135 9027
rect 5077 8987 5135 8993
rect 6178 8984 6184 9036
rect 6236 9024 6242 9036
rect 6236 8996 7420 9024
rect 6236 8984 6242 8996
rect 2878 8959 2936 8965
rect 2878 8956 2890 8959
rect 2648 8928 2890 8956
rect 2648 8916 2654 8928
rect 2878 8925 2890 8928
rect 2924 8925 2936 8959
rect 2878 8919 2936 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3786 8956 3792 8968
rect 3145 8919 3203 8925
rect 3252 8928 3792 8956
rect 1302 8848 1308 8900
rect 1360 8888 1366 8900
rect 1360 8860 1900 8888
rect 1360 8848 1366 8860
rect 1762 8820 1768 8832
rect 1723 8792 1768 8820
rect 1762 8780 1768 8792
rect 1820 8780 1826 8832
rect 1872 8820 1900 8860
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 3252 8888 3280 8928
rect 3786 8916 3792 8928
rect 3844 8916 3850 8968
rect 5350 8965 5356 8968
rect 5344 8956 5356 8965
rect 4985 8935 5043 8941
rect 4985 8932 4997 8935
rect 4908 8904 4997 8932
rect 2188 8860 3280 8888
rect 3329 8891 3387 8897
rect 2188 8848 2194 8860
rect 3329 8857 3341 8891
rect 3375 8888 3387 8891
rect 3510 8888 3516 8900
rect 3375 8860 3516 8888
rect 3375 8857 3387 8860
rect 3329 8851 3387 8857
rect 3344 8820 3372 8851
rect 3510 8848 3516 8860
rect 3568 8888 3574 8900
rect 3970 8888 3976 8900
rect 3568 8860 3976 8888
rect 3568 8848 3574 8860
rect 3970 8848 3976 8860
rect 4028 8848 4034 8900
rect 4430 8888 4436 8900
rect 4391 8860 4436 8888
rect 4430 8848 4436 8860
rect 4488 8848 4494 8900
rect 1872 8792 3372 8820
rect 3421 8823 3479 8829
rect 3421 8789 3433 8823
rect 3467 8820 3479 8823
rect 3694 8820 3700 8832
rect 3467 8792 3700 8820
rect 3467 8789 3479 8792
rect 3421 8783 3479 8789
rect 3694 8780 3700 8792
rect 3752 8780 3758 8832
rect 3786 8780 3792 8832
rect 3844 8820 3850 8832
rect 4154 8820 4160 8832
rect 3844 8792 4160 8820
rect 3844 8780 3850 8792
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4396 8792 4441 8820
rect 4396 8780 4402 8792
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4801 8823 4859 8829
rect 4801 8820 4813 8823
rect 4580 8792 4813 8820
rect 4580 8780 4586 8792
rect 4801 8789 4813 8792
rect 4847 8789 4859 8823
rect 4908 8820 4936 8904
rect 4985 8901 4997 8904
rect 5031 8901 5043 8935
rect 5311 8928 5356 8956
rect 5344 8919 5356 8928
rect 5350 8916 5356 8919
rect 5408 8916 5414 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6730 8956 6736 8968
rect 6595 8928 6736 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 6730 8916 6736 8928
rect 6788 8916 6794 8968
rect 7285 8959 7343 8965
rect 7285 8925 7297 8959
rect 7331 8925 7343 8959
rect 7392 8956 7420 8996
rect 8386 8956 8392 8968
rect 7392 8928 8392 8956
rect 7285 8919 7343 8925
rect 4985 8895 5043 8901
rect 5718 8848 5724 8900
rect 5776 8888 5782 8900
rect 6822 8888 6828 8900
rect 5776 8860 6828 8888
rect 5776 8848 5782 8860
rect 6822 8848 6828 8860
rect 6880 8888 6886 8900
rect 7300 8888 7328 8919
rect 8386 8916 8392 8928
rect 8444 8916 8450 8968
rect 7558 8897 7564 8900
rect 7552 8888 7564 8897
rect 6880 8860 7328 8888
rect 7519 8860 7564 8888
rect 6880 8848 6886 8860
rect 7552 8851 7564 8860
rect 7558 8848 7564 8851
rect 7616 8848 7622 8900
rect 5074 8820 5080 8832
rect 4908 8792 5080 8820
rect 4801 8783 4859 8789
rect 5074 8780 5080 8792
rect 5132 8780 5138 8832
rect 6270 8780 6276 8832
rect 6328 8820 6334 8832
rect 8496 8820 8524 9132
rect 9490 9120 9496 9132
rect 9548 9120 9554 9172
rect 9674 9120 9680 9172
rect 9732 9160 9738 9172
rect 10781 9163 10839 9169
rect 10781 9160 10793 9163
rect 9732 9132 10793 9160
rect 9732 9120 9738 9132
rect 10781 9129 10793 9132
rect 10827 9129 10839 9163
rect 10781 9123 10839 9129
rect 11238 9120 11244 9172
rect 11296 9160 11302 9172
rect 11698 9160 11704 9172
rect 11296 9132 11704 9160
rect 11296 9120 11302 9132
rect 11698 9120 11704 9132
rect 11756 9120 11762 9172
rect 13173 9163 13231 9169
rect 13173 9129 13185 9163
rect 13219 9160 13231 9163
rect 13354 9160 13360 9172
rect 13219 9132 13360 9160
rect 13219 9129 13231 9132
rect 13173 9123 13231 9129
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 13909 9163 13967 9169
rect 13909 9129 13921 9163
rect 13955 9160 13967 9163
rect 13998 9160 14004 9172
rect 13955 9132 14004 9160
rect 13955 9129 13967 9132
rect 13909 9123 13967 9129
rect 13998 9120 14004 9132
rect 14056 9120 14062 9172
rect 14090 9120 14096 9172
rect 14148 9160 14154 9172
rect 18138 9160 18144 9172
rect 14148 9132 14193 9160
rect 14568 9132 18144 9160
rect 14148 9120 14154 9132
rect 9306 9092 9312 9104
rect 8588 9064 9312 9092
rect 8588 8968 8616 9064
rect 9306 9052 9312 9064
rect 9364 9052 9370 9104
rect 10686 9092 10692 9104
rect 10599 9064 10692 9092
rect 10686 9052 10692 9064
rect 10744 9092 10750 9104
rect 10744 9064 12204 9092
rect 10744 9052 10750 9064
rect 10962 8984 10968 9036
rect 11020 9024 11026 9036
rect 12176 9033 12204 9064
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 14568 9092 14596 9132
rect 18138 9120 18144 9132
rect 18196 9120 18202 9172
rect 13872 9064 14596 9092
rect 13872 9052 13878 9064
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11020 8996 11345 9024
rect 11020 8984 11026 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11333 8987 11391 8993
rect 12161 9027 12219 9033
rect 12161 8993 12173 9027
rect 12207 8993 12219 9027
rect 12161 8987 12219 8993
rect 12618 8984 12624 9036
rect 12676 9024 12682 9036
rect 13446 9024 13452 9036
rect 12676 8996 13452 9024
rect 12676 8984 12682 8996
rect 13446 8984 13452 8996
rect 13504 8984 13510 9036
rect 15749 9027 15807 9033
rect 15749 8993 15761 9027
rect 15795 9024 15807 9027
rect 16114 9024 16120 9036
rect 15795 8996 16120 9024
rect 15795 8993 15807 8996
rect 15749 8987 15807 8993
rect 16114 8984 16120 8996
rect 16172 8984 16178 9036
rect 18690 8984 18696 9036
rect 18748 9024 18754 9036
rect 19334 9024 19340 9036
rect 18748 8996 19340 9024
rect 18748 8984 18754 8996
rect 19334 8984 19340 8996
rect 19392 8984 19398 9036
rect 8570 8916 8576 8968
rect 8628 8916 8634 8968
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 8941 8959 8999 8965
rect 8941 8956 8953 8959
rect 8812 8928 8953 8956
rect 8812 8916 8818 8928
rect 8941 8925 8953 8928
rect 8987 8925 8999 8959
rect 9306 8956 9312 8968
rect 9267 8928 9312 8956
rect 8941 8919 8999 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 9398 8916 9404 8968
rect 9456 8956 9462 8968
rect 9565 8959 9623 8965
rect 9565 8956 9577 8959
rect 9456 8928 9577 8956
rect 9456 8916 9462 8928
rect 9565 8925 9577 8928
rect 9611 8925 9623 8959
rect 9565 8919 9623 8925
rect 10318 8916 10324 8968
rect 10376 8956 10382 8968
rect 10870 8956 10876 8968
rect 10376 8928 10876 8956
rect 10376 8916 10382 8928
rect 10870 8916 10876 8928
rect 10928 8956 10934 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 10928 8928 11253 8956
rect 10928 8916 10934 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11977 8959 12035 8965
rect 11977 8925 11989 8959
rect 12023 8956 12035 8959
rect 12066 8956 12072 8968
rect 12023 8928 12072 8956
rect 12023 8925 12035 8928
rect 11977 8919 12035 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 12805 8959 12863 8965
rect 12805 8956 12817 8959
rect 12768 8928 12817 8956
rect 12768 8916 12774 8928
rect 12805 8925 12817 8928
rect 12851 8925 12863 8959
rect 12805 8919 12863 8925
rect 13265 8959 13323 8965
rect 13265 8925 13277 8959
rect 13311 8956 13323 8959
rect 13722 8956 13728 8968
rect 13311 8928 13728 8956
rect 13311 8925 13323 8928
rect 13265 8919 13323 8925
rect 13722 8916 13728 8928
rect 13780 8916 13786 8968
rect 14182 8916 14188 8968
rect 14240 8956 14246 8968
rect 15473 8959 15531 8965
rect 15473 8956 15485 8959
rect 14240 8928 15485 8956
rect 14240 8916 14246 8928
rect 15473 8925 15485 8928
rect 15519 8956 15531 8959
rect 15838 8956 15844 8968
rect 15519 8928 15844 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 15838 8916 15844 8928
rect 15896 8956 15902 8968
rect 16206 8956 16212 8968
rect 15896 8928 16212 8956
rect 15896 8916 15902 8928
rect 16206 8916 16212 8928
rect 16264 8956 16270 8968
rect 16485 8959 16543 8965
rect 16485 8956 16497 8959
rect 16264 8928 16497 8956
rect 16264 8916 16270 8928
rect 16485 8925 16497 8928
rect 16531 8925 16543 8959
rect 16485 8919 16543 8925
rect 16752 8959 16810 8965
rect 16752 8925 16764 8959
rect 16798 8956 16810 8959
rect 17126 8956 17132 8968
rect 16798 8928 17132 8956
rect 16798 8925 16810 8928
rect 16752 8919 16810 8925
rect 17126 8916 17132 8928
rect 17184 8916 17190 8968
rect 18233 8959 18291 8965
rect 18233 8925 18245 8959
rect 18279 8956 18291 8959
rect 18322 8956 18328 8968
rect 18279 8928 18328 8956
rect 18279 8925 18291 8928
rect 18233 8919 18291 8925
rect 18322 8916 18328 8928
rect 18380 8916 18386 8968
rect 18506 8956 18512 8968
rect 18467 8928 18512 8956
rect 18506 8916 18512 8928
rect 18564 8916 18570 8968
rect 8846 8848 8852 8900
rect 8904 8888 8910 8900
rect 8904 8860 11652 8888
rect 8904 8848 8910 8860
rect 8662 8820 8668 8832
rect 6328 8792 8524 8820
rect 8623 8792 8668 8820
rect 6328 8780 6334 8792
rect 8662 8780 8668 8792
rect 8720 8780 8726 8832
rect 8754 8780 8760 8832
rect 8812 8820 8818 8832
rect 9125 8823 9183 8829
rect 9125 8820 9137 8823
rect 8812 8792 9137 8820
rect 8812 8780 8818 8792
rect 9125 8789 9137 8792
rect 9171 8789 9183 8823
rect 9125 8783 9183 8789
rect 9766 8780 9772 8832
rect 9824 8820 9830 8832
rect 10962 8820 10968 8832
rect 9824 8792 10968 8820
rect 9824 8780 9830 8792
rect 10962 8780 10968 8792
rect 11020 8820 11026 8832
rect 11624 8829 11652 8860
rect 13354 8848 13360 8900
rect 13412 8888 13418 8900
rect 13412 8860 13584 8888
rect 13412 8848 13418 8860
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 11020 8792 11161 8820
rect 11020 8780 11026 8792
rect 11149 8789 11161 8792
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8789 11667 8823
rect 12066 8820 12072 8832
rect 12027 8792 12072 8820
rect 11609 8783 11667 8789
rect 12066 8780 12072 8792
rect 12124 8780 12130 8832
rect 12618 8780 12624 8832
rect 12676 8820 12682 8832
rect 12713 8823 12771 8829
rect 12713 8820 12725 8823
rect 12676 8792 12725 8820
rect 12676 8780 12682 8792
rect 12713 8789 12725 8792
rect 12759 8789 12771 8823
rect 12713 8783 12771 8789
rect 13170 8780 13176 8832
rect 13228 8820 13234 8832
rect 13446 8820 13452 8832
rect 13228 8792 13452 8820
rect 13228 8780 13234 8792
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13556 8820 13584 8860
rect 15194 8848 15200 8900
rect 15252 8897 15258 8900
rect 15252 8888 15264 8897
rect 15252 8860 15297 8888
rect 15252 8851 15264 8860
rect 15252 8848 15258 8851
rect 15562 8848 15568 8900
rect 15620 8888 15626 8900
rect 16025 8891 16083 8897
rect 16025 8888 16037 8891
rect 15620 8860 16037 8888
rect 15620 8848 15626 8860
rect 16025 8857 16037 8860
rect 16071 8888 16083 8891
rect 16298 8888 16304 8900
rect 16071 8860 16304 8888
rect 16071 8857 16083 8860
rect 16025 8851 16083 8857
rect 16298 8848 16304 8860
rect 16356 8888 16362 8900
rect 16356 8860 18368 8888
rect 16356 8848 16362 8860
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 13556 8792 15945 8820
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 16393 8823 16451 8829
rect 16393 8789 16405 8823
rect 16439 8820 16451 8823
rect 17126 8820 17132 8832
rect 16439 8792 17132 8820
rect 16439 8789 16451 8792
rect 16393 8783 16451 8789
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17276 8792 17877 8820
rect 17276 8780 17282 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 18046 8820 18052 8832
rect 18007 8792 18052 8820
rect 17865 8783 17923 8789
rect 18046 8780 18052 8792
rect 18104 8780 18110 8832
rect 18340 8829 18368 8860
rect 18325 8823 18383 8829
rect 18325 8789 18337 8823
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 1104 8730 18860 8752
rect 1104 8678 5398 8730
rect 5450 8678 5462 8730
rect 5514 8678 5526 8730
rect 5578 8678 5590 8730
rect 5642 8678 5654 8730
rect 5706 8678 9846 8730
rect 9898 8678 9910 8730
rect 9962 8678 9974 8730
rect 10026 8678 10038 8730
rect 10090 8678 10102 8730
rect 10154 8678 14294 8730
rect 14346 8678 14358 8730
rect 14410 8678 14422 8730
rect 14474 8678 14486 8730
rect 14538 8678 14550 8730
rect 14602 8678 18860 8730
rect 1104 8656 18860 8678
rect 2774 8576 2780 8628
rect 2832 8616 2838 8628
rect 6181 8619 6239 8625
rect 2832 8588 4272 8616
rect 2832 8576 2838 8588
rect 1670 8548 1676 8560
rect 1504 8520 1676 8548
rect 1504 8489 1532 8520
rect 1670 8508 1676 8520
rect 1728 8508 1734 8560
rect 2498 8508 2504 8560
rect 2556 8548 2562 8560
rect 3234 8548 3240 8560
rect 2556 8520 3240 8548
rect 2556 8508 2562 8520
rect 3234 8508 3240 8520
rect 3292 8508 3298 8560
rect 3418 8548 3424 8560
rect 3344 8520 3424 8548
rect 1762 8489 1768 8492
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8449 1547 8483
rect 1756 8480 1768 8489
rect 1675 8452 1768 8480
rect 1489 8443 1547 8449
rect 1756 8443 1768 8452
rect 1820 8480 1826 8492
rect 2590 8480 2596 8492
rect 1820 8452 2596 8480
rect 1762 8440 1768 8443
rect 1820 8440 1826 8452
rect 2590 8440 2596 8452
rect 2648 8440 2654 8492
rect 3142 8372 3148 8424
rect 3200 8372 3206 8424
rect 3344 8412 3372 8520
rect 3418 8508 3424 8520
rect 3476 8508 3482 8560
rect 3786 8548 3792 8560
rect 3712 8520 3792 8548
rect 3513 8483 3571 8489
rect 3513 8449 3525 8483
rect 3559 8480 3571 8483
rect 3712 8480 3740 8520
rect 3786 8508 3792 8520
rect 3844 8508 3850 8560
rect 3878 8508 3884 8560
rect 3936 8508 3942 8560
rect 4244 8557 4272 8588
rect 6181 8585 6193 8619
rect 6227 8616 6239 8619
rect 8478 8616 8484 8628
rect 6227 8588 8484 8616
rect 6227 8585 6239 8588
rect 6181 8579 6239 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 10226 8616 10232 8628
rect 9232 8588 10232 8616
rect 4229 8551 4287 8557
rect 4229 8517 4241 8551
rect 4275 8517 4287 8551
rect 4229 8511 4287 8517
rect 6822 8508 6828 8560
rect 6880 8548 6886 8560
rect 9145 8551 9203 8557
rect 6880 8520 7880 8548
rect 6880 8508 6886 8520
rect 3559 8452 3740 8480
rect 3559 8449 3571 8452
rect 3513 8443 3571 8449
rect 3789 8415 3847 8421
rect 3789 8412 3801 8415
rect 3344 8384 3801 8412
rect 3789 8381 3801 8384
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 2958 8344 2964 8356
rect 2915 8316 2964 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 2958 8304 2964 8316
rect 3016 8304 3022 8356
rect 3160 8344 3188 8372
rect 3160 8316 3648 8344
rect 3620 8294 3648 8316
rect 3896 8306 3924 8508
rect 3970 8440 3976 8492
rect 4028 8480 4034 8492
rect 5810 8480 5816 8492
rect 4028 8452 4073 8480
rect 5771 8452 5816 8480
rect 4028 8440 4034 8452
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 7852 8489 7880 8520
rect 9145 8517 9157 8551
rect 9191 8548 9203 8551
rect 9232 8548 9260 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10778 8576 10784 8628
rect 10836 8616 10842 8628
rect 12434 8616 12440 8628
rect 10836 8588 11468 8616
rect 12395 8588 12440 8616
rect 10836 8576 10842 8588
rect 9191 8520 9260 8548
rect 9191 8517 9203 8520
rect 9145 8511 9203 8517
rect 9306 8508 9312 8560
rect 9364 8548 9370 8560
rect 11440 8548 11468 8588
rect 12434 8576 12440 8588
rect 12492 8576 12498 8628
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 12710 8576 12716 8628
rect 12768 8616 12774 8628
rect 13449 8619 13507 8625
rect 13449 8616 13461 8619
rect 12768 8588 13461 8616
rect 12768 8576 12774 8588
rect 13449 8585 13461 8588
rect 13495 8585 13507 8619
rect 13449 8579 13507 8585
rect 13722 8576 13728 8628
rect 13780 8616 13786 8628
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13780 8588 13829 8616
rect 13780 8576 13786 8588
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 13817 8579 13875 8585
rect 13906 8576 13912 8628
rect 13964 8616 13970 8628
rect 14277 8619 14335 8625
rect 14277 8616 14289 8619
rect 13964 8588 14289 8616
rect 13964 8576 13970 8588
rect 14277 8585 14289 8588
rect 14323 8585 14335 8619
rect 14277 8579 14335 8585
rect 15286 8576 15292 8628
rect 15344 8616 15350 8628
rect 16022 8616 16028 8628
rect 15344 8588 16028 8616
rect 15344 8576 15350 8588
rect 16022 8576 16028 8588
rect 16080 8616 16086 8628
rect 16301 8619 16359 8625
rect 16301 8616 16313 8619
rect 16080 8588 16313 8616
rect 16080 8576 16086 8588
rect 16301 8585 16313 8588
rect 16347 8585 16359 8619
rect 17126 8616 17132 8628
rect 17087 8588 17132 8616
rect 16301 8579 16359 8585
rect 17126 8576 17132 8588
rect 17184 8576 17190 8628
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17368 8588 17509 8616
rect 17368 8576 17374 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 18322 8616 18328 8628
rect 18283 8588 18328 8616
rect 17497 8579 17555 8585
rect 18322 8576 18328 8588
rect 18380 8576 18386 8628
rect 12989 8551 13047 8557
rect 9364 8520 11376 8548
rect 11440 8520 12434 8548
rect 9364 8508 9370 8520
rect 9416 8489 9444 8520
rect 7570 8483 7628 8489
rect 7570 8480 7582 8483
rect 6840 8452 7582 8480
rect 5629 8415 5687 8421
rect 5629 8381 5641 8415
rect 5675 8381 5687 8415
rect 5629 8375 5687 8381
rect 5721 8415 5779 8421
rect 5721 8381 5733 8415
rect 5767 8412 5779 8415
rect 6178 8412 6184 8424
rect 5767 8384 6184 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 5353 8347 5411 8353
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5644 8344 5672 8375
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 5994 8344 6000 8356
rect 5399 8316 6000 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 3694 8294 3700 8306
rect 1486 8236 1492 8288
rect 1544 8276 1550 8288
rect 2222 8276 2228 8288
rect 1544 8248 2228 8276
rect 1544 8236 1550 8248
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 3620 8266 3700 8294
rect 3694 8254 3700 8266
rect 3752 8254 3758 8306
rect 3878 8254 3884 8306
rect 3936 8254 3942 8306
rect 5994 8304 6000 8316
rect 6052 8304 6058 8356
rect 6457 8347 6515 8353
rect 6457 8313 6469 8347
rect 6503 8344 6515 8347
rect 6730 8344 6736 8356
rect 6503 8316 6736 8344
rect 6503 8313 6515 8316
rect 6457 8307 6515 8313
rect 6730 8304 6736 8316
rect 6788 8304 6794 8356
rect 4338 8236 4344 8288
rect 4396 8276 4402 8288
rect 6270 8276 6276 8288
rect 4396 8248 6276 8276
rect 4396 8236 4402 8248
rect 6270 8236 6276 8248
rect 6328 8236 6334 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 6840 8276 6868 8452
rect 7570 8449 7582 8452
rect 7616 8449 7628 8483
rect 7570 8443 7628 8449
rect 7837 8483 7895 8489
rect 7837 8449 7849 8483
rect 7883 8449 7895 8483
rect 9401 8483 9459 8489
rect 7837 8443 7895 8449
rect 8404 8452 9352 8480
rect 8404 8412 8432 8452
rect 7852 8384 8432 8412
rect 9324 8412 9352 8452
rect 9401 8449 9413 8483
rect 9447 8449 9459 8483
rect 9401 8443 9459 8449
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 9548 8452 9593 8480
rect 9548 8440 9554 8452
rect 9674 8440 9680 8492
rect 9732 8480 9738 8492
rect 10134 8480 10140 8492
rect 9732 8452 10140 8480
rect 9732 8440 9738 8452
rect 10134 8440 10140 8452
rect 10192 8440 10198 8492
rect 10686 8440 10692 8492
rect 10744 8480 10750 8492
rect 11066 8483 11124 8489
rect 11066 8480 11078 8483
rect 10744 8452 11078 8480
rect 10744 8440 10750 8452
rect 11066 8449 11078 8452
rect 11112 8449 11124 8483
rect 11066 8443 11124 8449
rect 11348 8424 11376 8520
rect 11790 8480 11796 8492
rect 11751 8452 11796 8480
rect 11790 8440 11796 8452
rect 11848 8440 11854 8492
rect 12406 8480 12434 8520
rect 12989 8517 13001 8551
rect 13035 8548 13047 8551
rect 15470 8548 15476 8560
rect 13035 8520 15476 8548
rect 13035 8517 13047 8520
rect 12989 8511 13047 8517
rect 15470 8508 15476 8520
rect 15528 8508 15534 8560
rect 15596 8551 15654 8557
rect 15596 8517 15608 8551
rect 15642 8548 15654 8551
rect 15642 8520 16804 8548
rect 15642 8517 15654 8520
rect 15596 8511 15654 8517
rect 15286 8480 15292 8492
rect 12406 8452 15292 8480
rect 15286 8440 15292 8452
rect 15344 8440 15350 8492
rect 15838 8480 15844 8492
rect 15799 8452 15844 8480
rect 15838 8440 15844 8452
rect 15896 8440 15902 8492
rect 15930 8440 15936 8492
rect 15988 8480 15994 8492
rect 15988 8452 16033 8480
rect 15988 8440 15994 8452
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 16485 8483 16543 8489
rect 16485 8480 16497 8483
rect 16356 8452 16497 8480
rect 16356 8440 16362 8452
rect 16485 8449 16497 8452
rect 16531 8449 16543 8483
rect 16485 8443 16543 8449
rect 11330 8412 11336 8424
rect 9324 8384 10364 8412
rect 11291 8384 11336 8412
rect 6420 8248 6868 8276
rect 6420 8236 6426 8248
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7852 8276 7880 8384
rect 9398 8304 9404 8356
rect 9456 8344 9462 8356
rect 9677 8347 9735 8353
rect 9677 8344 9689 8347
rect 9456 8316 9689 8344
rect 9456 8304 9462 8316
rect 9677 8313 9689 8316
rect 9723 8313 9735 8347
rect 10336 8344 10364 8384
rect 11330 8372 11336 8384
rect 11388 8372 11394 8424
rect 11517 8415 11575 8421
rect 11517 8381 11529 8415
rect 11563 8412 11575 8415
rect 12066 8412 12072 8424
rect 11563 8384 12072 8412
rect 11563 8381 11575 8384
rect 11517 8375 11575 8381
rect 11532 8344 11560 8375
rect 12066 8372 12072 8384
rect 12124 8372 12130 8424
rect 13078 8412 13084 8424
rect 13039 8384 13084 8412
rect 13078 8372 13084 8384
rect 13136 8372 13142 8424
rect 13265 8415 13323 8421
rect 13265 8381 13277 8415
rect 13311 8381 13323 8415
rect 13906 8412 13912 8424
rect 13867 8384 13912 8412
rect 13265 8375 13323 8381
rect 10336 8316 10456 8344
rect 9677 8307 9735 8313
rect 8018 8276 8024 8288
rect 7156 8248 7880 8276
rect 7979 8248 8024 8276
rect 7156 8236 7162 8248
rect 8018 8236 8024 8248
rect 8076 8236 8082 8288
rect 9766 8236 9772 8288
rect 9824 8276 9830 8288
rect 9953 8279 10011 8285
rect 9953 8276 9965 8279
rect 9824 8248 9965 8276
rect 9824 8236 9830 8248
rect 9953 8245 9965 8248
rect 9999 8245 10011 8279
rect 10428 8276 10456 8316
rect 11348 8316 11560 8344
rect 13280 8344 13308 8375
rect 13906 8372 13912 8384
rect 13964 8372 13970 8424
rect 14090 8412 14096 8424
rect 14051 8384 14096 8412
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 16776 8412 16804 8520
rect 16850 8508 16856 8560
rect 16908 8548 16914 8560
rect 17865 8551 17923 8557
rect 17865 8548 17877 8551
rect 16908 8520 17877 8548
rect 16908 8508 16914 8520
rect 17865 8517 17877 8520
rect 17911 8517 17923 8551
rect 17865 8511 17923 8517
rect 17957 8551 18015 8557
rect 17957 8517 17969 8551
rect 18003 8548 18015 8551
rect 18598 8548 18604 8560
rect 18003 8520 18604 8548
rect 18003 8517 18015 8520
rect 17957 8511 18015 8517
rect 18598 8508 18604 8520
rect 18656 8508 18662 8560
rect 17034 8480 17040 8492
rect 16995 8452 17040 8480
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 18230 8440 18236 8492
rect 18288 8480 18294 8492
rect 18509 8483 18567 8489
rect 18509 8480 18521 8483
rect 18288 8452 18521 8480
rect 18288 8440 18294 8452
rect 18509 8449 18521 8452
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 17218 8412 17224 8424
rect 16776 8384 17224 8412
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 14108 8344 14136 8372
rect 16114 8344 16120 8356
rect 13280 8316 14136 8344
rect 14384 8316 14688 8344
rect 16075 8316 16120 8344
rect 11348 8276 11376 8316
rect 10428 8248 11376 8276
rect 9953 8239 10011 8245
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 11882 8276 11888 8288
rect 11756 8248 11888 8276
rect 11756 8236 11762 8248
rect 11882 8236 11888 8248
rect 11940 8236 11946 8288
rect 13262 8236 13268 8288
rect 13320 8276 13326 8288
rect 14384 8276 14412 8316
rect 13320 8248 14412 8276
rect 14461 8279 14519 8285
rect 13320 8236 13326 8248
rect 14461 8245 14473 8279
rect 14507 8276 14519 8279
rect 14550 8276 14556 8288
rect 14507 8248 14556 8276
rect 14507 8245 14519 8248
rect 14461 8239 14519 8245
rect 14550 8236 14556 8248
rect 14608 8236 14614 8288
rect 14660 8276 14688 8316
rect 16114 8304 16120 8316
rect 16172 8304 16178 8356
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 16264 8316 16681 8344
rect 16264 8304 16270 8316
rect 16669 8313 16681 8316
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 17862 8304 17868 8356
rect 17920 8344 17926 8356
rect 18064 8344 18092 8375
rect 17920 8316 18092 8344
rect 17920 8304 17926 8316
rect 16298 8276 16304 8288
rect 14660 8248 16304 8276
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 1104 8186 18860 8208
rect 1104 8134 3174 8186
rect 3226 8134 3238 8186
rect 3290 8134 3302 8186
rect 3354 8134 3366 8186
rect 3418 8134 3430 8186
rect 3482 8134 7622 8186
rect 7674 8134 7686 8186
rect 7738 8134 7750 8186
rect 7802 8134 7814 8186
rect 7866 8134 7878 8186
rect 7930 8134 12070 8186
rect 12122 8134 12134 8186
rect 12186 8134 12198 8186
rect 12250 8134 12262 8186
rect 12314 8134 12326 8186
rect 12378 8134 16518 8186
rect 16570 8134 16582 8186
rect 16634 8134 16646 8186
rect 16698 8134 16710 8186
rect 16762 8134 16774 8186
rect 16826 8134 18860 8186
rect 1104 8112 18860 8134
rect 1762 8032 1768 8084
rect 1820 8072 1826 8084
rect 2958 8072 2964 8084
rect 1820 8044 2964 8072
rect 1820 8032 1826 8044
rect 2958 8032 2964 8044
rect 3016 8072 3022 8084
rect 4154 8072 4160 8084
rect 3016 8044 4160 8072
rect 3016 8032 3022 8044
rect 4154 8032 4160 8044
rect 4212 8072 4218 8084
rect 4341 8075 4399 8081
rect 4212 8044 4292 8072
rect 4212 8032 4218 8044
rect 1670 7964 1676 8016
rect 1728 8004 1734 8016
rect 1946 8004 1952 8016
rect 1728 7976 1952 8004
rect 1728 7964 1734 7976
rect 1946 7964 1952 7976
rect 2004 7964 2010 8016
rect 2682 7964 2688 8016
rect 2740 7964 2746 8016
rect 3050 7964 3056 8016
rect 3108 7964 3114 8016
rect 3326 7964 3332 8016
rect 3384 8004 3390 8016
rect 3513 8007 3571 8013
rect 3513 8004 3525 8007
rect 3384 7976 3525 8004
rect 3384 7964 3390 7976
rect 3513 7973 3525 7976
rect 3559 7973 3571 8007
rect 3513 7967 3571 7973
rect 2225 7939 2283 7945
rect 2225 7905 2237 7939
rect 2271 7936 2283 7939
rect 2498 7936 2504 7948
rect 2271 7908 2504 7936
rect 2271 7905 2283 7908
rect 2225 7899 2283 7905
rect 2498 7896 2504 7908
rect 2556 7896 2562 7948
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2590 7828 2596 7880
rect 2648 7868 2654 7880
rect 2700 7868 2728 7964
rect 2648 7840 2728 7868
rect 2648 7828 2654 7840
rect 2774 7828 2780 7880
rect 2832 7868 2838 7880
rect 3068 7868 3096 7964
rect 3234 7936 3240 7948
rect 3160 7908 3240 7936
rect 3160 7877 3188 7908
rect 3234 7896 3240 7908
rect 3292 7896 3298 7948
rect 4264 7936 4292 8044
rect 4341 8041 4353 8075
rect 4387 8072 4399 8075
rect 5718 8072 5724 8084
rect 4387 8044 5396 8072
rect 5679 8044 5724 8072
rect 4387 8041 4399 8044
rect 4341 8035 4399 8041
rect 4430 8004 4436 8016
rect 4391 7976 4436 8004
rect 4430 7964 4436 7976
rect 4488 7964 4494 8016
rect 5368 8004 5396 8044
rect 5718 8032 5724 8044
rect 5776 8032 5782 8084
rect 6270 8032 6276 8084
rect 6328 8072 6334 8084
rect 11238 8072 11244 8084
rect 6328 8044 7972 8072
rect 6328 8032 6334 8044
rect 7944 8016 7972 8044
rect 8067 8044 11244 8072
rect 5902 8004 5908 8016
rect 5368 7976 5908 8004
rect 5902 7964 5908 7976
rect 5960 7964 5966 8016
rect 7006 7964 7012 8016
rect 7064 8004 7070 8016
rect 7834 8004 7840 8016
rect 7064 7976 7840 8004
rect 7064 7964 7070 7976
rect 7834 7964 7840 7976
rect 7892 7964 7898 8016
rect 7926 7964 7932 8016
rect 7984 7964 7990 8016
rect 4985 7939 5043 7945
rect 4985 7936 4997 7939
rect 4264 7908 4997 7936
rect 4985 7905 4997 7908
rect 5031 7905 5043 7939
rect 6914 7936 6920 7948
rect 4985 7899 5043 7905
rect 5929 7908 6920 7936
rect 2832 7840 3096 7868
rect 3145 7871 3203 7877
rect 2832 7828 2838 7840
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3510 7868 3516 7880
rect 3145 7831 3203 7837
rect 3252 7840 3516 7868
rect 750 7760 756 7812
rect 808 7800 814 7812
rect 808 7772 2176 7800
rect 808 7760 814 7772
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 2038 7732 2044 7744
rect 1636 7704 2044 7732
rect 1636 7692 1642 7704
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2148 7732 2176 7772
rect 2915 7735 2973 7741
rect 2915 7732 2927 7735
rect 2148 7704 2927 7732
rect 2915 7701 2927 7704
rect 2961 7732 2973 7735
rect 3252 7732 3280 7840
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 3786 7828 3792 7880
rect 3844 7868 3850 7880
rect 4157 7871 4215 7877
rect 3844 7840 4016 7868
rect 3844 7828 3850 7840
rect 3329 7803 3387 7809
rect 3329 7769 3341 7803
rect 3375 7769 3387 7803
rect 3329 7763 3387 7769
rect 2961 7704 3280 7732
rect 3344 7732 3372 7763
rect 3602 7760 3608 7812
rect 3660 7800 3666 7812
rect 3881 7803 3939 7809
rect 3881 7800 3893 7803
rect 3660 7772 3893 7800
rect 3660 7760 3666 7772
rect 3881 7769 3893 7772
rect 3927 7769 3939 7803
rect 3988 7800 4016 7840
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4801 7871 4859 7877
rect 4203 7840 4384 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4356 7812 4384 7840
rect 4801 7837 4813 7871
rect 4847 7864 4859 7871
rect 5929 7868 5957 7908
rect 6914 7896 6920 7908
rect 6972 7896 6978 7948
rect 7742 7936 7748 7948
rect 7703 7908 7748 7936
rect 7742 7896 7748 7908
rect 7800 7896 7806 7948
rect 4899 7864 5957 7868
rect 4847 7840 5957 7864
rect 7009 7871 7067 7877
rect 4847 7837 4927 7840
rect 4801 7836 4927 7837
rect 7009 7837 7021 7871
rect 7055 7837 7067 7871
rect 4801 7831 4859 7836
rect 7009 7831 7067 7837
rect 4065 7803 4123 7809
rect 4065 7800 4077 7803
rect 3988 7772 4077 7800
rect 3881 7763 3939 7769
rect 4065 7769 4077 7772
rect 4111 7769 4123 7803
rect 4065 7763 4123 7769
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 4522 7760 4528 7812
rect 4580 7800 4586 7812
rect 4580 7772 5396 7800
rect 4580 7760 4586 7772
rect 4614 7732 4620 7744
rect 3344 7704 4620 7732
rect 2961 7701 2973 7704
rect 2915 7695 2973 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 4893 7735 4951 7741
rect 4893 7701 4905 7735
rect 4939 7732 4951 7735
rect 5258 7732 5264 7744
rect 4939 7704 5264 7732
rect 4939 7701 4951 7704
rect 4893 7695 4951 7701
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 5368 7732 5396 7772
rect 5902 7760 5908 7812
rect 5960 7800 5966 7812
rect 7024 7800 7052 7831
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7374 7868 7380 7880
rect 7156 7840 7380 7868
rect 7156 7828 7162 7840
rect 7374 7828 7380 7840
rect 7432 7868 7438 7880
rect 7469 7871 7527 7877
rect 7469 7868 7481 7871
rect 7432 7840 7481 7868
rect 7432 7828 7438 7840
rect 7469 7837 7481 7840
rect 7515 7837 7527 7871
rect 7469 7831 7527 7837
rect 7558 7828 7564 7880
rect 7616 7868 7622 7880
rect 7929 7871 7987 7877
rect 7929 7868 7941 7871
rect 7616 7840 7941 7868
rect 7616 7828 7622 7840
rect 7929 7837 7941 7840
rect 7975 7868 7987 7871
rect 8067 7868 8095 8044
rect 11238 8032 11244 8044
rect 11296 8032 11302 8084
rect 11698 8032 11704 8084
rect 11756 8072 11762 8084
rect 13814 8072 13820 8084
rect 11756 8044 13820 8072
rect 11756 8032 11762 8044
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 15841 8075 15899 8081
rect 15841 8041 15853 8075
rect 15887 8072 15899 8075
rect 17310 8072 17316 8084
rect 15887 8044 17316 8072
rect 15887 8041 15899 8044
rect 15841 8035 15899 8041
rect 17310 8032 17316 8044
rect 17368 8032 17374 8084
rect 10778 8004 10784 8016
rect 8956 7976 10784 8004
rect 8386 7896 8392 7948
rect 8444 7936 8450 7948
rect 8956 7945 8984 7976
rect 10778 7964 10784 7976
rect 10836 7964 10842 8016
rect 10873 8007 10931 8013
rect 10873 7973 10885 8007
rect 10919 8004 10931 8007
rect 10919 7976 11376 8004
rect 10919 7973 10931 7976
rect 10873 7967 10931 7973
rect 11348 7948 11376 7976
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 8444 7908 8953 7936
rect 8444 7896 8450 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 10226 7936 10232 7948
rect 8941 7899 8999 7905
rect 9508 7908 10232 7936
rect 7975 7840 8095 7868
rect 8251 7871 8309 7877
rect 7975 7837 7987 7840
rect 7929 7831 7987 7837
rect 8251 7837 8263 7871
rect 8297 7837 8309 7871
rect 9214 7868 9220 7880
rect 9175 7840 9220 7868
rect 8251 7831 8309 7837
rect 5960 7772 7052 7800
rect 5960 7760 5966 7772
rect 7190 7760 7196 7812
rect 7248 7800 7254 7812
rect 7248 7772 7532 7800
rect 7248 7760 7254 7772
rect 6454 7732 6460 7744
rect 5368 7704 6460 7732
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 7098 7732 7104 7744
rect 7059 7704 7104 7732
rect 7098 7692 7104 7704
rect 7156 7692 7162 7744
rect 7504 7732 7532 7772
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 8266 7800 8294 7831
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 7708 7772 8294 7800
rect 7708 7760 7714 7772
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7504 7704 7573 7732
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 7926 7692 7932 7744
rect 7984 7732 7990 7744
rect 9508 7732 9536 7908
rect 10226 7896 10232 7908
rect 10284 7896 10290 7948
rect 11330 7896 11336 7948
rect 11388 7936 11394 7948
rect 12345 7939 12403 7945
rect 12345 7936 12357 7939
rect 11388 7908 12357 7936
rect 11388 7896 11394 7908
rect 12345 7905 12357 7908
rect 12391 7905 12403 7939
rect 12345 7899 12403 7905
rect 16025 7939 16083 7945
rect 16025 7905 16037 7939
rect 16071 7905 16083 7939
rect 16206 7936 16212 7948
rect 16167 7908 16212 7936
rect 16025 7899 16083 7905
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7868 10379 7871
rect 10410 7868 10416 7880
rect 10367 7840 10416 7868
rect 10367 7837 10379 7840
rect 10321 7831 10379 7837
rect 10410 7828 10416 7840
rect 10468 7828 10474 7880
rect 12612 7871 12670 7877
rect 10989 7840 12204 7868
rect 9582 7760 9588 7812
rect 9640 7800 9646 7812
rect 10989 7800 11017 7840
rect 9640 7772 11017 7800
rect 9640 7760 9646 7772
rect 11054 7760 11060 7812
rect 11112 7800 11118 7812
rect 11330 7800 11336 7812
rect 11112 7772 11336 7800
rect 11112 7760 11118 7772
rect 11330 7760 11336 7772
rect 11388 7760 11394 7812
rect 12176 7809 12204 7840
rect 12612 7837 12624 7871
rect 12658 7868 12670 7871
rect 13538 7868 13544 7880
rect 12658 7840 13544 7868
rect 12658 7837 12670 7840
rect 12612 7831 12670 7837
rect 13538 7828 13544 7840
rect 13596 7828 13602 7880
rect 13998 7828 14004 7880
rect 14056 7868 14062 7880
rect 14093 7871 14151 7877
rect 14093 7868 14105 7871
rect 14056 7840 14105 7868
rect 14056 7828 14062 7840
rect 14093 7837 14105 7840
rect 14139 7837 14151 7871
rect 14093 7831 14151 7837
rect 14182 7828 14188 7880
rect 14240 7868 14246 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14240 7840 14473 7868
rect 14240 7828 14246 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14550 7828 14556 7880
rect 14608 7868 14614 7880
rect 14728 7871 14786 7877
rect 14728 7868 14740 7871
rect 14608 7840 14740 7868
rect 14608 7828 14614 7840
rect 14728 7837 14740 7840
rect 14774 7868 14786 7871
rect 16040 7868 16068 7899
rect 16206 7896 16212 7908
rect 16264 7896 16270 7948
rect 17218 7896 17224 7948
rect 17276 7936 17282 7948
rect 17313 7939 17371 7945
rect 17313 7936 17325 7939
rect 17276 7908 17325 7936
rect 17276 7896 17282 7908
rect 17313 7905 17325 7908
rect 17359 7936 17371 7939
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17359 7908 18153 7936
rect 17359 7905 17371 7908
rect 17313 7899 17371 7905
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 17494 7868 17500 7880
rect 14774 7840 17500 7868
rect 14774 7837 14786 7840
rect 14728 7831 14786 7837
rect 17494 7828 17500 7840
rect 17552 7828 17558 7880
rect 17954 7828 17960 7880
rect 18012 7868 18018 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 18012 7840 18061 7868
rect 18012 7828 18018 7840
rect 18049 7837 18061 7840
rect 18095 7868 18107 7871
rect 19426 7868 19432 7880
rect 18095 7840 19432 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 19426 7828 19432 7840
rect 19484 7828 19490 7880
rect 12161 7803 12219 7809
rect 12161 7769 12173 7803
rect 12207 7800 12219 7803
rect 12710 7800 12716 7812
rect 12207 7772 12716 7800
rect 12207 7769 12219 7772
rect 12161 7763 12219 7769
rect 12710 7760 12716 7772
rect 12768 7760 12774 7812
rect 16301 7803 16359 7809
rect 13556 7772 14136 7800
rect 9861 7735 9919 7741
rect 9861 7732 9873 7735
rect 7984 7704 9873 7732
rect 7984 7692 7990 7704
rect 9861 7701 9873 7704
rect 9907 7701 9919 7735
rect 9861 7695 9919 7701
rect 10137 7735 10195 7741
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 10870 7732 10876 7744
rect 10183 7704 10876 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 10870 7692 10876 7704
rect 10928 7692 10934 7744
rect 11238 7692 11244 7744
rect 11296 7732 11302 7744
rect 13556 7732 13584 7772
rect 14108 7744 14136 7772
rect 16301 7769 16313 7803
rect 16347 7800 16359 7803
rect 16347 7772 16804 7800
rect 16347 7769 16359 7772
rect 16301 7763 16359 7769
rect 13722 7732 13728 7744
rect 11296 7704 13584 7732
rect 13683 7704 13728 7732
rect 11296 7692 11302 7704
rect 13722 7692 13728 7704
rect 13780 7692 13786 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 13872 7704 13917 7732
rect 13872 7692 13878 7704
rect 14090 7692 14096 7744
rect 14148 7692 14154 7744
rect 14277 7735 14335 7741
rect 14277 7701 14289 7735
rect 14323 7732 14335 7735
rect 14734 7732 14740 7744
rect 14323 7704 14740 7732
rect 14323 7701 14335 7704
rect 14277 7695 14335 7701
rect 14734 7692 14740 7704
rect 14792 7692 14798 7744
rect 16666 7732 16672 7744
rect 16627 7704 16672 7732
rect 16666 7692 16672 7704
rect 16724 7692 16730 7744
rect 16776 7741 16804 7772
rect 16942 7760 16948 7812
rect 17000 7800 17006 7812
rect 17221 7803 17279 7809
rect 17221 7800 17233 7803
rect 17000 7772 17233 7800
rect 17000 7760 17006 7772
rect 17221 7769 17233 7772
rect 17267 7769 17279 7803
rect 17221 7763 17279 7769
rect 16761 7735 16819 7741
rect 16761 7701 16773 7735
rect 16807 7701 16819 7735
rect 16761 7695 16819 7701
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 17129 7735 17187 7741
rect 17129 7732 17141 7735
rect 16908 7704 17141 7732
rect 16908 7692 16914 7704
rect 17129 7701 17141 7704
rect 17175 7701 17187 7735
rect 17586 7732 17592 7744
rect 17547 7704 17592 7732
rect 17129 7695 17187 7701
rect 17586 7692 17592 7704
rect 17644 7692 17650 7744
rect 17954 7732 17960 7744
rect 17915 7704 17960 7732
rect 17954 7692 17960 7704
rect 18012 7692 18018 7744
rect 18509 7735 18567 7741
rect 18509 7701 18521 7735
rect 18555 7732 18567 7735
rect 18782 7732 18788 7744
rect 18555 7704 18788 7732
rect 18555 7701 18567 7704
rect 18509 7695 18567 7701
rect 18782 7692 18788 7704
rect 18840 7692 18846 7744
rect 1104 7642 18860 7664
rect 1104 7590 5398 7642
rect 5450 7590 5462 7642
rect 5514 7590 5526 7642
rect 5578 7590 5590 7642
rect 5642 7590 5654 7642
rect 5706 7590 9846 7642
rect 9898 7590 9910 7642
rect 9962 7590 9974 7642
rect 10026 7590 10038 7642
rect 10090 7590 10102 7642
rect 10154 7590 14294 7642
rect 14346 7590 14358 7642
rect 14410 7590 14422 7642
rect 14474 7590 14486 7642
rect 14538 7590 14550 7642
rect 14602 7590 18860 7642
rect 1104 7568 18860 7590
rect 934 7488 940 7540
rect 992 7528 998 7540
rect 1394 7528 1400 7540
rect 992 7500 1400 7528
rect 992 7488 998 7500
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 2130 7488 2136 7540
rect 2188 7528 2194 7540
rect 2314 7528 2320 7540
rect 2188 7500 2320 7528
rect 2188 7488 2194 7500
rect 2314 7488 2320 7500
rect 2372 7488 2378 7540
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 3050 7528 3056 7540
rect 2547 7500 3056 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 3050 7488 3056 7500
rect 3108 7488 3114 7540
rect 4246 7528 4252 7540
rect 3160 7500 4252 7528
rect 1946 7420 1952 7472
rect 2004 7460 2010 7472
rect 3160 7460 3188 7500
rect 4246 7488 4252 7500
rect 4304 7488 4310 7540
rect 4893 7531 4951 7537
rect 4893 7497 4905 7531
rect 4939 7528 4951 7531
rect 5258 7528 5264 7540
rect 4939 7500 5264 7528
rect 4939 7497 4951 7500
rect 4893 7491 4951 7497
rect 5258 7488 5264 7500
rect 5316 7488 5322 7540
rect 6362 7528 6368 7540
rect 5460 7500 6368 7528
rect 5460 7472 5488 7500
rect 6362 7488 6368 7500
rect 6420 7488 6426 7540
rect 6914 7488 6920 7540
rect 6972 7528 6978 7540
rect 8021 7531 8079 7537
rect 8021 7528 8033 7531
rect 6972 7500 8033 7528
rect 6972 7488 6978 7500
rect 8021 7497 8033 7500
rect 8067 7497 8079 7531
rect 8021 7491 8079 7497
rect 8205 7531 8263 7537
rect 8205 7497 8217 7531
rect 8251 7497 8263 7531
rect 8846 7528 8852 7540
rect 8807 7500 8852 7528
rect 8205 7491 8263 7497
rect 2004 7432 3188 7460
rect 2004 7420 2010 7432
rect 3970 7420 3976 7472
rect 4028 7460 4034 7472
rect 4028 7432 4936 7460
rect 4028 7420 4034 7432
rect 4908 7404 4936 7432
rect 5442 7420 5448 7472
rect 5500 7420 5506 7472
rect 5629 7463 5687 7469
rect 5629 7429 5641 7463
rect 5675 7460 5687 7463
rect 5718 7460 5724 7472
rect 5675 7432 5724 7460
rect 5675 7429 5687 7432
rect 5629 7423 5687 7429
rect 5718 7420 5724 7432
rect 5776 7420 5782 7472
rect 6822 7420 6828 7472
rect 6880 7460 6886 7472
rect 6880 7432 7788 7460
rect 6880 7420 6886 7432
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 2130 7392 2136 7404
rect 2091 7364 2136 7392
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2498 7352 2504 7404
rect 2556 7392 2562 7404
rect 2593 7395 2651 7401
rect 2593 7392 2605 7395
rect 2556 7364 2605 7392
rect 2556 7352 2562 7364
rect 2593 7361 2605 7364
rect 2639 7392 2651 7395
rect 2958 7392 2964 7404
rect 2639 7364 2964 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2958 7352 2964 7364
rect 3016 7352 3022 7404
rect 4338 7392 4344 7404
rect 4299 7364 4344 7392
rect 4338 7352 4344 7364
rect 4396 7352 4402 7404
rect 4801 7395 4859 7401
rect 4801 7361 4813 7395
rect 4847 7361 4859 7395
rect 4801 7355 4859 7361
rect 1762 7284 1768 7336
rect 1820 7324 1826 7336
rect 1857 7327 1915 7333
rect 1857 7324 1869 7327
rect 1820 7296 1869 7324
rect 1820 7284 1826 7296
rect 1857 7293 1869 7296
rect 1903 7293 1915 7327
rect 1857 7287 1915 7293
rect 2041 7327 2099 7333
rect 2041 7293 2053 7327
rect 2087 7324 2099 7327
rect 2682 7324 2688 7336
rect 2087 7296 2688 7324
rect 2087 7293 2099 7296
rect 2041 7287 2099 7293
rect 2682 7284 2688 7296
rect 2740 7284 2746 7336
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4430 7324 4436 7336
rect 4212 7296 4436 7324
rect 4212 7284 4218 7296
rect 4430 7284 4436 7296
rect 4488 7284 4494 7336
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 4816 7324 4844 7355
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 7489 7395 7547 7401
rect 7489 7392 7501 7395
rect 5092 7364 7501 7392
rect 5092 7333 5120 7364
rect 4672 7296 4844 7324
rect 5077 7327 5135 7333
rect 4672 7284 4678 7296
rect 5077 7293 5089 7327
rect 5123 7293 5135 7327
rect 5077 7287 5135 7293
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 5920 7333 5948 7364
rect 7489 7361 7501 7364
rect 7535 7392 7547 7395
rect 7650 7392 7656 7404
rect 7535 7364 7656 7392
rect 7535 7361 7547 7364
rect 7489 7355 7547 7361
rect 7650 7352 7656 7364
rect 7708 7352 7714 7404
rect 7760 7401 7788 7432
rect 7926 7420 7932 7472
rect 7984 7460 7990 7472
rect 8220 7460 8248 7491
rect 8846 7488 8852 7500
rect 8904 7488 8910 7540
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 11330 7528 11336 7540
rect 11072 7500 11336 7528
rect 11072 7469 11100 7500
rect 11330 7488 11336 7500
rect 11388 7488 11394 7540
rect 12894 7528 12900 7540
rect 12855 7500 12900 7528
rect 12894 7488 12900 7500
rect 12952 7488 12958 7540
rect 13906 7488 13912 7540
rect 13964 7528 13970 7540
rect 14829 7531 14887 7537
rect 14829 7528 14841 7531
rect 13964 7500 14841 7528
rect 13964 7488 13970 7500
rect 14829 7497 14841 7500
rect 14875 7497 14887 7531
rect 14829 7491 14887 7497
rect 15470 7488 15476 7540
rect 15528 7528 15534 7540
rect 15657 7531 15715 7537
rect 15657 7528 15669 7531
rect 15528 7500 15669 7528
rect 15528 7488 15534 7500
rect 15657 7497 15669 7500
rect 15703 7497 15715 7531
rect 16942 7528 16948 7540
rect 15657 7491 15715 7497
rect 16040 7500 16948 7528
rect 7984 7432 8248 7460
rect 11057 7463 11115 7469
rect 7984 7420 7990 7432
rect 11057 7429 11069 7463
rect 11103 7429 11115 7463
rect 11698 7460 11704 7472
rect 11057 7423 11115 7429
rect 11164 7432 11704 7460
rect 7745 7395 7803 7401
rect 7745 7361 7757 7395
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 7834 7352 7840 7404
rect 7892 7392 7898 7404
rect 8389 7395 8447 7401
rect 8389 7392 8401 7395
rect 7892 7364 7937 7392
rect 8036 7364 8401 7392
rect 7892 7352 7898 7364
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5684 7296 5733 7324
rect 5684 7284 5690 7296
rect 5721 7293 5733 7296
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 5905 7327 5963 7333
rect 5905 7293 5917 7327
rect 5951 7293 5963 7327
rect 7668 7324 7696 7352
rect 7926 7324 7932 7336
rect 7668 7296 7932 7324
rect 5905 7287 5963 7293
rect 7926 7284 7932 7296
rect 7984 7284 7990 7336
rect 382 7216 388 7268
rect 440 7256 446 7268
rect 6089 7259 6147 7265
rect 6089 7256 6101 7259
rect 440 7228 6101 7256
rect 440 7216 446 7228
rect 6089 7225 6101 7228
rect 6135 7225 6147 7259
rect 6089 7219 6147 7225
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 4430 7188 4436 7200
rect 4391 7160 4436 7188
rect 4430 7148 4436 7160
rect 4488 7148 4494 7200
rect 4522 7148 4528 7200
rect 4580 7188 4586 7200
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4580 7160 5273 7188
rect 4580 7148 4586 7160
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 6104 7188 6132 7219
rect 8036 7188 8064 7364
rect 8389 7361 8401 7364
rect 8435 7361 8447 7395
rect 8389 7355 8447 7361
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 10410 7392 10416 7404
rect 8987 7364 10416 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 11164 7401 11192 7432
rect 11698 7420 11704 7432
rect 11756 7420 11762 7472
rect 16040 7469 16068 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17037 7531 17095 7537
rect 17037 7497 17049 7531
rect 17083 7528 17095 7531
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 17083 7500 17509 7528
rect 17083 7497 17095 7500
rect 17037 7491 17095 7497
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 17497 7491 17555 7497
rect 17586 7488 17592 7540
rect 17644 7528 17650 7540
rect 17957 7531 18015 7537
rect 17957 7528 17969 7531
rect 17644 7500 17969 7528
rect 17644 7488 17650 7500
rect 17957 7497 17969 7500
rect 18003 7497 18015 7531
rect 17957 7491 18015 7497
rect 16025 7463 16083 7469
rect 16025 7460 16037 7463
rect 15120 7432 16037 7460
rect 11790 7401 11796 7404
rect 11149 7395 11207 7401
rect 11149 7361 11161 7395
rect 11195 7361 11207 7395
rect 11784 7392 11796 7401
rect 11751 7364 11796 7392
rect 11149 7355 11207 7361
rect 11784 7355 11796 7364
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7324 9183 7327
rect 9674 7324 9680 7336
rect 9171 7296 9680 7324
rect 9171 7293 9183 7296
rect 9125 7287 9183 7293
rect 9674 7284 9680 7296
rect 9732 7284 9738 7336
rect 9766 7284 9772 7336
rect 9824 7324 9830 7336
rect 11164 7324 11192 7355
rect 11790 7352 11796 7355
rect 11848 7352 11854 7404
rect 12710 7352 12716 7404
rect 12768 7392 12774 7404
rect 12989 7395 13047 7401
rect 12989 7392 13001 7395
rect 12768 7364 13001 7392
rect 12768 7352 12774 7364
rect 12989 7361 13001 7364
rect 13035 7361 13047 7395
rect 12989 7355 13047 7361
rect 13170 7352 13176 7404
rect 13228 7392 13234 7404
rect 15120 7392 15148 7432
rect 16025 7429 16037 7432
rect 16071 7429 16083 7463
rect 16025 7423 16083 7429
rect 16117 7463 16175 7469
rect 16117 7429 16129 7463
rect 16163 7460 16175 7463
rect 16206 7460 16212 7472
rect 16163 7432 16212 7460
rect 16163 7429 16175 7432
rect 16117 7423 16175 7429
rect 16206 7420 16212 7432
rect 16264 7420 16270 7472
rect 16666 7420 16672 7472
rect 16724 7460 16730 7472
rect 17129 7463 17187 7469
rect 17129 7460 17141 7463
rect 16724 7432 17141 7460
rect 16724 7420 16730 7432
rect 17129 7429 17141 7432
rect 17175 7429 17187 7463
rect 17129 7423 17187 7429
rect 13228 7364 15148 7392
rect 15197 7395 15255 7401
rect 13228 7352 13234 7364
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 15470 7392 15476 7404
rect 15243 7364 15476 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 15470 7352 15476 7364
rect 15528 7352 15534 7404
rect 17862 7392 17868 7404
rect 17823 7364 17868 7392
rect 17862 7352 17868 7364
rect 17920 7352 17926 7404
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 18509 7395 18567 7401
rect 18509 7392 18521 7395
rect 18012 7364 18521 7392
rect 18012 7352 18018 7364
rect 18509 7361 18521 7364
rect 18555 7361 18567 7395
rect 18509 7355 18567 7361
rect 9824 7296 11192 7324
rect 9824 7284 9830 7296
rect 11238 7284 11244 7336
rect 11296 7324 11302 7336
rect 11517 7327 11575 7333
rect 11517 7324 11529 7327
rect 11296 7296 11529 7324
rect 11296 7284 11302 7296
rect 11517 7293 11529 7296
rect 11563 7293 11575 7327
rect 15102 7324 15108 7336
rect 11517 7287 11575 7293
rect 13280 7296 15108 7324
rect 8478 7188 8484 7200
rect 6104 7160 8064 7188
rect 8439 7160 8484 7188
rect 5261 7151 5319 7157
rect 8478 7148 8484 7160
rect 8536 7148 8542 7200
rect 11333 7191 11391 7197
rect 11333 7157 11345 7191
rect 11379 7188 11391 7191
rect 13280 7188 13308 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15286 7324 15292 7336
rect 15247 7296 15292 7324
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 15381 7327 15439 7333
rect 15381 7293 15393 7327
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 16209 7327 16267 7333
rect 16209 7293 16221 7327
rect 16255 7293 16267 7327
rect 17310 7324 17316 7336
rect 17271 7296 17316 7324
rect 16209 7287 16267 7293
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 15194 7256 15200 7268
rect 13780 7228 15200 7256
rect 13780 7216 13786 7228
rect 15194 7216 15200 7228
rect 15252 7256 15258 7268
rect 15396 7256 15424 7287
rect 16224 7256 16252 7287
rect 17310 7284 17316 7296
rect 17368 7284 17374 7336
rect 17494 7284 17500 7336
rect 17552 7324 17558 7336
rect 18049 7327 18107 7333
rect 18049 7324 18061 7327
rect 17552 7296 18061 7324
rect 17552 7284 17558 7296
rect 18049 7293 18061 7296
rect 18095 7293 18107 7327
rect 18049 7287 18107 7293
rect 16666 7256 16672 7268
rect 15252 7228 16252 7256
rect 16627 7228 16672 7256
rect 15252 7216 15258 7228
rect 16666 7216 16672 7228
rect 16724 7216 16730 7268
rect 11379 7160 13308 7188
rect 11379 7157 11391 7160
rect 11333 7151 11391 7157
rect 13998 7148 14004 7200
rect 14056 7188 14062 7200
rect 14182 7188 14188 7200
rect 14056 7160 14188 7188
rect 14056 7148 14062 7160
rect 14182 7148 14188 7160
rect 14240 7188 14246 7200
rect 14277 7191 14335 7197
rect 14277 7188 14289 7191
rect 14240 7160 14289 7188
rect 14240 7148 14246 7160
rect 14277 7157 14289 7160
rect 14323 7157 14335 7191
rect 14277 7151 14335 7157
rect 18230 7148 18236 7200
rect 18288 7188 18294 7200
rect 18325 7191 18383 7197
rect 18325 7188 18337 7191
rect 18288 7160 18337 7188
rect 18288 7148 18294 7160
rect 18325 7157 18337 7160
rect 18371 7157 18383 7191
rect 18325 7151 18383 7157
rect 1104 7098 18860 7120
rect 1104 7046 3174 7098
rect 3226 7046 3238 7098
rect 3290 7046 3302 7098
rect 3354 7046 3366 7098
rect 3418 7046 3430 7098
rect 3482 7046 7622 7098
rect 7674 7046 7686 7098
rect 7738 7046 7750 7098
rect 7802 7046 7814 7098
rect 7866 7046 7878 7098
rect 7930 7046 12070 7098
rect 12122 7046 12134 7098
rect 12186 7046 12198 7098
rect 12250 7046 12262 7098
rect 12314 7046 12326 7098
rect 12378 7046 16518 7098
rect 16570 7046 16582 7098
rect 16634 7046 16646 7098
rect 16698 7046 16710 7098
rect 16762 7046 16774 7098
rect 16826 7046 18860 7098
rect 1104 7024 18860 7046
rect 4724 6956 5212 6984
rect 2869 6919 2927 6925
rect 2869 6885 2881 6919
rect 2915 6916 2927 6919
rect 3142 6916 3148 6928
rect 2915 6888 3148 6916
rect 2915 6885 2927 6888
rect 2869 6879 2927 6885
rect 3142 6876 3148 6888
rect 3200 6876 3206 6928
rect 4614 6916 4620 6928
rect 4172 6888 4620 6916
rect 14 6808 20 6860
rect 72 6848 78 6860
rect 934 6848 940 6860
rect 72 6820 940 6848
rect 72 6808 78 6820
rect 934 6808 940 6820
rect 992 6808 998 6860
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 4172 6857 4200 6888
rect 4614 6876 4620 6888
rect 4672 6876 4678 6928
rect 4724 6925 4752 6956
rect 4709 6919 4767 6925
rect 4709 6885 4721 6919
rect 4755 6885 4767 6919
rect 4709 6879 4767 6885
rect 4801 6919 4859 6925
rect 4801 6885 4813 6919
rect 4847 6916 4859 6919
rect 4982 6916 4988 6928
rect 4847 6888 4988 6916
rect 4847 6885 4859 6888
rect 4801 6879 4859 6885
rect 4982 6876 4988 6888
rect 5040 6876 5046 6928
rect 3789 6851 3847 6857
rect 3789 6848 3801 6851
rect 3476 6820 3801 6848
rect 3476 6808 3482 6820
rect 3789 6817 3801 6820
rect 3835 6817 3847 6851
rect 3789 6811 3847 6817
rect 4157 6851 4215 6857
rect 4157 6817 4169 6851
rect 4203 6817 4215 6851
rect 4157 6811 4215 6817
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4430 6848 4436 6860
rect 4295 6820 4436 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4430 6808 4436 6820
rect 4488 6808 4494 6860
rect 4632 6820 5120 6848
rect 1489 6783 1547 6789
rect 1489 6749 1501 6783
rect 1535 6780 1547 6783
rect 2498 6780 2504 6792
rect 1535 6752 2504 6780
rect 1535 6749 1547 6752
rect 1489 6743 1547 6749
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 3605 6783 3663 6789
rect 3605 6749 3617 6783
rect 3651 6749 3663 6783
rect 3605 6743 3663 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4522 6780 4528 6792
rect 4387 6752 4528 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 1578 6672 1584 6724
rect 1636 6712 1642 6724
rect 1734 6715 1792 6721
rect 1734 6712 1746 6715
rect 1636 6684 1746 6712
rect 1636 6672 1642 6684
rect 1734 6681 1746 6684
rect 1780 6681 1792 6715
rect 3620 6712 3648 6743
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4632 6712 4660 6820
rect 3620 6684 4660 6712
rect 1734 6675 1792 6681
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3418 6644 3424 6656
rect 3007 6616 3424 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3510 6604 3516 6656
rect 3568 6644 3574 6656
rect 4614 6644 4620 6656
rect 3568 6616 4620 6644
rect 3568 6604 3574 6616
rect 4614 6604 4620 6616
rect 4672 6604 4678 6656
rect 5092 6644 5120 6820
rect 5184 6780 5212 6956
rect 6638 6944 6644 6996
rect 6696 6984 6702 6996
rect 7190 6984 7196 6996
rect 6696 6956 7052 6984
rect 7151 6956 7196 6984
rect 6696 6944 6702 6956
rect 6270 6876 6276 6928
rect 6328 6916 6334 6928
rect 6365 6919 6423 6925
rect 6365 6916 6377 6919
rect 6328 6888 6377 6916
rect 6328 6876 6334 6888
rect 6365 6885 6377 6888
rect 6411 6885 6423 6919
rect 6365 6879 6423 6885
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 6788 6888 6960 6916
rect 6788 6876 6794 6888
rect 6181 6851 6239 6857
rect 6181 6817 6193 6851
rect 6227 6848 6239 6851
rect 6822 6848 6828 6860
rect 6227 6820 6828 6848
rect 6227 6817 6239 6820
rect 6181 6811 6239 6817
rect 6822 6808 6828 6820
rect 6880 6808 6886 6860
rect 6932 6857 6960 6888
rect 6917 6851 6975 6857
rect 6917 6817 6929 6851
rect 6963 6817 6975 6851
rect 7024 6848 7052 6956
rect 7190 6944 7196 6956
rect 7248 6944 7254 6996
rect 7585 6956 8156 6984
rect 7585 6928 7613 6956
rect 7558 6876 7564 6928
rect 7616 6876 7622 6928
rect 8128 6916 8156 6956
rect 8248 6944 8254 6996
rect 8306 6984 8312 6996
rect 10410 6984 10416 6996
rect 8306 6956 8892 6984
rect 10371 6956 10416 6984
rect 8306 6944 8312 6956
rect 8386 6916 8392 6928
rect 8128 6888 8392 6916
rect 8386 6876 8392 6888
rect 8444 6876 8450 6928
rect 7653 6851 7711 6857
rect 7653 6848 7665 6851
rect 7024 6820 7665 6848
rect 6917 6811 6975 6817
rect 7653 6817 7665 6820
rect 7699 6817 7711 6851
rect 7653 6811 7711 6817
rect 7837 6851 7895 6857
rect 7837 6817 7849 6851
rect 7883 6817 7895 6851
rect 7837 6811 7895 6817
rect 6733 6783 6791 6789
rect 6733 6780 6745 6783
rect 5184 6752 6745 6780
rect 6733 6749 6745 6752
rect 6779 6749 6791 6783
rect 7558 6780 7564 6792
rect 7519 6752 7564 6780
rect 6733 6743 6791 6749
rect 7558 6740 7564 6752
rect 7616 6740 7622 6792
rect 7852 6780 7880 6811
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 8113 6851 8171 6857
rect 8113 6848 8125 6851
rect 7984 6820 8125 6848
rect 7984 6808 7990 6820
rect 8113 6817 8125 6820
rect 8159 6817 8171 6851
rect 8113 6811 8171 6817
rect 8297 6851 8355 6857
rect 8297 6817 8309 6851
rect 8343 6848 8355 6851
rect 8478 6848 8484 6860
rect 8343 6820 8484 6848
rect 8343 6817 8355 6820
rect 8297 6811 8355 6817
rect 8478 6808 8484 6820
rect 8536 6808 8542 6860
rect 8864 6848 8892 6956
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 13170 6984 13176 6996
rect 12860 6956 13176 6984
rect 12860 6944 12866 6956
rect 13170 6944 13176 6956
rect 13228 6944 13234 6996
rect 13998 6984 14004 6996
rect 13464 6956 14004 6984
rect 8864 6820 9076 6848
rect 8662 6780 8668 6792
rect 7852 6752 8668 6780
rect 8662 6740 8668 6752
rect 8720 6740 8726 6792
rect 5936 6715 5994 6721
rect 5936 6681 5948 6715
rect 5982 6712 5994 6715
rect 6086 6712 6092 6724
rect 5982 6684 6092 6712
rect 5982 6681 5994 6684
rect 5936 6675 5994 6681
rect 6086 6672 6092 6684
rect 6144 6672 6150 6724
rect 7926 6712 7932 6724
rect 6380 6684 7932 6712
rect 6380 6644 6408 6684
rect 7926 6672 7932 6684
rect 7984 6672 7990 6724
rect 8281 6684 8984 6712
rect 5092 6616 6408 6644
rect 6454 6604 6460 6656
rect 6512 6644 6518 6656
rect 6825 6647 6883 6653
rect 6825 6644 6837 6647
rect 6512 6616 6837 6644
rect 6512 6604 6518 6616
rect 6825 6613 6837 6616
rect 6871 6613 6883 6647
rect 6825 6607 6883 6613
rect 7006 6604 7012 6656
rect 7064 6644 7070 6656
rect 7374 6644 7380 6656
rect 7064 6616 7380 6644
rect 7064 6604 7070 6616
rect 7374 6604 7380 6616
rect 7432 6604 7438 6656
rect 7944 6644 7972 6672
rect 8110 6644 8116 6656
rect 7944 6616 8116 6644
rect 8110 6604 8116 6616
rect 8168 6644 8174 6656
rect 8281 6644 8309 6684
rect 8386 6644 8392 6656
rect 8168 6616 8309 6644
rect 8347 6616 8392 6644
rect 8168 6604 8174 6616
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 8662 6604 8668 6656
rect 8720 6644 8726 6656
rect 8956 6653 8984 6684
rect 8757 6647 8815 6653
rect 8757 6644 8769 6647
rect 8720 6616 8769 6644
rect 8720 6604 8726 6616
rect 8757 6613 8769 6616
rect 8803 6613 8815 6647
rect 8757 6607 8815 6613
rect 8941 6647 8999 6653
rect 8941 6613 8953 6647
rect 8987 6613 8999 6647
rect 9048 6644 9076 6820
rect 10686 6808 10692 6860
rect 10744 6848 10750 6860
rect 10962 6848 10968 6860
rect 10744 6820 10968 6848
rect 10744 6808 10750 6820
rect 10962 6808 10968 6820
rect 11020 6808 11026 6860
rect 13354 6848 13360 6860
rect 12912 6820 13360 6848
rect 10321 6783 10379 6789
rect 10321 6749 10333 6783
rect 10367 6780 10379 6783
rect 11238 6780 11244 6792
rect 10367 6752 11244 6780
rect 10367 6749 10379 6752
rect 10321 6743 10379 6749
rect 11238 6740 11244 6752
rect 11296 6740 11302 6792
rect 11514 6780 11520 6792
rect 11475 6752 11520 6780
rect 11514 6740 11520 6752
rect 11572 6740 11578 6792
rect 12912 6780 12940 6820
rect 13354 6808 13360 6820
rect 13412 6808 13418 6860
rect 12406 6752 12940 6780
rect 12989 6783 13047 6789
rect 9674 6672 9680 6724
rect 9732 6712 9738 6724
rect 10054 6715 10112 6721
rect 10054 6712 10066 6715
rect 9732 6684 10066 6712
rect 9732 6672 9738 6684
rect 10054 6681 10066 6684
rect 10100 6681 10112 6715
rect 10778 6712 10784 6724
rect 10739 6684 10784 6712
rect 10054 6675 10112 6681
rect 10778 6672 10784 6684
rect 10836 6672 10842 6724
rect 12406 6712 12434 6752
rect 12989 6749 13001 6783
rect 13035 6780 13047 6783
rect 13464 6780 13492 6956
rect 13998 6944 14004 6956
rect 14056 6944 14062 6996
rect 15194 6944 15200 6996
rect 15252 6984 15258 6996
rect 15930 6984 15936 6996
rect 15252 6956 15936 6984
rect 15252 6944 15258 6956
rect 15930 6944 15936 6956
rect 15988 6944 15994 6996
rect 17862 6944 17868 6996
rect 17920 6984 17926 6996
rect 18233 6987 18291 6993
rect 18233 6984 18245 6987
rect 17920 6956 18245 6984
rect 17920 6944 17926 6956
rect 18233 6953 18245 6956
rect 18279 6953 18291 6987
rect 18233 6947 18291 6953
rect 17218 6876 17224 6928
rect 17276 6916 17282 6928
rect 17276 6888 17632 6916
rect 17276 6876 17282 6888
rect 13722 6848 13728 6860
rect 13683 6820 13728 6848
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 17604 6857 17632 6888
rect 17589 6851 17647 6857
rect 17589 6817 17601 6851
rect 17635 6817 17647 6851
rect 17770 6848 17776 6860
rect 17731 6820 17776 6848
rect 17589 6811 17647 6817
rect 17770 6808 17776 6820
rect 17828 6808 17834 6860
rect 13035 6752 13492 6780
rect 13541 6783 13599 6789
rect 13035 6749 13047 6752
rect 12989 6743 13047 6749
rect 13541 6749 13553 6783
rect 13587 6780 13599 6783
rect 13587 6752 15332 6780
rect 13587 6749 13599 6752
rect 13541 6743 13599 6749
rect 10888 6684 12434 6712
rect 12744 6715 12802 6721
rect 10888 6653 10916 6684
rect 12744 6681 12756 6715
rect 12790 6712 12802 6715
rect 13814 6712 13820 6724
rect 12790 6684 13820 6712
rect 12790 6681 12802 6684
rect 12744 6675 12802 6681
rect 13814 6672 13820 6684
rect 13872 6712 13878 6724
rect 13872 6684 14136 6712
rect 13872 6672 13878 6684
rect 10873 6647 10931 6653
rect 10873 6644 10885 6647
rect 9048 6616 10885 6644
rect 8941 6607 8999 6613
rect 10873 6613 10885 6616
rect 10919 6613 10931 6647
rect 10873 6607 10931 6613
rect 11333 6647 11391 6653
rect 11333 6613 11345 6647
rect 11379 6644 11391 6647
rect 11422 6644 11428 6656
rect 11379 6616 11428 6644
rect 11379 6613 11391 6616
rect 11333 6607 11391 6613
rect 11422 6604 11428 6616
rect 11480 6604 11486 6656
rect 11609 6647 11667 6653
rect 11609 6613 11621 6647
rect 11655 6644 11667 6647
rect 11698 6644 11704 6656
rect 11655 6616 11704 6644
rect 11655 6613 11667 6616
rect 11609 6607 11667 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 13078 6604 13084 6656
rect 13136 6644 13142 6656
rect 13173 6647 13231 6653
rect 13173 6644 13185 6647
rect 13136 6616 13185 6644
rect 13136 6604 13142 6616
rect 13173 6613 13185 6616
rect 13219 6613 13231 6647
rect 13173 6607 13231 6613
rect 13354 6604 13360 6656
rect 13412 6644 13418 6656
rect 14108 6653 14136 6684
rect 14826 6672 14832 6724
rect 14884 6712 14890 6724
rect 15206 6715 15264 6721
rect 15206 6712 15218 6715
rect 14884 6684 15218 6712
rect 14884 6672 14890 6684
rect 15206 6681 15218 6684
rect 15252 6681 15264 6715
rect 15304 6712 15332 6752
rect 15378 6740 15384 6792
rect 15436 6780 15442 6792
rect 15473 6783 15531 6789
rect 15473 6780 15485 6783
rect 15436 6752 15485 6780
rect 15436 6740 15442 6752
rect 15473 6749 15485 6752
rect 15519 6780 15531 6783
rect 15657 6783 15715 6789
rect 15657 6780 15669 6783
rect 15519 6752 15669 6780
rect 15519 6749 15531 6752
rect 15473 6743 15531 6749
rect 15657 6749 15669 6752
rect 15703 6780 15715 6783
rect 16666 6780 16672 6792
rect 15703 6752 16672 6780
rect 15703 6749 15715 6752
rect 15657 6743 15715 6749
rect 16666 6740 16672 6752
rect 16724 6740 16730 6792
rect 17126 6780 17132 6792
rect 17087 6752 17132 6780
rect 17126 6740 17132 6752
rect 17184 6740 17190 6792
rect 18966 6780 18972 6792
rect 17788 6752 18972 6780
rect 15562 6712 15568 6724
rect 15304 6684 15568 6712
rect 15206 6675 15264 6681
rect 15562 6672 15568 6684
rect 15620 6672 15626 6724
rect 15924 6715 15982 6721
rect 15924 6681 15936 6715
rect 15970 6712 15982 6715
rect 16390 6712 16396 6724
rect 15970 6684 16396 6712
rect 15970 6681 15982 6684
rect 15924 6675 15982 6681
rect 16390 6672 16396 6684
rect 16448 6672 16454 6724
rect 17788 6712 17816 6752
rect 18966 6740 18972 6752
rect 19024 6740 19030 6792
rect 16868 6684 17816 6712
rect 17865 6715 17923 6721
rect 16868 6656 16896 6684
rect 17865 6681 17877 6715
rect 17911 6712 17923 6715
rect 18325 6715 18383 6721
rect 18325 6712 18337 6715
rect 17911 6684 18337 6712
rect 17911 6681 17923 6684
rect 17865 6675 17923 6681
rect 18325 6681 18337 6684
rect 18371 6681 18383 6715
rect 18325 6675 18383 6681
rect 13633 6647 13691 6653
rect 13633 6644 13645 6647
rect 13412 6616 13645 6644
rect 13412 6604 13418 6616
rect 13633 6613 13645 6616
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 14093 6647 14151 6653
rect 14093 6613 14105 6647
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 15286 6604 15292 6656
rect 15344 6644 15350 6656
rect 16482 6644 16488 6656
rect 15344 6616 16488 6644
rect 15344 6604 15350 6616
rect 16482 6604 16488 6616
rect 16540 6604 16546 6656
rect 16850 6604 16856 6656
rect 16908 6604 16914 6656
rect 17034 6644 17040 6656
rect 16995 6616 17040 6644
rect 17034 6604 17040 6616
rect 17092 6604 17098 6656
rect 17313 6647 17371 6653
rect 17313 6613 17325 6647
rect 17359 6644 17371 6647
rect 17494 6644 17500 6656
rect 17359 6616 17500 6644
rect 17359 6613 17371 6616
rect 17313 6607 17371 6613
rect 17494 6604 17500 6616
rect 17552 6604 17558 6656
rect 1104 6554 18860 6576
rect 1104 6502 5398 6554
rect 5450 6502 5462 6554
rect 5514 6502 5526 6554
rect 5578 6502 5590 6554
rect 5642 6502 5654 6554
rect 5706 6502 9846 6554
rect 9898 6502 9910 6554
rect 9962 6502 9974 6554
rect 10026 6502 10038 6554
rect 10090 6502 10102 6554
rect 10154 6502 14294 6554
rect 14346 6502 14358 6554
rect 14410 6502 14422 6554
rect 14474 6502 14486 6554
rect 14538 6502 14550 6554
rect 14602 6502 18860 6554
rect 1104 6480 18860 6502
rect 1581 6443 1639 6449
rect 1581 6409 1593 6443
rect 1627 6440 1639 6443
rect 2130 6440 2136 6452
rect 1627 6412 2136 6440
rect 1627 6409 1639 6412
rect 1581 6403 1639 6409
rect 2130 6400 2136 6412
rect 2188 6400 2194 6452
rect 2958 6400 2964 6452
rect 3016 6440 3022 6452
rect 4525 6443 4583 6449
rect 4525 6440 4537 6443
rect 3016 6412 4537 6440
rect 3016 6400 3022 6412
rect 4525 6409 4537 6412
rect 4571 6409 4583 6443
rect 4798 6440 4804 6452
rect 4759 6412 4804 6440
rect 4525 6403 4583 6409
rect 4798 6400 4804 6412
rect 4856 6400 4862 6452
rect 4982 6400 4988 6452
rect 5040 6440 5046 6452
rect 5902 6440 5908 6452
rect 5040 6412 5908 6440
rect 5040 6400 5046 6412
rect 5902 6400 5908 6412
rect 5960 6400 5966 6452
rect 6365 6443 6423 6449
rect 6365 6409 6377 6443
rect 6411 6440 6423 6443
rect 6454 6440 6460 6452
rect 6411 6412 6460 6440
rect 6411 6409 6423 6412
rect 6365 6403 6423 6409
rect 6454 6400 6460 6412
rect 6512 6400 6518 6452
rect 6733 6443 6791 6449
rect 6733 6409 6745 6443
rect 6779 6440 6791 6443
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 6779 6412 7205 6440
rect 6779 6409 6791 6412
rect 6733 6403 6791 6409
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 7193 6403 7251 6409
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 7524 6412 7665 6440
rect 7524 6400 7530 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 8386 6400 8392 6452
rect 8444 6440 8450 6452
rect 9493 6443 9551 6449
rect 9493 6440 9505 6443
rect 8444 6412 9505 6440
rect 8444 6400 8450 6412
rect 9493 6409 9505 6412
rect 9539 6409 9551 6443
rect 9493 6403 9551 6409
rect 9766 6400 9772 6452
rect 9824 6440 9830 6452
rect 9861 6443 9919 6449
rect 9861 6440 9873 6443
rect 9824 6412 9873 6440
rect 9824 6400 9830 6412
rect 9861 6409 9873 6412
rect 9907 6409 9919 6443
rect 9861 6403 9919 6409
rect 9953 6443 10011 6449
rect 9953 6409 9965 6443
rect 9999 6440 10011 6443
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 9999 6412 10333 6440
rect 9999 6409 10011 6412
rect 9953 6403 10011 6409
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 10410 6400 10416 6452
rect 10468 6440 10474 6452
rect 10689 6443 10747 6449
rect 10689 6440 10701 6443
rect 10468 6412 10701 6440
rect 10468 6400 10474 6412
rect 10689 6409 10701 6412
rect 10735 6409 10747 6443
rect 11330 6440 11336 6452
rect 11291 6412 11336 6440
rect 10689 6403 10747 6409
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 11790 6440 11796 6452
rect 11751 6412 11796 6440
rect 11790 6400 11796 6412
rect 11848 6400 11854 6452
rect 12158 6400 12164 6452
rect 12216 6400 12222 6452
rect 12802 6440 12808 6452
rect 12656 6412 12808 6440
rect 2501 6375 2559 6381
rect 2501 6341 2513 6375
rect 2547 6372 2559 6375
rect 2866 6372 2872 6384
rect 2547 6344 2872 6372
rect 2547 6341 2559 6344
rect 2501 6335 2559 6341
rect 2866 6332 2872 6344
rect 2924 6332 2930 6384
rect 3418 6332 3424 6384
rect 3476 6372 3482 6384
rect 6825 6375 6883 6381
rect 3476 6344 6040 6372
rect 3476 6332 3482 6344
rect 1670 6264 1676 6316
rect 1728 6304 1734 6316
rect 1949 6307 2007 6313
rect 1949 6304 1961 6307
rect 1728 6276 1961 6304
rect 1728 6264 1734 6276
rect 1949 6273 1961 6276
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 2409 6307 2467 6313
rect 2409 6273 2421 6307
rect 2455 6304 2467 6307
rect 2682 6304 2688 6316
rect 2455 6276 2688 6304
rect 2455 6273 2467 6276
rect 2409 6267 2467 6273
rect 2682 6264 2688 6276
rect 2740 6264 2746 6316
rect 3142 6313 3148 6316
rect 3136 6304 3148 6313
rect 3103 6276 3148 6304
rect 3136 6267 3148 6276
rect 3142 6264 3148 6267
rect 3200 6264 3206 6316
rect 3510 6264 3516 6316
rect 3568 6304 3574 6316
rect 4341 6307 4399 6313
rect 4341 6304 4353 6307
rect 3568 6276 4353 6304
rect 3568 6264 3574 6276
rect 4341 6273 4353 6276
rect 4387 6273 4399 6307
rect 4341 6267 4399 6273
rect 4522 6264 4528 6316
rect 4580 6304 4586 6316
rect 5350 6304 5356 6316
rect 4580 6276 5356 6304
rect 4580 6264 4586 6276
rect 5350 6264 5356 6276
rect 5408 6264 5414 6316
rect 5902 6304 5908 6316
rect 5960 6313 5966 6316
rect 5872 6276 5908 6304
rect 5902 6264 5908 6276
rect 5960 6267 5972 6313
rect 6012 6304 6040 6344
rect 6825 6341 6837 6375
rect 6871 6372 6883 6375
rect 7098 6372 7104 6384
rect 6871 6344 7104 6372
rect 6871 6341 6883 6344
rect 6825 6335 6883 6341
rect 7098 6332 7104 6344
rect 7156 6332 7162 6384
rect 8266 6375 8324 6381
rect 8266 6372 8278 6375
rect 7208 6344 8278 6372
rect 7208 6304 7236 6344
rect 8266 6341 8278 6344
rect 8312 6341 8324 6375
rect 8266 6335 8324 6341
rect 7558 6304 7564 6316
rect 6012 6276 7236 6304
rect 7519 6276 7564 6304
rect 5960 6264 5966 6267
rect 7558 6264 7564 6276
rect 7616 6264 7622 6316
rect 11790 6304 11796 6316
rect 7760 6276 11796 6304
rect 1762 6196 1768 6248
rect 1820 6236 1826 6248
rect 2130 6236 2136 6248
rect 1820 6208 2136 6236
rect 1820 6196 1826 6208
rect 2130 6196 2136 6208
rect 2188 6236 2194 6248
rect 2593 6239 2651 6245
rect 2593 6236 2605 6239
rect 2188 6208 2605 6236
rect 2188 6196 2194 6208
rect 2593 6205 2605 6208
rect 2639 6205 2651 6239
rect 2593 6199 2651 6205
rect 2869 6239 2927 6245
rect 2869 6205 2881 6239
rect 2915 6205 2927 6239
rect 2869 6199 2927 6205
rect 1762 6100 1768 6112
rect 1723 6072 1768 6100
rect 1762 6060 1768 6072
rect 1820 6060 1826 6112
rect 2041 6103 2099 6109
rect 2041 6069 2053 6103
rect 2087 6100 2099 6103
rect 2406 6100 2412 6112
rect 2087 6072 2412 6100
rect 2087 6069 2099 6072
rect 2041 6063 2099 6069
rect 2406 6060 2412 6072
rect 2464 6060 2470 6112
rect 2884 6100 2912 6199
rect 4430 6196 4436 6248
rect 4488 6236 4494 6248
rect 6181 6239 6239 6245
rect 4488 6208 4568 6236
rect 4488 6196 4494 6208
rect 3970 6100 3976 6112
rect 2884 6072 3976 6100
rect 3970 6060 3976 6072
rect 4028 6060 4034 6112
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 4430 6100 4436 6112
rect 4295 6072 4436 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 4430 6060 4436 6072
rect 4488 6060 4494 6112
rect 4540 6100 4568 6208
rect 6181 6205 6193 6239
rect 6227 6205 6239 6239
rect 6181 6199 6239 6205
rect 4706 6128 4712 6180
rect 4764 6168 4770 6180
rect 5074 6168 5080 6180
rect 4764 6140 5080 6168
rect 4764 6128 4770 6140
rect 5074 6128 5080 6140
rect 5132 6128 5138 6180
rect 6196 6168 6224 6199
rect 6362 6196 6368 6248
rect 6420 6236 6426 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6420 6208 6929 6236
rect 6420 6196 6426 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 7006 6196 7012 6248
rect 7064 6236 7070 6248
rect 7760 6236 7788 6276
rect 11790 6264 11796 6276
rect 11848 6264 11854 6316
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6304 11943 6307
rect 12066 6304 12072 6316
rect 11931 6276 12072 6304
rect 11931 6273 11943 6276
rect 11885 6267 11943 6273
rect 12066 6264 12072 6276
rect 12124 6264 12130 6316
rect 7064 6208 7788 6236
rect 7064 6196 7070 6208
rect 7834 6196 7840 6248
rect 7892 6236 7898 6248
rect 8021 6239 8079 6245
rect 7892 6208 7937 6236
rect 7892 6196 7898 6208
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 8036 6168 8064 6199
rect 9674 6196 9680 6248
rect 9732 6236 9738 6248
rect 10045 6239 10103 6245
rect 10045 6236 10057 6239
rect 9732 6208 10057 6236
rect 9732 6196 9738 6208
rect 10045 6205 10057 6208
rect 10091 6205 10103 6239
rect 10045 6199 10103 6205
rect 10226 6196 10232 6248
rect 10284 6236 10290 6248
rect 10781 6239 10839 6245
rect 10781 6236 10793 6239
rect 10284 6208 10793 6236
rect 10284 6196 10290 6208
rect 10781 6205 10793 6208
rect 10827 6205 10839 6239
rect 10962 6236 10968 6248
rect 10923 6208 10968 6236
rect 10781 6199 10839 6205
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11698 6236 11704 6248
rect 11659 6208 11704 6236
rect 11698 6196 11704 6208
rect 11756 6196 11762 6248
rect 12176 6236 12204 6400
rect 12250 6264 12256 6316
rect 12308 6304 12314 6316
rect 12656 6304 12684 6412
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 13078 6400 13084 6452
rect 13136 6440 13142 6452
rect 13173 6443 13231 6449
rect 13173 6440 13185 6443
rect 13136 6412 13185 6440
rect 13136 6400 13142 6412
rect 13173 6409 13185 6412
rect 13219 6409 13231 6443
rect 13173 6403 13231 6409
rect 13280 6412 14596 6440
rect 12986 6332 12992 6384
rect 13044 6372 13050 6384
rect 13280 6372 13308 6412
rect 13044 6344 13308 6372
rect 13044 6332 13050 6344
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 14369 6375 14427 6381
rect 14369 6372 14381 6375
rect 14056 6344 14381 6372
rect 14056 6332 14062 6344
rect 14369 6341 14381 6344
rect 14415 6341 14427 6375
rect 14369 6335 14427 6341
rect 14461 6375 14519 6381
rect 14461 6341 14473 6375
rect 14507 6341 14519 6375
rect 14568 6372 14596 6412
rect 15010 6400 15016 6452
rect 15068 6440 15074 6452
rect 15105 6443 15163 6449
rect 15105 6440 15117 6443
rect 15068 6412 15117 6440
rect 15068 6400 15074 6412
rect 15105 6409 15117 6412
rect 15151 6440 15163 6443
rect 18322 6440 18328 6452
rect 15151 6412 17908 6440
rect 18283 6412 18328 6440
rect 15151 6409 15163 6412
rect 15105 6403 15163 6409
rect 15194 6372 15200 6384
rect 14568 6344 15200 6372
rect 14461 6335 14519 6341
rect 12308 6276 12684 6304
rect 12713 6307 12771 6313
rect 12308 6264 12314 6276
rect 12713 6273 12725 6307
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6304 12863 6307
rect 13446 6304 13452 6316
rect 12851 6276 13452 6304
rect 12851 6273 12863 6276
rect 12805 6267 12863 6273
rect 12176 6208 12388 6236
rect 6196 6140 8064 6168
rect 6914 6100 6920 6112
rect 4540 6072 6920 6100
rect 6914 6060 6920 6072
rect 6972 6060 6978 6112
rect 8036 6100 8064 6140
rect 9122 6128 9128 6180
rect 9180 6168 9186 6180
rect 9401 6171 9459 6177
rect 9401 6168 9413 6171
rect 9180 6140 9413 6168
rect 9180 6128 9186 6140
rect 9401 6137 9413 6140
rect 9447 6168 9459 6171
rect 11054 6168 11060 6180
rect 9447 6140 11060 6168
rect 9447 6137 9459 6140
rect 9401 6131 9459 6137
rect 11054 6128 11060 6140
rect 11112 6128 11118 6180
rect 12360 6177 12388 6208
rect 12345 6171 12403 6177
rect 12345 6137 12357 6171
rect 12391 6137 12403 6171
rect 12345 6131 12403 6137
rect 8294 6100 8300 6112
rect 8036 6072 8300 6100
rect 8294 6060 8300 6072
rect 8352 6060 8358 6112
rect 12253 6103 12311 6109
rect 12253 6069 12265 6103
rect 12299 6100 12311 6103
rect 12728 6100 12756 6267
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 13541 6307 13599 6313
rect 13541 6273 13553 6307
rect 13587 6304 13599 6307
rect 13722 6304 13728 6316
rect 13587 6276 13728 6304
rect 13587 6273 13599 6276
rect 13541 6267 13599 6273
rect 13722 6264 13728 6276
rect 13780 6264 13786 6316
rect 14476 6304 14504 6335
rect 15194 6332 15200 6344
rect 15252 6332 15258 6384
rect 15470 6332 15476 6384
rect 15528 6372 15534 6384
rect 16936 6375 16994 6381
rect 15528 6344 16252 6372
rect 15528 6332 15534 6344
rect 14476 6276 15700 6304
rect 12894 6236 12900 6248
rect 12855 6208 12900 6236
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13170 6196 13176 6248
rect 13228 6236 13234 6248
rect 13633 6239 13691 6245
rect 13633 6236 13645 6239
rect 13228 6208 13645 6236
rect 13228 6196 13234 6208
rect 13633 6205 13645 6208
rect 13679 6205 13691 6239
rect 13814 6236 13820 6248
rect 13775 6208 13820 6236
rect 13633 6199 13691 6205
rect 13814 6196 13820 6208
rect 13872 6236 13878 6248
rect 14553 6239 14611 6245
rect 14553 6236 14565 6239
rect 13872 6208 14565 6236
rect 13872 6196 13878 6208
rect 14553 6205 14565 6208
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 12802 6128 12808 6180
rect 12860 6168 12866 6180
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 12860 6140 14013 6168
rect 12860 6128 12866 6140
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14568 6168 14596 6199
rect 14826 6196 14832 6248
rect 14884 6236 14890 6248
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14884 6208 14933 6236
rect 14884 6196 14890 6208
rect 14921 6205 14933 6208
rect 14967 6205 14979 6239
rect 15470 6236 15476 6248
rect 14921 6199 14979 6205
rect 15304 6208 15476 6236
rect 15304 6168 15332 6208
rect 15470 6196 15476 6208
rect 15528 6196 15534 6248
rect 15672 6236 15700 6276
rect 15746 6264 15752 6316
rect 15804 6304 15810 6316
rect 16025 6307 16083 6313
rect 16025 6304 16037 6307
rect 15804 6276 16037 6304
rect 15804 6264 15810 6276
rect 16025 6273 16037 6276
rect 16071 6273 16083 6307
rect 16025 6267 16083 6273
rect 16114 6236 16120 6248
rect 15672 6208 15884 6236
rect 16075 6208 16120 6236
rect 15657 6171 15715 6177
rect 15657 6168 15669 6171
rect 14568 6140 15332 6168
rect 15387 6140 15669 6168
rect 14001 6131 14059 6137
rect 12299 6072 12756 6100
rect 12299 6069 12311 6072
rect 12253 6063 12311 6069
rect 14550 6060 14556 6112
rect 14608 6100 14614 6112
rect 15387 6100 15415 6140
rect 15657 6137 15669 6140
rect 15703 6137 15715 6171
rect 15657 6131 15715 6137
rect 15562 6100 15568 6112
rect 14608 6072 15415 6100
rect 15523 6072 15568 6100
rect 14608 6060 14614 6072
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 15856 6100 15884 6208
rect 16114 6196 16120 6208
rect 16172 6196 16178 6248
rect 16224 6245 16252 6344
rect 16936 6341 16948 6375
rect 16982 6372 16994 6375
rect 17034 6372 17040 6384
rect 16982 6344 17040 6372
rect 16982 6341 16994 6344
rect 16936 6335 16994 6341
rect 17034 6332 17040 6344
rect 17092 6372 17098 6384
rect 17770 6372 17776 6384
rect 17092 6344 17776 6372
rect 17092 6332 17098 6344
rect 17770 6332 17776 6344
rect 17828 6332 17834 6384
rect 17880 6372 17908 6412
rect 18322 6400 18328 6412
rect 18380 6400 18386 6452
rect 18966 6372 18972 6384
rect 17880 6344 18972 6372
rect 18966 6332 18972 6344
rect 19024 6332 19030 6384
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6304 18199 6307
rect 19702 6304 19708 6316
rect 18187 6276 19708 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 16209 6239 16267 6245
rect 16209 6205 16221 6239
rect 16255 6205 16267 6239
rect 16666 6236 16672 6248
rect 16627 6208 16672 6236
rect 16209 6199 16267 6205
rect 16666 6196 16672 6208
rect 16724 6196 16730 6248
rect 19610 6168 19616 6180
rect 17604 6140 19616 6168
rect 17604 6100 17632 6140
rect 19610 6128 19616 6140
rect 19668 6128 19674 6180
rect 15856 6072 17632 6100
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 18049 6103 18107 6109
rect 18049 6100 18061 6103
rect 17736 6072 18061 6100
rect 17736 6060 17742 6072
rect 18049 6069 18061 6072
rect 18095 6069 18107 6103
rect 18049 6063 18107 6069
rect 1104 6010 18860 6032
rect 1104 5958 3174 6010
rect 3226 5958 3238 6010
rect 3290 5958 3302 6010
rect 3354 5958 3366 6010
rect 3418 5958 3430 6010
rect 3482 5958 7622 6010
rect 7674 5958 7686 6010
rect 7738 5958 7750 6010
rect 7802 5958 7814 6010
rect 7866 5958 7878 6010
rect 7930 5958 12070 6010
rect 12122 5958 12134 6010
rect 12186 5958 12198 6010
rect 12250 5958 12262 6010
rect 12314 5958 12326 6010
rect 12378 5958 16518 6010
rect 16570 5958 16582 6010
rect 16634 5958 16646 6010
rect 16698 5958 16710 6010
rect 16762 5958 16774 6010
rect 16826 5958 18860 6010
rect 1104 5936 18860 5958
rect 1949 5899 2007 5905
rect 1949 5865 1961 5899
rect 1995 5896 2007 5899
rect 3510 5896 3516 5908
rect 1995 5868 3516 5896
rect 1995 5865 2007 5868
rect 1949 5859 2007 5865
rect 3510 5856 3516 5868
rect 3568 5856 3574 5908
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 3651 5868 5028 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 1673 5831 1731 5837
rect 1673 5797 1685 5831
rect 1719 5828 1731 5831
rect 2314 5828 2320 5840
rect 1719 5800 2320 5828
rect 1719 5797 1731 5800
rect 1673 5791 1731 5797
rect 2314 5788 2320 5800
rect 2372 5788 2378 5840
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5828 2835 5831
rect 5000 5828 5028 5868
rect 5166 5856 5172 5908
rect 5224 5896 5230 5908
rect 5445 5899 5503 5905
rect 5445 5896 5457 5899
rect 5224 5868 5457 5896
rect 5224 5856 5230 5868
rect 5445 5865 5457 5868
rect 5491 5865 5503 5899
rect 5445 5859 5503 5865
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 6972 5868 9996 5896
rect 6972 5856 6978 5868
rect 5810 5828 5816 5840
rect 2823 5800 4108 5828
rect 5000 5800 5816 5828
rect 2823 5797 2835 5800
rect 2777 5791 2835 5797
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 2958 5760 2964 5772
rect 2271 5732 2964 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 2958 5720 2964 5732
rect 3016 5720 3022 5772
rect 4080 5760 4108 5800
rect 5810 5788 5816 5800
rect 5868 5788 5874 5840
rect 8570 5788 8576 5840
rect 8628 5828 8634 5840
rect 8757 5831 8815 5837
rect 8757 5828 8769 5831
rect 8628 5800 8769 5828
rect 8628 5788 8634 5800
rect 8757 5797 8769 5800
rect 8803 5797 8815 5831
rect 8757 5791 8815 5797
rect 6178 5760 6184 5772
rect 4080 5732 4200 5760
rect 1765 5695 1823 5701
rect 1765 5661 1777 5695
rect 1811 5692 1823 5695
rect 1946 5692 1952 5704
rect 1811 5664 1952 5692
rect 1811 5661 1823 5664
rect 1765 5655 1823 5661
rect 1946 5652 1952 5664
rect 2004 5652 2010 5704
rect 2406 5692 2412 5704
rect 2367 5664 2412 5692
rect 2406 5652 2412 5664
rect 2464 5652 2470 5704
rect 3050 5652 3056 5704
rect 3108 5692 3114 5704
rect 3237 5695 3295 5701
rect 3237 5692 3249 5695
rect 3108 5664 3249 5692
rect 3108 5652 3114 5664
rect 3237 5661 3249 5664
rect 3283 5661 3295 5695
rect 3237 5655 3295 5661
rect 3970 5652 3976 5704
rect 4028 5692 4034 5704
rect 4065 5695 4123 5701
rect 4065 5692 4077 5695
rect 4028 5664 4077 5692
rect 4028 5652 4034 5664
rect 4065 5661 4077 5664
rect 4111 5661 4123 5695
rect 4172 5692 4200 5732
rect 5092 5732 6184 5760
rect 5092 5692 5120 5732
rect 6178 5720 6184 5732
rect 6236 5720 6242 5772
rect 8110 5760 8116 5772
rect 8071 5732 8116 5760
rect 8110 5720 8116 5732
rect 8168 5720 8174 5772
rect 9968 5760 9996 5868
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 11756 5868 14688 5896
rect 11756 5856 11762 5868
rect 13725 5831 13783 5837
rect 13725 5828 13737 5831
rect 13372 5800 13737 5828
rect 9968 5732 12388 5760
rect 4172 5664 5120 5692
rect 5537 5695 5595 5701
rect 4065 5655 4123 5661
rect 5537 5661 5549 5695
rect 5583 5661 5595 5695
rect 5537 5655 5595 5661
rect 5813 5695 5871 5701
rect 5813 5661 5825 5695
rect 5859 5692 5871 5695
rect 6638 5692 6644 5704
rect 5859 5664 6644 5692
rect 5859 5661 5871 5664
rect 5813 5655 5871 5661
rect 1489 5627 1547 5633
rect 1489 5593 1501 5627
rect 1535 5624 1547 5627
rect 1670 5624 1676 5636
rect 1535 5596 1676 5624
rect 1535 5593 1547 5596
rect 1489 5587 1547 5593
rect 1670 5584 1676 5596
rect 1728 5584 1734 5636
rect 3145 5627 3203 5633
rect 3145 5593 3157 5627
rect 3191 5624 3203 5627
rect 4154 5624 4160 5636
rect 3191 5596 4160 5624
rect 3191 5593 3203 5596
rect 3145 5587 3203 5593
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 4332 5627 4390 5633
rect 4332 5593 4344 5627
rect 4378 5624 4390 5627
rect 4430 5624 4436 5636
rect 4378 5596 4436 5624
rect 4378 5593 4390 5596
rect 4332 5587 4390 5593
rect 4430 5584 4436 5596
rect 4488 5584 4494 5636
rect 4890 5584 4896 5636
rect 4948 5624 4954 5636
rect 5552 5624 5580 5655
rect 6638 5652 6644 5664
rect 6696 5652 6702 5704
rect 7929 5695 7987 5701
rect 7929 5661 7941 5695
rect 7975 5692 7987 5695
rect 8294 5692 8300 5704
rect 7975 5664 8300 5692
rect 7975 5661 7987 5664
rect 7929 5655 7987 5661
rect 8294 5652 8300 5664
rect 8352 5692 8358 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8352 5664 8953 5692
rect 8352 5652 8358 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 9208 5695 9266 5701
rect 9208 5661 9220 5695
rect 9254 5692 9266 5695
rect 10502 5692 10508 5704
rect 9254 5664 10508 5692
rect 9254 5661 9266 5664
rect 9208 5655 9266 5661
rect 10502 5652 10508 5664
rect 10560 5652 10566 5704
rect 12253 5695 12311 5701
rect 12253 5692 12265 5695
rect 11716 5664 12265 5692
rect 4948 5596 5580 5624
rect 7684 5627 7742 5633
rect 4948 5584 4954 5596
rect 7684 5593 7696 5627
rect 7730 5624 7742 5627
rect 8110 5624 8116 5636
rect 7730 5596 8116 5624
rect 7730 5593 7742 5596
rect 7684 5587 7742 5593
rect 8110 5584 8116 5596
rect 8168 5584 8174 5636
rect 9030 5624 9036 5636
rect 8312 5596 9036 5624
rect 2222 5516 2228 5568
rect 2280 5556 2286 5568
rect 2317 5559 2375 5565
rect 2317 5556 2329 5559
rect 2280 5528 2329 5556
rect 2280 5516 2286 5528
rect 2317 5525 2329 5528
rect 2363 5525 2375 5559
rect 2317 5519 2375 5525
rect 3973 5559 4031 5565
rect 3973 5525 3985 5559
rect 4019 5556 4031 5559
rect 5718 5556 5724 5568
rect 4019 5528 5724 5556
rect 4019 5525 4031 5528
rect 3973 5519 4031 5525
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 5902 5516 5908 5568
rect 5960 5556 5966 5568
rect 6086 5556 6092 5568
rect 5960 5528 6092 5556
rect 5960 5516 5966 5528
rect 6086 5516 6092 5528
rect 6144 5556 6150 5568
rect 8312 5565 8340 5596
rect 9030 5584 9036 5596
rect 9088 5584 9094 5636
rect 9582 5584 9588 5636
rect 9640 5624 9646 5636
rect 10413 5627 10471 5633
rect 10413 5624 10425 5627
rect 9640 5596 10425 5624
rect 9640 5584 9646 5596
rect 10413 5593 10425 5596
rect 10459 5624 10471 5627
rect 11330 5624 11336 5636
rect 10459 5596 11336 5624
rect 10459 5593 10471 5596
rect 10413 5587 10471 5593
rect 11330 5584 11336 5596
rect 11388 5584 11394 5636
rect 6549 5559 6607 5565
rect 6549 5556 6561 5559
rect 6144 5528 6561 5556
rect 6144 5516 6150 5528
rect 6549 5525 6561 5528
rect 6595 5525 6607 5559
rect 6549 5519 6607 5525
rect 8297 5559 8355 5565
rect 8297 5525 8309 5559
rect 8343 5525 8355 5559
rect 8297 5519 8355 5525
rect 8389 5559 8447 5565
rect 8389 5525 8401 5559
rect 8435 5556 8447 5559
rect 9766 5556 9772 5568
rect 8435 5528 9772 5556
rect 8435 5525 8447 5528
rect 8389 5519 8447 5525
rect 9766 5516 9772 5528
rect 9824 5516 9830 5568
rect 10321 5559 10379 5565
rect 10321 5525 10333 5559
rect 10367 5556 10379 5559
rect 10502 5556 10508 5568
rect 10367 5528 10508 5556
rect 10367 5525 10379 5528
rect 10321 5519 10379 5525
rect 10502 5516 10508 5528
rect 10560 5516 10566 5568
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11716 5565 11744 5664
rect 12253 5661 12265 5664
rect 12299 5661 12311 5695
rect 12360 5692 12388 5732
rect 12509 5695 12567 5701
rect 12509 5692 12521 5695
rect 12360 5664 12521 5692
rect 12253 5655 12311 5661
rect 12509 5661 12521 5664
rect 12555 5661 12567 5695
rect 12509 5655 12567 5661
rect 11790 5584 11796 5636
rect 11848 5624 11854 5636
rect 13372 5624 13400 5800
rect 13725 5797 13737 5800
rect 13771 5797 13783 5831
rect 14093 5831 14151 5837
rect 14093 5828 14105 5831
rect 13725 5791 13783 5797
rect 13832 5800 14105 5828
rect 13446 5652 13452 5704
rect 13504 5692 13510 5704
rect 13832 5692 13860 5800
rect 14093 5797 14105 5800
rect 14139 5797 14151 5831
rect 14093 5791 14151 5797
rect 14550 5760 14556 5772
rect 14511 5732 14556 5760
rect 14550 5720 14556 5732
rect 14608 5720 14614 5772
rect 14660 5769 14688 5868
rect 14826 5856 14832 5908
rect 14884 5896 14890 5908
rect 14884 5868 15700 5896
rect 14884 5856 14890 5868
rect 15562 5828 15568 5840
rect 15396 5800 15568 5828
rect 15396 5769 15424 5800
rect 15562 5788 15568 5800
rect 15620 5788 15626 5840
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 15381 5763 15439 5769
rect 15381 5729 15393 5763
rect 15427 5729 15439 5763
rect 15381 5723 15439 5729
rect 15470 5720 15476 5772
rect 15528 5760 15534 5772
rect 15672 5760 15700 5868
rect 16114 5856 16120 5908
rect 16172 5896 16178 5908
rect 16577 5899 16635 5905
rect 16577 5896 16589 5899
rect 16172 5868 16589 5896
rect 16172 5856 16178 5868
rect 16577 5865 16589 5868
rect 16623 5865 16635 5899
rect 16577 5859 16635 5865
rect 15930 5788 15936 5840
rect 15988 5828 15994 5840
rect 17405 5831 17463 5837
rect 17405 5828 17417 5831
rect 15988 5800 17417 5828
rect 15988 5788 15994 5800
rect 17405 5797 17417 5800
rect 17451 5797 17463 5831
rect 17405 5791 17463 5797
rect 16301 5763 16359 5769
rect 16301 5760 16313 5763
rect 15528 5732 15573 5760
rect 15672 5732 16313 5760
rect 15528 5720 15534 5732
rect 16301 5729 16313 5732
rect 16347 5760 16359 5763
rect 17129 5763 17187 5769
rect 17129 5760 17141 5763
rect 16347 5732 17141 5760
rect 16347 5729 16359 5732
rect 16301 5723 16359 5729
rect 17129 5729 17141 5732
rect 17175 5729 17187 5763
rect 17129 5723 17187 5729
rect 17678 5720 17684 5772
rect 17736 5760 17742 5772
rect 17957 5763 18015 5769
rect 17957 5760 17969 5763
rect 17736 5732 17969 5760
rect 17736 5720 17742 5732
rect 17957 5729 17969 5732
rect 18003 5729 18015 5763
rect 17957 5723 18015 5729
rect 13504 5664 13860 5692
rect 13504 5652 13510 5664
rect 13906 5652 13912 5704
rect 13964 5692 13970 5704
rect 13964 5664 14009 5692
rect 13964 5652 13970 5664
rect 16114 5652 16120 5704
rect 16172 5692 16178 5704
rect 16209 5695 16267 5701
rect 16209 5692 16221 5695
rect 16172 5664 16221 5692
rect 16172 5652 16178 5664
rect 16209 5661 16221 5664
rect 16255 5661 16267 5695
rect 16209 5655 16267 5661
rect 17402 5652 17408 5704
rect 17460 5692 17466 5704
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 17460 5664 17877 5692
rect 17460 5652 17466 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18233 5695 18291 5701
rect 18233 5661 18245 5695
rect 18279 5692 18291 5695
rect 19058 5692 19064 5704
rect 18279 5664 19064 5692
rect 18279 5661 18291 5664
rect 18233 5655 18291 5661
rect 19058 5652 19064 5664
rect 19116 5652 19122 5704
rect 11848 5596 13400 5624
rect 14461 5627 14519 5633
rect 11848 5584 11854 5596
rect 14461 5593 14473 5627
rect 14507 5624 14519 5627
rect 14507 5596 14964 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 11701 5559 11759 5565
rect 11701 5556 11713 5559
rect 11296 5528 11713 5556
rect 11296 5516 11302 5528
rect 11701 5525 11713 5528
rect 11747 5525 11759 5559
rect 11701 5519 11759 5525
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 14826 5556 14832 5568
rect 13679 5528 14832 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 14826 5516 14832 5528
rect 14884 5516 14890 5568
rect 14936 5565 14964 5596
rect 15010 5584 15016 5636
rect 15068 5624 15074 5636
rect 16945 5627 17003 5633
rect 16945 5624 16957 5627
rect 15068 5596 16957 5624
rect 15068 5584 15074 5596
rect 16945 5593 16957 5596
rect 16991 5593 17003 5627
rect 16945 5587 17003 5593
rect 17586 5584 17592 5636
rect 17644 5624 17650 5636
rect 17773 5627 17831 5633
rect 17773 5624 17785 5627
rect 17644 5596 17785 5624
rect 17644 5584 17650 5596
rect 17773 5593 17785 5596
rect 17819 5593 17831 5627
rect 17773 5587 17831 5593
rect 14921 5559 14979 5565
rect 14921 5525 14933 5559
rect 14967 5525 14979 5559
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 14921 5519 14979 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 15746 5556 15752 5568
rect 15707 5528 15752 5556
rect 15746 5516 15752 5528
rect 15804 5516 15810 5568
rect 16117 5559 16175 5565
rect 16117 5525 16129 5559
rect 16163 5556 16175 5559
rect 16850 5556 16856 5568
rect 16163 5528 16856 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 16850 5516 16856 5528
rect 16908 5516 16914 5568
rect 17037 5559 17095 5565
rect 17037 5525 17049 5559
rect 17083 5556 17095 5559
rect 18046 5556 18052 5568
rect 17083 5528 18052 5556
rect 17083 5525 17095 5528
rect 17037 5519 17095 5525
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18414 5556 18420 5568
rect 18375 5528 18420 5556
rect 18414 5516 18420 5528
rect 18472 5516 18478 5568
rect 1104 5466 18860 5488
rect 1104 5414 5398 5466
rect 5450 5414 5462 5466
rect 5514 5414 5526 5466
rect 5578 5414 5590 5466
rect 5642 5414 5654 5466
rect 5706 5414 9846 5466
rect 9898 5414 9910 5466
rect 9962 5414 9974 5466
rect 10026 5414 10038 5466
rect 10090 5414 10102 5466
rect 10154 5414 14294 5466
rect 14346 5414 14358 5466
rect 14410 5414 14422 5466
rect 14474 5414 14486 5466
rect 14538 5414 14550 5466
rect 14602 5414 18860 5466
rect 1104 5392 18860 5414
rect 2038 5352 2044 5364
rect 1999 5324 2044 5352
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 4522 5352 4528 5364
rect 3988 5324 4528 5352
rect 1949 5287 2007 5293
rect 1949 5253 1961 5287
rect 1995 5284 2007 5287
rect 3988 5284 4016 5324
rect 4522 5312 4528 5324
rect 4580 5312 4586 5364
rect 4614 5312 4620 5364
rect 4672 5352 4678 5364
rect 4982 5352 4988 5364
rect 4672 5324 4988 5352
rect 4672 5312 4678 5324
rect 4982 5312 4988 5324
rect 5040 5352 5046 5364
rect 6089 5355 6147 5361
rect 6089 5352 6101 5355
rect 5040 5324 6101 5352
rect 5040 5312 5046 5324
rect 6089 5321 6101 5324
rect 6135 5352 6147 5355
rect 6178 5352 6184 5364
rect 6135 5324 6184 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 6825 5355 6883 5361
rect 6825 5321 6837 5355
rect 6871 5352 6883 5355
rect 7282 5352 7288 5364
rect 6871 5324 7288 5352
rect 6871 5321 6883 5324
rect 6825 5315 6883 5321
rect 7282 5312 7288 5324
rect 7340 5312 7346 5364
rect 8570 5352 8576 5364
rect 8531 5324 8576 5352
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 9030 5352 9036 5364
rect 8991 5324 9036 5352
rect 9030 5312 9036 5324
rect 9088 5312 9094 5364
rect 9306 5312 9312 5364
rect 9364 5352 9370 5364
rect 9401 5355 9459 5361
rect 9401 5352 9413 5355
rect 9364 5324 9413 5352
rect 9364 5312 9370 5324
rect 9401 5321 9413 5324
rect 9447 5321 9459 5355
rect 9401 5315 9459 5321
rect 9493 5355 9551 5361
rect 9493 5321 9505 5355
rect 9539 5352 9551 5355
rect 12618 5352 12624 5364
rect 9539 5324 12624 5352
rect 9539 5321 9551 5324
rect 9493 5315 9551 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 12768 5324 13032 5352
rect 12768 5312 12774 5324
rect 1995 5256 4016 5284
rect 1995 5253 2007 5256
rect 1949 5247 2007 5253
rect 1397 5219 1455 5225
rect 1397 5185 1409 5219
rect 1443 5216 1455 5219
rect 1670 5216 1676 5228
rect 1443 5188 1676 5216
rect 1443 5185 1455 5188
rect 1397 5179 1455 5185
rect 1670 5176 1676 5188
rect 1728 5176 1734 5228
rect 2682 5176 2688 5228
rect 2740 5216 2746 5228
rect 3988 5225 4016 5256
rect 4884 5287 4942 5293
rect 4884 5253 4896 5287
rect 4930 5284 4942 5287
rect 5810 5284 5816 5296
rect 4930 5256 5816 5284
rect 4930 5253 4942 5256
rect 4884 5247 4942 5253
rect 5810 5244 5816 5256
rect 5868 5244 5874 5296
rect 8478 5284 8484 5296
rect 6748 5256 8484 5284
rect 3614 5219 3672 5225
rect 3614 5216 3626 5219
rect 2740 5188 3626 5216
rect 2740 5176 2746 5188
rect 3614 5185 3626 5188
rect 3660 5185 3672 5219
rect 3614 5179 3672 5185
rect 3973 5219 4031 5225
rect 3973 5185 3985 5219
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4154 5176 4160 5228
rect 4212 5216 4218 5228
rect 4249 5219 4307 5225
rect 4249 5216 4261 5219
rect 4212 5188 4261 5216
rect 4212 5176 4218 5188
rect 4249 5185 4261 5188
rect 4295 5185 4307 5219
rect 4249 5179 4307 5185
rect 4706 5176 4712 5228
rect 4764 5216 4770 5228
rect 4764 5188 6500 5216
rect 4764 5176 4770 5188
rect 6472 5160 6500 5188
rect 1578 5108 1584 5160
rect 1636 5148 1642 5160
rect 1857 5151 1915 5157
rect 1857 5148 1869 5151
rect 1636 5120 1869 5148
rect 1636 5108 1642 5120
rect 1857 5117 1869 5120
rect 1903 5148 1915 5151
rect 3881 5151 3939 5157
rect 1903 5120 2360 5148
rect 1903 5117 1915 5120
rect 1857 5111 1915 5117
rect 1581 5015 1639 5021
rect 1581 4981 1593 5015
rect 1627 5012 1639 5015
rect 2038 5012 2044 5024
rect 1627 4984 2044 5012
rect 1627 4981 1639 4984
rect 1581 4975 1639 4981
rect 2038 4972 2044 4984
rect 2096 4972 2102 5024
rect 2332 5012 2360 5120
rect 3881 5117 3893 5151
rect 3927 5148 3939 5151
rect 4617 5151 4675 5157
rect 4617 5148 4629 5151
rect 3927 5120 4629 5148
rect 3927 5117 3939 5120
rect 3881 5111 3939 5117
rect 4617 5117 4629 5120
rect 4663 5117 4675 5151
rect 6454 5148 6460 5160
rect 6415 5120 6460 5148
rect 4617 5111 4675 5117
rect 2409 5083 2467 5089
rect 2409 5049 2421 5083
rect 2455 5080 2467 5083
rect 2774 5080 2780 5092
rect 2455 5052 2780 5080
rect 2455 5049 2467 5052
rect 2409 5043 2467 5049
rect 2774 5040 2780 5052
rect 2832 5040 2838 5092
rect 3896 5080 3924 5111
rect 6454 5108 6460 5120
rect 6512 5108 6518 5160
rect 6748 5157 6776 5256
rect 8478 5244 8484 5256
rect 8536 5244 8542 5296
rect 8662 5284 8668 5296
rect 8623 5256 8668 5284
rect 8662 5244 8668 5256
rect 8720 5244 8726 5296
rect 10134 5244 10140 5296
rect 10192 5284 10198 5296
rect 10192 5256 11100 5284
rect 10192 5244 10198 5256
rect 6822 5176 6828 5228
rect 6880 5216 6886 5228
rect 6917 5219 6975 5225
rect 6917 5216 6929 5219
rect 6880 5188 6929 5216
rect 6880 5176 6886 5188
rect 6917 5185 6929 5188
rect 6963 5185 6975 5219
rect 6917 5179 6975 5185
rect 7745 5219 7803 5225
rect 7745 5185 7757 5219
rect 7791 5216 7803 5219
rect 9306 5216 9312 5228
rect 7791 5188 9312 5216
rect 7791 5185 7803 5188
rect 7745 5179 7803 5185
rect 9306 5176 9312 5188
rect 9364 5176 9370 5228
rect 9858 5176 9864 5228
rect 9916 5216 9922 5228
rect 10502 5216 10508 5228
rect 9916 5188 10508 5216
rect 9916 5176 9922 5188
rect 10502 5176 10508 5188
rect 10560 5176 10566 5228
rect 10962 5216 10968 5228
rect 11020 5225 11026 5228
rect 10932 5188 10968 5216
rect 10962 5176 10968 5188
rect 11020 5179 11032 5225
rect 11072 5216 11100 5256
rect 11330 5244 11336 5296
rect 11388 5284 11394 5296
rect 12728 5284 12756 5312
rect 13004 5293 13032 5324
rect 13998 5312 14004 5364
rect 14056 5352 14062 5364
rect 18417 5355 18475 5361
rect 14056 5324 17816 5352
rect 14056 5312 14062 5324
rect 11388 5256 12756 5284
rect 12989 5287 13047 5293
rect 11388 5244 11394 5256
rect 12989 5253 13001 5287
rect 13035 5253 13047 5287
rect 12989 5247 13047 5253
rect 13078 5244 13084 5296
rect 13136 5284 13142 5296
rect 14921 5287 14979 5293
rect 14921 5284 14933 5287
rect 13136 5256 14933 5284
rect 13136 5244 13142 5256
rect 14921 5253 14933 5256
rect 14967 5284 14979 5287
rect 15010 5284 15016 5296
rect 14967 5256 15016 5284
rect 14967 5253 14979 5256
rect 14921 5247 14979 5253
rect 15010 5244 15016 5256
rect 15068 5244 15074 5296
rect 15280 5287 15338 5293
rect 15280 5253 15292 5287
rect 15326 5284 15338 5287
rect 17034 5284 17040 5296
rect 15326 5256 17040 5284
rect 15326 5253 15338 5256
rect 15280 5247 15338 5253
rect 17034 5244 17040 5256
rect 17092 5284 17098 5296
rect 17678 5284 17684 5296
rect 17092 5256 17684 5284
rect 17092 5244 17098 5256
rect 17678 5244 17684 5256
rect 17736 5244 17742 5296
rect 12641 5219 12699 5225
rect 11072 5188 11376 5216
rect 11020 5176 11026 5179
rect 6733 5151 6791 5157
rect 6733 5117 6745 5151
rect 6779 5117 6791 5151
rect 6733 5111 6791 5117
rect 7466 5108 7472 5160
rect 7524 5148 7530 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 7524 5120 7849 5148
rect 7524 5108 7530 5120
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 8021 5151 8079 5157
rect 8021 5117 8033 5151
rect 8067 5148 8079 5151
rect 8110 5148 8116 5160
rect 8067 5120 8116 5148
rect 8067 5117 8079 5120
rect 8021 5111 8079 5117
rect 8110 5108 8116 5120
rect 8168 5108 8174 5160
rect 8849 5151 8907 5157
rect 8849 5117 8861 5151
rect 8895 5148 8907 5151
rect 9122 5148 9128 5160
rect 8895 5120 9128 5148
rect 8895 5117 8907 5120
rect 8849 5111 8907 5117
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10042 5148 10048 5160
rect 9732 5120 10048 5148
rect 9732 5108 9738 5120
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 11238 5148 11244 5160
rect 11199 5120 11244 5148
rect 11238 5108 11244 5120
rect 11296 5108 11302 5160
rect 3970 5080 3976 5092
rect 3896 5052 3976 5080
rect 3970 5040 3976 5052
rect 4028 5040 4034 5092
rect 4154 5080 4160 5092
rect 4115 5052 4160 5080
rect 4154 5040 4160 5052
rect 4212 5040 4218 5092
rect 7285 5083 7343 5089
rect 7285 5049 7297 5083
rect 7331 5080 7343 5083
rect 9030 5080 9036 5092
rect 7331 5052 9036 5080
rect 7331 5049 7343 5052
rect 7285 5043 7343 5049
rect 9030 5040 9036 5052
rect 9088 5040 9094 5092
rect 11348 5080 11376 5188
rect 12641 5185 12653 5219
rect 12687 5216 12699 5219
rect 13538 5216 13544 5228
rect 12687 5188 13544 5216
rect 12687 5185 12699 5188
rect 12641 5179 12699 5185
rect 13538 5176 13544 5188
rect 13596 5176 13602 5228
rect 13814 5176 13820 5228
rect 13872 5216 13878 5228
rect 16758 5216 16764 5228
rect 13872 5188 16068 5216
rect 16719 5188 16764 5216
rect 13872 5176 13878 5188
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5148 12955 5151
rect 15013 5151 15071 5157
rect 15013 5148 15025 5151
rect 12943 5120 15025 5148
rect 12943 5117 12955 5120
rect 12897 5111 12955 5117
rect 14292 5089 14320 5120
rect 15013 5117 15025 5120
rect 15059 5117 15071 5151
rect 16040 5148 16068 5188
rect 16758 5176 16764 5188
rect 16816 5176 16822 5228
rect 17497 5219 17555 5225
rect 17497 5216 17509 5219
rect 16868 5188 17509 5216
rect 16868 5148 16896 5188
rect 17497 5185 17509 5188
rect 17543 5185 17555 5219
rect 17497 5179 17555 5185
rect 17586 5148 17592 5160
rect 16040 5120 16896 5148
rect 17547 5120 17592 5148
rect 15013 5111 15071 5117
rect 14277 5083 14335 5089
rect 11348 5052 11560 5080
rect 11532 5024 11560 5052
rect 14277 5049 14289 5083
rect 14323 5049 14335 5083
rect 14277 5043 14335 5049
rect 2498 5012 2504 5024
rect 2332 4984 2504 5012
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 3510 4972 3516 5024
rect 3568 5012 3574 5024
rect 4433 5015 4491 5021
rect 4433 5012 4445 5015
rect 3568 4984 4445 5012
rect 3568 4972 3574 4984
rect 4433 4981 4445 4984
rect 4479 4981 4491 5015
rect 4433 4975 4491 4981
rect 4522 4972 4528 5024
rect 4580 5012 4586 5024
rect 5350 5012 5356 5024
rect 4580 4984 5356 5012
rect 4580 4972 4586 4984
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5994 5012 6000 5024
rect 5955 4984 6000 5012
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 7432 4984 7477 5012
rect 7432 4972 7438 4984
rect 8018 4972 8024 5024
rect 8076 5012 8082 5024
rect 8205 5015 8263 5021
rect 8205 5012 8217 5015
rect 8076 4984 8217 5012
rect 8076 4972 8082 4984
rect 8205 4981 8217 4984
rect 8251 4981 8263 5015
rect 8205 4975 8263 4981
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 9861 5015 9919 5021
rect 9861 5012 9873 5015
rect 8536 4984 9873 5012
rect 8536 4972 8542 4984
rect 9861 4981 9873 4984
rect 9907 5012 9919 5015
rect 11330 5012 11336 5024
rect 9907 4984 11336 5012
rect 9907 4981 9919 4984
rect 9861 4975 9919 4981
rect 11330 4972 11336 4984
rect 11388 4972 11394 5024
rect 11514 4972 11520 5024
rect 11572 5012 11578 5024
rect 11572 4984 11665 5012
rect 11572 4972 11578 4984
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 13078 5012 13084 5024
rect 11848 4984 13084 5012
rect 11848 4972 11854 4984
rect 13078 4972 13084 4984
rect 13136 4972 13142 5024
rect 15028 5012 15056 5111
rect 17586 5108 17592 5120
rect 17644 5108 17650 5160
rect 17696 5157 17724 5244
rect 17788 5216 17816 5324
rect 18417 5321 18429 5355
rect 18463 5352 18475 5355
rect 18690 5352 18696 5364
rect 18463 5324 18696 5352
rect 18463 5321 18475 5324
rect 18417 5315 18475 5321
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 17957 5219 18015 5225
rect 17957 5216 17969 5219
rect 17788 5188 17969 5216
rect 17957 5185 17969 5188
rect 18003 5185 18015 5219
rect 18230 5216 18236 5228
rect 18191 5188 18236 5216
rect 17957 5179 18015 5185
rect 18230 5176 18236 5188
rect 18288 5176 18294 5228
rect 17681 5151 17739 5157
rect 17681 5117 17693 5151
rect 17727 5117 17739 5151
rect 17681 5111 17739 5117
rect 15378 5012 15384 5024
rect 15028 4984 15384 5012
rect 15378 4972 15384 4984
rect 15436 4972 15442 5024
rect 16298 4972 16304 5024
rect 16356 5012 16362 5024
rect 16393 5015 16451 5021
rect 16393 5012 16405 5015
rect 16356 4984 16405 5012
rect 16356 4972 16362 4984
rect 16393 4981 16405 4984
rect 16439 4981 16451 5015
rect 16942 5012 16948 5024
rect 16903 4984 16948 5012
rect 16393 4975 16451 4981
rect 16942 4972 16948 4984
rect 17000 4972 17006 5024
rect 17126 5012 17132 5024
rect 17087 4984 17132 5012
rect 17126 4972 17132 4984
rect 17184 4972 17190 5024
rect 18141 5015 18199 5021
rect 18141 4981 18153 5015
rect 18187 5012 18199 5015
rect 18230 5012 18236 5024
rect 18187 4984 18236 5012
rect 18187 4981 18199 4984
rect 18141 4975 18199 4981
rect 18230 4972 18236 4984
rect 18288 4972 18294 5024
rect 1104 4922 18860 4944
rect 1104 4870 3174 4922
rect 3226 4870 3238 4922
rect 3290 4870 3302 4922
rect 3354 4870 3366 4922
rect 3418 4870 3430 4922
rect 3482 4870 7622 4922
rect 7674 4870 7686 4922
rect 7738 4870 7750 4922
rect 7802 4870 7814 4922
rect 7866 4870 7878 4922
rect 7930 4870 12070 4922
rect 12122 4870 12134 4922
rect 12186 4870 12198 4922
rect 12250 4870 12262 4922
rect 12314 4870 12326 4922
rect 12378 4870 16518 4922
rect 16570 4870 16582 4922
rect 16634 4870 16646 4922
rect 16698 4870 16710 4922
rect 16762 4870 16774 4922
rect 16826 4870 18860 4922
rect 1104 4848 18860 4870
rect 1857 4811 1915 4817
rect 1857 4777 1869 4811
rect 1903 4808 1915 4811
rect 1946 4808 1952 4820
rect 1903 4780 1952 4808
rect 1903 4777 1915 4780
rect 1857 4771 1915 4777
rect 1946 4768 1952 4780
rect 2004 4768 2010 4820
rect 2498 4808 2504 4820
rect 2148 4780 2504 4808
rect 1946 4632 1952 4684
rect 2004 4672 2010 4684
rect 2148 4681 2176 4780
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 2866 4808 2872 4820
rect 2827 4780 2872 4808
rect 2866 4768 2872 4780
rect 2924 4768 2930 4820
rect 3786 4808 3792 4820
rect 3747 4780 3792 4808
rect 3786 4768 3792 4780
rect 3844 4768 3850 4820
rect 8018 4808 8024 4820
rect 5460 4780 8024 4808
rect 5460 4740 5488 4780
rect 8018 4768 8024 4780
rect 8076 4768 8082 4820
rect 9766 4768 9772 4820
rect 9824 4808 9830 4820
rect 10413 4811 10471 4817
rect 10413 4808 10425 4811
rect 9824 4780 10425 4808
rect 9824 4768 9830 4780
rect 10413 4777 10425 4780
rect 10459 4777 10471 4811
rect 10413 4771 10471 4777
rect 11974 4768 11980 4820
rect 12032 4808 12038 4820
rect 12069 4811 12127 4817
rect 12069 4808 12081 4811
rect 12032 4780 12081 4808
rect 12032 4768 12038 4780
rect 12069 4777 12081 4780
rect 12115 4777 12127 4811
rect 12069 4771 12127 4777
rect 15102 4768 15108 4820
rect 15160 4808 15166 4820
rect 15160 4780 16988 4808
rect 15160 4768 15166 4780
rect 2516 4712 5488 4740
rect 6181 4743 6239 4749
rect 2133 4675 2191 4681
rect 2133 4672 2145 4675
rect 2004 4644 2145 4672
rect 2004 4632 2010 4644
rect 2133 4641 2145 4644
rect 2179 4641 2191 4675
rect 2314 4672 2320 4684
rect 2275 4644 2320 4672
rect 2133 4635 2191 4641
rect 2314 4632 2320 4644
rect 2372 4632 2378 4684
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4573 1455 4607
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1397 4567 1455 4573
rect 1412 4536 1440 4567
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2406 4604 2412 4616
rect 2367 4576 2412 4604
rect 2406 4564 2412 4576
rect 2464 4564 2470 4616
rect 2516 4536 2544 4712
rect 6181 4709 6193 4743
rect 6227 4740 6239 4743
rect 6914 4740 6920 4752
rect 6227 4712 6920 4740
rect 6227 4709 6239 4712
rect 6181 4703 6239 4709
rect 6914 4700 6920 4712
rect 6972 4700 6978 4752
rect 10134 4740 10140 4752
rect 8588 4712 10140 4740
rect 3418 4672 3424 4684
rect 3379 4644 3424 4672
rect 3418 4632 3424 4644
rect 3476 4632 3482 4684
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 4985 4675 5043 4681
rect 4985 4672 4997 4675
rect 4856 4644 4997 4672
rect 4856 4632 4862 4644
rect 4985 4641 4997 4644
rect 5031 4641 5043 4675
rect 4985 4635 5043 4641
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 5261 4675 5319 4681
rect 5261 4672 5273 4675
rect 5132 4644 5273 4672
rect 5132 4632 5138 4644
rect 5261 4641 5273 4644
rect 5307 4641 5319 4675
rect 8294 4672 8300 4684
rect 8255 4644 8300 4672
rect 5261 4635 5319 4641
rect 8294 4632 8300 4644
rect 8352 4632 8358 4684
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4341 4607 4399 4613
rect 4341 4573 4353 4607
rect 4387 4604 4399 4607
rect 5166 4604 5172 4616
rect 4387 4576 5172 4604
rect 4387 4573 4399 4576
rect 4341 4567 4399 4573
rect 3050 4536 3056 4548
rect 1412 4508 2544 4536
rect 2792 4508 3056 4536
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2406 4428 2412 4480
rect 2464 4468 2470 4480
rect 2682 4468 2688 4480
rect 2464 4440 2688 4468
rect 2464 4428 2470 4440
rect 2682 4428 2688 4440
rect 2740 4428 2746 4480
rect 2792 4477 2820 4508
rect 3050 4496 3056 4508
rect 3108 4496 3114 4548
rect 3694 4496 3700 4548
rect 3752 4496 3758 4548
rect 3988 4536 4016 4567
rect 5166 4564 5172 4576
rect 5224 4564 5230 4616
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 5537 4607 5595 4613
rect 5537 4604 5549 4607
rect 5408 4576 5549 4604
rect 5408 4564 5414 4576
rect 5537 4573 5549 4576
rect 5583 4604 5595 4607
rect 6825 4607 6883 4613
rect 5583 4576 6776 4604
rect 5583 4573 5595 4576
rect 5537 4567 5595 4573
rect 4801 4539 4859 4545
rect 3988 4508 4476 4536
rect 2777 4471 2835 4477
rect 2777 4437 2789 4471
rect 2823 4437 2835 4471
rect 3234 4468 3240 4480
rect 3195 4440 3240 4468
rect 2777 4431 2835 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4468 3387 4471
rect 3602 4468 3608 4480
rect 3375 4440 3608 4468
rect 3375 4437 3387 4440
rect 3329 4431 3387 4437
rect 3602 4428 3608 4440
rect 3660 4428 3666 4480
rect 3712 4468 3740 4496
rect 3878 4468 3884 4480
rect 3712 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 4154 4468 4160 4480
rect 4115 4440 4160 4468
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 4448 4477 4476 4508
rect 4801 4505 4813 4539
rect 4847 4536 4859 4539
rect 6546 4536 6552 4548
rect 4847 4508 6552 4536
rect 4847 4505 4859 4508
rect 4801 4499 4859 4505
rect 6546 4496 6552 4508
rect 6604 4496 6610 4548
rect 6748 4536 6776 4576
rect 6825 4573 6837 4607
rect 6871 4604 6883 4607
rect 8588 4604 8616 4712
rect 10134 4700 10140 4712
rect 10192 4700 10198 4752
rect 10318 4700 10324 4752
rect 10376 4740 10382 4752
rect 10376 4712 10421 4740
rect 10376 4700 10382 4712
rect 10594 4700 10600 4752
rect 10652 4740 10658 4752
rect 10652 4712 11284 4740
rect 10652 4700 10658 4712
rect 9122 4672 9128 4684
rect 8680 4644 9128 4672
rect 8680 4613 8708 4644
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 9306 4672 9312 4684
rect 9267 4644 9312 4672
rect 9306 4632 9312 4644
rect 9364 4632 9370 4684
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 9858 4672 9864 4684
rect 9815 4644 9864 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 9858 4632 9864 4644
rect 9916 4672 9922 4684
rect 10410 4672 10416 4684
rect 9916 4644 10416 4672
rect 9916 4632 9922 4644
rect 10410 4632 10416 4644
rect 10468 4632 10474 4684
rect 10686 4632 10692 4684
rect 10744 4672 10750 4684
rect 10873 4675 10931 4681
rect 10873 4672 10885 4675
rect 10744 4644 10885 4672
rect 10744 4632 10750 4644
rect 10873 4641 10885 4644
rect 10919 4641 10931 4675
rect 10873 4635 10931 4641
rect 10965 4675 11023 4681
rect 10965 4641 10977 4675
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 6871 4576 8616 4604
rect 8665 4607 8723 4613
rect 6871 4573 6883 4576
rect 6825 4567 6883 4573
rect 8665 4573 8677 4607
rect 8711 4573 8723 4607
rect 8938 4604 8944 4616
rect 8899 4576 8944 4604
rect 8665 4567 8723 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9953 4607 10011 4613
rect 9953 4604 9965 4607
rect 9416 4576 9965 4604
rect 8052 4539 8110 4545
rect 6748 4508 7972 4536
rect 4433 4471 4491 4477
rect 4433 4437 4445 4471
rect 4479 4437 4491 4471
rect 4433 4431 4491 4437
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 5166 4468 5172 4480
rect 4939 4440 5172 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 6917 4471 6975 4477
rect 6917 4437 6929 4471
rect 6963 4468 6975 4471
rect 7282 4468 7288 4480
rect 6963 4440 7288 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 7944 4468 7972 4508
rect 8052 4505 8064 4539
rect 8098 4536 8110 4539
rect 8202 4536 8208 4548
rect 8098 4508 8208 4536
rect 8098 4505 8110 4508
rect 8052 4499 8110 4505
rect 8202 4496 8208 4508
rect 8260 4496 8266 4548
rect 8312 4508 9260 4536
rect 8312 4468 8340 4508
rect 7944 4440 8340 4468
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 8481 4471 8539 4477
rect 8481 4468 8493 4471
rect 8444 4440 8493 4468
rect 8444 4428 8450 4440
rect 8481 4437 8493 4440
rect 8527 4437 8539 4471
rect 8481 4431 8539 4437
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9125 4471 9183 4477
rect 9125 4468 9137 4471
rect 8904 4440 9137 4468
rect 8904 4428 8910 4440
rect 9125 4437 9137 4440
rect 9171 4437 9183 4471
rect 9232 4468 9260 4508
rect 9306 4496 9312 4548
rect 9364 4536 9370 4548
rect 9416 4536 9444 4576
rect 9953 4573 9965 4576
rect 9999 4604 10011 4607
rect 9999 4576 10180 4604
rect 9999 4573 10011 4576
rect 9953 4567 10011 4573
rect 9766 4536 9772 4548
rect 9364 4508 9444 4536
rect 9646 4508 9772 4536
rect 9364 4496 9370 4508
rect 9646 4468 9674 4508
rect 9766 4496 9772 4508
rect 9824 4496 9830 4548
rect 9858 4496 9864 4548
rect 9916 4536 9922 4548
rect 10152 4536 10180 4576
rect 10226 4564 10232 4616
rect 10284 4604 10290 4616
rect 10980 4604 11008 4635
rect 10284 4576 11008 4604
rect 11256 4604 11284 4712
rect 11514 4700 11520 4752
rect 11572 4740 11578 4752
rect 14093 4743 14151 4749
rect 11572 4712 12434 4740
rect 11572 4700 11578 4712
rect 11330 4632 11336 4684
rect 11388 4672 11394 4684
rect 11793 4675 11851 4681
rect 11793 4672 11805 4675
rect 11388 4644 11805 4672
rect 11388 4632 11394 4644
rect 11793 4641 11805 4644
rect 11839 4641 11851 4675
rect 12406 4672 12434 4712
rect 14093 4709 14105 4743
rect 14139 4709 14151 4743
rect 14093 4703 14151 4709
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 12406 4644 12633 4672
rect 11793 4635 11851 4641
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 13538 4672 13544 4684
rect 13499 4644 13544 4672
rect 12621 4635 12679 4641
rect 13538 4632 13544 4644
rect 13596 4672 13602 4684
rect 14108 4672 14136 4703
rect 13596 4644 14136 4672
rect 16209 4675 16267 4681
rect 13596 4632 13602 4644
rect 16209 4641 16221 4675
rect 16255 4672 16267 4675
rect 16298 4672 16304 4684
rect 16255 4644 16304 4672
rect 16255 4641 16267 4644
rect 16209 4635 16267 4641
rect 16298 4632 16304 4644
rect 16356 4632 16362 4684
rect 11514 4604 11520 4616
rect 11256 4576 11520 4604
rect 10284 4564 10290 4576
rect 11514 4564 11520 4576
rect 11572 4564 11578 4616
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4604 11667 4607
rect 13449 4607 13507 4613
rect 11655 4576 13400 4604
rect 11655 4573 11667 4576
rect 11609 4567 11667 4573
rect 11790 4536 11796 4548
rect 9916 4508 9961 4536
rect 10152 4508 11796 4536
rect 9916 4496 9922 4508
rect 11790 4496 11796 4508
rect 11848 4496 11854 4548
rect 12437 4539 12495 4545
rect 12437 4505 12449 4539
rect 12483 4536 12495 4539
rect 13372 4536 13400 4576
rect 13449 4573 13461 4607
rect 13495 4604 13507 4607
rect 13814 4604 13820 4616
rect 13495 4576 13820 4604
rect 13495 4573 13507 4576
rect 13449 4567 13507 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 15378 4564 15384 4616
rect 15436 4604 15442 4616
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 15436 4576 15485 4604
rect 15436 4564 15442 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15930 4604 15936 4616
rect 15891 4576 15936 4604
rect 15473 4567 15531 4573
rect 15930 4564 15936 4576
rect 15988 4564 15994 4616
rect 16960 4613 16988 4780
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 18417 4811 18475 4817
rect 18012 4780 18276 4808
rect 18012 4768 18018 4780
rect 17034 4632 17040 4684
rect 17092 4672 17098 4684
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 17092 4644 17141 4672
rect 17092 4632 17098 4644
rect 17129 4641 17141 4644
rect 17175 4672 17187 4675
rect 17957 4675 18015 4681
rect 17957 4672 17969 4675
rect 17175 4644 17969 4672
rect 17175 4641 17187 4644
rect 17129 4635 17187 4641
rect 17957 4641 17969 4644
rect 18003 4641 18015 4675
rect 17957 4635 18015 4641
rect 18248 4613 18276 4780
rect 18417 4777 18429 4811
rect 18463 4808 18475 4811
rect 18506 4808 18512 4820
rect 18463 4780 18512 4808
rect 18463 4777 18475 4780
rect 18417 4771 18475 4777
rect 18506 4768 18512 4780
rect 18564 4768 18570 4820
rect 16945 4607 17003 4613
rect 16945 4573 16957 4607
rect 16991 4573 17003 4607
rect 18233 4607 18291 4613
rect 16945 4567 17003 4573
rect 17052 4576 18092 4604
rect 12483 4508 13032 4536
rect 13372 4508 14688 4536
rect 12483 4505 12495 4508
rect 12437 4499 12495 4505
rect 10778 4468 10784 4480
rect 9232 4440 9674 4468
rect 10739 4440 10784 4468
rect 9125 4431 9183 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 10870 4428 10876 4480
rect 10928 4468 10934 4480
rect 11241 4471 11299 4477
rect 11241 4468 11253 4471
rect 10928 4440 11253 4468
rect 10928 4428 10934 4440
rect 11241 4437 11253 4440
rect 11287 4437 11299 4471
rect 11241 4431 11299 4437
rect 11701 4471 11759 4477
rect 11701 4437 11713 4471
rect 11747 4468 11759 4471
rect 11882 4468 11888 4480
rect 11747 4440 11888 4468
rect 11747 4437 11759 4440
rect 11701 4431 11759 4437
rect 11882 4428 11888 4440
rect 11940 4468 11946 4480
rect 12342 4468 12348 4480
rect 11940 4440 12348 4468
rect 11940 4428 11946 4440
rect 12342 4428 12348 4440
rect 12400 4428 12406 4480
rect 12526 4468 12532 4480
rect 12487 4440 12532 4468
rect 12526 4428 12532 4440
rect 12584 4428 12590 4480
rect 13004 4477 13032 4508
rect 12989 4471 13047 4477
rect 12989 4437 13001 4471
rect 13035 4437 13047 4471
rect 13354 4468 13360 4480
rect 13315 4440 13360 4468
rect 12989 4431 13047 4437
rect 13354 4428 13360 4440
rect 13412 4428 13418 4480
rect 13906 4468 13912 4480
rect 13867 4440 13912 4468
rect 13906 4428 13912 4440
rect 13964 4428 13970 4480
rect 14660 4468 14688 4508
rect 14734 4496 14740 4548
rect 14792 4536 14798 4548
rect 17052 4545 17080 4576
rect 15206 4539 15264 4545
rect 15206 4536 15218 4539
rect 14792 4508 15218 4536
rect 14792 4496 14798 4508
rect 15206 4505 15218 4508
rect 15252 4505 15264 4539
rect 15206 4499 15264 4505
rect 16025 4539 16083 4545
rect 16025 4505 16037 4539
rect 16071 4536 16083 4539
rect 17037 4539 17095 4545
rect 16071 4508 16620 4536
rect 16071 4505 16083 4508
rect 16025 4499 16083 4505
rect 15286 4468 15292 4480
rect 14660 4440 15292 4468
rect 15286 4428 15292 4440
rect 15344 4428 15350 4480
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 16206 4428 16212 4480
rect 16264 4468 16270 4480
rect 16592 4477 16620 4508
rect 17037 4505 17049 4539
rect 17083 4505 17095 4539
rect 17037 4499 17095 4505
rect 17773 4539 17831 4545
rect 17773 4505 17785 4539
rect 17819 4536 17831 4539
rect 17954 4536 17960 4548
rect 17819 4508 17960 4536
rect 17819 4505 17831 4508
rect 17773 4499 17831 4505
rect 17954 4496 17960 4508
rect 18012 4496 18018 4548
rect 18064 4536 18092 4576
rect 18233 4573 18245 4607
rect 18279 4573 18291 4607
rect 18233 4567 18291 4573
rect 18414 4536 18420 4548
rect 18064 4508 18420 4536
rect 18414 4496 18420 4508
rect 18472 4536 18478 4548
rect 19610 4536 19616 4548
rect 18472 4508 19616 4536
rect 18472 4496 18478 4508
rect 19610 4496 19616 4508
rect 19668 4496 19674 4548
rect 16393 4471 16451 4477
rect 16393 4468 16405 4471
rect 16264 4440 16405 4468
rect 16264 4428 16270 4440
rect 16393 4437 16405 4440
rect 16439 4437 16451 4471
rect 16393 4431 16451 4437
rect 16577 4471 16635 4477
rect 16577 4437 16589 4471
rect 16623 4437 16635 4471
rect 17402 4468 17408 4480
rect 17363 4440 17408 4468
rect 16577 4431 16635 4437
rect 17402 4428 17408 4440
rect 17460 4428 17466 4480
rect 17862 4428 17868 4480
rect 17920 4468 17926 4480
rect 17920 4440 17965 4468
rect 17920 4428 17926 4440
rect 1104 4378 18860 4400
rect 1104 4326 5398 4378
rect 5450 4326 5462 4378
rect 5514 4326 5526 4378
rect 5578 4326 5590 4378
rect 5642 4326 5654 4378
rect 5706 4326 9846 4378
rect 9898 4326 9910 4378
rect 9962 4326 9974 4378
rect 10026 4326 10038 4378
rect 10090 4326 10102 4378
rect 10154 4326 14294 4378
rect 14346 4326 14358 4378
rect 14410 4326 14422 4378
rect 14474 4326 14486 4378
rect 14538 4326 14550 4378
rect 14602 4326 18860 4378
rect 1104 4304 18860 4326
rect 2958 4264 2964 4276
rect 2536 4236 2964 4264
rect 2536 4137 2564 4236
rect 2958 4224 2964 4236
rect 3016 4224 3022 4276
rect 4062 4224 4068 4276
rect 4120 4224 4126 4276
rect 5074 4224 5080 4276
rect 5132 4264 5138 4276
rect 5445 4267 5503 4273
rect 5132 4236 5177 4264
rect 5132 4224 5138 4236
rect 5445 4233 5457 4267
rect 5491 4233 5503 4267
rect 9214 4264 9220 4276
rect 5445 4227 5503 4233
rect 5644 4236 9220 4264
rect 4080 4196 4108 4224
rect 4430 4196 4436 4208
rect 2792 4168 4436 4196
rect 2521 4131 2579 4137
rect 2521 4097 2533 4131
rect 2567 4097 2579 4131
rect 2521 4091 2579 4097
rect 2792 4072 2820 4168
rect 4062 4128 4068 4140
rect 4120 4137 4126 4140
rect 4356 4137 4384 4168
rect 4430 4156 4436 4168
rect 4488 4156 4494 4208
rect 4985 4199 5043 4205
rect 4985 4165 4997 4199
rect 5031 4196 5043 4199
rect 5031 4168 5120 4196
rect 5031 4165 5043 4168
rect 4985 4159 5043 4165
rect 4120 4131 4143 4137
rect 3995 4100 4068 4128
rect 4062 4088 4068 4100
rect 4131 4128 4143 4131
rect 4341 4131 4399 4137
rect 4131 4100 4292 4128
rect 4131 4097 4143 4100
rect 4120 4091 4143 4097
rect 4120 4088 4126 4091
rect 2774 4060 2780 4072
rect 2735 4032 2780 4060
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 4264 4060 4292 4100
rect 4341 4097 4353 4131
rect 4387 4097 4399 4131
rect 4522 4128 4528 4140
rect 4483 4100 4528 4128
rect 4341 4091 4399 4097
rect 4522 4088 4528 4100
rect 4580 4088 4586 4140
rect 4614 4088 4620 4140
rect 4672 4128 4678 4140
rect 5092 4128 5120 4168
rect 5166 4156 5172 4208
rect 5224 4196 5230 4208
rect 5460 4196 5488 4227
rect 5224 4168 5488 4196
rect 5224 4156 5230 4168
rect 5644 4128 5672 4236
rect 9214 4224 9220 4236
rect 9272 4224 9278 4276
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9766 4264 9772 4276
rect 9548 4236 9772 4264
rect 9548 4224 9554 4236
rect 9766 4224 9772 4236
rect 9824 4224 9830 4276
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10226 4264 10232 4276
rect 10091 4236 10232 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10226 4224 10232 4236
rect 10284 4224 10290 4276
rect 10965 4267 11023 4273
rect 10965 4233 10977 4267
rect 11011 4264 11023 4267
rect 11011 4236 12480 4264
rect 11011 4233 11023 4236
rect 10965 4227 11023 4233
rect 8938 4196 8944 4208
rect 8128 4168 8944 4196
rect 4672 4100 5028 4128
rect 5092 4100 5672 4128
rect 5813 4131 5871 4137
rect 4672 4088 4678 4100
rect 4264 4032 4927 4060
rect 1397 3927 1455 3933
rect 1397 3893 1409 3927
rect 1443 3924 1455 3927
rect 2406 3924 2412 3936
rect 1443 3896 2412 3924
rect 1443 3893 1455 3896
rect 1397 3887 1455 3893
rect 2406 3884 2412 3896
rect 2464 3884 2470 3936
rect 2590 3884 2596 3936
rect 2648 3924 2654 3936
rect 2961 3927 3019 3933
rect 2961 3924 2973 3927
rect 2648 3896 2973 3924
rect 2648 3884 2654 3896
rect 2961 3893 2973 3896
rect 3007 3893 3019 3927
rect 2961 3887 3019 3893
rect 3694 3884 3700 3936
rect 3752 3924 3758 3936
rect 4522 3924 4528 3936
rect 3752 3896 4528 3924
rect 3752 3884 3758 3896
rect 4522 3884 4528 3896
rect 4580 3884 4586 3936
rect 4617 3927 4675 3933
rect 4617 3893 4629 3927
rect 4663 3924 4675 3927
rect 4798 3924 4804 3936
rect 4663 3896 4804 3924
rect 4663 3893 4675 3896
rect 4617 3887 4675 3893
rect 4798 3884 4804 3896
rect 4856 3884 4862 3936
rect 4899 3924 4927 4032
rect 5000 3992 5028 4100
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 6730 4128 6736 4140
rect 5859 4100 6736 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 6730 4088 6736 4100
rect 6788 4088 6794 4140
rect 7489 4131 7547 4137
rect 7489 4097 7501 4131
rect 7535 4128 7547 4131
rect 8018 4128 8024 4140
rect 7535 4100 8024 4128
rect 7535 4097 7547 4100
rect 7489 4091 7547 4097
rect 8018 4088 8024 4100
rect 8076 4088 8082 4140
rect 8128 4137 8156 4168
rect 8938 4156 8944 4168
rect 8996 4156 9002 4208
rect 9306 4156 9312 4208
rect 9364 4196 9370 4208
rect 9950 4196 9956 4208
rect 9364 4168 9956 4196
rect 9364 4156 9370 4168
rect 9950 4156 9956 4168
rect 10008 4156 10014 4208
rect 8113 4131 8171 4137
rect 8113 4097 8125 4131
rect 8159 4097 8171 4131
rect 8294 4128 8300 4140
rect 8113 4091 8171 4097
rect 8220 4100 8300 4128
rect 5258 4060 5264 4072
rect 5219 4032 5264 4060
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5902 4060 5908 4072
rect 5863 4032 5908 4060
rect 5902 4020 5908 4032
rect 5960 4020 5966 4072
rect 6086 4060 6092 4072
rect 6047 4032 6092 4060
rect 6086 4020 6092 4032
rect 6144 4020 6150 4072
rect 8220 4069 8248 4100
rect 8294 4088 8300 4100
rect 8352 4088 8358 4140
rect 8478 4137 8484 4140
rect 8472 4128 8484 4137
rect 8439 4100 8484 4128
rect 8472 4091 8484 4100
rect 8478 4088 8484 4091
rect 8536 4088 8542 4140
rect 10226 4088 10232 4140
rect 10284 4128 10290 4140
rect 10873 4131 10931 4137
rect 10873 4128 10885 4131
rect 10284 4100 10885 4128
rect 10284 4088 10290 4100
rect 10873 4097 10885 4100
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 7745 4063 7803 4069
rect 7745 4029 7757 4063
rect 7791 4060 7803 4063
rect 8205 4063 8263 4069
rect 8205 4060 8217 4063
rect 7791 4032 8217 4060
rect 7791 4029 7803 4032
rect 7745 4023 7803 4029
rect 8205 4029 8217 4032
rect 8251 4029 8263 4063
rect 9769 4063 9827 4069
rect 9769 4060 9781 4063
rect 8205 4023 8263 4029
rect 9600 4032 9781 4060
rect 5000 3964 6500 3992
rect 5994 3924 6000 3936
rect 4899 3896 6000 3924
rect 5994 3884 6000 3896
rect 6052 3884 6058 3936
rect 6362 3924 6368 3936
rect 6323 3896 6368 3924
rect 6362 3884 6368 3896
rect 6420 3884 6426 3936
rect 6472 3924 6500 3964
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 6472 3896 7941 3924
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 9214 3884 9220 3936
rect 9272 3924 9278 3936
rect 9600 3933 9628 4032
rect 9769 4029 9781 4032
rect 9815 4029 9827 4063
rect 9769 4023 9827 4029
rect 9950 4020 9956 4072
rect 10008 4060 10014 4072
rect 10008 4032 10053 4060
rect 10008 4020 10014 4032
rect 10134 4020 10140 4072
rect 10192 4060 10198 4072
rect 10980 4060 11008 4227
rect 11514 4156 11520 4208
rect 11572 4156 11578 4208
rect 11882 4196 11888 4208
rect 11843 4168 11888 4196
rect 11882 4156 11888 4168
rect 11940 4156 11946 4208
rect 12452 4196 12480 4236
rect 12526 4224 12532 4276
rect 12584 4264 12590 4276
rect 12621 4267 12679 4273
rect 12621 4264 12633 4267
rect 12584 4236 12633 4264
rect 12584 4224 12590 4236
rect 12621 4233 12633 4236
rect 12667 4233 12679 4267
rect 13814 4264 13820 4276
rect 13775 4236 13820 4264
rect 12621 4227 12679 4233
rect 13814 4224 13820 4236
rect 13872 4224 13878 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14185 4267 14243 4273
rect 14185 4264 14197 4267
rect 14056 4236 14197 4264
rect 14056 4224 14062 4236
rect 14185 4233 14197 4236
rect 14231 4233 14243 4267
rect 17405 4267 17463 4273
rect 14185 4227 14243 4233
rect 14292 4236 16528 4264
rect 12894 4196 12900 4208
rect 12452 4168 12900 4196
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 12989 4199 13047 4205
rect 12989 4165 13001 4199
rect 13035 4196 13047 4199
rect 14090 4196 14096 4208
rect 13035 4168 14096 4196
rect 13035 4165 13047 4168
rect 12989 4159 13047 4165
rect 14090 4156 14096 4168
rect 14148 4156 14154 4208
rect 11330 4128 11336 4140
rect 11164 4100 11336 4128
rect 11164 4072 11192 4100
rect 11330 4088 11336 4100
rect 11388 4088 11394 4140
rect 11532 4128 11560 4156
rect 11440 4100 11560 4128
rect 10192 4032 11008 4060
rect 10192 4020 10198 4032
rect 11146 4020 11152 4072
rect 11204 4060 11210 4072
rect 11204 4032 11297 4060
rect 11204 4020 11210 4032
rect 10413 3995 10471 4001
rect 10413 3961 10425 3995
rect 10459 3992 10471 3995
rect 10459 3964 10640 3992
rect 10459 3961 10471 3964
rect 10413 3955 10471 3961
rect 9585 3927 9643 3933
rect 9585 3924 9597 3927
rect 9272 3896 9597 3924
rect 9272 3884 9278 3896
rect 9585 3893 9597 3896
rect 9631 3893 9643 3927
rect 9585 3887 9643 3893
rect 9950 3884 9956 3936
rect 10008 3924 10014 3936
rect 10505 3927 10563 3933
rect 10505 3924 10517 3927
rect 10008 3896 10517 3924
rect 10008 3884 10014 3896
rect 10505 3893 10517 3896
rect 10551 3893 10563 3927
rect 10612 3924 10640 3964
rect 10870 3924 10876 3936
rect 10612 3896 10876 3924
rect 10505 3887 10563 3893
rect 10870 3884 10876 3896
rect 10928 3884 10934 3936
rect 11440 3924 11468 4100
rect 11606 4088 11612 4140
rect 11664 4128 11670 4140
rect 12529 4131 12587 4137
rect 11664 4100 12112 4128
rect 11664 4088 11670 4100
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 12084 4069 12112 4100
rect 12529 4097 12541 4131
rect 12575 4128 12587 4131
rect 12618 4128 12624 4140
rect 12575 4100 12624 4128
rect 12575 4097 12587 4100
rect 12529 4091 12587 4097
rect 12618 4088 12624 4100
rect 12676 4088 12682 4140
rect 13446 4128 13452 4140
rect 13407 4100 13452 4128
rect 13446 4088 13452 4100
rect 13504 4088 13510 4140
rect 13722 4088 13728 4140
rect 13780 4128 13786 4140
rect 14292 4128 14320 4236
rect 15378 4156 15384 4208
rect 15436 4196 15442 4208
rect 16500 4196 16528 4236
rect 17405 4233 17417 4267
rect 17451 4264 17463 4267
rect 17586 4264 17592 4276
rect 17451 4236 17592 4264
rect 17451 4233 17463 4236
rect 17405 4227 17463 4233
rect 17586 4224 17592 4236
rect 17644 4224 17650 4276
rect 18046 4264 18052 4276
rect 17696 4236 18052 4264
rect 17696 4196 17724 4236
rect 18046 4224 18052 4236
rect 18104 4224 18110 4276
rect 15436 4168 16436 4196
rect 16500 4168 17724 4196
rect 17773 4199 17831 4205
rect 15436 4156 15442 4168
rect 13780 4100 14320 4128
rect 14645 4131 14703 4137
rect 13780 4088 13786 4100
rect 14645 4097 14657 4131
rect 14691 4128 14703 4131
rect 15102 4128 15108 4140
rect 14691 4100 15108 4128
rect 14691 4097 14703 4100
rect 14645 4091 14703 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 16137 4131 16195 4137
rect 16137 4097 16149 4131
rect 16183 4128 16195 4131
rect 16298 4128 16304 4140
rect 16183 4100 16304 4128
rect 16183 4097 16195 4100
rect 16137 4091 16195 4097
rect 16298 4088 16304 4100
rect 16356 4088 16362 4140
rect 16408 4137 16436 4168
rect 17773 4165 17785 4199
rect 17819 4196 17831 4199
rect 18690 4196 18696 4208
rect 17819 4168 18696 4196
rect 17819 4165 17831 4168
rect 17773 4159 17831 4165
rect 18690 4156 18696 4168
rect 18748 4156 18754 4208
rect 16393 4131 16451 4137
rect 16393 4097 16405 4131
rect 16439 4097 16451 4131
rect 17310 4128 17316 4140
rect 17271 4100 17316 4128
rect 16393 4091 16451 4097
rect 17310 4088 17316 4100
rect 17368 4088 17374 4140
rect 17865 4131 17923 4137
rect 17865 4097 17877 4131
rect 17911 4128 17923 4131
rect 18230 4128 18236 4140
rect 17911 4100 18092 4128
rect 18191 4100 18236 4128
rect 17911 4097 17923 4100
rect 17865 4091 17923 4097
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11572 4032 11989 4060
rect 11572 4020 11578 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 11977 4023 12035 4029
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4029 12127 4063
rect 13078 4060 13084 4072
rect 13039 4032 13084 4060
rect 12069 4023 12127 4029
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13265 4063 13323 4069
rect 13265 4029 13277 4063
rect 13311 4060 13323 4063
rect 13538 4060 13544 4072
rect 13311 4032 13544 4060
rect 13311 4029 13323 4032
rect 13265 4023 13323 4029
rect 13538 4020 13544 4032
rect 13596 4020 13602 4072
rect 13998 4020 14004 4072
rect 14056 4060 14062 4072
rect 14277 4063 14335 4069
rect 14277 4060 14289 4063
rect 14056 4032 14289 4060
rect 14056 4020 14062 4032
rect 14277 4029 14289 4032
rect 14323 4029 14335 4063
rect 14277 4023 14335 4029
rect 14461 4063 14519 4069
rect 14461 4029 14473 4063
rect 14507 4060 14519 4063
rect 14734 4060 14740 4072
rect 14507 4032 14740 4060
rect 14507 4029 14519 4032
rect 14461 4023 14519 4029
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 16316 4060 16344 4088
rect 17218 4060 17224 4072
rect 16316 4032 17224 4060
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 17770 4020 17776 4072
rect 17828 4060 17834 4072
rect 17957 4063 18015 4069
rect 17957 4060 17969 4063
rect 17828 4032 17969 4060
rect 17828 4020 17834 4032
rect 17957 4029 17969 4032
rect 18003 4029 18015 4063
rect 18064 4060 18092 4100
rect 18230 4088 18236 4100
rect 18288 4088 18294 4140
rect 19518 4060 19524 4072
rect 18064 4032 19524 4060
rect 17957 4023 18015 4029
rect 19518 4020 19524 4032
rect 19576 4020 19582 4072
rect 12802 3952 12808 4004
rect 12860 3992 12866 4004
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 12860 3964 13645 3992
rect 12860 3952 12866 3964
rect 13633 3961 13645 3964
rect 13679 3961 13691 3995
rect 13633 3955 13691 3961
rect 13814 3952 13820 4004
rect 13872 3992 13878 4004
rect 14829 3995 14887 4001
rect 14829 3992 14841 3995
rect 13872 3964 14841 3992
rect 13872 3952 13878 3964
rect 14829 3961 14841 3964
rect 14875 3961 14887 3995
rect 15378 3992 15384 4004
rect 14829 3955 14887 3961
rect 14936 3964 15384 3992
rect 11517 3927 11575 3933
rect 11517 3924 11529 3927
rect 11440 3896 11529 3924
rect 11517 3893 11529 3896
rect 11563 3893 11575 3927
rect 11517 3887 11575 3893
rect 11790 3884 11796 3936
rect 11848 3924 11854 3936
rect 12345 3927 12403 3933
rect 12345 3924 12357 3927
rect 11848 3896 12357 3924
rect 11848 3884 11854 3896
rect 12345 3893 12357 3896
rect 12391 3893 12403 3927
rect 12345 3887 12403 3893
rect 12894 3884 12900 3936
rect 12952 3924 12958 3936
rect 14936 3924 14964 3964
rect 15378 3952 15384 3964
rect 15436 3952 15442 4004
rect 16390 3952 16396 4004
rect 16448 3992 16454 4004
rect 16669 3995 16727 4001
rect 16669 3992 16681 3995
rect 16448 3964 16681 3992
rect 16448 3952 16454 3964
rect 16669 3961 16681 3964
rect 16715 3961 16727 3995
rect 16669 3955 16727 3961
rect 18417 3995 18475 4001
rect 18417 3961 18429 3995
rect 18463 3992 18475 3995
rect 18598 3992 18604 4004
rect 18463 3964 18604 3992
rect 18463 3961 18475 3964
rect 18417 3955 18475 3961
rect 18598 3952 18604 3964
rect 18656 3952 18662 4004
rect 12952 3896 14964 3924
rect 12952 3884 12958 3896
rect 15010 3884 15016 3936
rect 15068 3924 15074 3936
rect 15068 3896 15113 3924
rect 15068 3884 15074 3896
rect 17678 3884 17684 3936
rect 17736 3924 17742 3936
rect 18138 3924 18144 3936
rect 17736 3896 18144 3924
rect 17736 3884 17742 3896
rect 18138 3884 18144 3896
rect 18196 3884 18202 3936
rect 1104 3834 18860 3856
rect 1104 3782 3174 3834
rect 3226 3782 3238 3834
rect 3290 3782 3302 3834
rect 3354 3782 3366 3834
rect 3418 3782 3430 3834
rect 3482 3782 7622 3834
rect 7674 3782 7686 3834
rect 7738 3782 7750 3834
rect 7802 3782 7814 3834
rect 7866 3782 7878 3834
rect 7930 3782 12070 3834
rect 12122 3782 12134 3834
rect 12186 3782 12198 3834
rect 12250 3782 12262 3834
rect 12314 3782 12326 3834
rect 12378 3782 16518 3834
rect 16570 3782 16582 3834
rect 16634 3782 16646 3834
rect 16698 3782 16710 3834
rect 16762 3782 16774 3834
rect 16826 3782 18860 3834
rect 1104 3760 18860 3782
rect 1578 3680 1584 3732
rect 1636 3720 1642 3732
rect 1636 3692 7696 3720
rect 1636 3680 1642 3692
rect 1489 3655 1547 3661
rect 1489 3621 1501 3655
rect 1535 3652 1547 3655
rect 3602 3652 3608 3664
rect 1535 3624 3608 3652
rect 1535 3621 1547 3624
rect 1489 3615 1547 3621
rect 3602 3612 3608 3624
rect 3660 3612 3666 3664
rect 6546 3652 6552 3664
rect 6507 3624 6552 3652
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 2498 3584 2504 3596
rect 2459 3556 2504 3584
rect 2498 3544 2504 3556
rect 2556 3584 2562 3596
rect 3329 3587 3387 3593
rect 3329 3584 3341 3587
rect 2556 3556 3341 3584
rect 2556 3544 2562 3556
rect 3329 3553 3341 3556
rect 3375 3553 3387 3587
rect 3970 3584 3976 3596
rect 3931 3556 3976 3584
rect 3329 3547 3387 3553
rect 3970 3544 3976 3556
rect 4028 3544 4034 3596
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 4488 3556 4629 3584
rect 4488 3544 4494 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 6086 3544 6092 3596
rect 6144 3584 6150 3596
rect 7101 3587 7159 3593
rect 7101 3584 7113 3587
rect 6144 3556 7113 3584
rect 6144 3544 6150 3556
rect 7101 3553 7113 3556
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 1854 3516 1860 3528
rect 1815 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4706 3516 4712 3528
rect 4203 3488 4712 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 4706 3476 4712 3488
rect 4764 3476 4770 3528
rect 4873 3519 4931 3525
rect 4873 3485 4885 3519
rect 4919 3516 4931 3519
rect 6457 3519 6515 3525
rect 4919 3488 5028 3516
rect 4919 3485 4931 3488
rect 4873 3479 4931 3485
rect 1302 3408 1308 3460
rect 1360 3448 1366 3460
rect 2409 3451 2467 3457
rect 2409 3448 2421 3451
rect 1360 3420 2421 3448
rect 1360 3408 1366 3420
rect 2409 3417 2421 3420
rect 2455 3417 2467 3451
rect 2409 3411 2467 3417
rect 4430 3408 4436 3460
rect 4488 3448 4494 3460
rect 4488 3420 4844 3448
rect 4488 3408 4494 3420
rect 1486 3340 1492 3392
rect 1544 3380 1550 3392
rect 1673 3383 1731 3389
rect 1673 3380 1685 3383
rect 1544 3352 1685 3380
rect 1544 3340 1550 3352
rect 1673 3349 1685 3352
rect 1719 3349 1731 3383
rect 1946 3380 1952 3392
rect 1907 3352 1952 3380
rect 1673 3343 1731 3349
rect 1946 3340 1952 3352
rect 2004 3340 2010 3392
rect 2314 3380 2320 3392
rect 2275 3352 2320 3380
rect 2314 3340 2320 3352
rect 2372 3340 2378 3392
rect 2498 3340 2504 3392
rect 2556 3380 2562 3392
rect 2777 3383 2835 3389
rect 2777 3380 2789 3383
rect 2556 3352 2789 3380
rect 2556 3340 2562 3352
rect 2777 3349 2789 3352
rect 2823 3349 2835 3383
rect 3142 3380 3148 3392
rect 3103 3352 3148 3380
rect 2777 3343 2835 3349
rect 3142 3340 3148 3352
rect 3200 3340 3206 3392
rect 3237 3383 3295 3389
rect 3237 3349 3249 3383
rect 3283 3380 3295 3383
rect 3510 3380 3516 3392
rect 3283 3352 3516 3380
rect 3283 3349 3295 3352
rect 3237 3343 3295 3349
rect 3510 3340 3516 3352
rect 3568 3380 3574 3392
rect 3786 3380 3792 3392
rect 3568 3352 3792 3380
rect 3568 3340 3574 3352
rect 3786 3340 3792 3352
rect 3844 3340 3850 3392
rect 3970 3340 3976 3392
rect 4028 3380 4034 3392
rect 4065 3383 4123 3389
rect 4065 3380 4077 3383
rect 4028 3352 4077 3380
rect 4028 3340 4034 3352
rect 4065 3349 4077 3352
rect 4111 3349 4123 3383
rect 4065 3343 4123 3349
rect 4246 3340 4252 3392
rect 4304 3380 4310 3392
rect 4525 3383 4583 3389
rect 4525 3380 4537 3383
rect 4304 3352 4537 3380
rect 4304 3340 4310 3352
rect 4525 3349 4537 3352
rect 4571 3349 4583 3383
rect 4816 3380 4844 3420
rect 5000 3380 5028 3488
rect 6457 3485 6469 3519
rect 6503 3485 6515 3519
rect 6457 3479 6515 3485
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3516 6975 3519
rect 7374 3516 7380 3528
rect 6963 3488 7380 3516
rect 6963 3485 6975 3488
rect 6917 3479 6975 3485
rect 5074 3408 5080 3460
rect 5132 3448 5138 3460
rect 6472 3448 6500 3479
rect 7374 3476 7380 3488
rect 7432 3476 7438 3528
rect 7668 3516 7696 3692
rect 8478 3680 8484 3732
rect 8536 3720 8542 3732
rect 10778 3720 10784 3732
rect 8536 3692 10784 3720
rect 8536 3680 8542 3692
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 10962 3680 10968 3732
rect 11020 3720 11026 3732
rect 11057 3723 11115 3729
rect 11057 3720 11069 3723
rect 11020 3692 11069 3720
rect 11020 3680 11026 3692
rect 11057 3689 11069 3692
rect 11103 3689 11115 3723
rect 11790 3720 11796 3732
rect 11057 3683 11115 3689
rect 11164 3692 11796 3720
rect 8202 3652 8208 3664
rect 7852 3624 8208 3652
rect 7852 3593 7880 3624
rect 8202 3612 8208 3624
rect 8260 3612 8266 3664
rect 7837 3587 7895 3593
rect 7837 3553 7849 3587
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 8021 3587 8079 3593
rect 8021 3553 8033 3587
rect 8067 3584 8079 3587
rect 8110 3584 8116 3596
rect 8067 3556 8116 3584
rect 8067 3553 8079 3556
rect 8021 3547 8079 3553
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 8294 3544 8300 3596
rect 8352 3584 8358 3596
rect 8941 3587 8999 3593
rect 8941 3584 8953 3587
rect 8352 3556 8953 3584
rect 8352 3544 8358 3556
rect 8941 3553 8953 3556
rect 8987 3553 8999 3587
rect 11164 3584 11192 3692
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 12406 3692 13032 3720
rect 12158 3612 12164 3664
rect 12216 3652 12222 3664
rect 12406 3652 12434 3692
rect 12216 3624 12434 3652
rect 12529 3655 12587 3661
rect 12216 3612 12222 3624
rect 12529 3621 12541 3655
rect 12575 3652 12587 3655
rect 12894 3652 12900 3664
rect 12575 3624 12900 3652
rect 12575 3621 12587 3624
rect 12529 3615 12587 3621
rect 12894 3612 12900 3624
rect 12952 3612 12958 3664
rect 8941 3547 8999 3553
rect 9968 3556 11192 3584
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 7668 3488 8493 3516
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 9968 3516 9996 3556
rect 10410 3516 10416 3528
rect 8481 3479 8539 3485
rect 8588 3488 9996 3516
rect 10371 3488 10416 3516
rect 8588 3448 8616 3488
rect 10410 3476 10416 3488
rect 10468 3476 10474 3528
rect 11149 3519 11207 3525
rect 11149 3485 11161 3519
rect 11195 3516 11207 3519
rect 11238 3516 11244 3528
rect 11195 3488 11244 3516
rect 11195 3485 11207 3488
rect 11149 3479 11207 3485
rect 11238 3476 11244 3488
rect 11296 3516 11302 3528
rect 12158 3516 12164 3528
rect 11296 3488 12164 3516
rect 11296 3476 11302 3488
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12618 3516 12624 3528
rect 12579 3488 12624 3516
rect 12618 3476 12624 3488
rect 12676 3476 12682 3528
rect 13004 3516 13032 3692
rect 13078 3680 13084 3732
rect 13136 3680 13142 3732
rect 13354 3680 13360 3732
rect 13412 3720 13418 3732
rect 13725 3723 13783 3729
rect 13725 3720 13737 3723
rect 13412 3692 13737 3720
rect 13412 3680 13418 3692
rect 13725 3689 13737 3692
rect 13771 3689 13783 3723
rect 13725 3683 13783 3689
rect 14642 3680 14648 3732
rect 14700 3720 14706 3732
rect 15470 3720 15476 3732
rect 14700 3692 15476 3720
rect 14700 3680 14706 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 17402 3720 17408 3732
rect 16776 3692 17408 3720
rect 13096 3652 13124 3680
rect 14093 3655 14151 3661
rect 14093 3652 14105 3655
rect 13096 3624 14105 3652
rect 14093 3621 14105 3624
rect 14139 3621 14151 3655
rect 14093 3615 14151 3621
rect 15286 3612 15292 3664
rect 15344 3652 15350 3664
rect 15344 3624 16160 3652
rect 15344 3612 15350 3624
rect 13173 3587 13231 3593
rect 13173 3553 13185 3587
rect 13219 3584 13231 3587
rect 14734 3584 14740 3596
rect 13219 3556 14740 3584
rect 13219 3553 13231 3556
rect 13173 3547 13231 3553
rect 14734 3544 14740 3556
rect 14792 3544 14798 3596
rect 15378 3544 15384 3596
rect 15436 3584 15442 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 15436 3556 15485 3584
rect 15436 3544 15442 3556
rect 15473 3553 15485 3556
rect 15519 3584 15531 3587
rect 15654 3584 15660 3596
rect 15519 3556 15660 3584
rect 15519 3553 15531 3556
rect 15473 3547 15531 3553
rect 15654 3544 15660 3556
rect 15712 3544 15718 3596
rect 16132 3593 16160 3624
rect 16117 3587 16175 3593
rect 16117 3553 16129 3587
rect 16163 3553 16175 3587
rect 16776 3584 16804 3692
rect 17402 3680 17408 3692
rect 17460 3680 17466 3732
rect 17589 3723 17647 3729
rect 17589 3689 17601 3723
rect 17635 3720 17647 3723
rect 17862 3720 17868 3732
rect 17635 3692 17868 3720
rect 17635 3689 17647 3692
rect 17589 3683 17647 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18509 3723 18567 3729
rect 18509 3689 18521 3723
rect 18555 3720 18567 3723
rect 18966 3720 18972 3732
rect 18555 3692 18972 3720
rect 18555 3689 18567 3692
rect 18509 3683 18567 3689
rect 18966 3680 18972 3692
rect 19024 3680 19030 3732
rect 17218 3612 17224 3664
rect 17276 3612 17282 3664
rect 19150 3652 19156 3664
rect 17512 3624 19156 3652
rect 16853 3587 16911 3593
rect 16853 3584 16865 3587
rect 16776 3556 16865 3584
rect 16117 3547 16175 3553
rect 16853 3553 16865 3556
rect 16899 3553 16911 3587
rect 16853 3547 16911 3553
rect 16991 3587 17049 3593
rect 16991 3553 17003 3587
rect 17037 3584 17049 3587
rect 17236 3584 17264 3612
rect 17037 3556 17264 3584
rect 17037 3553 17049 3556
rect 16991 3547 17049 3553
rect 13817 3519 13875 3525
rect 13817 3516 13829 3519
rect 13004 3488 13829 3516
rect 13817 3485 13829 3488
rect 13863 3485 13875 3519
rect 14458 3516 14464 3528
rect 14419 3488 14464 3516
rect 13817 3479 13875 3485
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15194 3476 15200 3528
rect 15252 3516 15258 3528
rect 15749 3519 15807 3525
rect 15749 3516 15761 3519
rect 15252 3488 15761 3516
rect 15252 3476 15258 3488
rect 15749 3485 15761 3488
rect 15795 3485 15807 3519
rect 15749 3479 15807 3485
rect 16761 3519 16819 3525
rect 16761 3485 16773 3519
rect 16807 3516 16819 3519
rect 17126 3516 17132 3528
rect 16807 3488 17132 3516
rect 16807 3485 16819 3488
rect 16761 3479 16819 3485
rect 17126 3476 17132 3488
rect 17184 3476 17190 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17276 3488 17321 3516
rect 17276 3476 17282 3488
rect 9214 3457 9220 3460
rect 9208 3448 9220 3457
rect 5132 3420 6316 3448
rect 6472 3420 8616 3448
rect 9175 3420 9220 3448
rect 5132 3408 5138 3420
rect 4816 3352 5028 3380
rect 5997 3383 6055 3389
rect 4525 3343 4583 3349
rect 5997 3349 6009 3383
rect 6043 3380 6055 3383
rect 6086 3380 6092 3392
rect 6043 3352 6092 3380
rect 6043 3349 6055 3352
rect 5997 3343 6055 3349
rect 6086 3340 6092 3352
rect 6144 3340 6150 3392
rect 6288 3389 6316 3420
rect 9208 3411 9220 3420
rect 9214 3408 9220 3411
rect 9272 3408 9278 3460
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 10134 3448 10140 3460
rect 9732 3420 10140 3448
rect 9732 3408 9738 3420
rect 10134 3408 10140 3420
rect 10192 3408 10198 3460
rect 10226 3408 10232 3460
rect 10284 3448 10290 3460
rect 11416 3451 11474 3457
rect 10284 3420 10916 3448
rect 10284 3408 10290 3420
rect 6273 3383 6331 3389
rect 6273 3349 6285 3383
rect 6319 3349 6331 3383
rect 6273 3343 6331 3349
rect 7009 3383 7067 3389
rect 7009 3349 7021 3383
rect 7055 3380 7067 3383
rect 7377 3383 7435 3389
rect 7377 3380 7389 3383
rect 7055 3352 7389 3380
rect 7055 3349 7067 3352
rect 7009 3343 7067 3349
rect 7377 3349 7389 3352
rect 7423 3349 7435 3383
rect 7377 3343 7435 3349
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 7745 3383 7803 3389
rect 7745 3380 7757 3383
rect 7616 3352 7757 3380
rect 7616 3340 7622 3352
rect 7745 3349 7757 3352
rect 7791 3349 7803 3383
rect 7745 3343 7803 3349
rect 8389 3383 8447 3389
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8478 3380 8484 3392
rect 8435 3352 8484 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8478 3340 8484 3352
rect 8536 3340 8542 3392
rect 8665 3383 8723 3389
rect 8665 3349 8677 3383
rect 8711 3380 8723 3383
rect 9306 3380 9312 3392
rect 8711 3352 9312 3380
rect 8711 3349 8723 3352
rect 8665 3343 8723 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 10321 3383 10379 3389
rect 10321 3349 10333 3383
rect 10367 3380 10379 3383
rect 10778 3380 10784 3392
rect 10367 3352 10784 3380
rect 10367 3349 10379 3352
rect 10321 3343 10379 3349
rect 10778 3340 10784 3352
rect 10836 3340 10842 3392
rect 10888 3380 10916 3420
rect 11416 3417 11428 3451
rect 11462 3448 11474 3451
rect 13722 3448 13728 3460
rect 11462 3420 13728 3448
rect 11462 3417 11474 3420
rect 11416 3411 11474 3417
rect 13722 3408 13728 3420
rect 13780 3408 13786 3460
rect 16114 3448 16120 3460
rect 14384 3420 16120 3448
rect 12805 3383 12863 3389
rect 12805 3380 12817 3383
rect 10888 3352 12817 3380
rect 12805 3349 12817 3352
rect 12851 3349 12863 3383
rect 12805 3343 12863 3349
rect 13170 3340 13176 3392
rect 13228 3380 13234 3392
rect 13265 3383 13323 3389
rect 13265 3380 13277 3383
rect 13228 3352 13277 3380
rect 13228 3340 13234 3352
rect 13265 3349 13277 3352
rect 13311 3349 13323 3383
rect 13265 3343 13323 3349
rect 13354 3340 13360 3392
rect 13412 3380 13418 3392
rect 13412 3352 13457 3380
rect 13412 3340 13418 3352
rect 13538 3340 13544 3392
rect 13596 3380 13602 3392
rect 14384 3380 14412 3420
rect 16114 3408 16120 3420
rect 16172 3448 16178 3460
rect 16482 3448 16488 3460
rect 16172 3420 16488 3448
rect 16172 3408 16178 3420
rect 16482 3408 16488 3420
rect 16540 3408 16546 3460
rect 16850 3408 16856 3460
rect 16908 3448 16914 3460
rect 17512 3448 17540 3624
rect 19150 3612 19156 3624
rect 19208 3612 19214 3664
rect 17770 3544 17776 3596
rect 17828 3584 17834 3596
rect 18141 3587 18199 3593
rect 18141 3584 18153 3587
rect 17828 3556 18153 3584
rect 17828 3544 17834 3556
rect 18141 3553 18153 3556
rect 18187 3553 18199 3587
rect 18141 3547 18199 3553
rect 18046 3516 18052 3528
rect 18007 3488 18052 3516
rect 18046 3476 18052 3488
rect 18104 3476 18110 3528
rect 16908 3420 17540 3448
rect 17957 3451 18015 3457
rect 16908 3408 16914 3420
rect 17957 3417 17969 3451
rect 18003 3448 18015 3451
rect 18322 3448 18328 3460
rect 18003 3420 18328 3448
rect 18003 3417 18015 3420
rect 17957 3411 18015 3417
rect 18322 3408 18328 3420
rect 18380 3408 18386 3460
rect 13596 3352 14412 3380
rect 14553 3383 14611 3389
rect 13596 3340 13602 3352
rect 14553 3349 14565 3383
rect 14599 3380 14611 3383
rect 14921 3383 14979 3389
rect 14921 3380 14933 3383
rect 14599 3352 14933 3380
rect 14599 3349 14611 3352
rect 14553 3343 14611 3349
rect 14921 3349 14933 3352
rect 14967 3349 14979 3383
rect 15286 3380 15292 3392
rect 15247 3352 15292 3380
rect 14921 3343 14979 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15381 3383 15439 3389
rect 15381 3349 15393 3383
rect 15427 3380 15439 3383
rect 15746 3380 15752 3392
rect 15427 3352 15752 3380
rect 15427 3349 15439 3352
rect 15381 3343 15439 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 15930 3380 15936 3392
rect 15891 3352 15936 3380
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16390 3380 16396 3392
rect 16351 3352 16396 3380
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 17405 3383 17463 3389
rect 17405 3349 17417 3383
rect 17451 3380 17463 3383
rect 17586 3380 17592 3392
rect 17451 3352 17592 3380
rect 17451 3349 17463 3352
rect 17405 3343 17463 3349
rect 17586 3340 17592 3352
rect 17644 3340 17650 3392
rect 1104 3290 18860 3312
rect 1104 3238 5398 3290
rect 5450 3238 5462 3290
rect 5514 3238 5526 3290
rect 5578 3238 5590 3290
rect 5642 3238 5654 3290
rect 5706 3238 9846 3290
rect 9898 3238 9910 3290
rect 9962 3238 9974 3290
rect 10026 3238 10038 3290
rect 10090 3238 10102 3290
rect 10154 3238 14294 3290
rect 14346 3238 14358 3290
rect 14410 3238 14422 3290
rect 14474 3238 14486 3290
rect 14538 3238 14550 3290
rect 14602 3238 18860 3290
rect 1104 3216 18860 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 1670 3176 1676 3188
rect 1627 3148 1676 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1670 3136 1676 3148
rect 1728 3136 1734 3188
rect 1946 3176 1952 3188
rect 1907 3148 1952 3176
rect 1946 3136 1952 3148
rect 2004 3136 2010 3188
rect 2041 3179 2099 3185
rect 2041 3145 2053 3179
rect 2087 3176 2099 3179
rect 2498 3176 2504 3188
rect 2087 3148 2504 3176
rect 2087 3145 2099 3148
rect 2041 3139 2099 3145
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 3142 3136 3148 3188
rect 3200 3176 3206 3188
rect 6730 3176 6736 3188
rect 3200 3148 6592 3176
rect 6691 3148 6736 3176
rect 3200 3136 3206 3148
rect 2774 3108 2780 3120
rect 2735 3080 2780 3108
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 4338 3108 4344 3120
rect 4299 3080 4344 3108
rect 4338 3068 4344 3080
rect 4396 3068 4402 3120
rect 4985 3111 5043 3117
rect 4985 3108 4997 3111
rect 4724 3080 4997 3108
rect 4724 3052 4752 3080
rect 4985 3077 4997 3080
rect 5031 3077 5043 3111
rect 5810 3108 5816 3120
rect 4985 3071 5043 3077
rect 5092 3080 5816 3108
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 4062 3040 4068 3052
rect 1504 3012 4068 3040
rect 1302 2932 1308 2984
rect 1360 2972 1366 2984
rect 1504 2972 1532 3012
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4706 3000 4712 3052
rect 4764 3000 4770 3052
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 4948 3012 4993 3040
rect 4948 3000 4954 3012
rect 1360 2944 1532 2972
rect 1857 2975 1915 2981
rect 1360 2932 1366 2944
rect 1857 2941 1869 2975
rect 1903 2972 1915 2975
rect 2130 2972 2136 2984
rect 1903 2944 2136 2972
rect 1903 2941 1915 2944
rect 1857 2935 1915 2941
rect 2130 2932 2136 2944
rect 2188 2932 2194 2984
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 5092 2972 5120 3080
rect 5810 3068 5816 3080
rect 5868 3068 5874 3120
rect 5258 3000 5264 3052
rect 5316 3040 5322 3052
rect 5721 3043 5779 3049
rect 5721 3040 5733 3043
rect 5316 3012 5733 3040
rect 5316 3000 5322 3012
rect 5721 3009 5733 3012
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 4028 2944 5120 2972
rect 5169 2975 5227 2981
rect 4028 2932 4034 2944
rect 5169 2941 5181 2975
rect 5215 2972 5227 2975
rect 5442 2972 5448 2984
rect 5215 2944 5448 2972
rect 5215 2941 5227 2944
rect 5169 2935 5227 2941
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5810 2972 5816 2984
rect 5771 2944 5816 2972
rect 5810 2932 5816 2944
rect 5868 2932 5874 2984
rect 5994 2972 6000 2984
rect 5955 2944 6000 2972
rect 5994 2932 6000 2944
rect 6052 2932 6058 2984
rect 2222 2864 2228 2916
rect 2280 2904 2286 2916
rect 2409 2907 2467 2913
rect 2409 2904 2421 2907
rect 2280 2876 2421 2904
rect 2280 2864 2286 2876
rect 2409 2873 2421 2876
rect 2455 2873 2467 2907
rect 2409 2867 2467 2873
rect 2958 2864 2964 2916
rect 3016 2904 3022 2916
rect 6457 2907 6515 2913
rect 6457 2904 6469 2907
rect 3016 2876 6469 2904
rect 3016 2864 3022 2876
rect 6457 2873 6469 2876
rect 6503 2873 6515 2907
rect 6457 2867 6515 2873
rect 1210 2796 1216 2848
rect 1268 2836 1274 2848
rect 2130 2836 2136 2848
rect 1268 2808 2136 2836
rect 1268 2796 1274 2808
rect 2130 2796 2136 2808
rect 2188 2796 2194 2848
rect 2498 2796 2504 2848
rect 2556 2836 2562 2848
rect 4062 2836 4068 2848
rect 2556 2808 4068 2836
rect 2556 2796 2562 2808
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 4522 2836 4528 2848
rect 4483 2808 4528 2836
rect 4522 2796 4528 2808
rect 4580 2796 4586 2848
rect 4614 2796 4620 2848
rect 4672 2836 4678 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 4672 2808 5365 2836
rect 4672 2796 4678 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 5442 2796 5448 2848
rect 5500 2836 5506 2848
rect 5994 2836 6000 2848
rect 5500 2808 6000 2836
rect 5500 2796 5506 2808
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6564 2836 6592 3148
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 6914 3136 6920 3188
rect 6972 3136 6978 3188
rect 7190 3136 7196 3188
rect 7248 3176 7254 3188
rect 8294 3176 8300 3188
rect 7248 3148 7613 3176
rect 8255 3148 8300 3176
rect 7248 3136 7254 3148
rect 6932 3108 6960 3136
rect 7101 3111 7159 3117
rect 7101 3108 7113 3111
rect 6932 3080 7113 3108
rect 7101 3077 7113 3080
rect 7147 3077 7159 3111
rect 7101 3071 7159 3077
rect 7585 3053 7613 3148
rect 8294 3136 8300 3148
rect 8352 3136 8358 3188
rect 8478 3136 8484 3188
rect 8536 3176 8542 3188
rect 9398 3176 9404 3188
rect 8536 3148 9404 3176
rect 8536 3136 8542 3148
rect 9398 3136 9404 3148
rect 9456 3136 9462 3188
rect 10137 3179 10195 3185
rect 10137 3145 10149 3179
rect 10183 3176 10195 3179
rect 10318 3176 10324 3188
rect 10183 3148 10324 3176
rect 10183 3145 10195 3148
rect 10137 3139 10195 3145
rect 10318 3136 10324 3148
rect 10376 3136 10382 3188
rect 10870 3176 10876 3188
rect 10831 3148 10876 3176
rect 10870 3136 10876 3148
rect 10928 3136 10934 3188
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 11698 3136 11704 3188
rect 11756 3176 11762 3188
rect 13814 3176 13820 3188
rect 11756 3148 13820 3176
rect 11756 3136 11762 3148
rect 13814 3136 13820 3148
rect 13872 3136 13878 3188
rect 14090 3176 14096 3188
rect 14051 3148 14096 3176
rect 14090 3136 14096 3148
rect 14148 3136 14154 3188
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 14553 3179 14611 3185
rect 14553 3176 14565 3179
rect 14240 3148 14565 3176
rect 14240 3136 14246 3148
rect 14553 3145 14565 3148
rect 14599 3145 14611 3179
rect 14553 3139 14611 3145
rect 15105 3179 15163 3185
rect 15105 3145 15117 3179
rect 15151 3145 15163 3179
rect 15378 3176 15384 3188
rect 15339 3148 15384 3176
rect 15105 3139 15163 3145
rect 9582 3108 9588 3120
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 7006 3040 7012 3052
rect 6687 3012 7012 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 7006 3000 7012 3012
rect 7064 3000 7070 3052
rect 7553 3047 7613 3053
rect 7553 3013 7565 3047
rect 7599 3016 7613 3047
rect 7760 3080 9588 3108
rect 7599 3013 7611 3016
rect 7553 3007 7611 3013
rect 7190 2972 7196 2984
rect 7151 2944 7196 2972
rect 7190 2932 7196 2944
rect 7248 2932 7254 2984
rect 7374 2972 7380 2984
rect 7335 2944 7380 2972
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7760 2972 7788 3080
rect 9582 3068 9588 3080
rect 9640 3068 9646 3120
rect 10045 3111 10103 3117
rect 10045 3077 10057 3111
rect 10091 3108 10103 3111
rect 10594 3108 10600 3120
rect 10091 3080 10600 3108
rect 10091 3077 10103 3080
rect 10045 3071 10103 3077
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 10060 3040 10088 3071
rect 10594 3068 10600 3080
rect 10652 3068 10658 3120
rect 10686 3068 10692 3120
rect 10744 3108 10750 3120
rect 11885 3111 11943 3117
rect 11885 3108 11897 3111
rect 10744 3080 11897 3108
rect 10744 3068 10750 3080
rect 11885 3077 11897 3080
rect 11931 3077 11943 3111
rect 11885 3071 11943 3077
rect 11977 3111 12035 3117
rect 11977 3077 11989 3111
rect 12023 3108 12035 3111
rect 12888 3111 12946 3117
rect 12023 3080 12848 3108
rect 12023 3077 12035 3080
rect 11977 3071 12035 3077
rect 10502 3040 10508 3052
rect 7984 3012 10088 3040
rect 10244 3012 10508 3040
rect 7984 3000 7990 3012
rect 7484 2944 7788 2972
rect 6638 2864 6644 2916
rect 6696 2904 6702 2916
rect 7484 2904 7512 2944
rect 7834 2932 7840 2984
rect 7892 2972 7898 2984
rect 8478 2972 8484 2984
rect 7892 2944 8484 2972
rect 7892 2932 7898 2944
rect 8478 2932 8484 2944
rect 8536 2932 8542 2984
rect 10244 2981 10272 3012
rect 10502 3000 10508 3012
rect 10560 3000 10566 3052
rect 10778 3000 10784 3052
rect 10836 3040 10842 3052
rect 12526 3040 12532 3052
rect 10836 3012 11100 3040
rect 12487 3012 12532 3040
rect 10836 3000 10842 3012
rect 10229 2975 10287 2981
rect 10229 2941 10241 2975
rect 10275 2941 10287 2975
rect 10962 2972 10968 2984
rect 10229 2935 10287 2941
rect 10336 2944 10824 2972
rect 10923 2944 10968 2972
rect 6696 2876 7512 2904
rect 7745 2907 7803 2913
rect 6696 2864 6702 2876
rect 7745 2873 7757 2907
rect 7791 2904 7803 2907
rect 7791 2876 8095 2904
rect 7791 2873 7803 2876
rect 7745 2867 7803 2873
rect 7190 2836 7196 2848
rect 6564 2808 7196 2836
rect 7190 2796 7196 2808
rect 7248 2796 7254 2848
rect 8067 2836 8095 2876
rect 8248 2864 8254 2916
rect 8306 2904 8312 2916
rect 10336 2904 10364 2944
rect 10502 2904 10508 2916
rect 8306 2876 10364 2904
rect 10463 2876 10508 2904
rect 8306 2864 8312 2876
rect 10502 2864 10508 2876
rect 10560 2864 10566 2916
rect 10796 2904 10824 2944
rect 10962 2932 10968 2944
rect 11020 2932 11026 2984
rect 11072 2981 11100 3012
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12820 3040 12848 3080
rect 12888 3077 12900 3111
rect 12934 3108 12946 3111
rect 14734 3108 14740 3120
rect 12934 3080 14740 3108
rect 12934 3077 12946 3080
rect 12888 3071 12946 3077
rect 14734 3068 14740 3080
rect 14792 3068 14798 3120
rect 15120 3108 15148 3139
rect 15378 3136 15384 3148
rect 15436 3136 15442 3188
rect 15562 3136 15568 3188
rect 15620 3176 15626 3188
rect 15749 3179 15807 3185
rect 15749 3176 15761 3179
rect 15620 3148 15761 3176
rect 15620 3136 15626 3148
rect 15749 3145 15761 3148
rect 15795 3145 15807 3179
rect 15749 3139 15807 3145
rect 15841 3179 15899 3185
rect 15841 3145 15853 3179
rect 15887 3176 15899 3179
rect 16390 3176 16396 3188
rect 15887 3148 16396 3176
rect 15887 3145 15899 3148
rect 15841 3139 15899 3145
rect 16390 3136 16396 3148
rect 16448 3136 16454 3188
rect 16482 3136 16488 3188
rect 16540 3176 16546 3188
rect 17497 3179 17555 3185
rect 17497 3176 17509 3179
rect 16540 3148 17509 3176
rect 16540 3136 16546 3148
rect 17497 3145 17509 3148
rect 17543 3145 17555 3179
rect 17954 3176 17960 3188
rect 17915 3148 17960 3176
rect 17497 3139 17555 3145
rect 17954 3136 17960 3148
rect 18012 3136 18018 3188
rect 18322 3136 18328 3188
rect 18380 3176 18386 3188
rect 19334 3176 19340 3188
rect 18380 3148 19340 3176
rect 18380 3136 18386 3148
rect 19334 3136 19340 3148
rect 19392 3136 19398 3188
rect 16022 3108 16028 3120
rect 15120 3080 16028 3108
rect 16022 3068 16028 3080
rect 16080 3068 16086 3120
rect 17034 3108 17040 3120
rect 16995 3080 17040 3108
rect 17034 3068 17040 3080
rect 17092 3068 17098 3120
rect 18414 3108 18420 3120
rect 18375 3080 18420 3108
rect 18414 3068 18420 3080
rect 18472 3068 18478 3120
rect 13906 3040 13912 3052
rect 12820 3012 13912 3040
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14458 3040 14464 3052
rect 14419 3012 14464 3040
rect 14458 3000 14464 3012
rect 14516 3000 14522 3052
rect 14918 3040 14924 3052
rect 14879 3012 14924 3040
rect 14918 3000 14924 3012
rect 14976 3000 14982 3052
rect 15286 3000 15292 3052
rect 15344 3040 15350 3052
rect 15838 3040 15844 3052
rect 15344 3012 15844 3040
rect 15344 3000 15350 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 16114 3000 16120 3052
rect 16172 3040 16178 3052
rect 16209 3043 16267 3049
rect 16209 3040 16221 3043
rect 16172 3012 16221 3040
rect 16172 3000 16178 3012
rect 16209 3009 16221 3012
rect 16255 3009 16267 3043
rect 16666 3040 16672 3052
rect 16627 3012 16672 3040
rect 16209 3003 16267 3009
rect 16666 3000 16672 3012
rect 16724 3000 16730 3052
rect 16758 3000 16764 3052
rect 16816 3040 16822 3052
rect 17589 3043 17647 3049
rect 17589 3040 17601 3043
rect 16816 3012 17601 3040
rect 16816 3000 16822 3012
rect 17589 3009 17601 3012
rect 17635 3009 17647 3043
rect 17589 3003 17647 3009
rect 18049 3043 18107 3049
rect 18049 3009 18061 3043
rect 18095 3040 18107 3043
rect 19886 3040 19892 3052
rect 18095 3012 19892 3040
rect 18095 3009 18107 3012
rect 18049 3003 18107 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 11057 2975 11115 2981
rect 11057 2941 11069 2975
rect 11103 2941 11115 2975
rect 12066 2972 12072 2984
rect 12027 2944 12072 2972
rect 11057 2935 11115 2941
rect 12066 2932 12072 2944
rect 12124 2932 12130 2984
rect 12158 2932 12164 2984
rect 12216 2972 12222 2984
rect 12621 2975 12679 2981
rect 12621 2972 12633 2975
rect 12216 2944 12633 2972
rect 12216 2932 12222 2944
rect 12621 2941 12633 2944
rect 12667 2941 12679 2975
rect 12621 2935 12679 2941
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 14366 2972 14372 2984
rect 13780 2944 14372 2972
rect 13780 2932 13786 2944
rect 14366 2932 14372 2944
rect 14424 2932 14430 2984
rect 14642 2972 14648 2984
rect 14603 2944 14648 2972
rect 14642 2932 14648 2944
rect 14700 2932 14706 2984
rect 15010 2932 15016 2984
rect 15068 2972 15074 2984
rect 15933 2975 15991 2981
rect 15933 2972 15945 2975
rect 15068 2944 15945 2972
rect 15068 2932 15074 2944
rect 15933 2941 15945 2944
rect 15979 2941 15991 2975
rect 15933 2935 15991 2941
rect 17405 2975 17463 2981
rect 17405 2941 17417 2975
rect 17451 2972 17463 2975
rect 17770 2972 17776 2984
rect 17451 2944 17776 2972
rect 17451 2941 17463 2944
rect 17405 2935 17463 2941
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18506 2972 18512 2984
rect 18012 2944 18512 2972
rect 18012 2932 18018 2944
rect 18506 2932 18512 2944
rect 18564 2932 18570 2984
rect 10796 2876 11008 2904
rect 9122 2836 9128 2848
rect 8067 2808 9128 2836
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9677 2839 9735 2845
rect 9677 2836 9689 2839
rect 9456 2808 9689 2836
rect 9456 2796 9462 2808
rect 9677 2805 9689 2808
rect 9723 2805 9735 2839
rect 10980 2836 11008 2876
rect 11606 2864 11612 2916
rect 11664 2904 11670 2916
rect 12345 2907 12403 2913
rect 12345 2904 12357 2907
rect 11664 2876 12357 2904
rect 11664 2864 11670 2876
rect 12345 2873 12357 2876
rect 12391 2873 12403 2907
rect 16393 2907 16451 2913
rect 16393 2904 16405 2907
rect 12345 2867 12403 2873
rect 13556 2876 16405 2904
rect 12894 2836 12900 2848
rect 10980 2808 12900 2836
rect 9677 2799 9735 2805
rect 12894 2796 12900 2808
rect 12952 2796 12958 2848
rect 13262 2796 13268 2848
rect 13320 2836 13326 2848
rect 13556 2836 13584 2876
rect 16393 2873 16405 2876
rect 16439 2873 16451 2907
rect 16393 2867 16451 2873
rect 16853 2907 16911 2913
rect 16853 2873 16865 2907
rect 16899 2904 16911 2907
rect 19426 2904 19432 2916
rect 16899 2876 19432 2904
rect 16899 2873 16911 2876
rect 16853 2867 16911 2873
rect 19426 2864 19432 2876
rect 19484 2864 19490 2916
rect 13320 2808 13584 2836
rect 14001 2839 14059 2845
rect 13320 2796 13326 2808
rect 14001 2805 14013 2839
rect 14047 2836 14059 2839
rect 14642 2836 14648 2848
rect 14047 2808 14648 2836
rect 14047 2805 14059 2808
rect 14001 2799 14059 2805
rect 14642 2796 14648 2808
rect 14700 2796 14706 2848
rect 14918 2796 14924 2848
rect 14976 2836 14982 2848
rect 17954 2836 17960 2848
rect 14976 2808 17960 2836
rect 14976 2796 14982 2808
rect 17954 2796 17960 2808
rect 18012 2796 18018 2848
rect 18230 2836 18236 2848
rect 18191 2808 18236 2836
rect 18230 2796 18236 2808
rect 18288 2796 18294 2848
rect 1104 2746 18860 2768
rect 1104 2694 3174 2746
rect 3226 2694 3238 2746
rect 3290 2694 3302 2746
rect 3354 2694 3366 2746
rect 3418 2694 3430 2746
rect 3482 2694 7622 2746
rect 7674 2694 7686 2746
rect 7738 2694 7750 2746
rect 7802 2694 7814 2746
rect 7866 2694 7878 2746
rect 7930 2694 12070 2746
rect 12122 2694 12134 2746
rect 12186 2694 12198 2746
rect 12250 2694 12262 2746
rect 12314 2694 12326 2746
rect 12378 2694 16518 2746
rect 16570 2694 16582 2746
rect 16634 2694 16646 2746
rect 16698 2694 16710 2746
rect 16762 2694 16774 2746
rect 16826 2694 18860 2746
rect 1104 2672 18860 2694
rect 2590 2632 2596 2644
rect 2056 2604 2596 2632
rect 2056 2505 2084 2604
rect 2590 2592 2596 2604
rect 2648 2632 2654 2644
rect 2958 2632 2964 2644
rect 2648 2604 2964 2632
rect 2648 2592 2654 2604
rect 2958 2592 2964 2604
rect 3016 2592 3022 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3878 2632 3884 2644
rect 3651 2604 3884 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3878 2592 3884 2604
rect 3936 2592 3942 2644
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 4617 2635 4675 2641
rect 4617 2632 4629 2635
rect 4120 2604 4629 2632
rect 4120 2592 4126 2604
rect 4617 2601 4629 2604
rect 4663 2601 4675 2635
rect 4617 2595 4675 2601
rect 5902 2592 5908 2644
rect 5960 2632 5966 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 5960 2604 7573 2632
rect 5960 2592 5966 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7561 2595 7619 2601
rect 9122 2592 9128 2644
rect 9180 2632 9186 2644
rect 10410 2632 10416 2644
rect 9180 2604 10416 2632
rect 9180 2592 9186 2604
rect 10410 2592 10416 2604
rect 10468 2592 10474 2644
rect 10686 2632 10692 2644
rect 10647 2604 10692 2632
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 13906 2592 13912 2644
rect 13964 2632 13970 2644
rect 14093 2635 14151 2641
rect 14093 2632 14105 2635
rect 13964 2604 14105 2632
rect 13964 2592 13970 2604
rect 14093 2601 14105 2604
rect 14139 2601 14151 2635
rect 14093 2595 14151 2601
rect 14182 2592 14188 2644
rect 14240 2592 14246 2644
rect 14366 2592 14372 2644
rect 14424 2632 14430 2644
rect 15565 2635 15623 2641
rect 15565 2632 15577 2635
rect 14424 2604 15577 2632
rect 14424 2592 14430 2604
rect 15565 2601 15577 2604
rect 15611 2601 15623 2635
rect 15565 2595 15623 2601
rect 3418 2524 3424 2576
rect 3476 2564 3482 2576
rect 6178 2564 6184 2576
rect 3476 2536 3521 2564
rect 6139 2536 6184 2564
rect 3476 2524 3482 2536
rect 6178 2524 6184 2536
rect 6236 2524 6242 2576
rect 7190 2524 7196 2576
rect 7248 2564 7254 2576
rect 8202 2564 8208 2576
rect 7248 2536 8208 2564
rect 7248 2524 7254 2536
rect 8202 2524 8208 2536
rect 8260 2524 8266 2576
rect 9674 2564 9680 2576
rect 8956 2536 9680 2564
rect 2041 2499 2099 2505
rect 2041 2465 2053 2499
rect 2087 2465 2099 2499
rect 2041 2459 2099 2465
rect 2133 2499 2191 2505
rect 2133 2465 2145 2499
rect 2179 2496 2191 2499
rect 2498 2496 2504 2508
rect 2179 2468 2504 2496
rect 2179 2465 2191 2468
rect 2133 2459 2191 2465
rect 2498 2456 2504 2468
rect 2556 2456 2562 2508
rect 2777 2499 2835 2505
rect 2777 2465 2789 2499
rect 2823 2465 2835 2499
rect 2777 2459 2835 2465
rect 1762 2428 1768 2440
rect 1723 2400 1768 2428
rect 1762 2388 1768 2400
rect 1820 2388 1826 2440
rect 2792 2428 2820 2459
rect 2866 2456 2872 2508
rect 2924 2496 2930 2508
rect 2961 2499 3019 2505
rect 2961 2496 2973 2499
rect 2924 2468 2973 2496
rect 2924 2456 2930 2468
rect 2961 2465 2973 2468
rect 3007 2465 3019 2499
rect 2961 2459 3019 2465
rect 3142 2456 3148 2508
rect 3200 2496 3206 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3200 2468 3893 2496
rect 3200 2456 3206 2468
rect 3881 2465 3893 2468
rect 3927 2496 3939 2499
rect 4430 2496 4436 2508
rect 3927 2468 4436 2496
rect 3927 2465 3939 2468
rect 3881 2459 3939 2465
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 5261 2499 5319 2505
rect 4632 2468 5120 2496
rect 3050 2428 3056 2440
rect 2792 2400 2912 2428
rect 3011 2400 3056 2428
rect 2884 2360 2912 2400
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3786 2428 3792 2440
rect 3160 2400 3792 2428
rect 3160 2360 3188 2400
rect 3786 2388 3792 2400
rect 3844 2388 3850 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4246 2428 4252 2440
rect 4203 2400 4252 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4632 2428 4660 2468
rect 4982 2428 4988 2440
rect 4448 2400 4660 2428
rect 4943 2400 4988 2428
rect 2608 2332 2774 2360
rect 2884 2332 3188 2360
rect 4065 2363 4123 2369
rect 1578 2292 1584 2304
rect 1539 2264 1584 2292
rect 1578 2252 1584 2264
rect 1636 2252 1642 2304
rect 2222 2292 2228 2304
rect 2183 2264 2228 2292
rect 2222 2252 2228 2264
rect 2280 2252 2286 2304
rect 2608 2301 2636 2332
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2261 2651 2295
rect 2746 2292 2774 2332
rect 4065 2329 4077 2363
rect 4111 2360 4123 2363
rect 4338 2360 4344 2372
rect 4111 2332 4344 2360
rect 4111 2329 4123 2332
rect 4065 2323 4123 2329
rect 4338 2320 4344 2332
rect 4396 2320 4402 2372
rect 4448 2292 4476 2400
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5092 2428 5120 2468
rect 5261 2465 5273 2499
rect 5307 2496 5319 2499
rect 5442 2496 5448 2508
rect 5307 2468 5448 2496
rect 5307 2465 5319 2468
rect 5261 2459 5319 2465
rect 5442 2456 5448 2468
rect 5500 2456 5506 2508
rect 5629 2499 5687 2505
rect 5629 2465 5641 2499
rect 5675 2496 5687 2499
rect 6086 2496 6092 2508
rect 5675 2468 6092 2496
rect 5675 2465 5687 2468
rect 5629 2459 5687 2465
rect 6086 2456 6092 2468
rect 6144 2456 6150 2508
rect 6362 2456 6368 2508
rect 6420 2496 6426 2508
rect 6822 2496 6828 2508
rect 6420 2468 6828 2496
rect 6420 2456 6426 2468
rect 6822 2456 6828 2468
rect 6880 2496 6886 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6880 2468 6929 2496
rect 6880 2456 6886 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7374 2456 7380 2508
rect 7432 2496 7438 2508
rect 8110 2496 8116 2508
rect 7432 2468 8116 2496
rect 7432 2456 7438 2468
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 8956 2505 8984 2536
rect 9674 2524 9680 2536
rect 9732 2524 9738 2576
rect 10502 2524 10508 2576
rect 10560 2564 10566 2576
rect 10962 2564 10968 2576
rect 10560 2536 10968 2564
rect 10560 2524 10566 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 14200 2564 14228 2592
rect 11440 2536 14228 2564
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 8220 2468 8953 2496
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5092 2400 5825 2428
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 6638 2428 6644 2440
rect 6599 2400 6644 2428
rect 5813 2391 5871 2397
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 8220 2428 8248 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 9214 2496 9220 2508
rect 9175 2468 9220 2496
rect 8941 2459 8999 2465
rect 9214 2456 9220 2468
rect 9272 2456 9278 2508
rect 9398 2496 9404 2508
rect 9359 2468 9404 2496
rect 9398 2456 9404 2468
rect 9456 2456 9462 2508
rect 10137 2499 10195 2505
rect 10137 2496 10149 2499
rect 9600 2468 10149 2496
rect 8478 2428 8484 2440
rect 7392 2400 8248 2428
rect 8439 2400 8484 2428
rect 5721 2363 5779 2369
rect 5721 2360 5733 2363
rect 4540 2332 5733 2360
rect 4540 2301 4568 2332
rect 5721 2329 5733 2332
rect 5767 2329 5779 2363
rect 7392 2360 7420 2400
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 9030 2388 9036 2440
rect 9088 2428 9094 2440
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9088 2400 9505 2428
rect 9088 2388 9094 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9493 2391 9551 2397
rect 8021 2363 8079 2369
rect 8021 2360 8033 2363
rect 5721 2323 5779 2329
rect 6288 2332 7420 2360
rect 7484 2332 8033 2360
rect 2746 2264 4476 2292
rect 4525 2295 4583 2301
rect 2593 2255 2651 2261
rect 4525 2261 4537 2295
rect 4571 2261 4583 2295
rect 4525 2255 4583 2261
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2292 5135 2295
rect 6288 2292 6316 2332
rect 6454 2292 6460 2304
rect 5123 2264 6316 2292
rect 6415 2264 6460 2292
rect 5123 2261 5135 2264
rect 5077 2255 5135 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 7006 2292 7012 2304
rect 6967 2264 7012 2292
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7098 2252 7104 2304
rect 7156 2292 7162 2304
rect 7484 2301 7512 2332
rect 8021 2329 8033 2332
rect 8067 2329 8079 2363
rect 8021 2323 8079 2329
rect 9398 2320 9404 2372
rect 9456 2360 9462 2372
rect 9600 2360 9628 2468
rect 10137 2465 10149 2468
rect 10183 2496 10195 2499
rect 11440 2496 11468 2536
rect 14734 2524 14740 2576
rect 14792 2564 14798 2576
rect 16301 2567 16359 2573
rect 16301 2564 16313 2567
rect 14792 2536 16313 2564
rect 14792 2524 14798 2536
rect 16301 2533 16313 2536
rect 16347 2533 16359 2567
rect 18046 2564 18052 2576
rect 18007 2536 18052 2564
rect 16301 2527 16359 2533
rect 18046 2524 18052 2536
rect 18104 2524 18110 2576
rect 12066 2496 12072 2508
rect 10183 2468 11468 2496
rect 12027 2468 12072 2496
rect 10183 2465 10195 2468
rect 10137 2459 10195 2465
rect 12066 2456 12072 2468
rect 12124 2496 12130 2508
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12124 2468 12541 2496
rect 12124 2456 12130 2468
rect 12529 2465 12541 2468
rect 12575 2496 12587 2499
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 12575 2468 13277 2496
rect 12575 2465 12587 2468
rect 12529 2459 12587 2465
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 13265 2459 13323 2465
rect 14366 2456 14372 2508
rect 14424 2496 14430 2508
rect 14645 2499 14703 2505
rect 14645 2496 14657 2499
rect 14424 2468 14657 2496
rect 14424 2456 14430 2468
rect 14645 2465 14657 2468
rect 14691 2465 14703 2499
rect 14645 2459 14703 2465
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 10321 2431 10379 2437
rect 10321 2428 10333 2431
rect 9824 2400 10333 2428
rect 9824 2388 9830 2400
rect 10321 2397 10333 2400
rect 10367 2397 10379 2431
rect 10321 2391 10379 2397
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10781 2431 10839 2437
rect 10468 2424 10732 2428
rect 10781 2424 10793 2431
rect 10468 2400 10793 2424
rect 10468 2388 10474 2400
rect 10704 2397 10793 2400
rect 10827 2397 10839 2431
rect 10704 2396 10839 2397
rect 10781 2391 10839 2396
rect 11333 2431 11391 2437
rect 11333 2397 11345 2431
rect 11379 2428 11391 2431
rect 11885 2431 11943 2437
rect 11379 2400 11836 2428
rect 11379 2397 11391 2400
rect 11333 2391 11391 2397
rect 9456 2332 9628 2360
rect 10229 2363 10287 2369
rect 9456 2320 9462 2332
rect 10229 2329 10241 2363
rect 10275 2360 10287 2363
rect 11808 2360 11836 2400
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 11974 2428 11980 2440
rect 11931 2400 11980 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 11974 2388 11980 2400
rect 12032 2388 12038 2440
rect 12250 2388 12256 2440
rect 12308 2428 12314 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 12308 2400 13461 2428
rect 12308 2388 12314 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 14553 2431 14611 2437
rect 14553 2428 14565 2431
rect 13449 2391 13507 2397
rect 13832 2400 14565 2428
rect 12342 2360 12348 2372
rect 10275 2332 11560 2360
rect 11808 2332 12348 2360
rect 10275 2329 10287 2332
rect 10229 2323 10287 2329
rect 7469 2295 7527 2301
rect 7156 2264 7201 2292
rect 7156 2252 7162 2264
rect 7469 2261 7481 2295
rect 7515 2261 7527 2295
rect 7926 2292 7932 2304
rect 7887 2264 7932 2292
rect 7469 2255 7527 2261
rect 7926 2252 7932 2264
rect 7984 2252 7990 2304
rect 8662 2292 8668 2304
rect 8623 2264 8668 2292
rect 8662 2252 8668 2264
rect 8720 2252 8726 2304
rect 9861 2295 9919 2301
rect 9861 2261 9873 2295
rect 9907 2292 9919 2295
rect 10502 2292 10508 2304
rect 9907 2264 10508 2292
rect 9907 2261 9919 2264
rect 9861 2255 9919 2261
rect 10502 2252 10508 2264
rect 10560 2252 10566 2304
rect 10962 2292 10968 2304
rect 10923 2264 10968 2292
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11146 2292 11152 2304
rect 11107 2264 11152 2292
rect 11146 2252 11152 2264
rect 11204 2252 11210 2304
rect 11532 2301 11560 2332
rect 12342 2320 12348 2332
rect 12400 2320 12406 2372
rect 12894 2320 12900 2372
rect 12952 2360 12958 2372
rect 13541 2363 13599 2369
rect 13541 2360 13553 2363
rect 12952 2332 13553 2360
rect 12952 2320 12958 2332
rect 13541 2329 13553 2332
rect 13587 2329 13599 2363
rect 13541 2323 13599 2329
rect 11517 2295 11575 2301
rect 11517 2261 11529 2295
rect 11563 2261 11575 2295
rect 11974 2292 11980 2304
rect 11935 2264 11980 2292
rect 11517 2255 11575 2261
rect 11974 2252 11980 2264
rect 12032 2252 12038 2304
rect 12618 2292 12624 2304
rect 12579 2264 12624 2292
rect 12618 2252 12624 2264
rect 12676 2252 12682 2304
rect 12710 2252 12716 2304
rect 12768 2292 12774 2304
rect 13081 2295 13139 2301
rect 12768 2264 12813 2292
rect 12768 2252 12774 2264
rect 13081 2261 13093 2295
rect 13127 2292 13139 2295
rect 13832 2292 13860 2400
rect 14553 2397 14565 2400
rect 14599 2397 14611 2431
rect 14918 2428 14924 2440
rect 14879 2400 14924 2428
rect 14553 2391 14611 2397
rect 14918 2388 14924 2400
rect 14976 2388 14982 2440
rect 15654 2428 15660 2440
rect 15615 2400 15660 2428
rect 15654 2388 15660 2400
rect 15712 2388 15718 2440
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 17402 2428 17408 2440
rect 17363 2400 17408 2428
rect 17402 2388 17408 2400
rect 17460 2388 17466 2440
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18141 2431 18199 2437
rect 18141 2428 18153 2431
rect 18012 2400 18153 2428
rect 18012 2388 18018 2400
rect 18141 2397 18153 2400
rect 18187 2397 18199 2431
rect 18141 2391 18199 2397
rect 14461 2363 14519 2369
rect 14461 2360 14473 2363
rect 13924 2332 14473 2360
rect 13924 2301 13952 2332
rect 14461 2329 14473 2332
rect 14507 2329 14519 2363
rect 14461 2323 14519 2329
rect 13127 2264 13860 2292
rect 13909 2295 13967 2301
rect 13127 2261 13139 2264
rect 13081 2255 13139 2261
rect 13909 2261 13921 2295
rect 13955 2261 13967 2295
rect 16390 2292 16396 2304
rect 16351 2264 16396 2292
rect 13909 2255 13967 2261
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 17310 2292 17316 2304
rect 17271 2264 17316 2292
rect 17310 2252 17316 2264
rect 17368 2252 17374 2304
rect 18138 2252 18144 2304
rect 18196 2292 18202 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18196 2264 18337 2292
rect 18196 2252 18202 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 1104 2202 18860 2224
rect 1104 2150 5398 2202
rect 5450 2150 5462 2202
rect 5514 2150 5526 2202
rect 5578 2150 5590 2202
rect 5642 2150 5654 2202
rect 5706 2150 9846 2202
rect 9898 2150 9910 2202
rect 9962 2150 9974 2202
rect 10026 2150 10038 2202
rect 10090 2150 10102 2202
rect 10154 2150 14294 2202
rect 14346 2150 14358 2202
rect 14410 2150 14422 2202
rect 14474 2150 14486 2202
rect 14538 2150 14550 2202
rect 14602 2150 18860 2202
rect 1104 2128 18860 2150
rect 4062 2048 4068 2100
rect 4120 2088 4126 2100
rect 8662 2088 8668 2100
rect 4120 2060 8668 2088
rect 4120 2048 4126 2060
rect 8662 2048 8668 2060
rect 8720 2048 8726 2100
rect 8938 2048 8944 2100
rect 8996 2088 9002 2100
rect 8996 2060 10824 2088
rect 8996 2048 9002 2060
rect 2222 1980 2228 2032
rect 2280 2020 2286 2032
rect 4614 2020 4620 2032
rect 2280 1992 4620 2020
rect 2280 1980 2286 1992
rect 4614 1980 4620 1992
rect 4672 1980 4678 2032
rect 6086 1980 6092 2032
rect 6144 2020 6150 2032
rect 10796 2020 10824 2060
rect 10870 2048 10876 2100
rect 10928 2088 10934 2100
rect 14918 2088 14924 2100
rect 10928 2060 14924 2088
rect 10928 2048 10934 2060
rect 14918 2048 14924 2060
rect 14976 2048 14982 2100
rect 11146 2020 11152 2032
rect 6144 1992 9904 2020
rect 10796 1992 11152 2020
rect 6144 1980 6150 1992
rect 3050 1912 3056 1964
rect 3108 1952 3114 1964
rect 5166 1952 5172 1964
rect 3108 1924 5172 1952
rect 3108 1912 3114 1924
rect 5166 1912 5172 1924
rect 5224 1912 5230 1964
rect 6822 1912 6828 1964
rect 6880 1952 6886 1964
rect 6880 1924 9720 1952
rect 6880 1912 6886 1924
rect 2406 1844 2412 1896
rect 2464 1884 2470 1896
rect 2464 1856 9628 1884
rect 2464 1844 2470 1856
rect 2038 1776 2044 1828
rect 2096 1816 2102 1828
rect 9398 1816 9404 1828
rect 2096 1788 9404 1816
rect 2096 1776 2102 1788
rect 9398 1776 9404 1788
rect 9456 1776 9462 1828
rect 4062 1708 4068 1760
rect 4120 1748 4126 1760
rect 8386 1748 8392 1760
rect 4120 1720 8392 1748
rect 4120 1708 4126 1720
rect 8386 1708 8392 1720
rect 8444 1708 8450 1760
rect 9600 1748 9628 1856
rect 9692 1816 9720 1924
rect 9876 1884 9904 1992
rect 11146 1980 11152 1992
rect 11204 1980 11210 2032
rect 12526 1980 12532 2032
rect 12584 2020 12590 2032
rect 16390 2020 16396 2032
rect 12584 1992 16396 2020
rect 12584 1980 12590 1992
rect 16390 1980 16396 1992
rect 16448 1980 16454 2032
rect 12342 1912 12348 1964
rect 12400 1952 12406 1964
rect 18690 1952 18696 1964
rect 12400 1924 18696 1952
rect 12400 1912 12406 1924
rect 18690 1912 18696 1924
rect 18748 1912 18754 1964
rect 17402 1884 17408 1896
rect 9876 1856 17408 1884
rect 17402 1844 17408 1856
rect 17460 1844 17466 1896
rect 16666 1816 16672 1828
rect 9692 1788 16672 1816
rect 16666 1776 16672 1788
rect 16724 1776 16730 1828
rect 12066 1748 12072 1760
rect 9600 1720 12072 1748
rect 12066 1708 12072 1720
rect 12124 1708 12130 1760
rect 12158 1708 12164 1760
rect 12216 1748 12222 1760
rect 18138 1748 18144 1760
rect 12216 1720 18144 1748
rect 12216 1708 12222 1720
rect 18138 1708 18144 1720
rect 18196 1708 18202 1760
rect 7006 1640 7012 1692
rect 7064 1680 7070 1692
rect 12618 1680 12624 1692
rect 7064 1652 12624 1680
rect 7064 1640 7070 1652
rect 12618 1640 12624 1652
rect 12676 1680 12682 1692
rect 15746 1680 15752 1692
rect 12676 1652 15752 1680
rect 12676 1640 12682 1652
rect 15746 1640 15752 1652
rect 15804 1640 15810 1692
rect 2314 1572 2320 1624
rect 2372 1612 2378 1624
rect 2372 1584 2774 1612
rect 2372 1572 2378 1584
rect 2746 1544 2774 1584
rect 3510 1572 3516 1624
rect 3568 1612 3574 1624
rect 7926 1612 7932 1624
rect 3568 1584 7932 1612
rect 3568 1572 3574 1584
rect 7926 1572 7932 1584
rect 7984 1612 7990 1624
rect 12250 1612 12256 1624
rect 7984 1584 12256 1612
rect 7984 1572 7990 1584
rect 12250 1572 12256 1584
rect 12308 1572 12314 1624
rect 12710 1612 12716 1624
rect 12406 1584 12716 1612
rect 7098 1544 7104 1556
rect 2746 1516 7104 1544
rect 7098 1504 7104 1516
rect 7156 1544 7162 1556
rect 12406 1544 12434 1584
rect 12710 1572 12716 1584
rect 12768 1572 12774 1624
rect 7156 1516 12434 1544
rect 7156 1504 7162 1516
rect 11238 1436 11244 1488
rect 11296 1476 11302 1488
rect 12802 1476 12808 1488
rect 11296 1448 12808 1476
rect 11296 1436 11302 1448
rect 12802 1436 12808 1448
rect 12860 1436 12866 1488
rect 4062 1300 4068 1352
rect 4120 1340 4126 1352
rect 10962 1340 10968 1352
rect 4120 1312 10968 1340
rect 4120 1300 4126 1312
rect 10962 1300 10968 1312
rect 11020 1300 11026 1352
rect 11974 1340 11980 1352
rect 11348 1312 11980 1340
rect 3602 1232 3608 1284
rect 3660 1272 3666 1284
rect 11348 1272 11376 1312
rect 11974 1300 11980 1312
rect 12032 1300 12038 1352
rect 13630 1300 13636 1352
rect 13688 1340 13694 1352
rect 15194 1340 15200 1352
rect 13688 1312 15200 1340
rect 13688 1300 13694 1312
rect 15194 1300 15200 1312
rect 15252 1300 15258 1352
rect 3660 1244 11376 1272
rect 3660 1232 3666 1244
rect 11422 1232 11428 1284
rect 11480 1272 11486 1284
rect 15930 1272 15936 1284
rect 11480 1244 15936 1272
rect 11480 1232 11486 1244
rect 15930 1232 15936 1244
rect 15988 1232 15994 1284
rect 11054 1164 11060 1216
rect 11112 1204 11118 1216
rect 15838 1204 15844 1216
rect 11112 1176 15844 1204
rect 11112 1164 11118 1176
rect 15838 1164 15844 1176
rect 15896 1164 15902 1216
rect 3418 824 3424 876
rect 3476 864 3482 876
rect 8846 864 8852 876
rect 3476 836 8852 864
rect 3476 824 3482 836
rect 8846 824 8852 836
rect 8904 824 8910 876
rect 3694 620 3700 672
rect 3752 660 3758 672
rect 6454 660 6460 672
rect 3752 632 6460 660
rect 3752 620 3758 632
rect 6454 620 6460 632
rect 6512 620 6518 672
rect 1578 8 1584 60
rect 1636 48 1642 60
rect 15654 48 15660 60
rect 1636 20 15660 48
rect 1636 8 1642 20
rect 15654 8 15660 20
rect 15712 8 15718 60
<< via1 >>
rect 6552 15784 6604 15836
rect 14832 15784 14884 15836
rect 4252 15648 4304 15700
rect 14556 15648 14608 15700
rect 2688 15580 2740 15632
rect 14648 15580 14700 15632
rect 5264 15512 5316 15564
rect 17960 15512 18012 15564
rect 756 15444 808 15496
rect 8116 15444 8168 15496
rect 13360 15444 13412 15496
rect 13912 15444 13964 15496
rect 20 15376 72 15428
rect 8484 15376 8536 15428
rect 10324 15376 10376 15428
rect 19892 15376 19944 15428
rect 2320 15308 2372 15360
rect 6460 15308 6512 15360
rect 11980 15308 12032 15360
rect 18512 15308 18564 15360
rect 2044 15240 2096 15292
rect 5816 15240 5868 15292
rect 12440 15240 12492 15292
rect 15476 15240 15528 15292
rect 2136 15172 2188 15224
rect 6644 15172 6696 15224
rect 12624 15172 12676 15224
rect 2504 15036 2556 15088
rect 7196 15104 7248 15156
rect 10508 15104 10560 15156
rect 3792 15036 3844 15088
rect 6920 15036 6972 15088
rect 11612 15036 11664 15088
rect 15016 15036 15068 15088
rect 17592 15104 17644 15156
rect 15292 15036 15344 15088
rect 15476 15036 15528 15088
rect 17684 15036 17736 15088
rect 4068 14968 4120 15020
rect 6736 14968 6788 15020
rect 12808 14968 12860 15020
rect 16304 14968 16356 15020
rect 4344 14900 4396 14952
rect 6092 14900 6144 14952
rect 7104 14900 7156 14952
rect 10600 14900 10652 14952
rect 12900 14900 12952 14952
rect 13176 14900 13228 14952
rect 15660 14900 15712 14952
rect 3884 14832 3936 14884
rect 6000 14832 6052 14884
rect 6184 14832 6236 14884
rect 11428 14832 11480 14884
rect 12532 14832 12584 14884
rect 16396 14832 16448 14884
rect 2872 14764 2924 14816
rect 4436 14764 4488 14816
rect 12992 14764 13044 14816
rect 16028 14764 16080 14816
rect 3174 14662 3226 14714
rect 3238 14662 3290 14714
rect 3302 14662 3354 14714
rect 3366 14662 3418 14714
rect 3430 14662 3482 14714
rect 7622 14662 7674 14714
rect 7686 14662 7738 14714
rect 7750 14662 7802 14714
rect 7814 14662 7866 14714
rect 7878 14662 7930 14714
rect 12070 14662 12122 14714
rect 12134 14662 12186 14714
rect 12198 14662 12250 14714
rect 12262 14662 12314 14714
rect 12326 14662 12378 14714
rect 16518 14662 16570 14714
rect 16582 14662 16634 14714
rect 16646 14662 16698 14714
rect 16710 14662 16762 14714
rect 16774 14662 16826 14714
rect 2780 14603 2832 14612
rect 2780 14569 2789 14603
rect 2789 14569 2823 14603
rect 2823 14569 2832 14603
rect 2780 14560 2832 14569
rect 2964 14560 3016 14612
rect 2228 14492 2280 14544
rect 4252 14603 4304 14612
rect 4252 14569 4261 14603
rect 4261 14569 4295 14603
rect 4295 14569 4304 14603
rect 4252 14560 4304 14569
rect 4528 14560 4580 14612
rect 4712 14560 4764 14612
rect 4804 14560 4856 14612
rect 5908 14560 5960 14612
rect 6644 14560 6696 14612
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 11888 14560 11940 14612
rect 11980 14560 12032 14612
rect 12440 14603 12492 14612
rect 12440 14569 12449 14603
rect 12449 14569 12483 14603
rect 12483 14569 12492 14603
rect 12624 14603 12676 14612
rect 12440 14560 12492 14569
rect 12624 14569 12633 14603
rect 12633 14569 12667 14603
rect 12667 14569 12676 14603
rect 12624 14560 12676 14569
rect 12808 14603 12860 14612
rect 12808 14569 12817 14603
rect 12817 14569 12851 14603
rect 12851 14569 12860 14603
rect 12808 14560 12860 14569
rect 12992 14603 13044 14612
rect 12992 14569 13001 14603
rect 13001 14569 13035 14603
rect 13035 14569 13044 14603
rect 12992 14560 13044 14569
rect 13176 14603 13228 14612
rect 13176 14569 13185 14603
rect 13185 14569 13219 14603
rect 13219 14569 13228 14603
rect 13176 14560 13228 14569
rect 1952 14467 2004 14476
rect 1952 14433 1961 14467
rect 1961 14433 1995 14467
rect 1995 14433 2004 14467
rect 1952 14424 2004 14433
rect 2136 14356 2188 14408
rect 2872 14424 2924 14476
rect 3240 14356 3292 14408
rect 3976 14424 4028 14476
rect 3424 14356 3476 14408
rect 3792 14399 3844 14408
rect 3792 14365 3801 14399
rect 3801 14365 3835 14399
rect 3835 14365 3844 14399
rect 3792 14356 3844 14365
rect 4068 14399 4120 14408
rect 4068 14365 4077 14399
rect 4077 14365 4111 14399
rect 4111 14365 4120 14399
rect 4068 14356 4120 14365
rect 4344 14399 4396 14408
rect 4344 14365 4353 14399
rect 4353 14365 4387 14399
rect 4387 14365 4396 14399
rect 4344 14356 4396 14365
rect 4620 14356 4672 14408
rect 5356 14492 5408 14544
rect 6000 14535 6052 14544
rect 6000 14501 6009 14535
rect 6009 14501 6043 14535
rect 6043 14501 6052 14535
rect 6000 14492 6052 14501
rect 6092 14535 6144 14544
rect 6092 14501 6101 14535
rect 6101 14501 6135 14535
rect 6135 14501 6144 14535
rect 6736 14535 6788 14544
rect 6092 14492 6144 14501
rect 6736 14501 6745 14535
rect 6745 14501 6779 14535
rect 6779 14501 6788 14535
rect 6736 14492 6788 14501
rect 6920 14535 6972 14544
rect 6920 14501 6929 14535
rect 6929 14501 6963 14535
rect 6963 14501 6972 14535
rect 6920 14492 6972 14501
rect 7012 14492 7064 14544
rect 11612 14492 11664 14544
rect 11796 14492 11848 14544
rect 14004 14560 14056 14612
rect 17868 14560 17920 14612
rect 6368 14399 6420 14408
rect 6368 14365 6377 14399
rect 6377 14365 6411 14399
rect 6411 14365 6420 14399
rect 6368 14356 6420 14365
rect 13176 14424 13228 14476
rect 9772 14356 9824 14408
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 2596 14220 2648 14272
rect 9680 14288 9732 14340
rect 15016 14492 15068 14544
rect 15108 14535 15160 14544
rect 15108 14501 15117 14535
rect 15117 14501 15151 14535
rect 15151 14501 15160 14535
rect 15108 14492 15160 14501
rect 13912 14424 13964 14476
rect 4620 14220 4672 14272
rect 4896 14220 4948 14272
rect 8576 14220 8628 14272
rect 9036 14220 9088 14272
rect 13820 14331 13872 14340
rect 13820 14297 13829 14331
rect 13829 14297 13863 14331
rect 13863 14297 13872 14331
rect 13820 14288 13872 14297
rect 14096 14288 14148 14340
rect 10416 14220 10468 14272
rect 11980 14263 12032 14272
rect 11980 14229 11989 14263
rect 11989 14229 12023 14263
rect 12023 14229 12032 14263
rect 11980 14220 12032 14229
rect 14556 14399 14608 14408
rect 14556 14365 14565 14399
rect 14565 14365 14599 14399
rect 14599 14365 14608 14399
rect 14556 14356 14608 14365
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 16948 14424 17000 14476
rect 17316 14467 17368 14476
rect 17316 14433 17325 14467
rect 17325 14433 17359 14467
rect 17359 14433 17368 14467
rect 17316 14424 17368 14433
rect 17592 14467 17644 14476
rect 17592 14433 17601 14467
rect 17601 14433 17635 14467
rect 17635 14433 17644 14467
rect 17592 14424 17644 14433
rect 18512 14467 18564 14476
rect 18512 14433 18521 14467
rect 18521 14433 18555 14467
rect 18555 14433 18564 14467
rect 18512 14424 18564 14433
rect 15016 14356 15068 14365
rect 15660 14399 15712 14408
rect 15660 14365 15669 14399
rect 15669 14365 15703 14399
rect 15703 14365 15712 14399
rect 15660 14356 15712 14365
rect 15844 14399 15896 14408
rect 15844 14365 15853 14399
rect 15853 14365 15887 14399
rect 15887 14365 15896 14399
rect 15844 14356 15896 14365
rect 16028 14399 16080 14408
rect 16028 14365 16037 14399
rect 16037 14365 16071 14399
rect 16071 14365 16080 14399
rect 16028 14356 16080 14365
rect 16304 14356 16356 14408
rect 18236 14399 18288 14408
rect 18236 14365 18245 14399
rect 18245 14365 18279 14399
rect 18279 14365 18288 14399
rect 18236 14356 18288 14365
rect 19616 14356 19668 14408
rect 15108 14288 15160 14340
rect 15200 14288 15252 14340
rect 17408 14288 17460 14340
rect 14740 14263 14792 14272
rect 14740 14229 14749 14263
rect 14749 14229 14783 14263
rect 14783 14229 14792 14263
rect 14740 14220 14792 14229
rect 15016 14220 15068 14272
rect 15292 14220 15344 14272
rect 17592 14220 17644 14272
rect 5398 14118 5450 14170
rect 5462 14118 5514 14170
rect 5526 14118 5578 14170
rect 5590 14118 5642 14170
rect 5654 14118 5706 14170
rect 9846 14118 9898 14170
rect 9910 14118 9962 14170
rect 9974 14118 10026 14170
rect 10038 14118 10090 14170
rect 10102 14118 10154 14170
rect 14294 14118 14346 14170
rect 14358 14118 14410 14170
rect 14422 14118 14474 14170
rect 14486 14118 14538 14170
rect 14550 14118 14602 14170
rect 2780 14059 2832 14068
rect 2780 14025 2789 14059
rect 2789 14025 2823 14059
rect 2823 14025 2832 14059
rect 2780 14016 2832 14025
rect 3424 14059 3476 14068
rect 3424 14025 3433 14059
rect 3433 14025 3467 14059
rect 3467 14025 3476 14059
rect 3424 14016 3476 14025
rect 1584 13948 1636 14000
rect 1124 13880 1176 13932
rect 2228 13923 2280 13932
rect 2228 13889 2237 13923
rect 2237 13889 2271 13923
rect 2271 13889 2280 13923
rect 2228 13880 2280 13889
rect 2688 13948 2740 14000
rect 2044 13812 2096 13864
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 3332 13880 3384 13932
rect 4436 14059 4488 14068
rect 4436 14025 4445 14059
rect 4445 14025 4479 14059
rect 4479 14025 4488 14059
rect 4436 14016 4488 14025
rect 4712 14016 4764 14068
rect 4988 14016 5040 14068
rect 5816 14016 5868 14068
rect 6368 14059 6420 14068
rect 6368 14025 6377 14059
rect 6377 14025 6411 14059
rect 6411 14025 6420 14059
rect 6368 14016 6420 14025
rect 6460 14016 6512 14068
rect 5172 13991 5224 14000
rect 5172 13957 5181 13991
rect 5181 13957 5215 13991
rect 5215 13957 5224 13991
rect 5172 13948 5224 13957
rect 5632 13948 5684 14000
rect 5724 13948 5776 14000
rect 7012 14016 7064 14068
rect 7196 14059 7248 14068
rect 7196 14025 7205 14059
rect 7205 14025 7239 14059
rect 7239 14025 7248 14059
rect 7196 14016 7248 14025
rect 8116 14059 8168 14068
rect 8116 14025 8125 14059
rect 8125 14025 8159 14059
rect 8159 14025 8168 14059
rect 8116 14016 8168 14025
rect 9312 14016 9364 14068
rect 9772 14059 9824 14068
rect 6920 13991 6972 14000
rect 6920 13957 6929 13991
rect 6929 13957 6963 13991
rect 6963 13957 6972 13991
rect 6920 13948 6972 13957
rect 7104 13991 7156 14000
rect 7104 13957 7113 13991
rect 7113 13957 7147 13991
rect 7147 13957 7156 13991
rect 7104 13948 7156 13957
rect 9404 13948 9456 14000
rect 9772 14025 9781 14059
rect 9781 14025 9815 14059
rect 9815 14025 9824 14059
rect 9772 14016 9824 14025
rect 10232 13948 10284 14000
rect 3884 13923 3936 13932
rect 3884 13889 3893 13923
rect 3893 13889 3927 13923
rect 3927 13889 3936 13923
rect 3884 13880 3936 13889
rect 4528 13880 4580 13932
rect 4712 13880 4764 13932
rect 5080 13880 5132 13932
rect 6000 13923 6052 13932
rect 4160 13812 4212 13864
rect 6000 13889 6009 13923
rect 6009 13889 6043 13923
rect 6043 13889 6052 13923
rect 6000 13880 6052 13889
rect 6552 13923 6604 13932
rect 6552 13889 6561 13923
rect 6561 13889 6595 13923
rect 6595 13889 6604 13923
rect 6552 13880 6604 13889
rect 6828 13880 6880 13932
rect 9312 13880 9364 13932
rect 9772 13880 9824 13932
rect 13636 14016 13688 14068
rect 13728 14059 13780 14068
rect 13728 14025 13737 14059
rect 13737 14025 13771 14059
rect 13771 14025 13780 14059
rect 13728 14016 13780 14025
rect 13912 14016 13964 14068
rect 14832 14059 14884 14068
rect 14832 14025 14841 14059
rect 14841 14025 14875 14059
rect 14875 14025 14884 14059
rect 14832 14016 14884 14025
rect 14924 14016 14976 14068
rect 8024 13812 8076 13864
rect 9404 13812 9456 13864
rect 4528 13744 4580 13796
rect 8576 13744 8628 13796
rect 12348 13991 12400 14000
rect 12348 13957 12357 13991
rect 12357 13957 12391 13991
rect 12391 13957 12400 13991
rect 12348 13948 12400 13957
rect 12532 13991 12584 14000
rect 12532 13957 12541 13991
rect 12541 13957 12575 13991
rect 12575 13957 12584 13991
rect 12532 13948 12584 13957
rect 12716 13991 12768 14000
rect 12716 13957 12725 13991
rect 12725 13957 12759 13991
rect 12759 13957 12768 13991
rect 12716 13948 12768 13957
rect 12164 13880 12216 13932
rect 13084 13923 13136 13932
rect 13084 13889 13093 13923
rect 13093 13889 13127 13923
rect 13127 13889 13136 13923
rect 13084 13880 13136 13889
rect 13176 13880 13228 13932
rect 13636 13880 13688 13932
rect 10784 13812 10836 13864
rect 11152 13744 11204 13796
rect 12072 13812 12124 13864
rect 13636 13744 13688 13796
rect 14648 13812 14700 13864
rect 14372 13787 14424 13796
rect 14372 13753 14381 13787
rect 14381 13753 14415 13787
rect 14415 13753 14424 13787
rect 14372 13744 14424 13753
rect 15660 14016 15712 14068
rect 19432 14016 19484 14068
rect 15108 13948 15160 14000
rect 15292 13923 15344 13932
rect 15292 13889 15301 13923
rect 15301 13889 15335 13923
rect 15335 13889 15344 13923
rect 15292 13880 15344 13889
rect 15384 13923 15436 13932
rect 15384 13889 15393 13923
rect 15393 13889 15427 13923
rect 15427 13889 15436 13923
rect 15844 13923 15896 13932
rect 15384 13880 15436 13889
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16120 13880 16172 13932
rect 16396 13812 16448 13864
rect 4068 13719 4120 13728
rect 4068 13685 4077 13719
rect 4077 13685 4111 13719
rect 4111 13685 4120 13719
rect 4068 13676 4120 13685
rect 5080 13676 5132 13728
rect 5356 13676 5408 13728
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 5908 13676 5960 13728
rect 6644 13676 6696 13728
rect 6828 13676 6880 13728
rect 11336 13676 11388 13728
rect 11612 13676 11664 13728
rect 11888 13719 11940 13728
rect 11888 13685 11897 13719
rect 11897 13685 11931 13719
rect 11931 13685 11940 13719
rect 11888 13676 11940 13685
rect 13176 13676 13228 13728
rect 14556 13676 14608 13728
rect 14924 13676 14976 13728
rect 15108 13719 15160 13728
rect 15108 13685 15117 13719
rect 15117 13685 15151 13719
rect 15151 13685 15160 13719
rect 15108 13676 15160 13685
rect 19064 13880 19116 13932
rect 17132 13812 17184 13864
rect 17684 13855 17736 13864
rect 17684 13821 17693 13855
rect 17693 13821 17727 13855
rect 17727 13821 17736 13855
rect 17684 13812 17736 13821
rect 18604 13812 18656 13864
rect 17040 13676 17092 13728
rect 3174 13574 3226 13626
rect 3238 13574 3290 13626
rect 3302 13574 3354 13626
rect 3366 13574 3418 13626
rect 3430 13574 3482 13626
rect 7622 13574 7674 13626
rect 7686 13574 7738 13626
rect 7750 13574 7802 13626
rect 7814 13574 7866 13626
rect 7878 13574 7930 13626
rect 12070 13574 12122 13626
rect 12134 13574 12186 13626
rect 12198 13574 12250 13626
rect 12262 13574 12314 13626
rect 12326 13574 12378 13626
rect 16518 13574 16570 13626
rect 16582 13574 16634 13626
rect 16646 13574 16698 13626
rect 16710 13574 16762 13626
rect 16774 13574 16826 13626
rect 848 13472 900 13524
rect 1216 13404 1268 13456
rect 2504 13336 2556 13388
rect 4252 13472 4304 13524
rect 5356 13472 5408 13524
rect 6644 13515 6696 13524
rect 6644 13481 6653 13515
rect 6653 13481 6687 13515
rect 6687 13481 6696 13515
rect 6644 13472 6696 13481
rect 7288 13472 7340 13524
rect 8024 13515 8076 13524
rect 8024 13481 8033 13515
rect 8033 13481 8067 13515
rect 8067 13481 8076 13515
rect 8024 13472 8076 13481
rect 8300 13515 8352 13524
rect 8300 13481 8309 13515
rect 8309 13481 8343 13515
rect 8343 13481 8352 13515
rect 8300 13472 8352 13481
rect 8576 13515 8628 13524
rect 8576 13481 8585 13515
rect 8585 13481 8619 13515
rect 8619 13481 8628 13515
rect 8576 13472 8628 13481
rect 9036 13515 9088 13524
rect 9036 13481 9045 13515
rect 9045 13481 9079 13515
rect 9079 13481 9088 13515
rect 9036 13472 9088 13481
rect 10416 13472 10468 13524
rect 10876 13472 10928 13524
rect 11428 13515 11480 13524
rect 11428 13481 11437 13515
rect 11437 13481 11471 13515
rect 11471 13481 11480 13515
rect 11428 13472 11480 13481
rect 11612 13472 11664 13524
rect 12808 13515 12860 13524
rect 4804 13404 4856 13456
rect 12808 13481 12817 13515
rect 12817 13481 12851 13515
rect 12851 13481 12860 13515
rect 12808 13472 12860 13481
rect 13544 13472 13596 13524
rect 15660 13472 15712 13524
rect 16120 13515 16172 13524
rect 16120 13481 16129 13515
rect 16129 13481 16163 13515
rect 16163 13481 16172 13515
rect 16120 13472 16172 13481
rect 16212 13472 16264 13524
rect 2136 13268 2188 13320
rect 2596 13311 2648 13320
rect 2596 13277 2605 13311
rect 2605 13277 2639 13311
rect 2639 13277 2648 13311
rect 2596 13268 2648 13277
rect 3332 13311 3384 13320
rect 3332 13277 3341 13311
rect 3341 13277 3375 13311
rect 3375 13277 3384 13311
rect 3332 13268 3384 13277
rect 3424 13311 3476 13320
rect 3424 13277 3433 13311
rect 3433 13277 3467 13311
rect 3467 13277 3476 13311
rect 3424 13268 3476 13277
rect 3884 13268 3936 13320
rect 4068 13311 4120 13320
rect 4068 13277 4077 13311
rect 4077 13277 4111 13311
rect 4111 13277 4120 13311
rect 5540 13336 5592 13388
rect 5632 13336 5684 13388
rect 6736 13336 6788 13388
rect 7196 13379 7248 13388
rect 7196 13345 7205 13379
rect 7205 13345 7239 13379
rect 7239 13345 7248 13379
rect 7196 13336 7248 13345
rect 8300 13336 8352 13388
rect 11520 13379 11572 13388
rect 11520 13345 11529 13379
rect 11529 13345 11563 13379
rect 11563 13345 11572 13379
rect 11520 13336 11572 13345
rect 12072 13404 12124 13456
rect 13084 13404 13136 13456
rect 13820 13404 13872 13456
rect 14924 13404 14976 13456
rect 15568 13404 15620 13456
rect 12348 13336 12400 13388
rect 12532 13336 12584 13388
rect 12992 13379 13044 13388
rect 12992 13345 13001 13379
rect 13001 13345 13035 13379
rect 13035 13345 13044 13379
rect 12992 13336 13044 13345
rect 14280 13336 14332 13388
rect 4068 13268 4120 13277
rect 4620 13268 4672 13320
rect 4804 13311 4856 13320
rect 4804 13277 4813 13311
rect 4813 13277 4847 13311
rect 4847 13277 4856 13311
rect 4804 13268 4856 13277
rect 4896 13311 4948 13320
rect 4896 13277 4905 13311
rect 4905 13277 4939 13311
rect 4939 13277 4948 13311
rect 4896 13268 4948 13277
rect 5080 13268 5132 13320
rect 5264 13268 5316 13320
rect 5816 13268 5868 13320
rect 10232 13268 10284 13320
rect 11060 13311 11112 13320
rect 11060 13277 11069 13311
rect 11069 13277 11103 13311
rect 11103 13277 11112 13311
rect 11060 13268 11112 13277
rect 12072 13268 12124 13320
rect 12440 13268 12492 13320
rect 12900 13268 12952 13320
rect 1308 13200 1360 13252
rect 2412 13175 2464 13184
rect 2412 13141 2421 13175
rect 2421 13141 2455 13175
rect 2455 13141 2464 13175
rect 2412 13132 2464 13141
rect 2780 13175 2832 13184
rect 2780 13141 2789 13175
rect 2789 13141 2823 13175
rect 2823 13141 2832 13175
rect 3792 13200 3844 13252
rect 6552 13200 6604 13252
rect 7288 13200 7340 13252
rect 10692 13200 10744 13252
rect 10968 13200 11020 13252
rect 11152 13243 11204 13252
rect 11152 13209 11161 13243
rect 11161 13209 11195 13243
rect 11195 13209 11204 13243
rect 11152 13200 11204 13209
rect 11244 13200 11296 13252
rect 12532 13243 12584 13252
rect 2780 13132 2832 13141
rect 3700 13132 3752 13184
rect 4068 13132 4120 13184
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 4436 13132 4488 13184
rect 5264 13132 5316 13184
rect 5908 13175 5960 13184
rect 5908 13141 5917 13175
rect 5917 13141 5951 13175
rect 5951 13141 5960 13175
rect 5908 13132 5960 13141
rect 6184 13175 6236 13184
rect 6184 13141 6193 13175
rect 6193 13141 6227 13175
rect 6227 13141 6236 13175
rect 6184 13132 6236 13141
rect 6920 13175 6972 13184
rect 6920 13141 6929 13175
rect 6929 13141 6963 13175
rect 6963 13141 6972 13175
rect 6920 13132 6972 13141
rect 7380 13175 7432 13184
rect 7380 13141 7389 13175
rect 7389 13141 7423 13175
rect 7423 13141 7432 13175
rect 7380 13132 7432 13141
rect 7472 13132 7524 13184
rect 7748 13175 7800 13184
rect 7748 13141 7757 13175
rect 7757 13141 7791 13175
rect 7791 13141 7800 13175
rect 7748 13132 7800 13141
rect 8024 13132 8076 13184
rect 10600 13175 10652 13184
rect 10600 13141 10609 13175
rect 10609 13141 10643 13175
rect 10643 13141 10652 13175
rect 10600 13132 10652 13141
rect 12072 13175 12124 13184
rect 12072 13141 12081 13175
rect 12081 13141 12115 13175
rect 12115 13141 12124 13175
rect 12072 13132 12124 13141
rect 12532 13209 12541 13243
rect 12541 13209 12575 13243
rect 12575 13209 12584 13243
rect 12532 13200 12584 13209
rect 13636 13268 13688 13320
rect 14188 13268 14240 13320
rect 15200 13336 15252 13388
rect 16856 13336 16908 13388
rect 17868 13336 17920 13388
rect 15384 13311 15436 13320
rect 15384 13277 15393 13311
rect 15393 13277 15427 13311
rect 15427 13277 15436 13311
rect 15384 13268 15436 13277
rect 15476 13268 15528 13320
rect 14924 13200 14976 13252
rect 16396 13200 16448 13252
rect 18052 13268 18104 13320
rect 17776 13200 17828 13252
rect 13452 13132 13504 13184
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 14004 13132 14056 13184
rect 14188 13132 14240 13184
rect 15384 13132 15436 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 15752 13132 15804 13184
rect 19156 13132 19208 13184
rect 5398 13030 5450 13082
rect 5462 13030 5514 13082
rect 5526 13030 5578 13082
rect 5590 13030 5642 13082
rect 5654 13030 5706 13082
rect 9846 13030 9898 13082
rect 9910 13030 9962 13082
rect 9974 13030 10026 13082
rect 10038 13030 10090 13082
rect 10102 13030 10154 13082
rect 14294 13030 14346 13082
rect 14358 13030 14410 13082
rect 14422 13030 14474 13082
rect 14486 13030 14538 13082
rect 14550 13030 14602 13082
rect 2320 12928 2372 12980
rect 4344 12971 4396 12980
rect 1768 12860 1820 12912
rect 4344 12937 4353 12971
rect 4353 12937 4387 12971
rect 4387 12937 4396 12971
rect 4344 12928 4396 12937
rect 5816 12971 5868 12980
rect 5816 12937 5825 12971
rect 5825 12937 5859 12971
rect 5859 12937 5868 12971
rect 5816 12928 5868 12937
rect 6552 12928 6604 12980
rect 6920 12928 6972 12980
rect 9496 12971 9548 12980
rect 9496 12937 9505 12971
rect 9505 12937 9539 12971
rect 9539 12937 9548 12971
rect 9496 12928 9548 12937
rect 10324 12928 10376 12980
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10692 12928 10744 12980
rect 11428 12928 11480 12980
rect 3056 12792 3108 12844
rect 3700 12792 3752 12844
rect 4252 12792 4304 12844
rect 6092 12860 6144 12912
rect 7288 12860 7340 12912
rect 8116 12903 8168 12912
rect 8116 12869 8125 12903
rect 8125 12869 8159 12903
rect 8159 12869 8168 12903
rect 8116 12860 8168 12869
rect 8300 12903 8352 12912
rect 8300 12869 8309 12903
rect 8309 12869 8343 12903
rect 8343 12869 8352 12903
rect 8300 12860 8352 12869
rect 8760 12903 8812 12912
rect 8760 12869 8769 12903
rect 8769 12869 8803 12903
rect 8803 12869 8812 12903
rect 9036 12903 9088 12912
rect 8760 12860 8812 12869
rect 9036 12869 9045 12903
rect 9045 12869 9079 12903
rect 9079 12869 9088 12903
rect 9036 12860 9088 12869
rect 9588 12860 9640 12912
rect 12164 12860 12216 12912
rect 12716 12928 12768 12980
rect 13176 12971 13228 12980
rect 13176 12937 13185 12971
rect 13185 12937 13219 12971
rect 13219 12937 13228 12971
rect 13176 12928 13228 12937
rect 13820 12971 13872 12980
rect 13820 12937 13829 12971
rect 13829 12937 13863 12971
rect 13863 12937 13872 12971
rect 13820 12928 13872 12937
rect 14096 12928 14148 12980
rect 4988 12835 5040 12844
rect 4988 12801 4997 12835
rect 4997 12801 5031 12835
rect 5031 12801 5040 12835
rect 4988 12792 5040 12801
rect 5172 12792 5224 12844
rect 5356 12835 5408 12844
rect 5356 12801 5365 12835
rect 5365 12801 5399 12835
rect 5399 12801 5408 12835
rect 5356 12792 5408 12801
rect 1492 12724 1544 12776
rect 2780 12724 2832 12776
rect 2964 12724 3016 12776
rect 3240 12724 3292 12776
rect 3608 12699 3660 12708
rect 3608 12665 3617 12699
rect 3617 12665 3651 12699
rect 3651 12665 3660 12699
rect 3608 12656 3660 12665
rect 2964 12588 3016 12640
rect 4068 12588 4120 12640
rect 4344 12656 4396 12708
rect 6276 12792 6328 12844
rect 6736 12792 6788 12844
rect 8392 12792 8444 12844
rect 6460 12724 6512 12776
rect 7196 12767 7248 12776
rect 7196 12733 7205 12767
rect 7205 12733 7239 12767
rect 7239 12733 7248 12767
rect 7196 12724 7248 12733
rect 8116 12724 8168 12776
rect 8852 12792 8904 12844
rect 9404 12792 9456 12844
rect 10692 12792 10744 12844
rect 9956 12724 10008 12776
rect 10600 12724 10652 12776
rect 5172 12656 5224 12708
rect 6276 12656 6328 12708
rect 6828 12656 6880 12708
rect 6920 12699 6972 12708
rect 6920 12665 6929 12699
rect 6929 12665 6963 12699
rect 6963 12665 6972 12699
rect 6920 12656 6972 12665
rect 5908 12588 5960 12640
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 7012 12631 7064 12640
rect 7012 12597 7021 12631
rect 7021 12597 7055 12631
rect 7055 12597 7064 12631
rect 7012 12588 7064 12597
rect 10876 12699 10928 12708
rect 8484 12631 8536 12640
rect 8484 12597 8493 12631
rect 8493 12597 8527 12631
rect 8527 12597 8536 12631
rect 8484 12588 8536 12597
rect 10876 12665 10885 12699
rect 10885 12665 10919 12699
rect 10919 12665 10928 12699
rect 11980 12792 12032 12844
rect 11520 12724 11572 12776
rect 12164 12767 12216 12776
rect 10876 12656 10928 12665
rect 11612 12656 11664 12708
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 12348 12792 12400 12844
rect 12808 12792 12860 12844
rect 13084 12792 13136 12844
rect 13544 12835 13596 12844
rect 13544 12801 13553 12835
rect 13553 12801 13587 12835
rect 13587 12801 13596 12835
rect 13544 12792 13596 12801
rect 14096 12792 14148 12844
rect 15844 12928 15896 12980
rect 14556 12792 14608 12844
rect 12532 12656 12584 12708
rect 13360 12724 13412 12776
rect 14740 12835 14792 12844
rect 14740 12801 14749 12835
rect 14749 12801 14783 12835
rect 14783 12801 14792 12835
rect 14740 12792 14792 12801
rect 15476 12792 15528 12844
rect 15660 12835 15712 12844
rect 15660 12801 15669 12835
rect 15669 12801 15703 12835
rect 15703 12801 15712 12835
rect 15660 12792 15712 12801
rect 16028 12835 16080 12844
rect 16028 12801 16037 12835
rect 16037 12801 16071 12835
rect 16071 12801 16080 12835
rect 16028 12792 16080 12801
rect 16488 12792 16540 12844
rect 12992 12656 13044 12708
rect 11520 12588 11572 12640
rect 14188 12656 14240 12708
rect 14280 12656 14332 12708
rect 13268 12631 13320 12640
rect 13268 12597 13277 12631
rect 13277 12597 13311 12631
rect 13311 12597 13320 12631
rect 13268 12588 13320 12597
rect 13636 12588 13688 12640
rect 14096 12631 14148 12640
rect 14096 12597 14105 12631
rect 14105 12597 14139 12631
rect 14139 12597 14148 12631
rect 14096 12588 14148 12597
rect 18236 12724 18288 12776
rect 15384 12656 15436 12708
rect 16212 12699 16264 12708
rect 16212 12665 16221 12699
rect 16221 12665 16255 12699
rect 16255 12665 16264 12699
rect 16212 12656 16264 12665
rect 18144 12656 18196 12708
rect 15200 12631 15252 12640
rect 15200 12597 15209 12631
rect 15209 12597 15243 12631
rect 15243 12597 15252 12631
rect 15200 12588 15252 12597
rect 16396 12588 16448 12640
rect 3174 12486 3226 12538
rect 3238 12486 3290 12538
rect 3302 12486 3354 12538
rect 3366 12486 3418 12538
rect 3430 12486 3482 12538
rect 7622 12486 7674 12538
rect 7686 12486 7738 12538
rect 7750 12486 7802 12538
rect 7814 12486 7866 12538
rect 7878 12486 7930 12538
rect 12070 12486 12122 12538
rect 12134 12486 12186 12538
rect 12198 12486 12250 12538
rect 12262 12486 12314 12538
rect 12326 12486 12378 12538
rect 16518 12486 16570 12538
rect 16582 12486 16634 12538
rect 16646 12486 16698 12538
rect 16710 12486 16762 12538
rect 16774 12486 16826 12538
rect 2780 12384 2832 12436
rect 7472 12384 7524 12436
rect 8576 12384 8628 12436
rect 2412 12291 2464 12300
rect 2412 12257 2421 12291
rect 2421 12257 2455 12291
rect 2455 12257 2464 12291
rect 2412 12248 2464 12257
rect 1952 12223 2004 12232
rect 1952 12189 1961 12223
rect 1961 12189 1995 12223
rect 1995 12189 2004 12223
rect 1952 12180 2004 12189
rect 2872 12316 2924 12368
rect 6736 12316 6788 12368
rect 6920 12316 6972 12368
rect 7196 12316 7248 12368
rect 3424 12291 3476 12300
rect 3424 12257 3433 12291
rect 3433 12257 3467 12291
rect 3467 12257 3476 12291
rect 3424 12248 3476 12257
rect 2964 12180 3016 12232
rect 4528 12248 4580 12300
rect 4620 12291 4672 12300
rect 4620 12257 4629 12291
rect 4629 12257 4663 12291
rect 4663 12257 4672 12291
rect 4620 12248 4672 12257
rect 5816 12248 5868 12300
rect 5908 12248 5960 12300
rect 6644 12248 6696 12300
rect 9588 12384 9640 12436
rect 9680 12384 9732 12436
rect 10140 12427 10192 12436
rect 10140 12393 10149 12427
rect 10149 12393 10183 12427
rect 10183 12393 10192 12427
rect 10140 12384 10192 12393
rect 10232 12384 10284 12436
rect 9404 12316 9456 12368
rect 10048 12316 10100 12368
rect 10416 12316 10468 12368
rect 10600 12316 10652 12368
rect 11244 12384 11296 12436
rect 11336 12384 11388 12436
rect 11796 12384 11848 12436
rect 11704 12316 11756 12368
rect 11888 12359 11940 12368
rect 11888 12325 11897 12359
rect 11897 12325 11931 12359
rect 11931 12325 11940 12359
rect 11888 12316 11940 12325
rect 14464 12384 14516 12436
rect 14924 12384 14976 12436
rect 7656 12248 7708 12300
rect 11060 12248 11112 12300
rect 11244 12248 11296 12300
rect 12440 12316 12492 12368
rect 13728 12316 13780 12368
rect 2504 12112 2556 12164
rect 2596 12087 2648 12096
rect 2596 12053 2605 12087
rect 2605 12053 2639 12087
rect 2639 12053 2648 12087
rect 2596 12044 2648 12053
rect 2688 12087 2740 12096
rect 2688 12053 2697 12087
rect 2697 12053 2731 12087
rect 2731 12053 2740 12087
rect 2688 12044 2740 12053
rect 3148 12044 3200 12096
rect 3332 12112 3384 12164
rect 4068 12112 4120 12164
rect 4804 12180 4856 12232
rect 5448 12223 5500 12232
rect 5448 12189 5457 12223
rect 5457 12189 5491 12223
rect 5491 12189 5500 12223
rect 5448 12180 5500 12189
rect 6000 12112 6052 12164
rect 6368 12180 6420 12232
rect 7288 12180 7340 12232
rect 7472 12223 7524 12232
rect 7472 12189 7481 12223
rect 7481 12189 7515 12223
rect 7515 12189 7524 12223
rect 7472 12180 7524 12189
rect 8300 12180 8352 12232
rect 8116 12155 8168 12164
rect 8116 12121 8125 12155
rect 8125 12121 8159 12155
rect 8159 12121 8168 12155
rect 8116 12112 8168 12121
rect 10968 12180 11020 12232
rect 12992 12248 13044 12300
rect 14832 12291 14884 12300
rect 11796 12180 11848 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 12900 12223 12952 12232
rect 12900 12189 12909 12223
rect 12909 12189 12943 12223
rect 12943 12189 12952 12223
rect 13176 12223 13228 12232
rect 12900 12180 12952 12189
rect 13176 12189 13185 12223
rect 13185 12189 13219 12223
rect 13219 12189 13228 12223
rect 13176 12180 13228 12189
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 4252 12087 4304 12096
rect 4252 12053 4261 12087
rect 4261 12053 4295 12087
rect 4295 12053 4304 12087
rect 4252 12044 4304 12053
rect 5816 12044 5868 12096
rect 6092 12087 6144 12096
rect 6092 12053 6101 12087
rect 6101 12053 6135 12087
rect 6135 12053 6144 12087
rect 6092 12044 6144 12053
rect 6184 12044 6236 12096
rect 6552 12044 6604 12096
rect 7104 12087 7156 12096
rect 7104 12053 7113 12087
rect 7113 12053 7147 12087
rect 7147 12053 7156 12087
rect 7104 12044 7156 12053
rect 7564 12044 7616 12096
rect 7748 12044 7800 12096
rect 10140 12112 10192 12164
rect 10692 12112 10744 12164
rect 11244 12112 11296 12164
rect 13728 12180 13780 12232
rect 14188 12180 14240 12232
rect 14832 12257 14841 12291
rect 14841 12257 14875 12291
rect 14875 12257 14884 12291
rect 14832 12248 14884 12257
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 9220 12044 9272 12096
rect 9496 12087 9548 12096
rect 9496 12053 9505 12087
rect 9505 12053 9539 12087
rect 9539 12053 9548 12087
rect 9496 12044 9548 12053
rect 9588 12044 9640 12096
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 10324 12044 10376 12053
rect 10416 12044 10468 12096
rect 11152 12044 11204 12096
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 11980 12087 12032 12096
rect 11980 12053 11989 12087
rect 11989 12053 12023 12087
rect 12023 12053 12032 12087
rect 11980 12044 12032 12053
rect 12164 12087 12216 12096
rect 12164 12053 12173 12087
rect 12173 12053 12207 12087
rect 12207 12053 12216 12087
rect 12164 12044 12216 12053
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 12532 12044 12584 12096
rect 13084 12087 13136 12096
rect 13084 12053 13093 12087
rect 13093 12053 13127 12087
rect 13127 12053 13136 12087
rect 13084 12044 13136 12053
rect 16212 12112 16264 12164
rect 16948 12384 17000 12436
rect 18972 12384 19024 12436
rect 18880 12316 18932 12368
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 17960 12291 18012 12300
rect 17960 12257 17969 12291
rect 17969 12257 18003 12291
rect 18003 12257 18012 12291
rect 17960 12248 18012 12257
rect 18052 12248 18104 12300
rect 18420 12248 18472 12300
rect 17224 12155 17276 12164
rect 17224 12121 17233 12155
rect 17233 12121 17267 12155
rect 17267 12121 17276 12155
rect 17224 12112 17276 12121
rect 17500 12180 17552 12232
rect 18052 12112 18104 12164
rect 13820 12087 13872 12096
rect 13820 12053 13829 12087
rect 13829 12053 13863 12087
rect 13863 12053 13872 12087
rect 13820 12044 13872 12053
rect 14924 12044 14976 12096
rect 15016 12044 15068 12096
rect 15292 12044 15344 12096
rect 15752 12087 15804 12096
rect 15752 12053 15761 12087
rect 15761 12053 15795 12087
rect 15795 12053 15804 12087
rect 15752 12044 15804 12053
rect 15936 12044 15988 12096
rect 16120 12044 16172 12096
rect 18328 12044 18380 12096
rect 5398 11942 5450 11994
rect 5462 11942 5514 11994
rect 5526 11942 5578 11994
rect 5590 11942 5642 11994
rect 5654 11942 5706 11994
rect 9846 11942 9898 11994
rect 9910 11942 9962 11994
rect 9974 11942 10026 11994
rect 10038 11942 10090 11994
rect 10102 11942 10154 11994
rect 14294 11942 14346 11994
rect 14358 11942 14410 11994
rect 14422 11942 14474 11994
rect 14486 11942 14538 11994
rect 14550 11942 14602 11994
rect 2596 11840 2648 11892
rect 2044 11772 2096 11824
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 3148 11772 3200 11824
rect 5908 11772 5960 11824
rect 3792 11704 3844 11756
rect 5724 11704 5776 11756
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 1124 11636 1176 11688
rect 2136 11636 2188 11688
rect 3056 11636 3108 11688
rect 2044 11568 2096 11620
rect 3976 11636 4028 11688
rect 1400 11500 1452 11552
rect 2596 11500 2648 11552
rect 4344 11636 4396 11688
rect 5356 11636 5408 11688
rect 6276 11772 6328 11824
rect 7012 11772 7064 11824
rect 7748 11815 7800 11824
rect 7748 11781 7757 11815
rect 7757 11781 7791 11815
rect 7791 11781 7800 11815
rect 7748 11772 7800 11781
rect 8024 11772 8076 11824
rect 6184 11704 6236 11756
rect 6460 11704 6512 11756
rect 6736 11704 6788 11756
rect 7656 11747 7708 11756
rect 6276 11636 6328 11688
rect 4160 11500 4212 11552
rect 4620 11500 4672 11552
rect 4896 11543 4948 11552
rect 4896 11509 4905 11543
rect 4905 11509 4939 11543
rect 4939 11509 4948 11543
rect 4896 11500 4948 11509
rect 5264 11500 5316 11552
rect 5908 11500 5960 11552
rect 6184 11500 6236 11552
rect 6460 11543 6512 11552
rect 6460 11509 6469 11543
rect 6469 11509 6503 11543
rect 6503 11509 6512 11543
rect 6460 11500 6512 11509
rect 6828 11568 6880 11620
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 9128 11772 9180 11824
rect 8852 11704 8904 11756
rect 7288 11636 7340 11688
rect 8024 11636 8076 11688
rect 8392 11679 8444 11688
rect 8392 11645 8401 11679
rect 8401 11645 8435 11679
rect 8435 11645 8444 11679
rect 8392 11636 8444 11645
rect 7932 11568 7984 11620
rect 10232 11704 10284 11756
rect 10416 11772 10468 11824
rect 11520 11840 11572 11892
rect 11980 11840 12032 11892
rect 12900 11772 12952 11824
rect 11060 11704 11112 11756
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 12532 11747 12584 11756
rect 12532 11713 12541 11747
rect 12541 11713 12575 11747
rect 12575 11713 12584 11747
rect 12532 11704 12584 11713
rect 13636 11704 13688 11756
rect 14004 11772 14056 11824
rect 14096 11713 14117 11740
rect 14117 11713 14148 11740
rect 14096 11688 14148 11713
rect 14924 11840 14976 11892
rect 15292 11840 15344 11892
rect 16120 11840 16172 11892
rect 16212 11840 16264 11892
rect 14556 11772 14608 11824
rect 15108 11772 15160 11824
rect 15752 11772 15804 11824
rect 19248 11772 19300 11824
rect 14648 11704 14700 11756
rect 14924 11747 14976 11756
rect 14924 11713 14933 11747
rect 14933 11713 14967 11747
rect 14967 11713 14976 11747
rect 14924 11704 14976 11713
rect 16304 11747 16356 11756
rect 16304 11713 16313 11747
rect 16313 11713 16347 11747
rect 16347 11713 16356 11747
rect 16304 11704 16356 11713
rect 11336 11636 11388 11688
rect 11520 11679 11572 11688
rect 11520 11645 11529 11679
rect 11529 11645 11563 11679
rect 11563 11645 11572 11679
rect 11520 11636 11572 11645
rect 12808 11611 12860 11620
rect 12808 11577 12817 11611
rect 12817 11577 12851 11611
rect 12851 11577 12860 11611
rect 12808 11568 12860 11577
rect 13084 11611 13136 11620
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 16120 11636 16172 11688
rect 18328 11704 18380 11756
rect 17684 11636 17736 11688
rect 17960 11679 18012 11688
rect 17960 11645 17969 11679
rect 17969 11645 18003 11679
rect 18003 11645 18012 11679
rect 17960 11636 18012 11645
rect 7288 11543 7340 11552
rect 7288 11509 7297 11543
rect 7297 11509 7331 11543
rect 7331 11509 7340 11543
rect 7288 11500 7340 11509
rect 9036 11500 9088 11552
rect 9404 11543 9456 11552
rect 9404 11509 9413 11543
rect 9413 11509 9447 11543
rect 9447 11509 9456 11543
rect 9404 11500 9456 11509
rect 10232 11500 10284 11552
rect 11888 11500 11940 11552
rect 12716 11543 12768 11552
rect 12716 11509 12725 11543
rect 12725 11509 12759 11543
rect 12759 11509 12768 11543
rect 12716 11500 12768 11509
rect 13636 11500 13688 11552
rect 13820 11500 13872 11552
rect 14372 11543 14424 11552
rect 14372 11509 14381 11543
rect 14381 11509 14415 11543
rect 14415 11509 14424 11543
rect 14372 11500 14424 11509
rect 14648 11543 14700 11552
rect 14648 11509 14657 11543
rect 14657 11509 14691 11543
rect 14691 11509 14700 11543
rect 14648 11500 14700 11509
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 15660 11543 15712 11552
rect 15660 11509 15669 11543
rect 15669 11509 15703 11543
rect 15703 11509 15712 11543
rect 15660 11500 15712 11509
rect 16028 11500 16080 11552
rect 17132 11500 17184 11552
rect 3174 11398 3226 11450
rect 3238 11398 3290 11450
rect 3302 11398 3354 11450
rect 3366 11398 3418 11450
rect 3430 11398 3482 11450
rect 7622 11398 7674 11450
rect 7686 11398 7738 11450
rect 7750 11398 7802 11450
rect 7814 11398 7866 11450
rect 7878 11398 7930 11450
rect 12070 11398 12122 11450
rect 12134 11398 12186 11450
rect 12198 11398 12250 11450
rect 12262 11398 12314 11450
rect 12326 11398 12378 11450
rect 16518 11398 16570 11450
rect 16582 11398 16634 11450
rect 16646 11398 16698 11450
rect 16710 11398 16762 11450
rect 16774 11398 16826 11450
rect 2688 11296 2740 11348
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 2044 11228 2096 11280
rect 2412 11228 2464 11280
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 3792 11160 3844 11212
rect 4160 11160 4212 11212
rect 4436 11203 4488 11212
rect 4436 11169 4445 11203
rect 4445 11169 4479 11203
rect 4479 11169 4488 11203
rect 4436 11160 4488 11169
rect 4528 11160 4580 11212
rect 1768 11135 1820 11144
rect 1768 11101 1777 11135
rect 1777 11101 1811 11135
rect 1811 11101 1820 11135
rect 1768 11092 1820 11101
rect 2872 11092 2924 11144
rect 2136 11024 2188 11076
rect 4436 11024 4488 11076
rect 5080 11024 5132 11076
rect 2504 10956 2556 11008
rect 3148 10956 3200 11008
rect 9312 11296 9364 11348
rect 8944 11228 8996 11280
rect 8024 11160 8076 11212
rect 10416 11160 10468 11212
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 8392 11092 8444 11144
rect 8484 11092 8536 11144
rect 8944 11092 8996 11144
rect 12808 11296 12860 11348
rect 13636 11296 13688 11348
rect 10692 11228 10744 11280
rect 13176 11228 13228 11280
rect 10968 11160 11020 11212
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 12256 11160 12308 11212
rect 14004 11296 14056 11348
rect 15016 11296 15068 11348
rect 15844 11296 15896 11348
rect 16304 11296 16356 11348
rect 11520 11092 11572 11144
rect 12440 11092 12492 11144
rect 12900 11135 12952 11144
rect 6184 11024 6236 11076
rect 6644 11024 6696 11076
rect 8116 11024 8168 11076
rect 9680 11024 9732 11076
rect 10232 11024 10284 11076
rect 11060 11024 11112 11076
rect 6828 10956 6880 11008
rect 7472 10999 7524 11008
rect 7472 10965 7481 10999
rect 7481 10965 7515 10999
rect 7515 10965 7524 10999
rect 7472 10956 7524 10965
rect 7564 10999 7616 11008
rect 7564 10965 7573 10999
rect 7573 10965 7607 10999
rect 7607 10965 7616 10999
rect 8392 10999 8444 11008
rect 7564 10956 7616 10965
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 8576 10999 8628 11008
rect 8576 10965 8585 10999
rect 8585 10965 8619 10999
rect 8619 10965 8628 10999
rect 8576 10956 8628 10965
rect 8852 10956 8904 11008
rect 10600 10956 10652 11008
rect 10784 10999 10836 11008
rect 10784 10965 10793 10999
rect 10793 10965 10827 10999
rect 10827 10965 10836 10999
rect 10784 10956 10836 10965
rect 12900 11101 12909 11135
rect 12909 11101 12943 11135
rect 12943 11101 12952 11135
rect 12900 11092 12952 11101
rect 13084 11092 13136 11144
rect 13452 11092 13504 11144
rect 16212 11092 16264 11144
rect 12164 10956 12216 11008
rect 12992 11024 13044 11076
rect 13544 11067 13596 11076
rect 13544 11033 13553 11067
rect 13553 11033 13587 11067
rect 13587 11033 13596 11067
rect 13544 11024 13596 11033
rect 14004 11024 14056 11076
rect 14556 11024 14608 11076
rect 15016 11024 15068 11076
rect 15660 11024 15712 11076
rect 12624 10956 12676 11008
rect 15384 10956 15436 11008
rect 17684 10956 17736 11008
rect 17960 10956 18012 11008
rect 5398 10854 5450 10906
rect 5462 10854 5514 10906
rect 5526 10854 5578 10906
rect 5590 10854 5642 10906
rect 5654 10854 5706 10906
rect 9846 10854 9898 10906
rect 9910 10854 9962 10906
rect 9974 10854 10026 10906
rect 10038 10854 10090 10906
rect 10102 10854 10154 10906
rect 14294 10854 14346 10906
rect 14358 10854 14410 10906
rect 14422 10854 14474 10906
rect 14486 10854 14538 10906
rect 14550 10854 14602 10906
rect 1400 10795 1452 10804
rect 1400 10761 1409 10795
rect 1409 10761 1443 10795
rect 1443 10761 1452 10795
rect 1400 10752 1452 10761
rect 1584 10752 1636 10804
rect 2044 10752 2096 10804
rect 3792 10752 3844 10804
rect 4528 10752 4580 10804
rect 6184 10795 6236 10804
rect 6184 10761 6193 10795
rect 6193 10761 6227 10795
rect 6227 10761 6236 10795
rect 6184 10752 6236 10761
rect 7288 10795 7340 10804
rect 7288 10761 7297 10795
rect 7297 10761 7331 10795
rect 7331 10761 7340 10795
rect 7288 10752 7340 10761
rect 9496 10752 9548 10804
rect 2412 10684 2464 10736
rect 2964 10727 3016 10736
rect 2964 10693 2973 10727
rect 2973 10693 3007 10727
rect 3007 10693 3016 10727
rect 2964 10684 3016 10693
rect 2872 10548 2924 10600
rect 4988 10684 5040 10736
rect 5908 10684 5960 10736
rect 7564 10684 7616 10736
rect 10784 10752 10836 10804
rect 12716 10752 12768 10804
rect 12992 10752 13044 10804
rect 14188 10752 14240 10804
rect 18144 10752 18196 10804
rect 10692 10727 10744 10736
rect 10692 10693 10701 10727
rect 10701 10693 10735 10727
rect 10735 10693 10744 10727
rect 10692 10684 10744 10693
rect 5724 10548 5776 10600
rect 6092 10548 6144 10600
rect 6552 10616 6604 10668
rect 6920 10616 6972 10668
rect 8760 10616 8812 10668
rect 9128 10616 9180 10668
rect 6828 10548 6880 10600
rect 8852 10548 8904 10600
rect 2780 10412 2832 10464
rect 3056 10455 3108 10464
rect 3056 10421 3065 10455
rect 3065 10421 3099 10455
rect 3099 10421 3108 10455
rect 3056 10412 3108 10421
rect 4436 10412 4488 10464
rect 7196 10480 7248 10532
rect 8484 10480 8536 10532
rect 9496 10548 9548 10600
rect 10140 10616 10192 10668
rect 14648 10684 14700 10736
rect 16396 10684 16448 10736
rect 16856 10684 16908 10736
rect 17592 10684 17644 10736
rect 11520 10659 11572 10668
rect 11520 10625 11529 10659
rect 11529 10625 11563 10659
rect 11563 10625 11572 10659
rect 11520 10616 11572 10625
rect 10232 10548 10284 10600
rect 10968 10548 11020 10600
rect 11152 10548 11204 10600
rect 11704 10548 11756 10600
rect 13268 10616 13320 10668
rect 17316 10659 17368 10668
rect 10508 10480 10560 10532
rect 12164 10523 12216 10532
rect 12164 10489 12173 10523
rect 12173 10489 12207 10523
rect 12207 10489 12216 10523
rect 12164 10480 12216 10489
rect 12256 10480 12308 10532
rect 13360 10548 13412 10600
rect 14096 10548 14148 10600
rect 15108 10548 15160 10600
rect 16212 10591 16264 10600
rect 16212 10557 16221 10591
rect 16221 10557 16255 10591
rect 16255 10557 16264 10591
rect 16212 10548 16264 10557
rect 16304 10591 16356 10600
rect 16304 10557 16313 10591
rect 16313 10557 16347 10591
rect 16347 10557 16356 10591
rect 16856 10591 16908 10600
rect 16304 10548 16356 10557
rect 16856 10557 16865 10591
rect 16865 10557 16899 10591
rect 16899 10557 16908 10591
rect 16856 10548 16908 10557
rect 17316 10625 17325 10659
rect 17325 10625 17359 10659
rect 17359 10625 17368 10659
rect 17316 10616 17368 10625
rect 18144 10659 18196 10668
rect 18144 10625 18153 10659
rect 18153 10625 18187 10659
rect 18187 10625 18196 10659
rect 18144 10616 18196 10625
rect 18788 10616 18840 10668
rect 17960 10548 18012 10600
rect 5540 10412 5592 10464
rect 6828 10455 6880 10464
rect 6828 10421 6837 10455
rect 6837 10421 6871 10455
rect 6871 10421 6880 10455
rect 6828 10412 6880 10421
rect 6920 10412 6972 10464
rect 8116 10412 8168 10464
rect 10048 10412 10100 10464
rect 10692 10412 10744 10464
rect 11704 10412 11756 10464
rect 12624 10412 12676 10464
rect 13176 10412 13228 10464
rect 14832 10455 14884 10464
rect 14832 10421 14841 10455
rect 14841 10421 14875 10455
rect 14875 10421 14884 10455
rect 14832 10412 14884 10421
rect 17500 10480 17552 10532
rect 17684 10480 17736 10532
rect 18512 10480 18564 10532
rect 19708 10480 19760 10532
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 3174 10310 3226 10362
rect 3238 10310 3290 10362
rect 3302 10310 3354 10362
rect 3366 10310 3418 10362
rect 3430 10310 3482 10362
rect 7622 10310 7674 10362
rect 7686 10310 7738 10362
rect 7750 10310 7802 10362
rect 7814 10310 7866 10362
rect 7878 10310 7930 10362
rect 12070 10310 12122 10362
rect 12134 10310 12186 10362
rect 12198 10310 12250 10362
rect 12262 10310 12314 10362
rect 12326 10310 12378 10362
rect 16518 10310 16570 10362
rect 16582 10310 16634 10362
rect 16646 10310 16698 10362
rect 16710 10310 16762 10362
rect 16774 10310 16826 10362
rect 1952 10208 2004 10260
rect 3792 10208 3844 10260
rect 6276 10208 6328 10260
rect 6736 10208 6788 10260
rect 2504 10140 2556 10192
rect 3608 10140 3660 10192
rect 3884 10140 3936 10192
rect 6552 10140 6604 10192
rect 8116 10208 8168 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 8852 10208 8904 10260
rect 9496 10251 9548 10260
rect 9496 10217 9505 10251
rect 9505 10217 9539 10251
rect 9539 10217 9548 10251
rect 9496 10208 9548 10217
rect 9588 10208 9640 10260
rect 10508 10208 10560 10260
rect 11336 10208 11388 10260
rect 2780 10072 2832 10124
rect 3056 10072 3108 10124
rect 3516 10072 3568 10124
rect 4988 10115 5040 10124
rect 4988 10081 4997 10115
rect 4997 10081 5031 10115
rect 5031 10081 5040 10115
rect 4988 10072 5040 10081
rect 5080 10072 5132 10124
rect 5816 10072 5868 10124
rect 6092 10072 6144 10124
rect 6460 10072 6512 10124
rect 7472 10072 7524 10124
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 8024 10072 8076 10124
rect 2136 10004 2188 10056
rect 1860 9936 1912 9988
rect 2688 10004 2740 10056
rect 3608 10047 3660 10056
rect 3608 10013 3617 10047
rect 3617 10013 3651 10047
rect 3651 10013 3660 10047
rect 3608 10004 3660 10013
rect 4068 10047 4120 10056
rect 4068 10013 4077 10047
rect 4077 10013 4111 10047
rect 4111 10013 4120 10047
rect 4068 10004 4120 10013
rect 4344 10047 4396 10056
rect 4344 10013 4353 10047
rect 4353 10013 4387 10047
rect 4387 10013 4396 10047
rect 4344 10004 4396 10013
rect 4252 9936 4304 9988
rect 5540 9936 5592 9988
rect 5816 9936 5868 9988
rect 6828 10004 6880 10056
rect 10232 10140 10284 10192
rect 8484 10072 8536 10124
rect 8392 10047 8444 10056
rect 8392 10013 8401 10047
rect 8401 10013 8435 10047
rect 8435 10013 8444 10047
rect 8392 10004 8444 10013
rect 9588 10072 9640 10124
rect 8668 9936 8720 9988
rect 3700 9868 3752 9920
rect 3884 9911 3936 9920
rect 3884 9877 3893 9911
rect 3893 9877 3927 9911
rect 3927 9877 3936 9911
rect 3884 9868 3936 9877
rect 4160 9911 4212 9920
rect 4160 9877 4169 9911
rect 4169 9877 4203 9911
rect 4203 9877 4212 9911
rect 4160 9868 4212 9877
rect 4344 9868 4396 9920
rect 6460 9868 6512 9920
rect 6920 9868 6972 9920
rect 7748 9868 7800 9920
rect 9312 10004 9364 10056
rect 9864 10047 9916 10056
rect 9864 10013 9873 10047
rect 9873 10013 9907 10047
rect 9907 10013 9916 10047
rect 9864 10004 9916 10013
rect 9496 9936 9548 9988
rect 11336 10004 11388 10056
rect 11704 10004 11756 10056
rect 14740 10208 14792 10260
rect 16028 10208 16080 10260
rect 17040 10208 17092 10260
rect 12624 9979 12676 9988
rect 9588 9868 9640 9920
rect 10232 9868 10284 9920
rect 12348 9868 12400 9920
rect 12624 9945 12658 9979
rect 12658 9945 12676 9979
rect 12624 9936 12676 9945
rect 14924 10140 14976 10192
rect 14096 10072 14148 10124
rect 15844 10115 15896 10124
rect 15844 10081 15853 10115
rect 15853 10081 15887 10115
rect 15887 10081 15896 10115
rect 15844 10072 15896 10081
rect 16028 10115 16080 10124
rect 16028 10081 16037 10115
rect 16037 10081 16071 10115
rect 16071 10081 16080 10115
rect 16028 10072 16080 10081
rect 17224 10140 17276 10192
rect 18420 10140 18472 10192
rect 17960 10115 18012 10124
rect 17960 10081 17969 10115
rect 17969 10081 18003 10115
rect 18003 10081 18012 10115
rect 17960 10072 18012 10081
rect 14372 10047 14424 10056
rect 14372 10013 14381 10047
rect 14381 10013 14415 10047
rect 14415 10013 14424 10047
rect 14372 10004 14424 10013
rect 16304 10004 16356 10056
rect 16948 10047 17000 10056
rect 16948 10013 16957 10047
rect 16957 10013 16991 10047
rect 16991 10013 17000 10047
rect 16948 10004 17000 10013
rect 18236 10047 18288 10056
rect 15200 9936 15252 9988
rect 15384 9979 15436 9988
rect 15384 9945 15393 9979
rect 15393 9945 15427 9979
rect 15427 9945 15436 9979
rect 15384 9936 15436 9945
rect 15660 9936 15712 9988
rect 17500 9936 17552 9988
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18328 9936 18380 9988
rect 13728 9911 13780 9920
rect 13728 9877 13737 9911
rect 13737 9877 13771 9911
rect 13771 9877 13780 9911
rect 13728 9868 13780 9877
rect 14832 9911 14884 9920
rect 14832 9877 14841 9911
rect 14841 9877 14875 9911
rect 14875 9877 14884 9911
rect 14832 9868 14884 9877
rect 14924 9911 14976 9920
rect 14924 9877 14933 9911
rect 14933 9877 14967 9911
rect 14967 9877 14976 9911
rect 16488 9911 16540 9920
rect 14924 9868 14976 9877
rect 16488 9877 16497 9911
rect 16497 9877 16531 9911
rect 16531 9877 16540 9911
rect 16488 9868 16540 9877
rect 17776 9911 17828 9920
rect 17776 9877 17785 9911
rect 17785 9877 17819 9911
rect 17819 9877 17828 9911
rect 17776 9868 17828 9877
rect 18420 9911 18472 9920
rect 18420 9877 18429 9911
rect 18429 9877 18463 9911
rect 18463 9877 18472 9911
rect 18420 9868 18472 9877
rect 5398 9766 5450 9818
rect 5462 9766 5514 9818
rect 5526 9766 5578 9818
rect 5590 9766 5642 9818
rect 5654 9766 5706 9818
rect 9846 9766 9898 9818
rect 9910 9766 9962 9818
rect 9974 9766 10026 9818
rect 10038 9766 10090 9818
rect 10102 9766 10154 9818
rect 14294 9766 14346 9818
rect 14358 9766 14410 9818
rect 14422 9766 14474 9818
rect 14486 9766 14538 9818
rect 14550 9766 14602 9818
rect 3792 9664 3844 9716
rect 2136 9596 2188 9648
rect 5080 9664 5132 9716
rect 7564 9664 7616 9716
rect 8116 9664 8168 9716
rect 8668 9664 8720 9716
rect 9680 9664 9732 9716
rect 9772 9664 9824 9716
rect 10416 9664 10468 9716
rect 11612 9664 11664 9716
rect 1952 9571 2004 9580
rect 1952 9537 1961 9571
rect 1961 9537 1995 9571
rect 1995 9537 2004 9571
rect 1952 9528 2004 9537
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 1400 9460 1452 9512
rect 2504 9528 2556 9580
rect 3884 9571 3936 9580
rect 3884 9537 3902 9571
rect 3902 9537 3936 9571
rect 3884 9528 3936 9537
rect 4068 9528 4120 9580
rect 1952 9392 2004 9444
rect 2228 9324 2280 9376
rect 2780 9367 2832 9376
rect 2780 9333 2789 9367
rect 2789 9333 2823 9367
rect 2823 9333 2832 9367
rect 2780 9324 2832 9333
rect 6552 9596 6604 9648
rect 7104 9596 7156 9648
rect 8484 9596 8536 9648
rect 7656 9528 7708 9580
rect 7840 9571 7892 9580
rect 7840 9537 7849 9571
rect 7849 9537 7883 9571
rect 7883 9537 7892 9571
rect 7840 9528 7892 9537
rect 8024 9528 8076 9580
rect 8668 9528 8720 9580
rect 10232 9528 10284 9580
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 12440 9596 12492 9648
rect 14096 9664 14148 9716
rect 14832 9664 14884 9716
rect 15292 9664 15344 9716
rect 17224 9664 17276 9716
rect 17500 9664 17552 9716
rect 17776 9664 17828 9716
rect 10784 9528 10836 9537
rect 4988 9503 5040 9512
rect 4988 9469 4997 9503
rect 4997 9469 5031 9503
rect 5031 9469 5040 9503
rect 4988 9460 5040 9469
rect 6368 9460 6420 9512
rect 10968 9503 11020 9512
rect 4160 9324 4212 9376
rect 4436 9367 4488 9376
rect 4436 9333 4445 9367
rect 4445 9333 4479 9367
rect 4479 9333 4488 9367
rect 4436 9324 4488 9333
rect 5080 9324 5132 9376
rect 5816 9392 5868 9444
rect 6184 9324 6236 9376
rect 6828 9324 6880 9376
rect 10968 9469 10977 9503
rect 10977 9469 11011 9503
rect 11011 9469 11020 9503
rect 10968 9460 11020 9469
rect 7932 9392 7984 9444
rect 9496 9435 9548 9444
rect 9496 9401 9505 9435
rect 9505 9401 9539 9435
rect 9539 9401 9548 9435
rect 9496 9392 9548 9401
rect 11704 9392 11756 9444
rect 12624 9528 12676 9580
rect 14188 9596 14240 9648
rect 13360 9460 13412 9512
rect 13728 9392 13780 9444
rect 14924 9528 14976 9580
rect 15568 9596 15620 9648
rect 16488 9596 16540 9648
rect 17040 9639 17092 9648
rect 17040 9605 17049 9639
rect 17049 9605 17083 9639
rect 17083 9605 17092 9639
rect 17040 9596 17092 9605
rect 18236 9596 18288 9648
rect 19524 9596 19576 9648
rect 16764 9528 16816 9580
rect 18972 9528 19024 9580
rect 14740 9503 14792 9512
rect 14740 9469 14749 9503
rect 14749 9469 14783 9503
rect 14783 9469 14792 9503
rect 14740 9460 14792 9469
rect 16120 9392 16172 9444
rect 17684 9392 17736 9444
rect 17868 9392 17920 9444
rect 9772 9324 9824 9376
rect 10232 9367 10284 9376
rect 10232 9333 10241 9367
rect 10241 9333 10275 9367
rect 10275 9333 10284 9367
rect 10232 9324 10284 9333
rect 11612 9367 11664 9376
rect 11612 9333 11621 9367
rect 11621 9333 11655 9367
rect 11655 9333 11664 9367
rect 11612 9324 11664 9333
rect 12532 9324 12584 9376
rect 13452 9324 13504 9376
rect 14740 9324 14792 9376
rect 3174 9222 3226 9274
rect 3238 9222 3290 9274
rect 3302 9222 3354 9274
rect 3366 9222 3418 9274
rect 3430 9222 3482 9274
rect 7622 9222 7674 9274
rect 7686 9222 7738 9274
rect 7750 9222 7802 9274
rect 7814 9222 7866 9274
rect 7878 9222 7930 9274
rect 12070 9222 12122 9274
rect 12134 9222 12186 9274
rect 12198 9222 12250 9274
rect 12262 9222 12314 9274
rect 12326 9222 12378 9274
rect 16518 9222 16570 9274
rect 16582 9222 16634 9274
rect 16646 9222 16698 9274
rect 16710 9222 16762 9274
rect 16774 9222 16826 9274
rect 2872 9120 2924 9172
rect 3976 9163 4028 9172
rect 1768 9052 1820 9104
rect 3976 9129 3985 9163
rect 3985 9129 4019 9163
rect 4019 9129 4028 9163
rect 3976 9120 4028 9129
rect 4160 9120 4212 9172
rect 1676 9027 1728 9036
rect 1676 8993 1685 9027
rect 1685 8993 1719 9027
rect 1719 8993 1728 9027
rect 1676 8984 1728 8993
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 2596 8916 2648 8968
rect 4068 9052 4120 9104
rect 6368 9120 6420 9172
rect 8024 9120 8076 9172
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 6644 9052 6696 9104
rect 4528 8984 4580 8993
rect 6184 8984 6236 9036
rect 3792 8959 3844 8968
rect 1308 8848 1360 8900
rect 1768 8823 1820 8832
rect 1768 8789 1777 8823
rect 1777 8789 1811 8823
rect 1811 8789 1820 8823
rect 1768 8780 1820 8789
rect 2136 8848 2188 8900
rect 3792 8925 3801 8959
rect 3801 8925 3835 8959
rect 3835 8925 3844 8959
rect 3792 8916 3844 8925
rect 5356 8959 5408 8968
rect 3516 8848 3568 8900
rect 3976 8848 4028 8900
rect 4436 8891 4488 8900
rect 4436 8857 4445 8891
rect 4445 8857 4479 8891
rect 4479 8857 4488 8891
rect 4436 8848 4488 8857
rect 3700 8780 3752 8832
rect 3792 8780 3844 8832
rect 4160 8780 4212 8832
rect 4344 8823 4396 8832
rect 4344 8789 4353 8823
rect 4353 8789 4387 8823
rect 4387 8789 4396 8823
rect 4344 8780 4396 8789
rect 4528 8780 4580 8832
rect 5356 8925 5390 8959
rect 5390 8925 5408 8959
rect 5356 8916 5408 8925
rect 6736 8916 6788 8968
rect 5724 8848 5776 8900
rect 6828 8848 6880 8900
rect 8392 8916 8444 8968
rect 7564 8891 7616 8900
rect 7564 8857 7598 8891
rect 7598 8857 7616 8891
rect 7564 8848 7616 8857
rect 5080 8780 5132 8832
rect 6276 8780 6328 8832
rect 9496 9120 9548 9172
rect 9680 9120 9732 9172
rect 11244 9120 11296 9172
rect 11704 9120 11756 9172
rect 13360 9120 13412 9172
rect 14004 9120 14056 9172
rect 14096 9163 14148 9172
rect 14096 9129 14105 9163
rect 14105 9129 14139 9163
rect 14139 9129 14148 9163
rect 14096 9120 14148 9129
rect 9312 9052 9364 9104
rect 10692 9095 10744 9104
rect 10692 9061 10701 9095
rect 10701 9061 10735 9095
rect 10735 9061 10744 9095
rect 10692 9052 10744 9061
rect 10968 8984 11020 9036
rect 13820 9052 13872 9104
rect 18144 9120 18196 9172
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 13452 8984 13504 9036
rect 16120 8984 16172 9036
rect 18696 8984 18748 9036
rect 19340 8984 19392 9036
rect 8576 8916 8628 8968
rect 8760 8916 8812 8968
rect 9312 8959 9364 8968
rect 9312 8925 9321 8959
rect 9321 8925 9355 8959
rect 9355 8925 9364 8959
rect 9312 8916 9364 8925
rect 9404 8916 9456 8968
rect 10324 8916 10376 8968
rect 10876 8916 10928 8968
rect 12072 8916 12124 8968
rect 12716 8916 12768 8968
rect 13728 8916 13780 8968
rect 14188 8916 14240 8968
rect 15844 8916 15896 8968
rect 16212 8916 16264 8968
rect 17132 8916 17184 8968
rect 18328 8916 18380 8968
rect 18512 8959 18564 8968
rect 18512 8925 18521 8959
rect 18521 8925 18555 8959
rect 18555 8925 18564 8959
rect 18512 8916 18564 8925
rect 8852 8848 8904 8900
rect 8668 8823 8720 8832
rect 8668 8789 8677 8823
rect 8677 8789 8711 8823
rect 8711 8789 8720 8823
rect 8668 8780 8720 8789
rect 8760 8780 8812 8832
rect 9772 8780 9824 8832
rect 10968 8780 11020 8832
rect 13360 8848 13412 8900
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 12624 8780 12676 8832
rect 13176 8780 13228 8832
rect 13452 8780 13504 8832
rect 15200 8891 15252 8900
rect 15200 8857 15218 8891
rect 15218 8857 15252 8891
rect 15200 8848 15252 8857
rect 15568 8848 15620 8900
rect 16304 8848 16356 8900
rect 17132 8780 17184 8832
rect 17224 8780 17276 8832
rect 18052 8823 18104 8832
rect 18052 8789 18061 8823
rect 18061 8789 18095 8823
rect 18095 8789 18104 8823
rect 18052 8780 18104 8789
rect 5398 8678 5450 8730
rect 5462 8678 5514 8730
rect 5526 8678 5578 8730
rect 5590 8678 5642 8730
rect 5654 8678 5706 8730
rect 9846 8678 9898 8730
rect 9910 8678 9962 8730
rect 9974 8678 10026 8730
rect 10038 8678 10090 8730
rect 10102 8678 10154 8730
rect 14294 8678 14346 8730
rect 14358 8678 14410 8730
rect 14422 8678 14474 8730
rect 14486 8678 14538 8730
rect 14550 8678 14602 8730
rect 2780 8576 2832 8628
rect 1676 8508 1728 8560
rect 2504 8508 2556 8560
rect 3240 8508 3292 8560
rect 1768 8483 1820 8492
rect 1768 8449 1802 8483
rect 1802 8449 1820 8483
rect 1768 8440 1820 8449
rect 2596 8440 2648 8492
rect 3148 8372 3200 8424
rect 3424 8508 3476 8560
rect 3792 8508 3844 8560
rect 3884 8508 3936 8560
rect 8484 8576 8536 8628
rect 6828 8508 6880 8560
rect 2964 8304 3016 8356
rect 3976 8483 4028 8492
rect 3976 8449 3985 8483
rect 3985 8449 4019 8483
rect 4019 8449 4028 8483
rect 5816 8483 5868 8492
rect 3976 8440 4028 8449
rect 5816 8449 5825 8483
rect 5825 8449 5859 8483
rect 5859 8449 5868 8483
rect 5816 8440 5868 8449
rect 10232 8576 10284 8628
rect 10784 8576 10836 8628
rect 12440 8619 12492 8628
rect 9312 8508 9364 8560
rect 12440 8585 12449 8619
rect 12449 8585 12483 8619
rect 12483 8585 12492 8619
rect 12440 8576 12492 8585
rect 12624 8619 12676 8628
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 12716 8576 12768 8628
rect 13728 8576 13780 8628
rect 13912 8576 13964 8628
rect 15292 8576 15344 8628
rect 16028 8576 16080 8628
rect 17132 8619 17184 8628
rect 17132 8585 17141 8619
rect 17141 8585 17175 8619
rect 17175 8585 17184 8619
rect 17132 8576 17184 8585
rect 17316 8576 17368 8628
rect 18328 8619 18380 8628
rect 18328 8585 18337 8619
rect 18337 8585 18371 8619
rect 18371 8585 18380 8619
rect 18328 8576 18380 8585
rect 6184 8372 6236 8424
rect 1492 8236 1544 8288
rect 2228 8236 2280 8288
rect 3700 8254 3752 8306
rect 3884 8254 3936 8306
rect 6000 8304 6052 8356
rect 6736 8304 6788 8356
rect 4344 8236 4396 8288
rect 6276 8236 6328 8288
rect 6368 8236 6420 8288
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9680 8440 9732 8492
rect 10140 8440 10192 8492
rect 10692 8440 10744 8492
rect 11796 8483 11848 8492
rect 11796 8449 11805 8483
rect 11805 8449 11839 8483
rect 11839 8449 11848 8483
rect 11796 8440 11848 8449
rect 15476 8508 15528 8560
rect 15292 8440 15344 8492
rect 15844 8483 15896 8492
rect 15844 8449 15853 8483
rect 15853 8449 15887 8483
rect 15887 8449 15896 8483
rect 15844 8440 15896 8449
rect 15936 8483 15988 8492
rect 15936 8449 15945 8483
rect 15945 8449 15979 8483
rect 15979 8449 15988 8483
rect 15936 8440 15988 8449
rect 16304 8440 16356 8492
rect 11336 8415 11388 8424
rect 7104 8236 7156 8288
rect 9404 8304 9456 8356
rect 11336 8381 11345 8415
rect 11345 8381 11379 8415
rect 11379 8381 11388 8415
rect 11336 8372 11388 8381
rect 12072 8372 12124 8424
rect 13084 8415 13136 8424
rect 13084 8381 13093 8415
rect 13093 8381 13127 8415
rect 13127 8381 13136 8415
rect 13084 8372 13136 8381
rect 13912 8415 13964 8424
rect 8024 8279 8076 8288
rect 8024 8245 8033 8279
rect 8033 8245 8067 8279
rect 8067 8245 8076 8279
rect 8024 8236 8076 8245
rect 9772 8236 9824 8288
rect 13912 8381 13921 8415
rect 13921 8381 13955 8415
rect 13955 8381 13964 8415
rect 13912 8372 13964 8381
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 16856 8508 16908 8560
rect 18604 8508 18656 8560
rect 17040 8483 17092 8492
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 18236 8440 18288 8492
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 16120 8347 16172 8356
rect 11704 8236 11756 8288
rect 11888 8236 11940 8288
rect 13268 8236 13320 8288
rect 14556 8236 14608 8288
rect 16120 8313 16129 8347
rect 16129 8313 16163 8347
rect 16163 8313 16172 8347
rect 16120 8304 16172 8313
rect 16212 8304 16264 8356
rect 17868 8304 17920 8356
rect 16304 8236 16356 8288
rect 3174 8134 3226 8186
rect 3238 8134 3290 8186
rect 3302 8134 3354 8186
rect 3366 8134 3418 8186
rect 3430 8134 3482 8186
rect 7622 8134 7674 8186
rect 7686 8134 7738 8186
rect 7750 8134 7802 8186
rect 7814 8134 7866 8186
rect 7878 8134 7930 8186
rect 12070 8134 12122 8186
rect 12134 8134 12186 8186
rect 12198 8134 12250 8186
rect 12262 8134 12314 8186
rect 12326 8134 12378 8186
rect 16518 8134 16570 8186
rect 16582 8134 16634 8186
rect 16646 8134 16698 8186
rect 16710 8134 16762 8186
rect 16774 8134 16826 8186
rect 1768 8032 1820 8084
rect 2964 8032 3016 8084
rect 4160 8032 4212 8084
rect 1676 7964 1728 8016
rect 1952 7964 2004 8016
rect 2688 7964 2740 8016
rect 3056 7964 3108 8016
rect 3332 7964 3384 8016
rect 2504 7896 2556 7948
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2596 7828 2648 7880
rect 2780 7828 2832 7880
rect 3240 7896 3292 7948
rect 5724 8075 5776 8084
rect 4436 8007 4488 8016
rect 4436 7973 4445 8007
rect 4445 7973 4479 8007
rect 4479 7973 4488 8007
rect 4436 7964 4488 7973
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6276 8032 6328 8084
rect 5908 7964 5960 8016
rect 7012 7964 7064 8016
rect 7840 7964 7892 8016
rect 7932 7964 7984 8016
rect 756 7760 808 7812
rect 1584 7692 1636 7744
rect 2044 7692 2096 7744
rect 3516 7828 3568 7880
rect 3792 7828 3844 7880
rect 3608 7760 3660 7812
rect 6920 7896 6972 7948
rect 7748 7939 7800 7948
rect 7748 7905 7757 7939
rect 7757 7905 7791 7939
rect 7791 7905 7800 7939
rect 7748 7896 7800 7905
rect 4344 7760 4396 7812
rect 4528 7760 4580 7812
rect 4620 7692 4672 7744
rect 5264 7692 5316 7744
rect 5908 7760 5960 7812
rect 7104 7828 7156 7880
rect 7380 7828 7432 7880
rect 7564 7828 7616 7880
rect 11244 8032 11296 8084
rect 11704 8032 11756 8084
rect 13820 8032 13872 8084
rect 17316 8032 17368 8084
rect 8392 7896 8444 7948
rect 10784 7964 10836 8016
rect 9220 7871 9272 7880
rect 7196 7760 7248 7812
rect 6460 7692 6512 7744
rect 7104 7735 7156 7744
rect 7104 7701 7113 7735
rect 7113 7701 7147 7735
rect 7147 7701 7156 7735
rect 7104 7692 7156 7701
rect 7656 7760 7708 7812
rect 9220 7837 9229 7871
rect 9229 7837 9263 7871
rect 9263 7837 9272 7871
rect 9220 7828 9272 7837
rect 7932 7692 7984 7744
rect 10232 7896 10284 7948
rect 11336 7896 11388 7948
rect 16212 7939 16264 7948
rect 10416 7828 10468 7880
rect 9588 7760 9640 7812
rect 11060 7760 11112 7812
rect 11336 7760 11388 7812
rect 13544 7828 13596 7880
rect 14004 7828 14056 7880
rect 14188 7828 14240 7880
rect 14556 7828 14608 7880
rect 16212 7905 16221 7939
rect 16221 7905 16255 7939
rect 16255 7905 16264 7939
rect 16212 7896 16264 7905
rect 17224 7896 17276 7948
rect 17500 7828 17552 7880
rect 17960 7828 18012 7880
rect 19432 7828 19484 7880
rect 12716 7760 12768 7812
rect 10876 7692 10928 7744
rect 11244 7692 11296 7744
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 13820 7735 13872 7744
rect 13820 7701 13829 7735
rect 13829 7701 13863 7735
rect 13863 7701 13872 7735
rect 13820 7692 13872 7701
rect 14096 7692 14148 7744
rect 14740 7692 14792 7744
rect 16672 7735 16724 7744
rect 16672 7701 16681 7735
rect 16681 7701 16715 7735
rect 16715 7701 16724 7735
rect 16672 7692 16724 7701
rect 16948 7760 17000 7812
rect 16856 7692 16908 7744
rect 17592 7735 17644 7744
rect 17592 7701 17601 7735
rect 17601 7701 17635 7735
rect 17635 7701 17644 7735
rect 17592 7692 17644 7701
rect 17960 7735 18012 7744
rect 17960 7701 17969 7735
rect 17969 7701 18003 7735
rect 18003 7701 18012 7735
rect 17960 7692 18012 7701
rect 18788 7692 18840 7744
rect 5398 7590 5450 7642
rect 5462 7590 5514 7642
rect 5526 7590 5578 7642
rect 5590 7590 5642 7642
rect 5654 7590 5706 7642
rect 9846 7590 9898 7642
rect 9910 7590 9962 7642
rect 9974 7590 10026 7642
rect 10038 7590 10090 7642
rect 10102 7590 10154 7642
rect 14294 7590 14346 7642
rect 14358 7590 14410 7642
rect 14422 7590 14474 7642
rect 14486 7590 14538 7642
rect 14550 7590 14602 7642
rect 940 7488 992 7540
rect 1400 7488 1452 7540
rect 2136 7488 2188 7540
rect 2320 7488 2372 7540
rect 3056 7488 3108 7540
rect 1952 7420 2004 7472
rect 4252 7488 4304 7540
rect 5264 7488 5316 7540
rect 6368 7531 6420 7540
rect 6368 7497 6377 7531
rect 6377 7497 6411 7531
rect 6411 7497 6420 7531
rect 6368 7488 6420 7497
rect 6920 7488 6972 7540
rect 8852 7531 8904 7540
rect 3976 7420 4028 7472
rect 5448 7420 5500 7472
rect 5724 7420 5776 7472
rect 6828 7420 6880 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2136 7395 2188 7404
rect 2136 7361 2145 7395
rect 2145 7361 2179 7395
rect 2179 7361 2188 7395
rect 2136 7352 2188 7361
rect 2504 7352 2556 7404
rect 2964 7352 3016 7404
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 1768 7284 1820 7336
rect 2688 7284 2740 7336
rect 4160 7284 4212 7336
rect 4436 7284 4488 7336
rect 4620 7284 4672 7336
rect 4896 7352 4948 7404
rect 5632 7284 5684 7336
rect 7656 7352 7708 7404
rect 7932 7420 7984 7472
rect 8852 7497 8861 7531
rect 8861 7497 8895 7531
rect 8895 7497 8904 7531
rect 8852 7488 8904 7497
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 11336 7488 11388 7540
rect 12900 7531 12952 7540
rect 12900 7497 12909 7531
rect 12909 7497 12943 7531
rect 12943 7497 12952 7531
rect 12900 7488 12952 7497
rect 13912 7488 13964 7540
rect 15476 7488 15528 7540
rect 7840 7395 7892 7404
rect 7840 7361 7849 7395
rect 7849 7361 7883 7395
rect 7883 7361 7892 7395
rect 7840 7352 7892 7361
rect 7932 7284 7984 7336
rect 388 7216 440 7268
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 4436 7191 4488 7200
rect 4436 7157 4445 7191
rect 4445 7157 4479 7191
rect 4479 7157 4488 7191
rect 4436 7148 4488 7157
rect 4528 7148 4580 7200
rect 10416 7352 10468 7404
rect 11704 7420 11756 7472
rect 16948 7488 17000 7540
rect 17592 7488 17644 7540
rect 11796 7395 11848 7404
rect 11796 7361 11830 7395
rect 11830 7361 11848 7395
rect 9680 7284 9732 7336
rect 9772 7284 9824 7336
rect 11796 7352 11848 7361
rect 12716 7352 12768 7404
rect 13176 7352 13228 7404
rect 16212 7420 16264 7472
rect 16672 7420 16724 7472
rect 15476 7352 15528 7404
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 17960 7352 18012 7404
rect 11244 7284 11296 7336
rect 8484 7191 8536 7200
rect 8484 7157 8493 7191
rect 8493 7157 8527 7191
rect 8527 7157 8536 7191
rect 8484 7148 8536 7157
rect 15108 7284 15160 7336
rect 15292 7327 15344 7336
rect 15292 7293 15301 7327
rect 15301 7293 15335 7327
rect 15335 7293 15344 7327
rect 15292 7284 15344 7293
rect 17316 7327 17368 7336
rect 13728 7216 13780 7268
rect 15200 7216 15252 7268
rect 17316 7293 17325 7327
rect 17325 7293 17359 7327
rect 17359 7293 17368 7327
rect 17316 7284 17368 7293
rect 17500 7284 17552 7336
rect 16672 7259 16724 7268
rect 16672 7225 16681 7259
rect 16681 7225 16715 7259
rect 16715 7225 16724 7259
rect 16672 7216 16724 7225
rect 14004 7148 14056 7200
rect 14188 7148 14240 7200
rect 18236 7148 18288 7200
rect 3174 7046 3226 7098
rect 3238 7046 3290 7098
rect 3302 7046 3354 7098
rect 3366 7046 3418 7098
rect 3430 7046 3482 7098
rect 7622 7046 7674 7098
rect 7686 7046 7738 7098
rect 7750 7046 7802 7098
rect 7814 7046 7866 7098
rect 7878 7046 7930 7098
rect 12070 7046 12122 7098
rect 12134 7046 12186 7098
rect 12198 7046 12250 7098
rect 12262 7046 12314 7098
rect 12326 7046 12378 7098
rect 16518 7046 16570 7098
rect 16582 7046 16634 7098
rect 16646 7046 16698 7098
rect 16710 7046 16762 7098
rect 16774 7046 16826 7098
rect 3148 6876 3200 6928
rect 20 6808 72 6860
rect 940 6808 992 6860
rect 3424 6808 3476 6860
rect 4620 6876 4672 6928
rect 4988 6876 5040 6928
rect 4436 6808 4488 6860
rect 2504 6740 2556 6792
rect 1584 6672 1636 6724
rect 4528 6740 4580 6792
rect 3424 6604 3476 6656
rect 3516 6604 3568 6656
rect 4620 6604 4672 6656
rect 6644 6944 6696 6996
rect 7196 6987 7248 6996
rect 6276 6876 6328 6928
rect 6736 6876 6788 6928
rect 6828 6808 6880 6860
rect 7196 6953 7205 6987
rect 7205 6953 7239 6987
rect 7239 6953 7248 6987
rect 7196 6944 7248 6953
rect 7564 6876 7616 6928
rect 8254 6944 8306 6996
rect 10416 6987 10468 6996
rect 8392 6876 8444 6928
rect 7564 6783 7616 6792
rect 7564 6749 7573 6783
rect 7573 6749 7607 6783
rect 7607 6749 7616 6783
rect 7564 6740 7616 6749
rect 7932 6808 7984 6860
rect 8484 6808 8536 6860
rect 10416 6953 10425 6987
rect 10425 6953 10459 6987
rect 10459 6953 10468 6987
rect 10416 6944 10468 6953
rect 12808 6944 12860 6996
rect 13176 6944 13228 6996
rect 8668 6740 8720 6792
rect 6092 6672 6144 6724
rect 7932 6672 7984 6724
rect 6460 6604 6512 6656
rect 7012 6604 7064 6656
rect 7380 6604 7432 6656
rect 8116 6604 8168 6656
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 8668 6604 8720 6656
rect 10692 6808 10744 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 11244 6740 11296 6792
rect 11520 6783 11572 6792
rect 11520 6749 11529 6783
rect 11529 6749 11563 6783
rect 11563 6749 11572 6783
rect 11520 6740 11572 6749
rect 13360 6808 13412 6860
rect 9680 6672 9732 6724
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 14004 6944 14056 6996
rect 15200 6944 15252 6996
rect 15936 6944 15988 6996
rect 17868 6944 17920 6996
rect 17224 6876 17276 6928
rect 13728 6851 13780 6860
rect 13728 6817 13737 6851
rect 13737 6817 13771 6851
rect 13771 6817 13780 6851
rect 13728 6808 13780 6817
rect 17776 6851 17828 6860
rect 17776 6817 17785 6851
rect 17785 6817 17819 6851
rect 17819 6817 17828 6851
rect 17776 6808 17828 6817
rect 13820 6672 13872 6724
rect 11428 6604 11480 6656
rect 11704 6604 11756 6656
rect 13084 6604 13136 6656
rect 13360 6604 13412 6656
rect 14832 6672 14884 6724
rect 15384 6740 15436 6792
rect 16672 6740 16724 6792
rect 17132 6783 17184 6792
rect 17132 6749 17141 6783
rect 17141 6749 17175 6783
rect 17175 6749 17184 6783
rect 17132 6740 17184 6749
rect 15568 6672 15620 6724
rect 16396 6672 16448 6724
rect 18972 6740 19024 6792
rect 15292 6604 15344 6656
rect 16488 6604 16540 6656
rect 16856 6604 16908 6656
rect 17040 6647 17092 6656
rect 17040 6613 17049 6647
rect 17049 6613 17083 6647
rect 17083 6613 17092 6647
rect 17040 6604 17092 6613
rect 17500 6604 17552 6656
rect 5398 6502 5450 6554
rect 5462 6502 5514 6554
rect 5526 6502 5578 6554
rect 5590 6502 5642 6554
rect 5654 6502 5706 6554
rect 9846 6502 9898 6554
rect 9910 6502 9962 6554
rect 9974 6502 10026 6554
rect 10038 6502 10090 6554
rect 10102 6502 10154 6554
rect 14294 6502 14346 6554
rect 14358 6502 14410 6554
rect 14422 6502 14474 6554
rect 14486 6502 14538 6554
rect 14550 6502 14602 6554
rect 2136 6400 2188 6452
rect 2964 6400 3016 6452
rect 4804 6443 4856 6452
rect 4804 6409 4813 6443
rect 4813 6409 4847 6443
rect 4847 6409 4856 6443
rect 4804 6400 4856 6409
rect 4988 6400 5040 6452
rect 5908 6400 5960 6452
rect 6460 6400 6512 6452
rect 7472 6400 7524 6452
rect 8392 6400 8444 6452
rect 9772 6400 9824 6452
rect 10416 6400 10468 6452
rect 11336 6443 11388 6452
rect 11336 6409 11345 6443
rect 11345 6409 11379 6443
rect 11379 6409 11388 6443
rect 11336 6400 11388 6409
rect 11796 6443 11848 6452
rect 11796 6409 11805 6443
rect 11805 6409 11839 6443
rect 11839 6409 11848 6443
rect 11796 6400 11848 6409
rect 12164 6400 12216 6452
rect 2872 6332 2924 6384
rect 3424 6332 3476 6384
rect 1676 6264 1728 6316
rect 2688 6264 2740 6316
rect 3148 6307 3200 6316
rect 3148 6273 3182 6307
rect 3182 6273 3200 6307
rect 3148 6264 3200 6273
rect 3516 6264 3568 6316
rect 4528 6264 4580 6316
rect 5356 6264 5408 6316
rect 5908 6307 5960 6316
rect 5908 6273 5926 6307
rect 5926 6273 5960 6307
rect 5908 6264 5960 6273
rect 7104 6332 7156 6384
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 1768 6196 1820 6248
rect 2136 6196 2188 6248
rect 1768 6103 1820 6112
rect 1768 6069 1777 6103
rect 1777 6069 1811 6103
rect 1811 6069 1820 6103
rect 1768 6060 1820 6069
rect 2412 6060 2464 6112
rect 4436 6196 4488 6248
rect 3976 6060 4028 6112
rect 4436 6060 4488 6112
rect 4712 6128 4764 6180
rect 5080 6128 5132 6180
rect 6368 6196 6420 6248
rect 7012 6196 7064 6248
rect 11796 6264 11848 6316
rect 12072 6264 12124 6316
rect 7840 6239 7892 6248
rect 7840 6205 7849 6239
rect 7849 6205 7883 6239
rect 7883 6205 7892 6239
rect 7840 6196 7892 6205
rect 9680 6196 9732 6248
rect 10232 6196 10284 6248
rect 10968 6239 11020 6248
rect 10968 6205 10977 6239
rect 10977 6205 11011 6239
rect 11011 6205 11020 6239
rect 10968 6196 11020 6205
rect 11704 6239 11756 6248
rect 11704 6205 11713 6239
rect 11713 6205 11747 6239
rect 11747 6205 11756 6239
rect 11704 6196 11756 6205
rect 12256 6264 12308 6316
rect 12808 6400 12860 6452
rect 13084 6400 13136 6452
rect 12992 6332 13044 6384
rect 14004 6332 14056 6384
rect 15016 6400 15068 6452
rect 18328 6443 18380 6452
rect 15200 6375 15252 6384
rect 6920 6060 6972 6112
rect 9128 6128 9180 6180
rect 11060 6128 11112 6180
rect 8300 6060 8352 6112
rect 13452 6264 13504 6316
rect 13728 6264 13780 6316
rect 15200 6341 15209 6375
rect 15209 6341 15243 6375
rect 15243 6341 15252 6375
rect 15200 6332 15252 6341
rect 15476 6332 15528 6384
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 13176 6196 13228 6248
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 12808 6128 12860 6180
rect 14832 6196 14884 6248
rect 15476 6196 15528 6248
rect 15752 6264 15804 6316
rect 16120 6239 16172 6248
rect 14556 6060 14608 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 16120 6205 16129 6239
rect 16129 6205 16163 6239
rect 16163 6205 16172 6239
rect 16120 6196 16172 6205
rect 17040 6332 17092 6384
rect 17776 6332 17828 6384
rect 18328 6409 18337 6443
rect 18337 6409 18371 6443
rect 18371 6409 18380 6443
rect 18328 6400 18380 6409
rect 18972 6332 19024 6384
rect 19708 6264 19760 6316
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 19616 6128 19668 6180
rect 17684 6060 17736 6112
rect 3174 5958 3226 6010
rect 3238 5958 3290 6010
rect 3302 5958 3354 6010
rect 3366 5958 3418 6010
rect 3430 5958 3482 6010
rect 7622 5958 7674 6010
rect 7686 5958 7738 6010
rect 7750 5958 7802 6010
rect 7814 5958 7866 6010
rect 7878 5958 7930 6010
rect 12070 5958 12122 6010
rect 12134 5958 12186 6010
rect 12198 5958 12250 6010
rect 12262 5958 12314 6010
rect 12326 5958 12378 6010
rect 16518 5958 16570 6010
rect 16582 5958 16634 6010
rect 16646 5958 16698 6010
rect 16710 5958 16762 6010
rect 16774 5958 16826 6010
rect 3516 5856 3568 5908
rect 2320 5788 2372 5840
rect 5172 5856 5224 5908
rect 6920 5856 6972 5908
rect 2964 5763 3016 5772
rect 2964 5729 2973 5763
rect 2973 5729 3007 5763
rect 3007 5729 3016 5763
rect 2964 5720 3016 5729
rect 5816 5788 5868 5840
rect 8576 5788 8628 5840
rect 1952 5652 2004 5704
rect 2412 5695 2464 5704
rect 2412 5661 2421 5695
rect 2421 5661 2455 5695
rect 2455 5661 2464 5695
rect 2412 5652 2464 5661
rect 3056 5652 3108 5704
rect 3976 5652 4028 5704
rect 6184 5720 6236 5772
rect 8116 5763 8168 5772
rect 8116 5729 8125 5763
rect 8125 5729 8159 5763
rect 8159 5729 8168 5763
rect 8116 5720 8168 5729
rect 11704 5856 11756 5908
rect 1676 5584 1728 5636
rect 4160 5584 4212 5636
rect 4436 5584 4488 5636
rect 4896 5584 4948 5636
rect 6644 5652 6696 5704
rect 8300 5652 8352 5704
rect 10508 5652 10560 5704
rect 8116 5584 8168 5636
rect 2228 5516 2280 5568
rect 5724 5516 5776 5568
rect 5908 5516 5960 5568
rect 6092 5516 6144 5568
rect 9036 5584 9088 5636
rect 9588 5584 9640 5636
rect 11336 5584 11388 5636
rect 9772 5516 9824 5568
rect 10508 5516 10560 5568
rect 11244 5516 11296 5568
rect 11796 5584 11848 5636
rect 13452 5652 13504 5704
rect 14556 5763 14608 5772
rect 14556 5729 14565 5763
rect 14565 5729 14599 5763
rect 14599 5729 14608 5763
rect 14556 5720 14608 5729
rect 14832 5856 14884 5908
rect 15568 5788 15620 5840
rect 15476 5763 15528 5772
rect 15476 5729 15485 5763
rect 15485 5729 15519 5763
rect 15519 5729 15528 5763
rect 16120 5856 16172 5908
rect 15936 5788 15988 5840
rect 15476 5720 15528 5729
rect 17684 5720 17736 5772
rect 13912 5695 13964 5704
rect 13912 5661 13921 5695
rect 13921 5661 13955 5695
rect 13955 5661 13964 5695
rect 13912 5652 13964 5661
rect 16120 5652 16172 5704
rect 17408 5652 17460 5704
rect 19064 5652 19116 5704
rect 14832 5516 14884 5568
rect 15016 5584 15068 5636
rect 17592 5584 17644 5636
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 15752 5559 15804 5568
rect 15752 5525 15761 5559
rect 15761 5525 15795 5559
rect 15795 5525 15804 5559
rect 15752 5516 15804 5525
rect 16856 5516 16908 5568
rect 18052 5516 18104 5568
rect 18420 5559 18472 5568
rect 18420 5525 18429 5559
rect 18429 5525 18463 5559
rect 18463 5525 18472 5559
rect 18420 5516 18472 5525
rect 5398 5414 5450 5466
rect 5462 5414 5514 5466
rect 5526 5414 5578 5466
rect 5590 5414 5642 5466
rect 5654 5414 5706 5466
rect 9846 5414 9898 5466
rect 9910 5414 9962 5466
rect 9974 5414 10026 5466
rect 10038 5414 10090 5466
rect 10102 5414 10154 5466
rect 14294 5414 14346 5466
rect 14358 5414 14410 5466
rect 14422 5414 14474 5466
rect 14486 5414 14538 5466
rect 14550 5414 14602 5466
rect 2044 5355 2096 5364
rect 2044 5321 2053 5355
rect 2053 5321 2087 5355
rect 2087 5321 2096 5355
rect 2044 5312 2096 5321
rect 4528 5312 4580 5364
rect 4620 5312 4672 5364
rect 4988 5312 5040 5364
rect 6184 5312 6236 5364
rect 7288 5312 7340 5364
rect 8576 5355 8628 5364
rect 8576 5321 8585 5355
rect 8585 5321 8619 5355
rect 8619 5321 8628 5355
rect 8576 5312 8628 5321
rect 9036 5355 9088 5364
rect 9036 5321 9045 5355
rect 9045 5321 9079 5355
rect 9079 5321 9088 5355
rect 9036 5312 9088 5321
rect 9312 5312 9364 5364
rect 12624 5312 12676 5364
rect 12716 5312 12768 5364
rect 1676 5176 1728 5228
rect 2688 5176 2740 5228
rect 5816 5244 5868 5296
rect 4160 5176 4212 5228
rect 4712 5176 4764 5228
rect 1584 5108 1636 5160
rect 2044 4972 2096 5024
rect 6460 5151 6512 5160
rect 2780 5040 2832 5092
rect 6460 5117 6469 5151
rect 6469 5117 6503 5151
rect 6503 5117 6512 5151
rect 6460 5108 6512 5117
rect 8484 5244 8536 5296
rect 8668 5287 8720 5296
rect 8668 5253 8677 5287
rect 8677 5253 8711 5287
rect 8711 5253 8720 5287
rect 8668 5244 8720 5253
rect 10140 5244 10192 5296
rect 6828 5176 6880 5228
rect 9312 5176 9364 5228
rect 9864 5176 9916 5228
rect 10508 5176 10560 5228
rect 10968 5219 11020 5228
rect 10968 5185 10986 5219
rect 10986 5185 11020 5219
rect 10968 5176 11020 5185
rect 11336 5244 11388 5296
rect 14004 5312 14056 5364
rect 13084 5244 13136 5296
rect 15016 5244 15068 5296
rect 17040 5244 17092 5296
rect 17684 5244 17736 5296
rect 7472 5108 7524 5160
rect 8116 5108 8168 5160
rect 9128 5108 9180 5160
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 10048 5108 10100 5160
rect 11244 5151 11296 5160
rect 11244 5117 11253 5151
rect 11253 5117 11287 5151
rect 11287 5117 11296 5151
rect 11244 5108 11296 5117
rect 3976 5040 4028 5092
rect 4160 5083 4212 5092
rect 4160 5049 4169 5083
rect 4169 5049 4203 5083
rect 4203 5049 4212 5083
rect 4160 5040 4212 5049
rect 9036 5040 9088 5092
rect 13544 5176 13596 5228
rect 13820 5176 13872 5228
rect 16764 5219 16816 5228
rect 16764 5185 16773 5219
rect 16773 5185 16807 5219
rect 16807 5185 16816 5219
rect 16764 5176 16816 5185
rect 17592 5151 17644 5160
rect 2504 5015 2556 5024
rect 2504 4981 2513 5015
rect 2513 4981 2547 5015
rect 2547 4981 2556 5015
rect 2504 4972 2556 4981
rect 3516 4972 3568 5024
rect 4528 4972 4580 5024
rect 5356 4972 5408 5024
rect 6000 5015 6052 5024
rect 6000 4981 6009 5015
rect 6009 4981 6043 5015
rect 6043 4981 6052 5015
rect 6000 4972 6052 4981
rect 7380 5015 7432 5024
rect 7380 4981 7389 5015
rect 7389 4981 7423 5015
rect 7423 4981 7432 5015
rect 7380 4972 7432 4981
rect 8024 4972 8076 5024
rect 8484 4972 8536 5024
rect 11336 4972 11388 5024
rect 11520 5015 11572 5024
rect 11520 4981 11529 5015
rect 11529 4981 11563 5015
rect 11563 4981 11572 5015
rect 11520 4972 11572 4981
rect 11796 4972 11848 5024
rect 13084 4972 13136 5024
rect 17592 5117 17601 5151
rect 17601 5117 17635 5151
rect 17635 5117 17644 5151
rect 17592 5108 17644 5117
rect 18696 5312 18748 5364
rect 18236 5219 18288 5228
rect 18236 5185 18245 5219
rect 18245 5185 18279 5219
rect 18279 5185 18288 5219
rect 18236 5176 18288 5185
rect 15384 4972 15436 5024
rect 16304 4972 16356 5024
rect 16948 5015 17000 5024
rect 16948 4981 16957 5015
rect 16957 4981 16991 5015
rect 16991 4981 17000 5015
rect 16948 4972 17000 4981
rect 17132 5015 17184 5024
rect 17132 4981 17141 5015
rect 17141 4981 17175 5015
rect 17175 4981 17184 5015
rect 17132 4972 17184 4981
rect 18236 4972 18288 5024
rect 3174 4870 3226 4922
rect 3238 4870 3290 4922
rect 3302 4870 3354 4922
rect 3366 4870 3418 4922
rect 3430 4870 3482 4922
rect 7622 4870 7674 4922
rect 7686 4870 7738 4922
rect 7750 4870 7802 4922
rect 7814 4870 7866 4922
rect 7878 4870 7930 4922
rect 12070 4870 12122 4922
rect 12134 4870 12186 4922
rect 12198 4870 12250 4922
rect 12262 4870 12314 4922
rect 12326 4870 12378 4922
rect 16518 4870 16570 4922
rect 16582 4870 16634 4922
rect 16646 4870 16698 4922
rect 16710 4870 16762 4922
rect 16774 4870 16826 4922
rect 1952 4768 2004 4820
rect 1952 4632 2004 4684
rect 2504 4768 2556 4820
rect 2872 4811 2924 4820
rect 2872 4777 2881 4811
rect 2881 4777 2915 4811
rect 2915 4777 2924 4811
rect 2872 4768 2924 4777
rect 3792 4811 3844 4820
rect 3792 4777 3801 4811
rect 3801 4777 3835 4811
rect 3835 4777 3844 4811
rect 3792 4768 3844 4777
rect 8024 4768 8076 4820
rect 9772 4768 9824 4820
rect 11980 4768 12032 4820
rect 15108 4768 15160 4820
rect 2320 4675 2372 4684
rect 2320 4641 2329 4675
rect 2329 4641 2363 4675
rect 2363 4641 2372 4675
rect 2320 4632 2372 4641
rect 1676 4607 1728 4616
rect 1676 4573 1685 4607
rect 1685 4573 1719 4607
rect 1719 4573 1728 4607
rect 1676 4564 1728 4573
rect 2412 4607 2464 4616
rect 2412 4573 2421 4607
rect 2421 4573 2455 4607
rect 2455 4573 2464 4607
rect 2412 4564 2464 4573
rect 6920 4700 6972 4752
rect 3424 4675 3476 4684
rect 3424 4641 3433 4675
rect 3433 4641 3467 4675
rect 3467 4641 3476 4675
rect 3424 4632 3476 4641
rect 4804 4632 4856 4684
rect 5080 4632 5132 4684
rect 8300 4675 8352 4684
rect 8300 4641 8309 4675
rect 8309 4641 8343 4675
rect 8343 4641 8352 4675
rect 8300 4632 8352 4641
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2412 4428 2464 4480
rect 2688 4428 2740 4480
rect 3056 4496 3108 4548
rect 3700 4496 3752 4548
rect 5172 4564 5224 4616
rect 5356 4564 5408 4616
rect 3240 4471 3292 4480
rect 3240 4437 3249 4471
rect 3249 4437 3283 4471
rect 3283 4437 3292 4471
rect 3240 4428 3292 4437
rect 3608 4428 3660 4480
rect 3884 4428 3936 4480
rect 4160 4471 4212 4480
rect 4160 4437 4169 4471
rect 4169 4437 4203 4471
rect 4203 4437 4212 4471
rect 4160 4428 4212 4437
rect 6552 4496 6604 4548
rect 10140 4700 10192 4752
rect 10324 4743 10376 4752
rect 10324 4709 10333 4743
rect 10333 4709 10367 4743
rect 10367 4709 10376 4743
rect 10324 4700 10376 4709
rect 10600 4700 10652 4752
rect 9128 4632 9180 4684
rect 9312 4675 9364 4684
rect 9312 4641 9321 4675
rect 9321 4641 9355 4675
rect 9355 4641 9364 4675
rect 9312 4632 9364 4641
rect 9864 4632 9916 4684
rect 10416 4632 10468 4684
rect 10692 4632 10744 4684
rect 8944 4607 8996 4616
rect 8944 4573 8953 4607
rect 8953 4573 8987 4607
rect 8987 4573 8996 4607
rect 8944 4564 8996 4573
rect 5172 4428 5224 4480
rect 7288 4428 7340 4480
rect 8208 4496 8260 4548
rect 8392 4428 8444 4480
rect 8852 4428 8904 4480
rect 9312 4496 9364 4548
rect 9772 4496 9824 4548
rect 9864 4539 9916 4548
rect 9864 4505 9873 4539
rect 9873 4505 9907 4539
rect 9907 4505 9916 4539
rect 10232 4564 10284 4616
rect 11520 4700 11572 4752
rect 11336 4632 11388 4684
rect 13544 4675 13596 4684
rect 13544 4641 13553 4675
rect 13553 4641 13587 4675
rect 13587 4641 13596 4675
rect 13544 4632 13596 4641
rect 16304 4632 16356 4684
rect 11520 4564 11572 4616
rect 9864 4496 9916 4505
rect 11796 4496 11848 4548
rect 13820 4564 13872 4616
rect 15384 4564 15436 4616
rect 15936 4607 15988 4616
rect 15936 4573 15945 4607
rect 15945 4573 15979 4607
rect 15979 4573 15988 4607
rect 15936 4564 15988 4573
rect 17960 4768 18012 4820
rect 17040 4632 17092 4684
rect 18512 4768 18564 4820
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 10876 4428 10928 4480
rect 11888 4428 11940 4480
rect 12348 4428 12400 4480
rect 12532 4471 12584 4480
rect 12532 4437 12541 4471
rect 12541 4437 12575 4471
rect 12575 4437 12584 4471
rect 12532 4428 12584 4437
rect 13360 4471 13412 4480
rect 13360 4437 13369 4471
rect 13369 4437 13403 4471
rect 13403 4437 13412 4471
rect 13360 4428 13412 4437
rect 13912 4471 13964 4480
rect 13912 4437 13921 4471
rect 13921 4437 13955 4471
rect 13955 4437 13964 4471
rect 13912 4428 13964 4437
rect 14740 4496 14792 4548
rect 15292 4428 15344 4480
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 16212 4428 16264 4480
rect 17960 4496 18012 4548
rect 18420 4496 18472 4548
rect 19616 4496 19668 4548
rect 17408 4471 17460 4480
rect 17408 4437 17417 4471
rect 17417 4437 17451 4471
rect 17451 4437 17460 4471
rect 17408 4428 17460 4437
rect 17868 4471 17920 4480
rect 17868 4437 17877 4471
rect 17877 4437 17911 4471
rect 17911 4437 17920 4471
rect 17868 4428 17920 4437
rect 5398 4326 5450 4378
rect 5462 4326 5514 4378
rect 5526 4326 5578 4378
rect 5590 4326 5642 4378
rect 5654 4326 5706 4378
rect 9846 4326 9898 4378
rect 9910 4326 9962 4378
rect 9974 4326 10026 4378
rect 10038 4326 10090 4378
rect 10102 4326 10154 4378
rect 14294 4326 14346 4378
rect 14358 4326 14410 4378
rect 14422 4326 14474 4378
rect 14486 4326 14538 4378
rect 14550 4326 14602 4378
rect 2964 4224 3016 4276
rect 4068 4224 4120 4276
rect 5080 4267 5132 4276
rect 5080 4233 5089 4267
rect 5089 4233 5123 4267
rect 5123 4233 5132 4267
rect 5080 4224 5132 4233
rect 4068 4131 4120 4140
rect 4436 4156 4488 4208
rect 4068 4097 4097 4131
rect 4097 4097 4120 4131
rect 4068 4088 4120 4097
rect 2780 4063 2832 4072
rect 2780 4029 2789 4063
rect 2789 4029 2823 4063
rect 2823 4029 2832 4063
rect 2780 4020 2832 4029
rect 4528 4131 4580 4140
rect 4528 4097 4537 4131
rect 4537 4097 4571 4131
rect 4571 4097 4580 4131
rect 4528 4088 4580 4097
rect 4620 4088 4672 4140
rect 5172 4156 5224 4208
rect 9220 4224 9272 4276
rect 9496 4224 9548 4276
rect 9772 4224 9824 4276
rect 10232 4224 10284 4276
rect 2412 3884 2464 3936
rect 2596 3884 2648 3936
rect 3700 3884 3752 3936
rect 4528 3884 4580 3936
rect 4804 3884 4856 3936
rect 6736 4088 6788 4140
rect 8024 4088 8076 4140
rect 8944 4156 8996 4208
rect 9312 4156 9364 4208
rect 9956 4156 10008 4208
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 5908 4063 5960 4072
rect 5908 4029 5917 4063
rect 5917 4029 5951 4063
rect 5951 4029 5960 4063
rect 5908 4020 5960 4029
rect 6092 4063 6144 4072
rect 6092 4029 6101 4063
rect 6101 4029 6135 4063
rect 6135 4029 6144 4063
rect 6092 4020 6144 4029
rect 8300 4088 8352 4140
rect 8484 4131 8536 4140
rect 8484 4097 8518 4131
rect 8518 4097 8536 4131
rect 8484 4088 8536 4097
rect 10232 4088 10284 4140
rect 6000 3884 6052 3936
rect 6368 3927 6420 3936
rect 6368 3893 6377 3927
rect 6377 3893 6411 3927
rect 6411 3893 6420 3927
rect 6368 3884 6420 3893
rect 9220 3884 9272 3936
rect 9956 4063 10008 4072
rect 9956 4029 9965 4063
rect 9965 4029 9999 4063
rect 9999 4029 10008 4063
rect 9956 4020 10008 4029
rect 10140 4020 10192 4072
rect 11520 4156 11572 4208
rect 11888 4199 11940 4208
rect 11888 4165 11897 4199
rect 11897 4165 11931 4199
rect 11931 4165 11940 4199
rect 11888 4156 11940 4165
rect 12532 4224 12584 4276
rect 13820 4267 13872 4276
rect 13820 4233 13829 4267
rect 13829 4233 13863 4267
rect 13863 4233 13872 4267
rect 13820 4224 13872 4233
rect 14004 4224 14056 4276
rect 12900 4156 12952 4208
rect 14096 4156 14148 4208
rect 11336 4088 11388 4140
rect 11152 4063 11204 4072
rect 11152 4029 11161 4063
rect 11161 4029 11195 4063
rect 11195 4029 11204 4063
rect 11152 4020 11204 4029
rect 9956 3884 10008 3936
rect 10876 3884 10928 3936
rect 11612 4088 11664 4140
rect 11520 4020 11572 4072
rect 12624 4088 12676 4140
rect 13452 4131 13504 4140
rect 13452 4097 13461 4131
rect 13461 4097 13495 4131
rect 13495 4097 13504 4131
rect 13452 4088 13504 4097
rect 13728 4088 13780 4140
rect 15384 4156 15436 4208
rect 17592 4224 17644 4276
rect 18052 4224 18104 4276
rect 15108 4088 15160 4140
rect 16304 4088 16356 4140
rect 18696 4156 18748 4208
rect 17316 4131 17368 4140
rect 17316 4097 17325 4131
rect 17325 4097 17359 4131
rect 17359 4097 17368 4131
rect 17316 4088 17368 4097
rect 18236 4131 18288 4140
rect 13084 4063 13136 4072
rect 13084 4029 13093 4063
rect 13093 4029 13127 4063
rect 13127 4029 13136 4063
rect 13084 4020 13136 4029
rect 13544 4020 13596 4072
rect 14004 4020 14056 4072
rect 14740 4020 14792 4072
rect 17224 4020 17276 4072
rect 17776 4020 17828 4072
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 19524 4020 19576 4072
rect 12808 3952 12860 4004
rect 13820 3952 13872 4004
rect 11796 3884 11848 3936
rect 12900 3884 12952 3936
rect 15384 3952 15436 4004
rect 16396 3952 16448 4004
rect 18604 3952 18656 4004
rect 15016 3927 15068 3936
rect 15016 3893 15025 3927
rect 15025 3893 15059 3927
rect 15059 3893 15068 3927
rect 15016 3884 15068 3893
rect 17684 3884 17736 3936
rect 18144 3884 18196 3936
rect 3174 3782 3226 3834
rect 3238 3782 3290 3834
rect 3302 3782 3354 3834
rect 3366 3782 3418 3834
rect 3430 3782 3482 3834
rect 7622 3782 7674 3834
rect 7686 3782 7738 3834
rect 7750 3782 7802 3834
rect 7814 3782 7866 3834
rect 7878 3782 7930 3834
rect 12070 3782 12122 3834
rect 12134 3782 12186 3834
rect 12198 3782 12250 3834
rect 12262 3782 12314 3834
rect 12326 3782 12378 3834
rect 16518 3782 16570 3834
rect 16582 3782 16634 3834
rect 16646 3782 16698 3834
rect 16710 3782 16762 3834
rect 16774 3782 16826 3834
rect 1584 3680 1636 3732
rect 3608 3612 3660 3664
rect 6552 3655 6604 3664
rect 6552 3621 6561 3655
rect 6561 3621 6595 3655
rect 6595 3621 6604 3655
rect 6552 3612 6604 3621
rect 2504 3587 2556 3596
rect 2504 3553 2513 3587
rect 2513 3553 2547 3587
rect 2547 3553 2556 3587
rect 2504 3544 2556 3553
rect 3976 3587 4028 3596
rect 3976 3553 3985 3587
rect 3985 3553 4019 3587
rect 4019 3553 4028 3587
rect 3976 3544 4028 3553
rect 4436 3544 4488 3596
rect 6092 3544 6144 3596
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 4712 3476 4764 3528
rect 1308 3408 1360 3460
rect 4436 3408 4488 3460
rect 1492 3340 1544 3392
rect 1952 3383 2004 3392
rect 1952 3349 1961 3383
rect 1961 3349 1995 3383
rect 1995 3349 2004 3383
rect 1952 3340 2004 3349
rect 2320 3383 2372 3392
rect 2320 3349 2329 3383
rect 2329 3349 2363 3383
rect 2363 3349 2372 3383
rect 2320 3340 2372 3349
rect 2504 3340 2556 3392
rect 3148 3383 3200 3392
rect 3148 3349 3157 3383
rect 3157 3349 3191 3383
rect 3191 3349 3200 3383
rect 3148 3340 3200 3349
rect 3516 3340 3568 3392
rect 3792 3340 3844 3392
rect 3976 3340 4028 3392
rect 4252 3340 4304 3392
rect 5080 3408 5132 3460
rect 7380 3476 7432 3528
rect 8484 3680 8536 3732
rect 10784 3680 10836 3732
rect 10968 3680 11020 3732
rect 8208 3612 8260 3664
rect 8116 3544 8168 3596
rect 8300 3544 8352 3596
rect 11796 3680 11848 3732
rect 12164 3612 12216 3664
rect 12900 3612 12952 3664
rect 10416 3519 10468 3528
rect 10416 3485 10425 3519
rect 10425 3485 10459 3519
rect 10459 3485 10468 3519
rect 10416 3476 10468 3485
rect 11244 3476 11296 3528
rect 12164 3476 12216 3528
rect 12624 3519 12676 3528
rect 12624 3485 12633 3519
rect 12633 3485 12667 3519
rect 12667 3485 12676 3519
rect 12624 3476 12676 3485
rect 13084 3680 13136 3732
rect 13360 3680 13412 3732
rect 14648 3680 14700 3732
rect 15476 3680 15528 3732
rect 15292 3612 15344 3664
rect 14740 3587 14792 3596
rect 14740 3553 14749 3587
rect 14749 3553 14783 3587
rect 14783 3553 14792 3587
rect 14740 3544 14792 3553
rect 15384 3544 15436 3596
rect 15660 3544 15712 3596
rect 17408 3680 17460 3732
rect 17868 3680 17920 3732
rect 18972 3680 19024 3732
rect 17224 3612 17276 3664
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 15200 3476 15252 3528
rect 17132 3476 17184 3528
rect 17224 3519 17276 3528
rect 17224 3485 17233 3519
rect 17233 3485 17267 3519
rect 17267 3485 17276 3519
rect 17224 3476 17276 3485
rect 9220 3451 9272 3460
rect 6092 3340 6144 3392
rect 9220 3417 9254 3451
rect 9254 3417 9272 3451
rect 9220 3408 9272 3417
rect 9680 3408 9732 3460
rect 10140 3408 10192 3460
rect 10232 3408 10284 3460
rect 7564 3340 7616 3392
rect 8484 3340 8536 3392
rect 9312 3340 9364 3392
rect 10784 3340 10836 3392
rect 13728 3408 13780 3460
rect 13176 3340 13228 3392
rect 13360 3383 13412 3392
rect 13360 3349 13369 3383
rect 13369 3349 13403 3383
rect 13403 3349 13412 3383
rect 13360 3340 13412 3349
rect 13544 3340 13596 3392
rect 16120 3408 16172 3460
rect 16488 3408 16540 3460
rect 16856 3408 16908 3460
rect 19156 3612 19208 3664
rect 17776 3544 17828 3596
rect 18052 3519 18104 3528
rect 18052 3485 18061 3519
rect 18061 3485 18095 3519
rect 18095 3485 18104 3519
rect 18052 3476 18104 3485
rect 18328 3408 18380 3460
rect 15292 3383 15344 3392
rect 15292 3349 15301 3383
rect 15301 3349 15335 3383
rect 15335 3349 15344 3383
rect 15292 3340 15344 3349
rect 15752 3340 15804 3392
rect 15936 3383 15988 3392
rect 15936 3349 15945 3383
rect 15945 3349 15979 3383
rect 15979 3349 15988 3383
rect 15936 3340 15988 3349
rect 16396 3383 16448 3392
rect 16396 3349 16405 3383
rect 16405 3349 16439 3383
rect 16439 3349 16448 3383
rect 16396 3340 16448 3349
rect 17592 3340 17644 3392
rect 5398 3238 5450 3290
rect 5462 3238 5514 3290
rect 5526 3238 5578 3290
rect 5590 3238 5642 3290
rect 5654 3238 5706 3290
rect 9846 3238 9898 3290
rect 9910 3238 9962 3290
rect 9974 3238 10026 3290
rect 10038 3238 10090 3290
rect 10102 3238 10154 3290
rect 14294 3238 14346 3290
rect 14358 3238 14410 3290
rect 14422 3238 14474 3290
rect 14486 3238 14538 3290
rect 14550 3238 14602 3290
rect 1676 3136 1728 3188
rect 1952 3179 2004 3188
rect 1952 3145 1961 3179
rect 1961 3145 1995 3179
rect 1995 3145 2004 3179
rect 1952 3136 2004 3145
rect 2504 3136 2556 3188
rect 3148 3136 3200 3188
rect 6736 3179 6788 3188
rect 2780 3111 2832 3120
rect 2780 3077 2789 3111
rect 2789 3077 2823 3111
rect 2823 3077 2832 3111
rect 2780 3068 2832 3077
rect 4344 3111 4396 3120
rect 4344 3077 4353 3111
rect 4353 3077 4387 3111
rect 4387 3077 4396 3111
rect 4344 3068 4396 3077
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 1308 2932 1360 2984
rect 4068 3000 4120 3052
rect 4712 3000 4764 3052
rect 4896 3043 4948 3052
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 2136 2932 2188 2984
rect 3976 2932 4028 2984
rect 5816 3068 5868 3120
rect 5264 3000 5316 3052
rect 5448 2932 5500 2984
rect 5816 2975 5868 2984
rect 5816 2941 5825 2975
rect 5825 2941 5859 2975
rect 5859 2941 5868 2975
rect 5816 2932 5868 2941
rect 6000 2975 6052 2984
rect 6000 2941 6009 2975
rect 6009 2941 6043 2975
rect 6043 2941 6052 2975
rect 6000 2932 6052 2941
rect 2228 2864 2280 2916
rect 2964 2864 3016 2916
rect 1216 2796 1268 2848
rect 2136 2796 2188 2848
rect 2504 2796 2556 2848
rect 4068 2796 4120 2848
rect 4528 2839 4580 2848
rect 4528 2805 4537 2839
rect 4537 2805 4571 2839
rect 4571 2805 4580 2839
rect 4528 2796 4580 2805
rect 4620 2796 4672 2848
rect 5448 2796 5500 2848
rect 6000 2796 6052 2848
rect 6736 3145 6745 3179
rect 6745 3145 6779 3179
rect 6779 3145 6788 3179
rect 6736 3136 6788 3145
rect 6920 3136 6972 3188
rect 7196 3136 7248 3188
rect 8300 3179 8352 3188
rect 8300 3145 8309 3179
rect 8309 3145 8343 3179
rect 8343 3145 8352 3179
rect 8300 3136 8352 3145
rect 8484 3136 8536 3188
rect 9404 3136 9456 3188
rect 10324 3136 10376 3188
rect 10876 3179 10928 3188
rect 10876 3145 10885 3179
rect 10885 3145 10919 3179
rect 10919 3145 10928 3179
rect 10876 3136 10928 3145
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 11704 3136 11756 3188
rect 13820 3136 13872 3188
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 14188 3136 14240 3188
rect 15384 3179 15436 3188
rect 9588 3111 9640 3120
rect 7012 3000 7064 3052
rect 7196 2975 7248 2984
rect 7196 2941 7205 2975
rect 7205 2941 7239 2975
rect 7239 2941 7248 2975
rect 7196 2932 7248 2941
rect 7380 2975 7432 2984
rect 7380 2941 7389 2975
rect 7389 2941 7423 2975
rect 7423 2941 7432 2975
rect 7380 2932 7432 2941
rect 9588 3077 9597 3111
rect 9597 3077 9631 3111
rect 9631 3077 9640 3111
rect 9588 3068 9640 3077
rect 7932 3000 7984 3052
rect 10600 3068 10652 3120
rect 10692 3068 10744 3120
rect 6644 2864 6696 2916
rect 7840 2932 7892 2984
rect 8484 2932 8536 2984
rect 10508 3000 10560 3052
rect 10784 3000 10836 3052
rect 12532 3043 12584 3052
rect 10968 2975 11020 2984
rect 7196 2796 7248 2848
rect 8254 2864 8306 2916
rect 10508 2907 10560 2916
rect 10508 2873 10517 2907
rect 10517 2873 10551 2907
rect 10551 2873 10560 2907
rect 10508 2864 10560 2873
rect 10968 2941 10977 2975
rect 10977 2941 11011 2975
rect 11011 2941 11020 2975
rect 10968 2932 11020 2941
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 14740 3068 14792 3120
rect 15384 3145 15393 3179
rect 15393 3145 15427 3179
rect 15427 3145 15436 3179
rect 15384 3136 15436 3145
rect 15568 3136 15620 3188
rect 16396 3136 16448 3188
rect 16488 3136 16540 3188
rect 17960 3179 18012 3188
rect 17960 3145 17969 3179
rect 17969 3145 18003 3179
rect 18003 3145 18012 3179
rect 17960 3136 18012 3145
rect 18328 3136 18380 3188
rect 19340 3136 19392 3188
rect 16028 3068 16080 3120
rect 17040 3111 17092 3120
rect 17040 3077 17049 3111
rect 17049 3077 17083 3111
rect 17083 3077 17092 3111
rect 17040 3068 17092 3077
rect 18420 3111 18472 3120
rect 18420 3077 18429 3111
rect 18429 3077 18463 3111
rect 18463 3077 18472 3111
rect 18420 3068 18472 3077
rect 13912 3000 13964 3052
rect 14464 3043 14516 3052
rect 14464 3009 14473 3043
rect 14473 3009 14507 3043
rect 14507 3009 14516 3043
rect 14464 3000 14516 3009
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15292 3000 15344 3052
rect 15844 3000 15896 3052
rect 16120 3000 16172 3052
rect 16672 3043 16724 3052
rect 16672 3009 16681 3043
rect 16681 3009 16715 3043
rect 16715 3009 16724 3043
rect 16672 3000 16724 3009
rect 16764 3000 16816 3052
rect 19892 3000 19944 3052
rect 12072 2975 12124 2984
rect 12072 2941 12081 2975
rect 12081 2941 12115 2975
rect 12115 2941 12124 2975
rect 12072 2932 12124 2941
rect 12164 2932 12216 2984
rect 13728 2932 13780 2984
rect 14372 2932 14424 2984
rect 14648 2975 14700 2984
rect 14648 2941 14657 2975
rect 14657 2941 14691 2975
rect 14691 2941 14700 2975
rect 14648 2932 14700 2941
rect 15016 2932 15068 2984
rect 17776 2932 17828 2984
rect 17960 2932 18012 2984
rect 18512 2932 18564 2984
rect 9128 2796 9180 2848
rect 9404 2796 9456 2848
rect 11612 2864 11664 2916
rect 12900 2796 12952 2848
rect 13268 2796 13320 2848
rect 19432 2864 19484 2916
rect 14648 2796 14700 2848
rect 14924 2796 14976 2848
rect 17960 2796 18012 2848
rect 18236 2839 18288 2848
rect 18236 2805 18245 2839
rect 18245 2805 18279 2839
rect 18279 2805 18288 2839
rect 18236 2796 18288 2805
rect 3174 2694 3226 2746
rect 3238 2694 3290 2746
rect 3302 2694 3354 2746
rect 3366 2694 3418 2746
rect 3430 2694 3482 2746
rect 7622 2694 7674 2746
rect 7686 2694 7738 2746
rect 7750 2694 7802 2746
rect 7814 2694 7866 2746
rect 7878 2694 7930 2746
rect 12070 2694 12122 2746
rect 12134 2694 12186 2746
rect 12198 2694 12250 2746
rect 12262 2694 12314 2746
rect 12326 2694 12378 2746
rect 16518 2694 16570 2746
rect 16582 2694 16634 2746
rect 16646 2694 16698 2746
rect 16710 2694 16762 2746
rect 16774 2694 16826 2746
rect 2596 2592 2648 2644
rect 2964 2592 3016 2644
rect 3884 2592 3936 2644
rect 4068 2592 4120 2644
rect 5908 2592 5960 2644
rect 9128 2592 9180 2644
rect 10416 2592 10468 2644
rect 10692 2635 10744 2644
rect 10692 2601 10701 2635
rect 10701 2601 10735 2635
rect 10735 2601 10744 2635
rect 10692 2592 10744 2601
rect 13912 2592 13964 2644
rect 14188 2592 14240 2644
rect 14372 2592 14424 2644
rect 3424 2567 3476 2576
rect 3424 2533 3433 2567
rect 3433 2533 3467 2567
rect 3467 2533 3476 2567
rect 6184 2567 6236 2576
rect 3424 2524 3476 2533
rect 6184 2533 6193 2567
rect 6193 2533 6227 2567
rect 6227 2533 6236 2567
rect 6184 2524 6236 2533
rect 7196 2524 7248 2576
rect 8208 2524 8260 2576
rect 2504 2456 2556 2508
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 2872 2456 2924 2508
rect 3148 2456 3200 2508
rect 4436 2456 4488 2508
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 3792 2388 3844 2440
rect 4252 2388 4304 2440
rect 4988 2431 5040 2440
rect 1584 2295 1636 2304
rect 1584 2261 1593 2295
rect 1593 2261 1627 2295
rect 1627 2261 1636 2295
rect 1584 2252 1636 2261
rect 2228 2295 2280 2304
rect 2228 2261 2237 2295
rect 2237 2261 2271 2295
rect 2271 2261 2280 2295
rect 2228 2252 2280 2261
rect 4344 2320 4396 2372
rect 4988 2397 4997 2431
rect 4997 2397 5031 2431
rect 5031 2397 5040 2431
rect 4988 2388 5040 2397
rect 5448 2456 5500 2508
rect 6092 2456 6144 2508
rect 6368 2456 6420 2508
rect 6828 2456 6880 2508
rect 7380 2456 7432 2508
rect 8116 2499 8168 2508
rect 8116 2465 8125 2499
rect 8125 2465 8159 2499
rect 8159 2465 8168 2499
rect 8116 2456 8168 2465
rect 9680 2524 9732 2576
rect 10508 2524 10560 2576
rect 10968 2524 11020 2576
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 9220 2499 9272 2508
rect 9220 2465 9229 2499
rect 9229 2465 9263 2499
rect 9263 2465 9272 2499
rect 9220 2456 9272 2465
rect 9404 2499 9456 2508
rect 9404 2465 9413 2499
rect 9413 2465 9447 2499
rect 9447 2465 9456 2499
rect 9404 2456 9456 2465
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 9036 2388 9088 2440
rect 6460 2295 6512 2304
rect 6460 2261 6469 2295
rect 6469 2261 6503 2295
rect 6503 2261 6512 2295
rect 6460 2252 6512 2261
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 7104 2295 7156 2304
rect 7104 2261 7113 2295
rect 7113 2261 7147 2295
rect 7147 2261 7156 2295
rect 9404 2320 9456 2372
rect 14740 2524 14792 2576
rect 18052 2567 18104 2576
rect 18052 2533 18061 2567
rect 18061 2533 18095 2567
rect 18095 2533 18104 2567
rect 18052 2524 18104 2533
rect 12072 2499 12124 2508
rect 12072 2465 12081 2499
rect 12081 2465 12115 2499
rect 12115 2465 12124 2499
rect 12072 2456 12124 2465
rect 14372 2456 14424 2508
rect 9772 2388 9824 2440
rect 10416 2388 10468 2440
rect 11980 2388 12032 2440
rect 12256 2388 12308 2440
rect 7104 2252 7156 2261
rect 7932 2295 7984 2304
rect 7932 2261 7941 2295
rect 7941 2261 7975 2295
rect 7975 2261 7984 2295
rect 7932 2252 7984 2261
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 10508 2252 10560 2304
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 11152 2295 11204 2304
rect 11152 2261 11161 2295
rect 11161 2261 11195 2295
rect 11195 2261 11204 2295
rect 11152 2252 11204 2261
rect 12348 2320 12400 2372
rect 12900 2320 12952 2372
rect 11980 2295 12032 2304
rect 11980 2261 11989 2295
rect 11989 2261 12023 2295
rect 12023 2261 12032 2295
rect 11980 2252 12032 2261
rect 12624 2295 12676 2304
rect 12624 2261 12633 2295
rect 12633 2261 12667 2295
rect 12667 2261 12676 2295
rect 12624 2252 12676 2261
rect 12716 2295 12768 2304
rect 12716 2261 12725 2295
rect 12725 2261 12759 2295
rect 12759 2261 12768 2295
rect 12716 2252 12768 2261
rect 14924 2431 14976 2440
rect 14924 2397 14933 2431
rect 14933 2397 14967 2431
rect 14967 2397 14976 2431
rect 14924 2388 14976 2397
rect 15660 2431 15712 2440
rect 15660 2397 15669 2431
rect 15669 2397 15703 2431
rect 15703 2397 15712 2431
rect 15660 2388 15712 2397
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 17408 2431 17460 2440
rect 17408 2397 17417 2431
rect 17417 2397 17451 2431
rect 17451 2397 17460 2431
rect 17408 2388 17460 2397
rect 17960 2388 18012 2440
rect 16396 2295 16448 2304
rect 16396 2261 16405 2295
rect 16405 2261 16439 2295
rect 16439 2261 16448 2295
rect 16396 2252 16448 2261
rect 17316 2295 17368 2304
rect 17316 2261 17325 2295
rect 17325 2261 17359 2295
rect 17359 2261 17368 2295
rect 17316 2252 17368 2261
rect 18144 2252 18196 2304
rect 5398 2150 5450 2202
rect 5462 2150 5514 2202
rect 5526 2150 5578 2202
rect 5590 2150 5642 2202
rect 5654 2150 5706 2202
rect 9846 2150 9898 2202
rect 9910 2150 9962 2202
rect 9974 2150 10026 2202
rect 10038 2150 10090 2202
rect 10102 2150 10154 2202
rect 14294 2150 14346 2202
rect 14358 2150 14410 2202
rect 14422 2150 14474 2202
rect 14486 2150 14538 2202
rect 14550 2150 14602 2202
rect 4068 2048 4120 2100
rect 8668 2048 8720 2100
rect 8944 2048 8996 2100
rect 2228 1980 2280 2032
rect 4620 1980 4672 2032
rect 6092 1980 6144 2032
rect 10876 2048 10928 2100
rect 14924 2048 14976 2100
rect 3056 1912 3108 1964
rect 5172 1912 5224 1964
rect 6828 1912 6880 1964
rect 2412 1844 2464 1896
rect 2044 1776 2096 1828
rect 9404 1776 9456 1828
rect 4068 1708 4120 1760
rect 8392 1708 8444 1760
rect 11152 1980 11204 2032
rect 12532 1980 12584 2032
rect 16396 1980 16448 2032
rect 12348 1912 12400 1964
rect 18696 1912 18748 1964
rect 17408 1844 17460 1896
rect 16672 1776 16724 1828
rect 12072 1708 12124 1760
rect 12164 1708 12216 1760
rect 18144 1708 18196 1760
rect 7012 1640 7064 1692
rect 12624 1640 12676 1692
rect 15752 1640 15804 1692
rect 2320 1572 2372 1624
rect 3516 1572 3568 1624
rect 7932 1572 7984 1624
rect 12256 1572 12308 1624
rect 7104 1504 7156 1556
rect 12716 1572 12768 1624
rect 11244 1436 11296 1488
rect 12808 1436 12860 1488
rect 4068 1300 4120 1352
rect 10968 1300 11020 1352
rect 3608 1232 3660 1284
rect 11980 1300 12032 1352
rect 13636 1300 13688 1352
rect 15200 1300 15252 1352
rect 11428 1232 11480 1284
rect 15936 1232 15988 1284
rect 11060 1164 11112 1216
rect 15844 1164 15896 1216
rect 3424 824 3476 876
rect 8852 824 8904 876
rect 3700 620 3752 672
rect 6460 620 6512 672
rect 1584 8 1636 60
rect 15660 8 15712 60
<< metal2 >>
rect 1950 16538 2006 17200
rect 3790 16960 3846 16969
rect 3790 16895 3846 16904
rect 1950 16510 2268 16538
rect 1950 16400 2006 16510
rect 2134 16008 2190 16017
rect 2134 15943 2190 15952
rect 756 15496 808 15502
rect 756 15438 808 15444
rect 20 15428 72 15434
rect 20 15370 72 15376
rect 32 6866 60 15370
rect 768 7818 796 15438
rect 2044 15292 2096 15298
rect 2044 15234 2096 15240
rect 1490 14920 1546 14929
rect 1490 14855 1546 14864
rect 1124 13932 1176 13938
rect 1124 13874 1176 13880
rect 848 13524 900 13530
rect 848 13466 900 13472
rect 860 7959 888 13466
rect 1136 13025 1164 13874
rect 1216 13456 1268 13462
rect 1216 13398 1268 13404
rect 1122 13016 1178 13025
rect 1122 12951 1178 12960
rect 938 12608 994 12617
rect 938 12543 994 12552
rect 846 7950 902 7959
rect 846 7885 902 7894
rect 756 7812 808 7818
rect 756 7754 808 7760
rect 952 7546 980 12543
rect 1030 12472 1086 12481
rect 1030 12407 1086 12416
rect 940 7540 992 7546
rect 940 7482 992 7488
rect 1044 7426 1072 12407
rect 1124 11688 1176 11694
rect 1124 11630 1176 11636
rect 1136 7449 1164 11630
rect 860 7398 1072 7426
rect 1122 7440 1178 7449
rect 388 7268 440 7274
rect 388 7210 440 7216
rect 20 6860 72 6866
rect 20 6802 72 6808
rect 400 800 428 7210
rect 860 7188 888 7398
rect 1122 7375 1178 7384
rect 860 7160 1072 7188
rect 940 6860 992 6866
rect 940 6802 992 6808
rect 952 6769 980 6802
rect 938 6760 994 6769
rect 938 6695 994 6704
rect 1044 3369 1072 7160
rect 1122 6216 1178 6225
rect 1122 6151 1178 6160
rect 1136 4729 1164 6151
rect 1122 4720 1178 4729
rect 1122 4655 1178 4664
rect 1030 3360 1086 3369
rect 1030 3295 1086 3304
rect 1228 2854 1256 13398
rect 1308 13252 1360 13258
rect 1308 13194 1360 13200
rect 1320 9489 1348 13194
rect 1504 12782 1532 14855
rect 1950 14512 2006 14521
rect 1950 14447 1952 14456
rect 2004 14447 2006 14456
rect 1952 14418 2004 14424
rect 1584 14000 1636 14006
rect 1584 13942 1636 13948
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 10810 1440 11494
rect 1400 10804 1452 10810
rect 1400 10746 1452 10752
rect 1504 10690 1532 12718
rect 1596 10810 1624 13942
rect 2056 13870 2084 15234
rect 2148 15230 2176 15943
rect 2136 15224 2188 15230
rect 2136 15166 2188 15172
rect 2148 14414 2176 15166
rect 2240 14550 2268 16510
rect 2688 15632 2740 15638
rect 2688 15574 2740 15580
rect 2320 15360 2372 15366
rect 2320 15302 2372 15308
rect 2228 14544 2280 14550
rect 2228 14486 2280 14492
rect 2136 14408 2188 14414
rect 2136 14350 2188 14356
rect 2226 14240 2282 14249
rect 2226 14175 2282 14184
rect 2240 13938 2268 14175
rect 2228 13932 2280 13938
rect 2228 13874 2280 13880
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 1858 13424 1914 13433
rect 1858 13359 1914 13368
rect 1768 12912 1820 12918
rect 1768 12854 1820 12860
rect 1674 12200 1730 12209
rect 1674 12135 1730 12144
rect 1688 11218 1716 12135
rect 1676 11212 1728 11218
rect 1676 11154 1728 11160
rect 1780 11150 1808 12854
rect 1768 11144 1820 11150
rect 1768 11086 1820 11092
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1504 10662 1624 10690
rect 1490 10024 1546 10033
rect 1490 9959 1546 9968
rect 1400 9512 1452 9518
rect 1306 9480 1362 9489
rect 1400 9454 1452 9460
rect 1306 9415 1362 9424
rect 1308 8900 1360 8906
rect 1308 8842 1360 8848
rect 1320 3466 1348 8842
rect 1412 8809 1440 9454
rect 1504 8974 1532 9959
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1492 8288 1544 8294
rect 1492 8230 1544 8236
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1412 4593 1440 7482
rect 1504 7290 1532 8230
rect 1596 7750 1624 10662
rect 1872 9994 1900 13359
rect 1952 12232 2004 12238
rect 1952 12174 2004 12180
rect 1964 11257 1992 12174
rect 2056 11830 2084 13806
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2044 11824 2096 11830
rect 2148 11801 2176 13262
rect 2332 13138 2360 15302
rect 2504 15088 2556 15094
rect 2504 15030 2556 15036
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 13977 2452 14214
rect 2410 13968 2466 13977
rect 2410 13903 2466 13912
rect 2516 13394 2544 15030
rect 2596 14272 2648 14278
rect 2596 14214 2648 14220
rect 2504 13388 2556 13394
rect 2504 13330 2556 13336
rect 2410 13288 2466 13297
rect 2410 13223 2466 13232
rect 2424 13190 2452 13223
rect 2240 13110 2360 13138
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2044 11766 2096 11772
rect 2134 11792 2190 11801
rect 2240 11762 2268 13110
rect 2320 12980 2372 12986
rect 2320 12922 2372 12928
rect 2134 11727 2190 11736
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2136 11688 2188 11694
rect 2136 11630 2188 11636
rect 2044 11620 2096 11626
rect 2044 11562 2096 11568
rect 2056 11286 2084 11562
rect 2044 11280 2096 11286
rect 1950 11248 2006 11257
rect 2044 11222 2096 11228
rect 1950 11183 2006 11192
rect 2148 11082 2176 11630
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 1964 10033 1992 10202
rect 1950 10024 2006 10033
rect 1860 9988 1912 9994
rect 1950 9959 2006 9968
rect 1860 9930 1912 9936
rect 1872 9353 1900 9930
rect 1950 9616 2006 9625
rect 1950 9551 1952 9560
rect 2004 9551 2006 9560
rect 1952 9522 2004 9528
rect 1952 9444 2004 9450
rect 1952 9386 2004 9392
rect 1858 9344 1914 9353
rect 1858 9279 1914 9288
rect 1768 9104 1820 9110
rect 1674 9072 1730 9081
rect 1768 9046 1820 9052
rect 1674 9007 1676 9016
rect 1728 9007 1730 9016
rect 1676 8978 1728 8984
rect 1780 8922 1808 9046
rect 1688 8894 1808 8922
rect 1688 8566 1716 8894
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1858 8800 1914 8809
rect 1676 8560 1728 8566
rect 1676 8502 1728 8508
rect 1780 8498 1808 8774
rect 1858 8735 1914 8744
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1768 8084 1820 8090
rect 1768 8026 1820 8032
rect 1676 8016 1728 8022
rect 1676 7958 1728 7964
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1688 7410 1716 7958
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1780 7342 1808 8026
rect 1768 7336 1820 7342
rect 1504 7262 1716 7290
rect 1768 7278 1820 7284
rect 1492 7200 1544 7206
rect 1492 7142 1544 7148
rect 1504 5137 1532 7142
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1596 5166 1624 6666
rect 1688 6322 1716 7262
rect 1676 6316 1728 6322
rect 1676 6258 1728 6264
rect 1780 6254 1808 7278
rect 1768 6248 1820 6254
rect 1768 6190 1820 6196
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1674 5672 1730 5681
rect 1674 5607 1676 5616
rect 1728 5607 1730 5616
rect 1676 5578 1728 5584
rect 1780 5409 1808 6054
rect 1766 5400 1822 5409
rect 1766 5335 1822 5344
rect 1676 5228 1728 5234
rect 1676 5170 1728 5176
rect 1584 5160 1636 5166
rect 1490 5128 1546 5137
rect 1584 5102 1636 5108
rect 1490 5063 1546 5072
rect 1688 4706 1716 5170
rect 1688 4678 1808 4706
rect 1676 4616 1728 4622
rect 1398 4584 1454 4593
rect 1676 4558 1728 4564
rect 1398 4519 1454 4528
rect 1584 4480 1636 4486
rect 1584 4422 1636 4428
rect 1596 3738 1624 4422
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1308 3460 1360 3466
rect 1308 3402 1360 3408
rect 1492 3392 1544 3398
rect 1492 3334 1544 3340
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1308 2984 1360 2990
rect 1412 2961 1440 2994
rect 1308 2926 1360 2932
rect 1398 2952 1454 2961
rect 1216 2848 1268 2854
rect 1216 2790 1268 2796
rect 1320 2258 1348 2926
rect 1398 2887 1454 2896
rect 1228 2230 1348 2258
rect 1228 800 1256 2230
rect 386 0 442 800
rect 1214 0 1270 800
rect 1504 241 1532 3334
rect 1688 3194 1716 4558
rect 1676 3188 1728 3194
rect 1676 3130 1728 3136
rect 1780 2961 1808 4678
rect 1872 3534 1900 8735
rect 1964 8022 1992 9386
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 1952 7880 2004 7886
rect 2056 7868 2084 10746
rect 2240 10713 2268 11698
rect 2226 10704 2282 10713
rect 2226 10639 2282 10648
rect 2226 10568 2282 10577
rect 2226 10503 2282 10512
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2148 9654 2176 9998
rect 2240 9761 2268 10503
rect 2226 9752 2282 9761
rect 2226 9687 2282 9696
rect 2136 9648 2188 9654
rect 2136 9590 2188 9596
rect 2240 9586 2268 9687
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2228 9376 2280 9382
rect 2228 9318 2280 9324
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2004 7840 2084 7868
rect 1952 7822 2004 7828
rect 1964 7478 1992 7822
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 1950 6760 2006 6769
rect 1950 6695 2006 6704
rect 1964 5710 1992 6695
rect 1952 5704 2004 5710
rect 1952 5646 2004 5652
rect 2056 5370 2084 7686
rect 2148 7546 2176 8842
rect 2240 8537 2268 9318
rect 2226 8528 2282 8537
rect 2226 8463 2282 8472
rect 2228 8288 2280 8294
rect 2332 8242 2360 12922
rect 2516 12345 2544 13330
rect 2608 13326 2636 14214
rect 2700 14006 2728 15574
rect 3804 15094 3832 16895
rect 4066 16688 4122 16697
rect 4066 16623 4122 16632
rect 3882 15328 3938 15337
rect 3882 15263 3938 15272
rect 3792 15088 3844 15094
rect 2778 15056 2834 15065
rect 3792 15030 3844 15036
rect 2778 14991 2834 15000
rect 2792 14618 2820 14991
rect 2872 14816 2924 14822
rect 2872 14758 2924 14764
rect 2780 14612 2832 14618
rect 2780 14554 2832 14560
rect 2884 14482 2912 14758
rect 3174 14716 3482 14736
rect 3174 14714 3180 14716
rect 3236 14714 3260 14716
rect 3316 14714 3340 14716
rect 3396 14714 3420 14716
rect 3476 14714 3482 14716
rect 3236 14662 3238 14714
rect 3418 14662 3420 14714
rect 3174 14660 3180 14662
rect 3236 14660 3260 14662
rect 3316 14660 3340 14662
rect 3396 14660 3420 14662
rect 3476 14660 3482 14662
rect 2962 14648 3018 14657
rect 3174 14640 3482 14660
rect 2962 14583 2964 14592
rect 3016 14583 3018 14592
rect 2964 14554 3016 14560
rect 2872 14476 2924 14482
rect 2872 14418 2924 14424
rect 3804 14414 3832 15030
rect 3896 14890 3924 15263
rect 4080 15026 4108 16623
rect 5906 16400 5962 17200
rect 9862 16538 9918 17200
rect 9862 16510 10456 16538
rect 9862 16400 9918 16510
rect 4342 16280 4398 16289
rect 4342 16215 4398 16224
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 3884 14884 3936 14890
rect 3884 14826 3936 14832
rect 3240 14408 3292 14414
rect 2778 14376 2834 14385
rect 3240 14350 3292 14356
rect 3424 14408 3476 14414
rect 3424 14350 3476 14356
rect 3792 14408 3844 14414
rect 3792 14350 3844 14356
rect 2778 14311 2834 14320
rect 2792 14074 2820 14311
rect 3054 14104 3110 14113
rect 2780 14068 2832 14074
rect 3252 14090 3280 14350
rect 3252 14062 3372 14090
rect 3436 14074 3464 14350
rect 3054 14039 3110 14048
rect 2780 14010 2832 14016
rect 2688 14000 2740 14006
rect 2688 13942 2740 13948
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12889 2820 13126
rect 3068 12968 3096 14039
rect 3238 13968 3294 13977
rect 3344 13938 3372 14062
rect 3424 14068 3476 14074
rect 3424 14010 3476 14016
rect 3896 13938 3924 14826
rect 3976 14476 4028 14482
rect 3976 14418 4028 14424
rect 3988 14260 4016 14418
rect 4080 14414 4108 14962
rect 4264 14618 4292 15642
rect 4356 14958 4384 16215
rect 4618 15600 4674 15609
rect 4618 15535 4674 15544
rect 5264 15564 5316 15570
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4252 14612 4304 14618
rect 4252 14554 4304 14560
rect 4356 14414 4384 14894
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4632 14770 4660 15535
rect 5264 15506 5316 15512
rect 4986 15056 5042 15065
rect 4986 14991 5042 15000
rect 4068 14408 4120 14414
rect 4068 14350 4120 14356
rect 4344 14408 4396 14414
rect 4344 14350 4396 14356
rect 3988 14232 4292 14260
rect 3238 13903 3240 13912
rect 3292 13903 3294 13912
rect 3332 13932 3384 13938
rect 3240 13874 3292 13880
rect 3332 13874 3384 13880
rect 3884 13932 3936 13938
rect 3884 13874 3936 13880
rect 4160 13864 4212 13870
rect 4066 13832 4122 13841
rect 4160 13806 4212 13812
rect 4066 13767 4122 13776
rect 4080 13734 4108 13767
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3174 13628 3482 13648
rect 3174 13626 3180 13628
rect 3236 13626 3260 13628
rect 3316 13626 3340 13628
rect 3396 13626 3420 13628
rect 3476 13626 3482 13628
rect 3236 13574 3238 13626
rect 3418 13574 3420 13626
rect 3174 13572 3180 13574
rect 3236 13572 3260 13574
rect 3316 13572 3340 13574
rect 3396 13572 3420 13574
rect 3476 13572 3482 13574
rect 3174 13552 3482 13572
rect 3606 13560 3662 13569
rect 3344 13504 3606 13512
rect 3344 13495 3662 13504
rect 3344 13484 3648 13495
rect 3344 13326 3372 13484
rect 3790 13424 3846 13433
rect 3790 13359 3846 13368
rect 4066 13424 4122 13433
rect 4066 13359 4122 13368
rect 3332 13320 3384 13326
rect 3424 13320 3476 13326
rect 3332 13262 3384 13268
rect 3422 13288 3424 13297
rect 3476 13288 3478 13297
rect 3804 13258 3832 13359
rect 4080 13326 4108 13359
rect 3884 13320 3936 13326
rect 3884 13262 3936 13268
rect 4068 13320 4120 13326
rect 4068 13262 4120 13268
rect 3422 13223 3478 13232
rect 3792 13252 3844 13258
rect 3792 13194 3844 13200
rect 3700 13184 3752 13190
rect 3528 13144 3700 13172
rect 3238 13016 3294 13025
rect 3068 12940 3188 12968
rect 3238 12951 3294 12960
rect 2778 12880 2834 12889
rect 2778 12815 2834 12824
rect 3054 12880 3110 12889
rect 3054 12815 3056 12824
rect 3108 12815 3110 12824
rect 3056 12786 3108 12792
rect 2780 12776 2832 12782
rect 2964 12776 3016 12782
rect 2780 12718 2832 12724
rect 2870 12744 2926 12753
rect 2792 12442 2820 12718
rect 2926 12724 2964 12730
rect 3160 12730 3188 12940
rect 3252 12782 3280 12951
rect 2926 12718 3016 12724
rect 2926 12702 3004 12718
rect 3068 12702 3188 12730
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 2870 12679 2926 12688
rect 2964 12640 3016 12646
rect 2964 12582 3016 12588
rect 2976 12481 3004 12582
rect 2962 12472 3018 12481
rect 2780 12436 2832 12442
rect 2962 12407 3018 12416
rect 2780 12378 2832 12384
rect 2502 12336 2558 12345
rect 2412 12300 2464 12306
rect 2502 12271 2558 12280
rect 2412 12242 2464 12248
rect 2424 11286 2452 12242
rect 2504 12164 2556 12170
rect 2504 12106 2556 12112
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2424 10742 2452 11222
rect 2516 11014 2544 12106
rect 2596 12096 2648 12102
rect 2596 12038 2648 12044
rect 2688 12096 2740 12102
rect 2792 12073 2820 12378
rect 2872 12368 2924 12374
rect 2872 12310 2924 12316
rect 2688 12038 2740 12044
rect 2778 12064 2834 12073
rect 2608 11898 2636 12038
rect 2596 11892 2648 11898
rect 2596 11834 2648 11840
rect 2596 11552 2648 11558
rect 2596 11494 2648 11500
rect 2504 11008 2556 11014
rect 2504 10950 2556 10956
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2516 9586 2544 10134
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2608 8974 2636 11494
rect 2700 11354 2728 12038
rect 2778 11999 2834 12008
rect 2884 11665 2912 12310
rect 2964 12232 3016 12238
rect 2964 12174 3016 12180
rect 2870 11656 2926 11665
rect 2870 11591 2926 11600
rect 2976 11393 3004 12174
rect 3068 11694 3096 12702
rect 3174 12540 3482 12560
rect 3174 12538 3180 12540
rect 3236 12538 3260 12540
rect 3316 12538 3340 12540
rect 3396 12538 3420 12540
rect 3476 12538 3482 12540
rect 3236 12486 3238 12538
rect 3418 12486 3420 12538
rect 3174 12484 3180 12486
rect 3236 12484 3260 12486
rect 3316 12484 3340 12486
rect 3396 12484 3420 12486
rect 3476 12484 3482 12486
rect 3174 12464 3482 12484
rect 3422 12336 3478 12345
rect 3422 12271 3424 12280
rect 3476 12271 3478 12280
rect 3424 12242 3476 12248
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3148 12096 3200 12102
rect 3148 12038 3200 12044
rect 3160 11830 3188 12038
rect 3148 11824 3200 11830
rect 3148 11766 3200 11772
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3344 11540 3372 12106
rect 3068 11512 3372 11540
rect 2962 11384 3018 11393
rect 2688 11348 2740 11354
rect 2962 11319 3018 11328
rect 2688 11290 2740 11296
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2884 10606 2912 11086
rect 2962 10976 3018 10985
rect 2962 10911 3018 10920
rect 2976 10742 3004 10911
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2872 10600 2924 10606
rect 3068 10554 3096 11512
rect 3174 11452 3482 11472
rect 3174 11450 3180 11452
rect 3236 11450 3260 11452
rect 3316 11450 3340 11452
rect 3396 11450 3420 11452
rect 3476 11450 3482 11452
rect 3236 11398 3238 11450
rect 3418 11398 3420 11450
rect 3174 11396 3180 11398
rect 3236 11396 3260 11398
rect 3316 11396 3340 11398
rect 3396 11396 3420 11398
rect 3476 11396 3482 11398
rect 3174 11376 3482 11396
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 2872 10542 2924 10548
rect 2780 10464 2832 10470
rect 2778 10432 2780 10441
rect 2832 10432 2834 10441
rect 2778 10367 2834 10376
rect 2792 10130 2820 10367
rect 2780 10124 2832 10130
rect 2780 10066 2832 10072
rect 2688 10056 2740 10062
rect 2688 9998 2740 10004
rect 2596 8968 2648 8974
rect 2502 8936 2558 8945
rect 2596 8910 2648 8916
rect 2502 8871 2558 8880
rect 2516 8566 2544 8871
rect 2504 8560 2556 8566
rect 2504 8502 2556 8508
rect 2280 8236 2360 8242
rect 2228 8230 2360 8236
rect 2240 8214 2360 8230
rect 2516 7954 2544 8502
rect 2596 8492 2648 8498
rect 2596 8434 2648 8440
rect 2608 8265 2636 8434
rect 2594 8256 2650 8265
rect 2594 8191 2650 8200
rect 2700 8022 2728 9998
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2792 8634 2820 9318
rect 2884 9178 2912 10542
rect 2976 10526 3096 10554
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2780 8628 2832 8634
rect 2780 8570 2832 8576
rect 2792 8265 2820 8570
rect 2778 8256 2834 8265
rect 2778 8191 2834 8200
rect 2688 8016 2740 8022
rect 2688 7958 2740 7964
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2596 7880 2648 7886
rect 2596 7822 2648 7828
rect 2780 7880 2832 7886
rect 2884 7868 2912 9114
rect 2976 8537 3004 10526
rect 3056 10464 3108 10470
rect 3160 10452 3188 10950
rect 3108 10424 3188 10452
rect 3056 10406 3108 10412
rect 3068 10248 3096 10406
rect 3174 10364 3482 10384
rect 3174 10362 3180 10364
rect 3236 10362 3260 10364
rect 3316 10362 3340 10364
rect 3396 10362 3420 10364
rect 3476 10362 3482 10364
rect 3236 10310 3238 10362
rect 3418 10310 3420 10362
rect 3174 10308 3180 10310
rect 3236 10308 3260 10310
rect 3316 10308 3340 10310
rect 3396 10308 3420 10310
rect 3476 10308 3482 10310
rect 3174 10288 3482 10308
rect 3068 10220 3464 10248
rect 3056 10124 3108 10130
rect 3056 10066 3108 10072
rect 2962 8528 3018 8537
rect 2962 8463 3018 8472
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2976 8090 3004 8298
rect 2964 8084 3016 8090
rect 2964 8026 3016 8032
rect 3068 8022 3096 10066
rect 3436 10010 3464 10220
rect 3528 10130 3556 13144
rect 3700 13126 3752 13132
rect 3790 12880 3846 12889
rect 3700 12844 3752 12850
rect 3790 12815 3846 12824
rect 3700 12786 3752 12792
rect 3608 12708 3660 12714
rect 3608 12650 3660 12656
rect 3620 12617 3648 12650
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 3712 12434 3740 12786
rect 3804 12617 3832 12815
rect 3790 12608 3846 12617
rect 3790 12543 3846 12552
rect 3620 12406 3740 12434
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 3620 10441 3648 12406
rect 3804 12356 3832 12407
rect 3712 12328 3832 12356
rect 3606 10432 3662 10441
rect 3606 10367 3662 10376
rect 3606 10296 3662 10305
rect 3606 10231 3662 10240
rect 3620 10198 3648 10231
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3608 10056 3660 10062
rect 3436 9982 3556 10010
rect 3608 9998 3660 10004
rect 3712 10010 3740 12328
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3804 11354 3832 11698
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3792 11212 3844 11218
rect 3792 11154 3844 11160
rect 3804 10810 3832 11154
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3790 10704 3846 10713
rect 3790 10639 3846 10648
rect 3804 10266 3832 10639
rect 3792 10260 3844 10266
rect 3792 10202 3844 10208
rect 3896 10198 3924 13262
rect 4080 13190 4108 13262
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4172 12866 4200 13806
rect 4264 13530 4292 14232
rect 4448 14074 4476 14758
rect 4632 14742 4844 14770
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4540 13938 4568 14554
rect 4632 14414 4660 14742
rect 4816 14618 4844 14742
rect 4712 14612 4764 14618
rect 4712 14554 4764 14560
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4620 14272 4672 14278
rect 4620 14214 4672 14220
rect 4528 13932 4580 13938
rect 4528 13874 4580 13880
rect 4528 13796 4580 13802
rect 4528 13738 4580 13744
rect 4252 13524 4304 13530
rect 4252 13466 4304 13472
rect 4252 13184 4304 13190
rect 4436 13184 4488 13190
rect 4252 13126 4304 13132
rect 4342 13152 4398 13161
rect 4264 13025 4292 13126
rect 4436 13126 4488 13132
rect 4342 13087 4398 13096
rect 4250 13016 4306 13025
rect 4356 12986 4384 13087
rect 4250 12951 4306 12960
rect 4344 12980 4396 12986
rect 4344 12922 4396 12928
rect 3988 12838 4200 12866
rect 4250 12880 4306 12889
rect 3988 12186 4016 12838
rect 4250 12815 4252 12824
rect 4304 12815 4306 12824
rect 4252 12786 4304 12792
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4068 12640 4120 12646
rect 4068 12582 4120 12588
rect 4080 12288 4108 12582
rect 4080 12260 4200 12288
rect 3988 12170 4108 12186
rect 3988 12164 4120 12170
rect 3988 12158 4068 12164
rect 4068 12106 4120 12112
rect 3976 12096 4028 12102
rect 3974 12064 3976 12073
rect 4028 12064 4030 12073
rect 4172 12050 4200 12260
rect 3974 11999 4030 12008
rect 4080 12022 4200 12050
rect 4252 12096 4304 12102
rect 4252 12038 4304 12044
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3884 10192 3936 10198
rect 3884 10134 3936 10140
rect 3174 9276 3482 9296
rect 3174 9274 3180 9276
rect 3236 9274 3260 9276
rect 3316 9274 3340 9276
rect 3396 9274 3420 9276
rect 3476 9274 3482 9276
rect 3236 9222 3238 9274
rect 3418 9222 3420 9274
rect 3174 9220 3180 9222
rect 3236 9220 3260 9222
rect 3316 9220 3340 9222
rect 3396 9220 3420 9222
rect 3476 9220 3482 9222
rect 3174 9200 3482 9220
rect 3528 9160 3556 9982
rect 3344 9132 3556 9160
rect 3146 8936 3202 8945
rect 3146 8871 3202 8880
rect 3160 8430 3188 8871
rect 3240 8560 3292 8566
rect 3238 8528 3240 8537
rect 3292 8528 3294 8537
rect 3238 8463 3294 8472
rect 3148 8424 3200 8430
rect 3344 8412 3372 9132
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3528 8786 3556 8842
rect 3436 8758 3556 8786
rect 3436 8566 3464 8758
rect 3620 8650 3648 9998
rect 3712 9982 3832 10010
rect 3700 9920 3752 9926
rect 3700 9862 3752 9868
rect 3712 9081 3740 9862
rect 3804 9722 3832 9982
rect 3884 9920 3936 9926
rect 3884 9862 3936 9868
rect 3896 9761 3924 9862
rect 3882 9752 3938 9761
rect 3792 9716 3844 9722
rect 3882 9687 3938 9696
rect 3792 9658 3844 9664
rect 3698 9072 3754 9081
rect 3698 9007 3754 9016
rect 3804 8974 3832 9658
rect 3884 9580 3936 9586
rect 3884 9522 3936 9528
rect 3792 8968 3844 8974
rect 3698 8936 3754 8945
rect 3792 8910 3844 8916
rect 3698 8871 3754 8880
rect 3712 8838 3740 8871
rect 3700 8832 3752 8838
rect 3700 8774 3752 8780
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3896 8786 3924 9522
rect 3988 9178 4016 11630
rect 4080 10962 4108 12022
rect 4160 11552 4212 11558
rect 4160 11494 4212 11500
rect 4172 11218 4200 11494
rect 4160 11212 4212 11218
rect 4160 11154 4212 11160
rect 4264 11121 4292 12038
rect 4356 11937 4384 12650
rect 4342 11928 4398 11937
rect 4342 11863 4398 11872
rect 4344 11688 4396 11694
rect 4344 11630 4396 11636
rect 4250 11112 4306 11121
rect 4250 11047 4306 11056
rect 4080 10934 4200 10962
rect 4066 10840 4122 10849
rect 4066 10775 4122 10784
rect 4080 10062 4108 10775
rect 4068 10056 4120 10062
rect 4172 10033 4200 10934
rect 4356 10062 4384 11630
rect 4448 11336 4476 13126
rect 4540 12306 4568 13738
rect 4632 13326 4660 14214
rect 4724 14074 4752 14554
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 4712 14068 4764 14074
rect 4712 14010 4764 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4724 13841 4752 13874
rect 4710 13832 4766 13841
rect 4710 13767 4766 13776
rect 4908 13705 4936 14214
rect 5000 14113 5028 14991
rect 5078 14240 5134 14249
rect 5078 14175 5134 14184
rect 4986 14104 5042 14113
rect 4986 14039 4988 14048
rect 5040 14039 5042 14048
rect 4988 14010 5040 14016
rect 5000 13979 5028 14010
rect 5092 13938 5120 14175
rect 5172 14000 5224 14006
rect 5172 13942 5224 13948
rect 5080 13932 5132 13938
rect 5080 13874 5132 13880
rect 5080 13728 5132 13734
rect 4894 13696 4950 13705
rect 4894 13631 4950 13640
rect 5000 13688 5080 13716
rect 4804 13456 4856 13462
rect 4804 13398 4856 13404
rect 4816 13326 4844 13398
rect 4620 13320 4672 13326
rect 4620 13262 4672 13268
rect 4804 13320 4856 13326
rect 4804 13262 4856 13268
rect 4896 13320 4948 13326
rect 4896 13262 4948 13268
rect 4710 13016 4766 13025
rect 4710 12951 4766 12960
rect 4528 12300 4580 12306
rect 4528 12242 4580 12248
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4632 11558 4660 12242
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4448 11308 4660 11336
rect 4436 11212 4488 11218
rect 4436 11154 4488 11160
rect 4528 11212 4580 11218
rect 4528 11154 4580 11160
rect 4448 11082 4476 11154
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4448 10470 4476 11018
rect 4540 10810 4568 11154
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4436 10464 4488 10470
rect 4488 10424 4568 10452
rect 4436 10406 4488 10412
rect 4344 10056 4396 10062
rect 4068 9998 4120 10004
rect 4158 10024 4214 10033
rect 4344 9998 4396 10004
rect 4158 9959 4214 9968
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9580 4120 9586
rect 4068 9522 4120 9528
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 4080 9110 4108 9522
rect 4172 9382 4200 9862
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4068 9104 4120 9110
rect 3974 9072 4030 9081
rect 4068 9046 4120 9052
rect 3974 9007 4030 9016
rect 3988 8906 4016 9007
rect 3976 8900 4028 8906
rect 3976 8842 4028 8848
rect 3620 8622 3740 8650
rect 3424 8560 3476 8566
rect 3712 8548 3740 8622
rect 3804 8566 3832 8774
rect 3896 8758 3933 8786
rect 3905 8566 3933 8758
rect 3424 8502 3476 8508
rect 3620 8520 3740 8548
rect 3792 8560 3844 8566
rect 3344 8384 3556 8412
rect 3148 8366 3200 8372
rect 3174 8188 3482 8208
rect 3174 8186 3180 8188
rect 3236 8186 3260 8188
rect 3316 8186 3340 8188
rect 3396 8186 3420 8188
rect 3476 8186 3482 8188
rect 3236 8134 3238 8186
rect 3418 8134 3420 8186
rect 3174 8132 3180 8134
rect 3236 8132 3260 8134
rect 3316 8132 3340 8134
rect 3396 8132 3420 8134
rect 3476 8132 3482 8134
rect 3174 8112 3482 8132
rect 3528 8072 3556 8384
rect 3620 8129 3648 8520
rect 3792 8502 3844 8508
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3976 8492 4028 8498
rect 4080 8480 4108 9046
rect 4172 8838 4200 9114
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4028 8452 4108 8480
rect 3976 8434 4028 8440
rect 3974 8392 4030 8401
rect 3974 8327 4030 8336
rect 3700 8306 3752 8312
rect 3884 8306 3936 8312
rect 3752 8254 3832 8294
rect 3700 8248 3832 8254
rect 3882 8256 3884 8265
rect 3988 8294 4016 8327
rect 3988 8266 4108 8294
rect 3936 8256 3938 8265
rect 3436 8044 3556 8072
rect 3606 8120 3662 8129
rect 3712 8106 3740 8248
rect 3882 8191 3938 8200
rect 3712 8078 3832 8106
rect 3606 8055 3662 8064
rect 3804 8072 3832 8078
rect 3804 8044 3924 8072
rect 3056 8016 3108 8022
rect 3332 8016 3384 8022
rect 3056 7958 3108 7964
rect 3238 7984 3294 7993
rect 3332 7958 3384 7964
rect 3238 7919 3240 7928
rect 3292 7919 3294 7928
rect 3240 7890 3292 7896
rect 2884 7840 3004 7868
rect 3344 7857 3372 7958
rect 2780 7822 2832 7828
rect 2136 7540 2188 7546
rect 2136 7482 2188 7488
rect 2320 7540 2372 7546
rect 2320 7482 2372 7488
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 2148 6458 2176 7346
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2136 6248 2188 6254
rect 2136 6190 2188 6196
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 1950 5264 2006 5273
rect 1950 5199 2006 5208
rect 1964 4826 1992 5199
rect 2044 5024 2096 5030
rect 2044 4966 2096 4972
rect 1952 4820 2004 4826
rect 1952 4762 2004 4768
rect 1952 4684 2004 4690
rect 1952 4626 2004 4632
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1964 3482 1992 4626
rect 2056 3641 2084 4966
rect 2042 3632 2098 3641
rect 2042 3567 2098 3576
rect 1964 3454 2084 3482
rect 1952 3392 2004 3398
rect 1952 3334 2004 3340
rect 1964 3194 1992 3334
rect 1952 3188 2004 3194
rect 1952 3130 2004 3136
rect 1766 2952 1822 2961
rect 1766 2887 1822 2896
rect 1766 2680 1822 2689
rect 1766 2615 1822 2624
rect 1780 2446 1808 2615
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 1584 2304 1636 2310
rect 1584 2246 1636 2252
rect 1490 232 1546 241
rect 1490 167 1546 176
rect 1596 66 1624 2246
rect 2056 1834 2084 3454
rect 2148 2990 2176 6190
rect 2332 5846 2360 7482
rect 2504 7404 2556 7410
rect 2504 7346 2556 7352
rect 2516 6798 2544 7346
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2608 6304 2636 7822
rect 2686 7576 2742 7585
rect 2686 7511 2742 7520
rect 2700 7342 2728 7511
rect 2688 7336 2740 7342
rect 2688 7278 2740 7284
rect 2792 7041 2820 7822
rect 2976 7410 3004 7840
rect 3330 7848 3386 7857
rect 3330 7783 3386 7792
rect 3056 7540 3108 7546
rect 3056 7482 3108 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2778 7032 2834 7041
rect 2778 6967 2834 6976
rect 2964 6452 3016 6458
rect 2964 6394 3016 6400
rect 2872 6384 2924 6390
rect 2872 6326 2924 6332
rect 2688 6316 2740 6322
rect 2608 6276 2688 6304
rect 2688 6258 2740 6264
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2320 5840 2372 5846
rect 2320 5782 2372 5788
rect 2424 5710 2452 6054
rect 2412 5704 2464 5710
rect 2412 5646 2464 5652
rect 2228 5568 2280 5574
rect 2700 5545 2728 6258
rect 2228 5510 2280 5516
rect 2686 5536 2742 5545
rect 2136 2984 2188 2990
rect 2136 2926 2188 2932
rect 2240 2922 2268 5510
rect 2686 5471 2742 5480
rect 2688 5228 2740 5234
rect 2688 5170 2740 5176
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2410 4856 2466 4865
rect 2516 4826 2544 4966
rect 2410 4791 2466 4800
rect 2504 4820 2556 4826
rect 2318 4720 2374 4729
rect 2318 4655 2320 4664
rect 2372 4655 2374 4664
rect 2320 4626 2372 4632
rect 2424 4622 2452 4791
rect 2504 4762 2556 4768
rect 2502 4720 2558 4729
rect 2502 4655 2558 4664
rect 2412 4616 2464 4622
rect 2412 4558 2464 4564
rect 2412 4480 2464 4486
rect 2412 4422 2464 4428
rect 2424 3942 2452 4422
rect 2412 3936 2464 3942
rect 2412 3878 2464 3884
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2228 2916 2280 2922
rect 2228 2858 2280 2864
rect 2136 2848 2188 2854
rect 2136 2790 2188 2796
rect 2044 1828 2096 1834
rect 2044 1770 2096 1776
rect 2148 800 2176 2790
rect 2228 2304 2280 2310
rect 2228 2246 2280 2252
rect 2240 2038 2268 2246
rect 2228 2032 2280 2038
rect 2228 1974 2280 1980
rect 2332 1630 2360 3334
rect 2424 1902 2452 3878
rect 2516 3602 2544 4655
rect 2700 4486 2728 5170
rect 2780 5092 2832 5098
rect 2780 5034 2832 5040
rect 2792 4706 2820 5034
rect 2884 4826 2912 6326
rect 2976 6089 3004 6394
rect 2962 6080 3018 6089
rect 2962 6015 3018 6024
rect 2962 5944 3018 5953
rect 2962 5879 3018 5888
rect 2976 5778 3004 5879
rect 2964 5772 3016 5778
rect 2964 5714 3016 5720
rect 3068 5710 3096 7482
rect 3436 7460 3464 8044
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3792 7880 3844 7886
rect 3896 7868 3924 8044
rect 3844 7840 3924 7868
rect 3792 7822 3844 7828
rect 3528 7562 3556 7822
rect 3608 7812 3660 7818
rect 3608 7754 3660 7760
rect 3620 7721 3648 7754
rect 3606 7712 3662 7721
rect 3606 7647 3662 7656
rect 3528 7534 3648 7562
rect 3436 7432 3556 7460
rect 3174 7100 3482 7120
rect 3174 7098 3180 7100
rect 3236 7098 3260 7100
rect 3316 7098 3340 7100
rect 3396 7098 3420 7100
rect 3476 7098 3482 7100
rect 3236 7046 3238 7098
rect 3418 7046 3420 7098
rect 3174 7044 3180 7046
rect 3236 7044 3260 7046
rect 3316 7044 3340 7046
rect 3396 7044 3420 7046
rect 3476 7044 3482 7046
rect 3174 7024 3482 7044
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 3422 6896 3478 6905
rect 3160 6361 3188 6870
rect 3422 6831 3424 6840
rect 3476 6831 3478 6840
rect 3424 6802 3476 6808
rect 3528 6662 3556 7432
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3436 6390 3464 6598
rect 3424 6384 3476 6390
rect 3146 6352 3202 6361
rect 3424 6326 3476 6332
rect 3146 6287 3148 6296
rect 3200 6287 3202 6296
rect 3516 6316 3568 6322
rect 3148 6258 3200 6264
rect 3516 6258 3568 6264
rect 3174 6012 3482 6032
rect 3174 6010 3180 6012
rect 3236 6010 3260 6012
rect 3316 6010 3340 6012
rect 3396 6010 3420 6012
rect 3476 6010 3482 6012
rect 3236 5958 3238 6010
rect 3418 5958 3420 6010
rect 3174 5956 3180 5958
rect 3236 5956 3260 5958
rect 3316 5956 3340 5958
rect 3396 5956 3420 5958
rect 3476 5956 3482 5958
rect 3174 5936 3482 5956
rect 3528 5914 3556 6258
rect 3516 5908 3568 5914
rect 3516 5850 3568 5856
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2962 5128 3018 5137
rect 2962 5063 3018 5072
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 2792 4678 2912 4706
rect 2688 4480 2740 4486
rect 2688 4422 2740 4428
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2596 3936 2648 3942
rect 2596 3878 2648 3884
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2504 3392 2556 3398
rect 2504 3334 2556 3340
rect 2516 3194 2544 3334
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2504 2848 2556 2854
rect 2504 2790 2556 2796
rect 2516 2514 2544 2790
rect 2608 2650 2636 3878
rect 2792 3126 2820 4014
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2884 2514 2912 4678
rect 2976 4282 3004 5063
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3174 4924 3482 4944
rect 3174 4922 3180 4924
rect 3236 4922 3260 4924
rect 3316 4922 3340 4924
rect 3396 4922 3420 4924
rect 3476 4922 3482 4924
rect 3236 4870 3238 4922
rect 3418 4870 3420 4922
rect 3174 4868 3180 4870
rect 3236 4868 3260 4870
rect 3316 4868 3340 4870
rect 3396 4868 3420 4870
rect 3476 4868 3482 4870
rect 3174 4848 3482 4868
rect 3422 4720 3478 4729
rect 3422 4655 3424 4664
rect 3476 4655 3478 4664
rect 3424 4626 3476 4632
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2976 2825 3004 2858
rect 2962 2816 3018 2825
rect 2962 2751 3018 2760
rect 2964 2644 3016 2650
rect 2964 2586 3016 2592
rect 2504 2508 2556 2514
rect 2504 2450 2556 2456
rect 2872 2508 2924 2514
rect 2872 2450 2924 2456
rect 2976 2292 3004 2586
rect 3068 2446 3096 4490
rect 3240 4480 3292 4486
rect 3240 4422 3292 4428
rect 3252 4321 3280 4422
rect 3238 4312 3294 4321
rect 3238 4247 3294 4256
rect 3174 3836 3482 3856
rect 3174 3834 3180 3836
rect 3236 3834 3260 3836
rect 3316 3834 3340 3836
rect 3396 3834 3420 3836
rect 3476 3834 3482 3836
rect 3236 3782 3238 3834
rect 3418 3782 3420 3834
rect 3174 3780 3180 3782
rect 3236 3780 3260 3782
rect 3316 3780 3340 3782
rect 3396 3780 3420 3782
rect 3476 3780 3482 3782
rect 3174 3760 3482 3780
rect 3528 3505 3556 4966
rect 3620 4486 3648 7534
rect 3698 7304 3754 7313
rect 3698 7239 3754 7248
rect 3712 4554 3740 7239
rect 3804 7177 3832 7822
rect 4080 7721 4108 8266
rect 4158 8256 4214 8265
rect 4158 8191 4214 8200
rect 4172 8090 4200 8191
rect 4264 8129 4292 9930
rect 4344 9920 4396 9926
rect 4344 9862 4396 9868
rect 4356 8838 4384 9862
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4448 8906 4476 9318
rect 4540 9042 4568 10424
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4436 8900 4488 8906
rect 4436 8842 4488 8848
rect 4344 8832 4396 8838
rect 4528 8832 4580 8838
rect 4344 8774 4396 8780
rect 4526 8800 4528 8809
rect 4580 8800 4582 8809
rect 4526 8735 4582 8744
rect 4344 8288 4396 8294
rect 4344 8230 4396 8236
rect 4250 8120 4306 8129
rect 4160 8084 4212 8090
rect 4250 8055 4306 8064
rect 4160 8026 4212 8032
rect 4356 7936 4384 8230
rect 4436 8016 4488 8022
rect 4436 7958 4488 7964
rect 4264 7908 4384 7936
rect 4066 7712 4122 7721
rect 4066 7647 4122 7656
rect 4264 7546 4292 7908
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4356 7721 4384 7754
rect 4342 7712 4398 7721
rect 4342 7647 4398 7656
rect 4252 7540 4304 7546
rect 4252 7482 4304 7488
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 3790 7168 3846 7177
rect 3790 7103 3846 7112
rect 3790 6624 3846 6633
rect 3790 6559 3846 6568
rect 3804 4826 3832 6559
rect 3988 6202 4016 7414
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3988 6174 4108 6202
rect 3976 6112 4028 6118
rect 3976 6054 4028 6060
rect 3988 5710 4016 6054
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3988 5098 4016 5646
rect 3976 5092 4028 5098
rect 3976 5034 4028 5040
rect 3792 4820 3844 4826
rect 3792 4762 3844 4768
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3608 4480 3660 4486
rect 3608 4422 3660 4428
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3620 3670 3648 4422
rect 3790 4040 3846 4049
rect 3790 3975 3846 3984
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3608 3664 3660 3670
rect 3608 3606 3660 3612
rect 3514 3496 3570 3505
rect 3514 3431 3570 3440
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3516 3392 3568 3398
rect 3516 3334 3568 3340
rect 3160 3194 3188 3334
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3174 2748 3482 2768
rect 3174 2746 3180 2748
rect 3236 2746 3260 2748
rect 3316 2746 3340 2748
rect 3396 2746 3420 2748
rect 3476 2746 3482 2748
rect 3236 2694 3238 2746
rect 3418 2694 3420 2746
rect 3174 2692 3180 2694
rect 3236 2692 3260 2694
rect 3316 2692 3340 2694
rect 3396 2692 3420 2694
rect 3476 2692 3482 2694
rect 3174 2672 3482 2692
rect 3424 2576 3476 2582
rect 3424 2518 3476 2524
rect 3148 2508 3200 2514
rect 3148 2450 3200 2456
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 3160 2292 3188 2450
rect 2976 2264 3188 2292
rect 3436 2009 3464 2518
rect 3422 2000 3478 2009
rect 3056 1964 3108 1970
rect 3422 1935 3478 1944
rect 3056 1906 3108 1912
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2320 1624 2372 1630
rect 2320 1566 2372 1572
rect 3068 800 3096 1906
rect 3528 1630 3556 3334
rect 3516 1624 3568 1630
rect 3516 1566 3568 1572
rect 3620 1290 3648 3606
rect 3712 3097 3740 3878
rect 3804 3398 3832 3975
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3698 3088 3754 3097
rect 3698 3023 3754 3032
rect 3896 2836 3924 4422
rect 3988 4264 4016 5034
rect 4080 4457 4108 6174
rect 4172 5642 4200 7278
rect 4356 6225 4384 7346
rect 4448 7342 4476 7958
rect 4526 7848 4582 7857
rect 4526 7783 4528 7792
rect 4580 7783 4582 7792
rect 4528 7754 4580 7760
rect 4632 7750 4660 11308
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4632 7585 4660 7686
rect 4618 7576 4674 7585
rect 4618 7511 4674 7520
rect 4436 7336 4488 7342
rect 4620 7336 4672 7342
rect 4436 7278 4488 7284
rect 4618 7304 4620 7313
rect 4672 7304 4674 7313
rect 4618 7239 4674 7248
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4448 6866 4476 7142
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 4540 6798 4568 7142
rect 4632 7041 4660 7239
rect 4618 7032 4674 7041
rect 4618 6967 4674 6976
rect 4620 6928 4672 6934
rect 4618 6896 4620 6905
rect 4672 6896 4674 6905
rect 4618 6831 4674 6840
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4620 6656 4672 6662
rect 4620 6598 4672 6604
rect 4434 6488 4490 6497
rect 4434 6423 4490 6432
rect 4448 6254 4476 6423
rect 4528 6316 4580 6322
rect 4528 6258 4580 6264
rect 4436 6248 4488 6254
rect 4342 6216 4398 6225
rect 4436 6190 4488 6196
rect 4342 6151 4398 6160
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4172 5098 4200 5170
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4250 4584 4306 4593
rect 4250 4519 4306 4528
rect 4160 4480 4212 4486
rect 4066 4448 4122 4457
rect 4160 4422 4212 4428
rect 4066 4383 4122 4392
rect 4068 4276 4120 4282
rect 3988 4236 4068 4264
rect 4068 4218 4120 4224
rect 4068 4140 4120 4146
rect 3988 4100 4068 4128
rect 3988 3602 4016 4100
rect 4068 4082 4120 4088
rect 3976 3596 4028 3602
rect 3976 3538 4028 3544
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3988 2990 4016 3334
rect 4172 3074 4200 4422
rect 4264 3777 4292 4519
rect 4250 3768 4306 3777
rect 4250 3703 4306 3712
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4080 3058 4200 3074
rect 4068 3052 4200 3058
rect 4120 3046 4200 3052
rect 4068 2994 4120 3000
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 4068 2848 4120 2854
rect 3790 2816 3846 2825
rect 3896 2808 4016 2836
rect 3790 2751 3846 2760
rect 3804 2446 3832 2751
rect 3882 2680 3938 2689
rect 3882 2615 3884 2624
rect 3936 2615 3938 2624
rect 3884 2586 3936 2592
rect 3792 2440 3844 2446
rect 3792 2382 3844 2388
rect 3608 1284 3660 1290
rect 3608 1226 3660 1232
rect 3424 876 3476 882
rect 3424 818 3476 824
rect 1584 60 1636 66
rect 1584 2 1636 8
rect 2134 0 2190 800
rect 3054 0 3110 800
rect 3436 785 3464 818
rect 3988 800 4016 2808
rect 4068 2790 4120 2796
rect 4080 2650 4108 2790
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4264 2446 4292 3334
rect 4356 3126 4384 6151
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4448 5642 4476 6054
rect 4436 5636 4488 5642
rect 4436 5578 4488 5584
rect 4448 4593 4476 5578
rect 4540 5370 4568 6258
rect 4632 5370 4660 6598
rect 4724 6186 4752 12951
rect 4908 12889 4936 13262
rect 4894 12880 4950 12889
rect 5000 12850 5028 13688
rect 5080 13670 5132 13676
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4894 12815 4950 12824
rect 4988 12844 5040 12850
rect 4988 12786 5040 12792
rect 5092 12434 5120 13262
rect 5184 12850 5212 13942
rect 5276 13705 5304 15506
rect 5816 15292 5868 15298
rect 5816 15234 5868 15240
rect 5722 14920 5778 14929
rect 5722 14855 5778 14864
rect 5354 14648 5410 14657
rect 5354 14583 5410 14592
rect 5368 14550 5396 14583
rect 5356 14544 5408 14550
rect 5356 14486 5408 14492
rect 5736 14385 5764 14855
rect 5722 14376 5778 14385
rect 5722 14311 5778 14320
rect 5828 14226 5856 15234
rect 5920 14618 5948 16400
rect 6552 15836 6604 15842
rect 6552 15778 6604 15784
rect 6460 15360 6512 15366
rect 6460 15302 6512 15308
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6000 14884 6052 14890
rect 6000 14826 6052 14832
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6012 14550 6040 14826
rect 6104 14550 6132 14894
rect 6184 14884 6236 14890
rect 6184 14826 6236 14832
rect 6000 14544 6052 14550
rect 6000 14486 6052 14492
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 6196 14362 6224 14826
rect 6368 14408 6420 14414
rect 6012 14334 6224 14362
rect 6274 14376 6330 14385
rect 5828 14198 5948 14226
rect 5398 14172 5706 14192
rect 5398 14170 5404 14172
rect 5460 14170 5484 14172
rect 5540 14170 5564 14172
rect 5620 14170 5644 14172
rect 5700 14170 5706 14172
rect 5460 14118 5462 14170
rect 5642 14118 5644 14170
rect 5398 14116 5404 14118
rect 5460 14116 5484 14118
rect 5540 14116 5564 14118
rect 5620 14116 5644 14118
rect 5700 14116 5706 14118
rect 5398 14096 5706 14116
rect 5814 14104 5870 14113
rect 5814 14039 5816 14048
rect 5868 14039 5870 14048
rect 5816 14010 5868 14016
rect 5632 14000 5684 14006
rect 5632 13942 5684 13948
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5356 13728 5408 13734
rect 5262 13696 5318 13705
rect 5540 13728 5592 13734
rect 5446 13696 5502 13705
rect 5408 13676 5446 13682
rect 5356 13670 5446 13676
rect 5368 13654 5446 13670
rect 5262 13631 5318 13640
rect 5540 13670 5592 13676
rect 5446 13631 5502 13640
rect 5276 13326 5304 13631
rect 5356 13524 5408 13530
rect 5356 13466 5408 13472
rect 5368 13433 5396 13466
rect 5354 13424 5410 13433
rect 5552 13394 5580 13670
rect 5644 13394 5672 13942
rect 5354 13359 5410 13368
rect 5540 13388 5592 13394
rect 5540 13330 5592 13336
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5264 13320 5316 13326
rect 5264 13262 5316 13268
rect 5264 13184 5316 13190
rect 5264 13126 5316 13132
rect 5172 12844 5224 12850
rect 5172 12786 5224 12792
rect 5170 12744 5226 12753
rect 5170 12679 5172 12688
rect 5224 12679 5226 12688
rect 5172 12650 5224 12656
rect 5000 12406 5120 12434
rect 4804 12232 4856 12238
rect 4804 12174 4856 12180
rect 4816 6458 4844 12174
rect 4896 11552 4948 11558
rect 4896 11494 4948 11500
rect 4908 7410 4936 11494
rect 5000 10985 5028 12406
rect 5276 12152 5304 13126
rect 5398 13084 5706 13104
rect 5398 13082 5404 13084
rect 5460 13082 5484 13084
rect 5540 13082 5564 13084
rect 5620 13082 5644 13084
rect 5700 13082 5706 13084
rect 5460 13030 5462 13082
rect 5642 13030 5644 13082
rect 5398 13028 5404 13030
rect 5460 13028 5484 13030
rect 5540 13028 5564 13030
rect 5620 13028 5644 13030
rect 5700 13028 5706 13030
rect 5398 13008 5706 13028
rect 5736 12900 5764 13942
rect 5920 13734 5948 14198
rect 6012 13938 6040 14334
rect 6368 14350 6420 14356
rect 6274 14311 6330 14320
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5816 13320 5868 13326
rect 5816 13262 5868 13268
rect 5828 12986 5856 13262
rect 5908 13184 5960 13190
rect 5908 13126 5960 13132
rect 5816 12980 5868 12986
rect 5816 12922 5868 12928
rect 5644 12872 5764 12900
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5368 12209 5396 12786
rect 5644 12345 5672 12872
rect 5920 12646 5948 13126
rect 5908 12640 5960 12646
rect 6012 12617 6040 13874
rect 6090 13424 6146 13433
rect 6090 13359 6146 13368
rect 6104 12918 6132 13359
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6092 12912 6144 12918
rect 6196 12889 6224 13126
rect 6092 12854 6144 12860
rect 6182 12880 6238 12889
rect 6288 12850 6316 14311
rect 6380 14074 6408 14350
rect 6472 14074 6500 15302
rect 6368 14068 6420 14074
rect 6368 14010 6420 14016
rect 6460 14068 6512 14074
rect 6460 14010 6512 14016
rect 6564 13938 6592 15778
rect 8116 15496 8168 15502
rect 8116 15438 8168 15444
rect 6644 15224 6696 15230
rect 6644 15166 6696 15172
rect 6656 14618 6684 15166
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 6920 15088 6972 15094
rect 6920 15030 6972 15036
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6748 14550 6776 14962
rect 6932 14550 6960 15030
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 14657 7144 14894
rect 7102 14648 7158 14657
rect 7102 14583 7158 14592
rect 6736 14544 6788 14550
rect 6736 14486 6788 14492
rect 6920 14544 6972 14550
rect 6920 14486 6972 14492
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7024 14362 7052 14486
rect 6748 14334 7052 14362
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6644 13728 6696 13734
rect 6644 13670 6696 13676
rect 6656 13530 6684 13670
rect 6644 13524 6696 13530
rect 6644 13466 6696 13472
rect 6748 13394 6776 14334
rect 6826 14240 6882 14249
rect 6826 14175 6882 14184
rect 6840 13938 6868 14175
rect 7012 14068 7064 14074
rect 7012 14010 7064 14016
rect 6920 14000 6972 14006
rect 6918 13968 6920 13977
rect 6972 13968 6974 13977
rect 6828 13932 6880 13938
rect 6918 13903 6974 13912
rect 6828 13874 6880 13880
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 6550 13288 6606 13297
rect 6550 13223 6552 13232
rect 6604 13223 6606 13232
rect 6552 13194 6604 13200
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6182 12815 6238 12824
rect 6276 12844 6328 12850
rect 6090 12744 6146 12753
rect 6090 12679 6146 12688
rect 6104 12646 6132 12679
rect 6092 12640 6144 12646
rect 5908 12582 5960 12588
rect 5998 12608 6054 12617
rect 5630 12336 5686 12345
rect 5920 12306 5948 12582
rect 6196 12617 6224 12815
rect 6276 12786 6328 12792
rect 6460 12776 6512 12782
rect 6460 12718 6512 12724
rect 6276 12708 6328 12714
rect 6276 12650 6328 12656
rect 6092 12582 6144 12588
rect 6182 12608 6238 12617
rect 5998 12543 6054 12552
rect 6182 12543 6238 12552
rect 6182 12472 6238 12481
rect 6182 12407 6238 12416
rect 5630 12271 5686 12280
rect 5816 12300 5868 12306
rect 5816 12242 5868 12248
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 5448 12232 5500 12238
rect 5092 12124 5304 12152
rect 5354 12200 5410 12209
rect 5448 12174 5500 12180
rect 5828 12186 5856 12242
rect 5998 12200 6054 12209
rect 5354 12135 5410 12144
rect 5092 11665 5120 12124
rect 5460 12084 5488 12174
rect 5828 12158 5948 12186
rect 5184 12056 5488 12084
rect 5816 12096 5868 12102
rect 5078 11656 5134 11665
rect 5078 11591 5134 11600
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 4986 10976 5042 10985
rect 4986 10911 5042 10920
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 5000 10130 5028 10678
rect 5092 10130 5120 11018
rect 4988 10124 5040 10130
rect 4988 10066 5040 10072
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 5000 9518 5028 10066
rect 5092 9722 5120 10066
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 5000 6934 5028 9454
rect 5080 9376 5132 9382
rect 5078 9344 5080 9353
rect 5132 9344 5134 9353
rect 5078 9279 5134 9288
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 5092 6769 5120 8774
rect 5078 6760 5134 6769
rect 5078 6695 5134 6704
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 4710 5536 4766 5545
rect 4710 5471 4766 5480
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4724 5234 4752 5471
rect 4712 5228 4764 5234
rect 4712 5170 4764 5176
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4434 4584 4490 4593
rect 4434 4519 4490 4528
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4448 3602 4476 4150
rect 4540 4146 4568 4966
rect 4816 4690 4844 6394
rect 5000 6225 5028 6394
rect 4986 6216 5042 6225
rect 4986 6151 5042 6160
rect 5080 6180 5132 6186
rect 5080 6122 5132 6128
rect 4894 6080 4950 6089
rect 4894 6015 4950 6024
rect 4908 5642 4936 6015
rect 5092 5681 5120 6122
rect 5184 5914 5212 12056
rect 5920 12073 5948 12158
rect 5998 12135 6000 12144
rect 6052 12135 6054 12144
rect 6000 12106 6052 12112
rect 6196 12102 6224 12407
rect 6092 12096 6144 12102
rect 5816 12038 5868 12044
rect 5906 12064 5962 12073
rect 5398 11996 5706 12016
rect 5398 11994 5404 11996
rect 5460 11994 5484 11996
rect 5540 11994 5564 11996
rect 5620 11994 5644 11996
rect 5700 11994 5706 11996
rect 5460 11942 5462 11994
rect 5642 11942 5644 11994
rect 5398 11940 5404 11942
rect 5460 11940 5484 11942
rect 5540 11940 5564 11942
rect 5620 11940 5644 11942
rect 5700 11940 5706 11942
rect 5398 11920 5706 11940
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5264 11552 5316 11558
rect 5368 11529 5396 11630
rect 5264 11494 5316 11500
rect 5354 11520 5410 11529
rect 5276 8956 5304 11494
rect 5354 11455 5410 11464
rect 5736 11393 5764 11698
rect 5722 11384 5778 11393
rect 5722 11319 5778 11328
rect 5398 10908 5706 10928
rect 5398 10906 5404 10908
rect 5460 10906 5484 10908
rect 5540 10906 5564 10908
rect 5620 10906 5644 10908
rect 5700 10906 5706 10908
rect 5460 10854 5462 10906
rect 5642 10854 5644 10906
rect 5398 10852 5404 10854
rect 5460 10852 5484 10854
rect 5540 10852 5564 10854
rect 5620 10852 5644 10854
rect 5700 10852 5706 10854
rect 5398 10832 5706 10852
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5540 10464 5592 10470
rect 5540 10406 5592 10412
rect 5552 9994 5580 10406
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5398 9820 5706 9840
rect 5398 9818 5404 9820
rect 5460 9818 5484 9820
rect 5540 9818 5564 9820
rect 5620 9818 5644 9820
rect 5700 9818 5706 9820
rect 5460 9766 5462 9818
rect 5642 9766 5644 9818
rect 5398 9764 5404 9766
rect 5460 9764 5484 9766
rect 5540 9764 5564 9766
rect 5620 9764 5644 9766
rect 5700 9764 5706 9766
rect 5398 9744 5706 9764
rect 5356 8968 5408 8974
rect 5276 8928 5356 8956
rect 5356 8910 5408 8916
rect 5736 8906 5764 10542
rect 5828 10130 5856 12038
rect 6092 12038 6144 12044
rect 6184 12096 6236 12102
rect 6184 12038 6236 12044
rect 5906 11999 5962 12008
rect 5908 11824 5960 11830
rect 5906 11792 5908 11801
rect 5960 11792 5962 11801
rect 5906 11727 5962 11736
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 10849 5948 11494
rect 5906 10840 5962 10849
rect 5906 10775 5962 10784
rect 5908 10736 5960 10742
rect 5908 10678 5960 10684
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5816 9988 5868 9994
rect 5816 9930 5868 9936
rect 5828 9450 5856 9930
rect 5816 9444 5868 9450
rect 5816 9386 5868 9392
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5398 8732 5706 8752
rect 5398 8730 5404 8732
rect 5460 8730 5484 8732
rect 5540 8730 5564 8732
rect 5620 8730 5644 8732
rect 5700 8730 5706 8732
rect 5460 8678 5462 8730
rect 5642 8678 5644 8730
rect 5398 8676 5404 8678
rect 5460 8676 5484 8678
rect 5540 8676 5564 8678
rect 5620 8676 5644 8678
rect 5700 8676 5706 8678
rect 5262 8664 5318 8673
rect 5398 8656 5706 8676
rect 5262 8599 5318 8608
rect 5276 8401 5304 8599
rect 5262 8392 5318 8401
rect 5262 8327 5318 8336
rect 5736 8090 5764 8842
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5262 7848 5318 7857
rect 5262 7783 5318 7792
rect 5276 7750 5304 7783
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5398 7644 5706 7664
rect 5398 7642 5404 7644
rect 5460 7642 5484 7644
rect 5540 7642 5564 7644
rect 5620 7642 5644 7644
rect 5700 7642 5706 7644
rect 5460 7590 5462 7642
rect 5642 7590 5644 7642
rect 5398 7588 5404 7590
rect 5460 7588 5484 7590
rect 5540 7588 5564 7590
rect 5620 7588 5644 7590
rect 5700 7588 5706 7590
rect 5398 7568 5706 7588
rect 5264 7540 5316 7546
rect 5264 7482 5316 7488
rect 5276 7041 5304 7482
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 5724 7472 5776 7478
rect 5724 7414 5776 7420
rect 5460 7177 5488 7414
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 7177 5672 7278
rect 5446 7168 5502 7177
rect 5446 7103 5502 7112
rect 5630 7168 5686 7177
rect 5630 7103 5686 7112
rect 5262 7032 5318 7041
rect 5262 6967 5318 6976
rect 5276 6304 5304 6967
rect 5398 6556 5706 6576
rect 5398 6554 5404 6556
rect 5460 6554 5484 6556
rect 5540 6554 5564 6556
rect 5620 6554 5644 6556
rect 5700 6554 5706 6556
rect 5460 6502 5462 6554
rect 5642 6502 5644 6554
rect 5398 6500 5404 6502
rect 5460 6500 5484 6502
rect 5540 6500 5564 6502
rect 5620 6500 5644 6502
rect 5700 6500 5706 6502
rect 5398 6480 5706 6500
rect 5356 6316 5408 6322
rect 5276 6276 5356 6304
rect 5356 6258 5408 6264
rect 5172 5908 5224 5914
rect 5224 5868 5304 5896
rect 5172 5850 5224 5856
rect 5078 5672 5134 5681
rect 4896 5636 4948 5642
rect 5078 5607 5134 5616
rect 4896 5578 4948 5584
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4908 4570 4936 5578
rect 4988 5364 5040 5370
rect 4988 5306 5040 5312
rect 4816 4542 4936 4570
rect 4816 4162 4844 4542
rect 4528 4140 4580 4146
rect 4528 4082 4580 4088
rect 4620 4140 4672 4146
rect 4816 4134 4936 4162
rect 4620 4082 4672 4088
rect 4528 3936 4580 3942
rect 4632 3924 4660 4082
rect 4580 3896 4660 3924
rect 4804 3936 4856 3942
rect 4710 3904 4766 3913
rect 4528 3878 4580 3884
rect 4804 3878 4856 3884
rect 4710 3839 4766 3848
rect 4436 3596 4488 3602
rect 4436 3538 4488 3544
rect 4724 3534 4752 3839
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4436 3460 4488 3466
rect 4436 3402 4488 3408
rect 4344 3120 4396 3126
rect 4344 3062 4396 3068
rect 4356 2689 4384 3062
rect 4342 2680 4398 2689
rect 4342 2615 4398 2624
rect 4448 2514 4476 3402
rect 4712 3052 4764 3058
rect 4816 3040 4844 3878
rect 4908 3058 4936 4134
rect 4764 3012 4844 3040
rect 4896 3052 4948 3058
rect 4712 2994 4764 3000
rect 4896 2994 4948 3000
rect 4528 2848 4580 2854
rect 4528 2790 4580 2796
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4252 2440 4304 2446
rect 4540 2394 4568 2790
rect 4252 2382 4304 2388
rect 4356 2378 4568 2394
rect 4344 2372 4568 2378
rect 4396 2366 4568 2372
rect 4344 2314 4396 2320
rect 4068 2100 4120 2106
rect 4068 2042 4120 2048
rect 4080 1873 4108 2042
rect 4632 2038 4660 2790
rect 5000 2446 5028 5306
rect 5092 4690 5120 5607
rect 5170 4720 5226 4729
rect 5080 4684 5132 4690
rect 5170 4655 5226 4664
rect 5080 4626 5132 4632
rect 5092 4282 5120 4626
rect 5184 4622 5212 4655
rect 5172 4616 5224 4622
rect 5172 4558 5224 4564
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 5184 4214 5212 4422
rect 5172 4208 5224 4214
rect 5078 4176 5134 4185
rect 5172 4150 5224 4156
rect 5078 4111 5134 4120
rect 5092 3466 5120 4111
rect 5276 4078 5304 5868
rect 5736 5574 5764 7414
rect 5828 5846 5856 8434
rect 5920 8022 5948 10678
rect 6012 8362 6040 11698
rect 6104 11257 6132 12038
rect 6288 11830 6316 12650
rect 6368 12232 6420 12238
rect 6368 12174 6420 12180
rect 6276 11824 6328 11830
rect 6276 11766 6328 11772
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6196 11558 6224 11698
rect 6276 11688 6328 11694
rect 6276 11630 6328 11636
rect 6184 11552 6236 11558
rect 6184 11494 6236 11500
rect 6090 11248 6146 11257
rect 6090 11183 6146 11192
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 10606 6132 11086
rect 6184 11076 6236 11082
rect 6184 11018 6236 11024
rect 6196 10810 6224 11018
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6092 10600 6144 10606
rect 6092 10542 6144 10548
rect 6288 10266 6316 11630
rect 6276 10260 6328 10266
rect 6276 10202 6328 10208
rect 6092 10124 6144 10130
rect 6092 10066 6144 10072
rect 6000 8356 6052 8362
rect 6000 8298 6052 8304
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5920 6458 5948 7754
rect 5998 7576 6054 7585
rect 5998 7511 6054 7520
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5816 5840 5868 5846
rect 5816 5782 5868 5788
rect 5920 5574 5948 6258
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5908 5568 5960 5574
rect 5908 5510 5960 5516
rect 5398 5468 5706 5488
rect 5398 5466 5404 5468
rect 5460 5466 5484 5468
rect 5540 5466 5564 5468
rect 5620 5466 5644 5468
rect 5700 5466 5706 5468
rect 5460 5414 5462 5466
rect 5642 5414 5644 5466
rect 5398 5412 5404 5414
rect 5460 5412 5484 5414
rect 5540 5412 5564 5414
rect 5620 5412 5644 5414
rect 5700 5412 5706 5414
rect 5398 5392 5706 5412
rect 5814 5400 5870 5409
rect 5814 5335 5870 5344
rect 5828 5302 5856 5335
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 6012 5137 6040 7511
rect 6104 6730 6132 10066
rect 6274 9616 6330 9625
rect 6274 9551 6330 9560
rect 6184 9376 6236 9382
rect 6184 9318 6236 9324
rect 6196 9042 6224 9318
rect 6184 9036 6236 9042
rect 6184 8978 6236 8984
rect 6288 8838 6316 9551
rect 6380 9518 6408 12174
rect 6472 11762 6500 12718
rect 6564 12345 6592 12922
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6748 12374 6776 12786
rect 6840 12714 6868 13670
rect 7024 13297 7052 14010
rect 7116 14006 7144 14583
rect 7208 14074 7236 15098
rect 7622 14716 7930 14736
rect 7622 14714 7628 14716
rect 7684 14714 7708 14716
rect 7764 14714 7788 14716
rect 7844 14714 7868 14716
rect 7924 14714 7930 14716
rect 7684 14662 7686 14714
rect 7866 14662 7868 14714
rect 7622 14660 7628 14662
rect 7684 14660 7708 14662
rect 7764 14660 7788 14662
rect 7844 14660 7868 14662
rect 7924 14660 7930 14662
rect 7622 14640 7930 14660
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 7196 14068 7248 14074
rect 7196 14010 7248 14016
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7392 13705 7420 14554
rect 8128 14074 8156 15438
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 10324 15428 10376 15434
rect 10324 15370 10376 15376
rect 8298 14104 8354 14113
rect 8116 14068 8168 14074
rect 8298 14039 8354 14048
rect 8116 14010 8168 14016
rect 8024 13864 8076 13870
rect 8128 13841 8156 14010
rect 8024 13806 8076 13812
rect 8114 13832 8170 13841
rect 7378 13696 7434 13705
rect 7378 13631 7434 13640
rect 7622 13628 7930 13648
rect 7622 13626 7628 13628
rect 7684 13626 7708 13628
rect 7764 13626 7788 13628
rect 7844 13626 7868 13628
rect 7924 13626 7930 13628
rect 7684 13574 7686 13626
rect 7866 13574 7868 13626
rect 7622 13572 7628 13574
rect 7684 13572 7708 13574
rect 7764 13572 7788 13574
rect 7844 13572 7868 13574
rect 7924 13572 7930 13574
rect 7622 13552 7930 13572
rect 8036 13530 8064 13806
rect 8114 13767 8170 13776
rect 8312 13530 8340 14039
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8300 13524 8352 13530
rect 8352 13484 8432 13512
rect 8300 13466 8352 13472
rect 7194 13424 7250 13433
rect 7194 13359 7196 13368
rect 7248 13359 7250 13368
rect 7196 13330 7248 13336
rect 7010 13288 7066 13297
rect 7300 13258 7328 13466
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8114 13288 8170 13297
rect 7010 13223 7066 13232
rect 7288 13252 7340 13258
rect 8114 13223 8170 13232
rect 7288 13194 7340 13200
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 7380 13184 7432 13190
rect 7380 13126 7432 13132
rect 7472 13184 7524 13190
rect 7748 13184 7800 13190
rect 7472 13126 7524 13132
rect 7746 13152 7748 13161
rect 8024 13184 8076 13190
rect 7800 13152 7802 13161
rect 6932 12986 6960 13126
rect 7010 13016 7066 13025
rect 6920 12980 6972 12986
rect 7010 12951 7066 12960
rect 6920 12922 6972 12928
rect 6828 12708 6880 12714
rect 6828 12650 6880 12656
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6840 12481 6868 12650
rect 6932 12617 6960 12650
rect 7024 12646 7052 12951
rect 7288 12912 7340 12918
rect 7116 12872 7288 12900
rect 7012 12640 7064 12646
rect 6918 12608 6974 12617
rect 7012 12582 7064 12588
rect 6918 12543 6974 12552
rect 7024 12481 7052 12582
rect 6826 12472 6882 12481
rect 6826 12407 6882 12416
rect 7010 12472 7066 12481
rect 7010 12407 7066 12416
rect 6736 12368 6788 12374
rect 6550 12336 6606 12345
rect 6736 12310 6788 12316
rect 6920 12368 6972 12374
rect 6920 12310 6972 12316
rect 6550 12271 6606 12280
rect 6644 12300 6696 12306
rect 6644 12242 6696 12248
rect 6552 12096 6604 12102
rect 6552 12038 6604 12044
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6460 11552 6512 11558
rect 6460 11494 6512 11500
rect 6472 10130 6500 11494
rect 6564 11121 6592 12038
rect 6550 11112 6606 11121
rect 6656 11082 6684 12242
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6550 11047 6606 11056
rect 6644 11076 6696 11082
rect 6644 11018 6696 11024
rect 6642 10840 6698 10849
rect 6642 10775 6698 10784
rect 6552 10668 6604 10674
rect 6552 10610 6604 10616
rect 6564 10305 6592 10610
rect 6550 10296 6606 10305
rect 6550 10231 6606 10240
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6472 9625 6500 9862
rect 6564 9654 6592 10134
rect 6552 9648 6604 9654
rect 6458 9616 6514 9625
rect 6552 9590 6604 9596
rect 6458 9551 6514 9560
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6380 9178 6408 9454
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6276 8832 6328 8838
rect 6276 8774 6328 8780
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6092 6724 6144 6730
rect 6092 6666 6144 6672
rect 6196 5778 6224 8366
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6288 8090 6316 8230
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6380 7546 6408 8230
rect 6472 7750 6500 9551
rect 6656 9500 6684 10775
rect 6748 10266 6776 11698
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6840 11014 6868 11562
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10606 6868 10950
rect 6932 10674 6960 12310
rect 7116 12186 7144 12872
rect 7288 12854 7340 12860
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 7208 12374 7236 12718
rect 7196 12368 7248 12374
rect 7392 12345 7420 13126
rect 7484 12442 7512 13126
rect 8024 13126 8076 13132
rect 7746 13087 7802 13096
rect 7622 12540 7930 12560
rect 7622 12538 7628 12540
rect 7684 12538 7708 12540
rect 7764 12538 7788 12540
rect 7844 12538 7868 12540
rect 7924 12538 7930 12540
rect 7684 12486 7686 12538
rect 7866 12486 7868 12538
rect 7622 12484 7628 12486
rect 7684 12484 7708 12486
rect 7764 12484 7788 12486
rect 7844 12484 7868 12486
rect 7924 12484 7930 12486
rect 7622 12464 7930 12484
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7196 12310 7248 12316
rect 7378 12336 7434 12345
rect 7378 12271 7434 12280
rect 7562 12336 7618 12345
rect 7562 12271 7618 12280
rect 7656 12300 7708 12306
rect 7288 12232 7340 12238
rect 7116 12158 7236 12186
rect 7288 12174 7340 12180
rect 7472 12232 7524 12238
rect 7472 12174 7524 12180
rect 7104 12096 7156 12102
rect 7104 12038 7156 12044
rect 7012 11824 7064 11830
rect 7012 11766 7064 11772
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 6828 10600 6880 10606
rect 6828 10542 6880 10548
rect 6828 10464 6880 10470
rect 6828 10406 6880 10412
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6840 10062 6868 10406
rect 6932 10169 6960 10406
rect 6918 10160 6974 10169
rect 6918 10095 6974 10104
rect 6828 10056 6880 10062
rect 6828 9998 6880 10004
rect 6920 9920 6972 9926
rect 6826 9888 6882 9897
rect 6920 9862 6972 9868
rect 6826 9823 6882 9832
rect 6564 9472 6684 9500
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6368 7540 6420 7546
rect 6368 7482 6420 7488
rect 6276 6928 6328 6934
rect 6274 6896 6276 6905
rect 6328 6896 6330 6905
rect 6274 6831 6330 6840
rect 6380 6254 6408 7482
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 6458 6500 6598
rect 6460 6452 6512 6458
rect 6460 6394 6512 6400
rect 6368 6248 6420 6254
rect 6368 6190 6420 6196
rect 6184 5772 6236 5778
rect 6184 5714 6236 5720
rect 6564 5692 6592 9472
rect 6840 9466 6868 9823
rect 6932 9761 6960 9862
rect 6918 9752 6974 9761
rect 6918 9687 6974 9696
rect 6840 9438 6960 9466
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6644 9104 6696 9110
rect 6644 9046 6696 9052
rect 6656 7721 6684 9046
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8362 6776 8910
rect 6840 8906 6868 9318
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6840 8566 6868 8842
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6736 8356 6788 8362
rect 6736 8298 6788 8304
rect 6642 7712 6698 7721
rect 6642 7647 6698 7656
rect 6656 7002 6684 7647
rect 6644 6996 6696 7002
rect 6644 6938 6696 6944
rect 6748 6934 6776 8298
rect 6840 7478 6868 8502
rect 6932 7954 6960 9438
rect 7024 8022 7052 11766
rect 7116 9654 7144 12038
rect 7208 10538 7236 12158
rect 7300 12073 7328 12174
rect 7286 12064 7342 12073
rect 7286 11999 7342 12008
rect 7286 11792 7342 11801
rect 7286 11727 7342 11736
rect 7300 11694 7328 11727
rect 7288 11688 7340 11694
rect 7288 11630 7340 11636
rect 7484 11608 7512 12174
rect 7576 12102 7604 12271
rect 7656 12242 7708 12248
rect 7564 12096 7616 12102
rect 7564 12038 7616 12044
rect 7668 11762 7696 12242
rect 7748 12096 7800 12102
rect 7748 12038 7800 12044
rect 7760 11830 7788 12038
rect 8036 11914 8064 13126
rect 8128 12918 8156 13223
rect 8312 12918 8340 13330
rect 8116 12912 8168 12918
rect 8116 12854 8168 12860
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8404 12850 8432 13484
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8116 12776 8168 12782
rect 8496 12730 8524 15370
rect 8758 15056 8814 15065
rect 8758 14991 8814 15000
rect 8576 14272 8628 14278
rect 8576 14214 8628 14220
rect 8588 13802 8616 14214
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13530 8616 13738
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8116 12718 8168 12724
rect 8128 12617 8156 12718
rect 8404 12702 8524 12730
rect 8114 12608 8170 12617
rect 8114 12543 8170 12552
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8128 11937 8156 12106
rect 7944 11886 8064 11914
rect 8114 11928 8170 11937
rect 7748 11824 7800 11830
rect 7748 11766 7800 11772
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7944 11626 7972 11886
rect 8114 11863 8170 11872
rect 8024 11824 8076 11830
rect 8022 11792 8024 11801
rect 8076 11792 8078 11801
rect 8022 11727 8078 11736
rect 8024 11688 8076 11694
rect 8024 11630 8076 11636
rect 7392 11580 7512 11608
rect 7932 11620 7984 11626
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 10810 7328 11494
rect 7392 11268 7420 11580
rect 7932 11562 7984 11568
rect 7622 11452 7930 11472
rect 7622 11450 7628 11452
rect 7684 11450 7708 11452
rect 7764 11450 7788 11452
rect 7844 11450 7868 11452
rect 7924 11450 7930 11452
rect 7684 11398 7686 11450
rect 7866 11398 7868 11450
rect 7622 11396 7628 11398
rect 7684 11396 7708 11398
rect 7764 11396 7788 11398
rect 7844 11396 7868 11398
rect 7924 11396 7930 11398
rect 7622 11376 7930 11396
rect 7392 11240 7512 11268
rect 7484 11014 7512 11240
rect 8036 11218 8064 11630
rect 8024 11212 8076 11218
rect 8024 11154 8076 11160
rect 7472 11008 7524 11014
rect 7472 10950 7524 10956
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7196 10532 7248 10538
rect 7196 10474 7248 10480
rect 7378 10432 7434 10441
rect 7378 10367 7434 10376
rect 7286 10296 7342 10305
rect 7286 10231 7342 10240
rect 7194 10160 7250 10169
rect 7194 10095 7250 10104
rect 7104 9648 7156 9654
rect 7104 9590 7156 9596
rect 7208 8294 7236 10095
rect 7300 8673 7328 10231
rect 7392 10010 7420 10367
rect 7484 10130 7512 10950
rect 7576 10742 7604 10950
rect 7564 10736 7616 10742
rect 7564 10678 7616 10684
rect 7622 10364 7930 10384
rect 7622 10362 7628 10364
rect 7684 10362 7708 10364
rect 7764 10362 7788 10364
rect 7844 10362 7868 10364
rect 7924 10362 7930 10364
rect 7684 10310 7686 10362
rect 7866 10310 7868 10362
rect 7622 10308 7628 10310
rect 7684 10308 7708 10310
rect 7764 10308 7788 10310
rect 7844 10308 7868 10310
rect 7924 10308 7930 10310
rect 7622 10288 7930 10308
rect 8036 10130 8064 11154
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10849 8156 11018
rect 8114 10840 8170 10849
rect 8114 10775 8170 10784
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8128 10266 8156 10406
rect 8116 10260 8168 10266
rect 8116 10202 8168 10208
rect 7472 10124 7524 10130
rect 7472 10066 7524 10072
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 7392 9982 7512 10010
rect 7378 9480 7434 9489
rect 7484 9466 7512 9982
rect 7576 9722 7604 10066
rect 7748 9920 7800 9926
rect 7654 9888 7710 9897
rect 7748 9862 7800 9868
rect 7654 9823 7710 9832
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7668 9586 7696 9823
rect 7760 9761 7788 9862
rect 7746 9752 7802 9761
rect 7746 9687 7802 9696
rect 7930 9752 7986 9761
rect 7930 9687 7986 9696
rect 8116 9716 8168 9722
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7562 9480 7618 9489
rect 7484 9438 7562 9466
rect 7378 9415 7434 9424
rect 7852 9466 7880 9522
rect 7562 9415 7618 9424
rect 7668 9438 7880 9466
rect 7944 9450 7972 9687
rect 8116 9658 8168 9664
rect 8024 9580 8076 9586
rect 8024 9522 8076 9528
rect 7932 9444 7984 9450
rect 7286 8664 7342 8673
rect 7286 8599 7342 8608
rect 7104 8288 7156 8294
rect 7208 8266 7328 8294
rect 7104 8230 7156 8236
rect 7012 8016 7064 8022
rect 7012 7958 7064 7964
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6932 7698 6960 7890
rect 7116 7886 7144 8230
rect 7104 7880 7156 7886
rect 7104 7822 7156 7828
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7104 7744 7156 7750
rect 6932 7670 7052 7698
rect 7104 7686 7156 7692
rect 6920 7540 6972 7546
rect 6920 7482 6972 7488
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6840 6866 6868 7414
rect 6828 6860 6880 6866
rect 6828 6802 6880 6808
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 6644 5704 6696 5710
rect 6564 5664 6644 5692
rect 6644 5646 6696 5652
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 5998 5128 6054 5137
rect 5998 5063 6054 5072
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5368 4622 5396 4966
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5398 4380 5706 4400
rect 5398 4378 5404 4380
rect 5460 4378 5484 4380
rect 5540 4378 5564 4380
rect 5620 4378 5644 4380
rect 5700 4378 5706 4380
rect 5460 4326 5462 4378
rect 5642 4326 5644 4378
rect 5398 4324 5404 4326
rect 5460 4324 5484 4326
rect 5540 4324 5564 4326
rect 5620 4324 5644 4326
rect 5700 4324 5706 4326
rect 5398 4304 5706 4324
rect 5264 4072 5316 4078
rect 5170 4040 5226 4049
rect 5264 4014 5316 4020
rect 5908 4072 5960 4078
rect 5908 4014 5960 4020
rect 5170 3975 5226 3984
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 4894 2272 4950 2281
rect 4894 2207 4950 2216
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 4066 1864 4122 1873
rect 4066 1799 4122 1808
rect 4068 1760 4120 1766
rect 4068 1702 4120 1708
rect 4080 1465 4108 1702
rect 4066 1456 4122 1465
rect 4066 1391 4122 1400
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 4080 1193 4108 1294
rect 4066 1184 4122 1193
rect 4066 1119 4122 1128
rect 4908 800 4936 2207
rect 5184 1970 5212 3975
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5276 3058 5304 3703
rect 5398 3292 5706 3312
rect 5398 3290 5404 3292
rect 5460 3290 5484 3292
rect 5540 3290 5564 3292
rect 5620 3290 5644 3292
rect 5700 3290 5706 3292
rect 5460 3238 5462 3290
rect 5642 3238 5644 3290
rect 5398 3236 5404 3238
rect 5460 3236 5484 3238
rect 5540 3236 5564 3238
rect 5620 3236 5644 3238
rect 5700 3236 5706 3238
rect 5398 3216 5706 3236
rect 5814 3224 5870 3233
rect 5814 3159 5870 3168
rect 5828 3126 5856 3159
rect 5816 3120 5868 3126
rect 5816 3062 5868 3068
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5816 2984 5868 2990
rect 5816 2926 5868 2932
rect 5460 2854 5488 2926
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5460 2514 5488 2790
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5398 2204 5706 2224
rect 5398 2202 5404 2204
rect 5460 2202 5484 2204
rect 5540 2202 5564 2204
rect 5620 2202 5644 2204
rect 5700 2202 5706 2204
rect 5460 2150 5462 2202
rect 5642 2150 5644 2202
rect 5398 2148 5404 2150
rect 5460 2148 5484 2150
rect 5540 2148 5564 2150
rect 5620 2148 5644 2150
rect 5700 2148 5706 2150
rect 5262 2136 5318 2145
rect 5398 2128 5706 2148
rect 5262 2071 5318 2080
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 5276 1737 5304 2071
rect 5262 1728 5318 1737
rect 5262 1663 5318 1672
rect 5828 1465 5856 2926
rect 5920 2650 5948 4014
rect 6012 3942 6040 4966
rect 6104 4078 6132 5510
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 6196 4457 6224 5306
rect 6460 5160 6512 5166
rect 6458 5128 6460 5137
rect 6512 5128 6514 5137
rect 6458 5063 6514 5072
rect 6552 4548 6604 4554
rect 6552 4490 6604 4496
rect 6182 4448 6238 4457
rect 6182 4383 6238 4392
rect 6092 4072 6144 4078
rect 6092 4014 6144 4020
rect 6000 3936 6052 3942
rect 6000 3878 6052 3884
rect 6012 2990 6040 3878
rect 6104 3602 6132 4014
rect 6368 3936 6420 3942
rect 6368 3878 6420 3884
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 6274 3496 6330 3505
rect 6274 3431 6330 3440
rect 6092 3392 6144 3398
rect 6092 3334 6144 3340
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 6012 2854 6040 2926
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5908 2644 5960 2650
rect 5908 2586 5960 2592
rect 6104 2514 6132 3334
rect 6184 2576 6236 2582
rect 6182 2544 6184 2553
rect 6236 2544 6238 2553
rect 6092 2508 6144 2514
rect 6182 2479 6238 2488
rect 6092 2450 6144 2456
rect 6104 2038 6132 2450
rect 6092 2032 6144 2038
rect 6092 1974 6144 1980
rect 5814 1456 5870 1465
rect 5814 1391 5870 1400
rect 5828 870 5948 898
rect 5828 800 5856 870
rect 3422 776 3478 785
rect 3422 711 3478 720
rect 3700 672 3752 678
rect 3700 614 3752 620
rect 3712 513 3740 614
rect 3698 504 3754 513
rect 3698 439 3754 448
rect 3974 0 4030 800
rect 4894 0 4950 800
rect 5814 0 5870 800
rect 5920 762 5948 870
rect 6288 762 6316 3431
rect 6380 2514 6408 3878
rect 6564 3670 6592 4490
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 6656 3369 6684 5646
rect 6840 5234 6868 6287
rect 6932 6118 6960 7482
rect 7024 6662 7052 7670
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7116 6390 7144 7686
rect 7208 7002 7236 7754
rect 7196 6996 7248 7002
rect 7196 6938 7248 6944
rect 7104 6384 7156 6390
rect 7104 6326 7156 6332
rect 7012 6248 7064 6254
rect 7012 6190 7064 6196
rect 6920 6112 6972 6118
rect 6920 6054 6972 6060
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6828 5228 6880 5234
rect 6828 5170 6880 5176
rect 6736 4140 6788 4146
rect 6736 4082 6788 4088
rect 6642 3360 6698 3369
rect 6642 3295 6698 3304
rect 6748 3194 6776 4082
rect 6840 3913 6868 5170
rect 6932 4758 6960 5850
rect 6920 4752 6972 4758
rect 6920 4694 6972 4700
rect 6826 3904 6882 3913
rect 6826 3839 6882 3848
rect 6918 3496 6974 3505
rect 6918 3431 6974 3440
rect 6932 3194 6960 3431
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6734 3088 6790 3097
rect 6734 3023 6790 3032
rect 6918 3088 6974 3097
rect 7024 3058 7052 6190
rect 7300 5370 7328 8266
rect 7392 7886 7420 9415
rect 7668 9364 7696 9438
rect 7932 9386 7984 9392
rect 7484 9353 7696 9364
rect 7470 9344 7696 9353
rect 7526 9336 7696 9344
rect 7470 9279 7526 9288
rect 7484 8809 7512 9279
rect 7622 9276 7930 9296
rect 7622 9274 7628 9276
rect 7684 9274 7708 9276
rect 7764 9274 7788 9276
rect 7844 9274 7868 9276
rect 7924 9274 7930 9276
rect 7684 9222 7686 9274
rect 7866 9222 7868 9274
rect 7622 9220 7628 9222
rect 7684 9220 7708 9222
rect 7764 9220 7788 9222
rect 7844 9220 7868 9222
rect 7924 9220 7930 9222
rect 7622 9200 7930 9220
rect 8036 9178 8064 9522
rect 8024 9172 8076 9178
rect 8024 9114 8076 9120
rect 8128 8945 8156 9658
rect 7746 8936 7802 8945
rect 7564 8900 7616 8906
rect 7746 8871 7802 8880
rect 8114 8936 8170 8945
rect 8114 8871 8170 8880
rect 7564 8842 7616 8848
rect 7470 8800 7526 8809
rect 7470 8735 7526 8744
rect 7576 8673 7604 8842
rect 7562 8664 7618 8673
rect 7562 8599 7618 8608
rect 7760 8276 7788 8871
rect 8114 8800 8170 8809
rect 8114 8735 8170 8744
rect 7484 8265 7788 8276
rect 7470 8256 7788 8265
rect 7526 8248 7788 8256
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7470 8191 7526 8200
rect 7484 7970 7512 8191
rect 7622 8188 7930 8208
rect 7622 8186 7628 8188
rect 7684 8186 7708 8188
rect 7764 8186 7788 8188
rect 7844 8186 7868 8188
rect 7924 8186 7930 8188
rect 7684 8134 7686 8186
rect 7866 8134 7868 8186
rect 7622 8132 7628 8134
rect 7684 8132 7708 8134
rect 7764 8132 7788 8134
rect 7844 8132 7868 8134
rect 7924 8132 7930 8134
rect 7622 8112 7930 8132
rect 7840 8016 7892 8022
rect 7484 7942 7696 7970
rect 7840 7958 7892 7964
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7380 7880 7432 7886
rect 7564 7880 7616 7886
rect 7380 7822 7432 7828
rect 7484 7840 7564 7868
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7392 5409 7420 6598
rect 7484 6458 7512 7840
rect 7564 7822 7616 7828
rect 7668 7818 7696 7942
rect 7748 7948 7800 7954
rect 7748 7890 7800 7896
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7656 7404 7708 7410
rect 7760 7392 7788 7890
rect 7852 7410 7880 7958
rect 7944 7750 7972 7958
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7930 7576 7986 7585
rect 7930 7511 7986 7520
rect 7944 7478 7972 7511
rect 7932 7472 7984 7478
rect 7932 7414 7984 7420
rect 7708 7364 7788 7392
rect 7840 7404 7892 7410
rect 7656 7346 7708 7352
rect 7840 7346 7892 7352
rect 7932 7336 7984 7342
rect 8036 7324 8064 8230
rect 7984 7296 8064 7324
rect 7932 7278 7984 7284
rect 7622 7100 7930 7120
rect 7622 7098 7628 7100
rect 7684 7098 7708 7100
rect 7764 7098 7788 7100
rect 7844 7098 7868 7100
rect 7924 7098 7930 7100
rect 7684 7046 7686 7098
rect 7866 7046 7868 7098
rect 7622 7044 7628 7046
rect 7684 7044 7708 7046
rect 7764 7044 7788 7046
rect 7844 7044 7868 7046
rect 7924 7044 7930 7046
rect 7622 7024 7930 7044
rect 8036 6984 8064 7296
rect 7852 6956 8064 6984
rect 7564 6928 7616 6934
rect 7564 6870 7616 6876
rect 7576 6798 7604 6870
rect 7564 6792 7616 6798
rect 7564 6734 7616 6740
rect 7562 6488 7618 6497
rect 7472 6452 7524 6458
rect 7562 6423 7618 6432
rect 7472 6394 7524 6400
rect 7576 6322 7604 6423
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7852 6254 7880 6956
rect 8128 6916 8156 8735
rect 8312 8537 8340 12174
rect 8404 12084 8432 12702
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12186 8524 12582
rect 8588 12442 8616 13466
rect 8772 12918 8800 14991
rect 9402 14648 9458 14657
rect 9402 14583 9458 14592
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 13530 9076 14214
rect 9312 14068 9364 14074
rect 9312 14010 9364 14016
rect 9324 13938 9352 14010
rect 9416 14006 9444 14583
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14340 9732 14346
rect 9680 14282 9732 14288
rect 9404 14000 9456 14006
rect 9404 13942 9456 13948
rect 9312 13932 9364 13938
rect 9692 13920 9720 14282
rect 9784 14074 9812 14350
rect 10230 14240 10286 14249
rect 9846 14172 10154 14192
rect 10230 14175 10286 14184
rect 9846 14170 9852 14172
rect 9908 14170 9932 14172
rect 9988 14170 10012 14172
rect 10068 14170 10092 14172
rect 10148 14170 10154 14172
rect 9908 14118 9910 14170
rect 10090 14118 10092 14170
rect 9846 14116 9852 14118
rect 9908 14116 9932 14118
rect 9988 14116 10012 14118
rect 10068 14116 10092 14118
rect 10148 14116 10154 14118
rect 9846 14096 10154 14116
rect 9772 14068 9824 14074
rect 9772 14010 9824 14016
rect 10244 14006 10272 14175
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 9772 13932 9824 13938
rect 9692 13892 9772 13920
rect 9312 13874 9364 13880
rect 9772 13874 9824 13880
rect 9404 13864 9456 13870
rect 9404 13806 9456 13812
rect 9416 13705 9444 13806
rect 9402 13696 9458 13705
rect 9402 13631 9458 13640
rect 9036 13524 9088 13530
rect 8956 13484 9036 13512
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8850 12880 8906 12889
rect 8850 12815 8852 12824
rect 8904 12815 8906 12824
rect 8852 12786 8904 12792
rect 8576 12436 8628 12442
rect 8576 12378 8628 12384
rect 8496 12158 8708 12186
rect 8484 12096 8536 12102
rect 8404 12056 8484 12084
rect 8484 12038 8536 12044
rect 8392 11688 8444 11694
rect 8392 11630 8444 11636
rect 8404 11150 8432 11630
rect 8496 11150 8524 12038
rect 8392 11144 8444 11150
rect 8392 11086 8444 11092
rect 8484 11144 8536 11150
rect 8484 11086 8536 11092
rect 8392 11008 8444 11014
rect 8390 10976 8392 10985
rect 8576 11008 8628 11014
rect 8444 10976 8446 10985
rect 8576 10950 8628 10956
rect 8390 10911 8446 10920
rect 8390 10568 8446 10577
rect 8390 10503 8446 10512
rect 8484 10532 8536 10538
rect 8404 10062 8432 10503
rect 8484 10474 8536 10480
rect 8496 10130 8524 10474
rect 8484 10124 8536 10130
rect 8484 10066 8536 10072
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8404 8974 8432 9998
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8496 8634 8524 9590
rect 8588 9081 8616 10950
rect 8680 10713 8708 12158
rect 8852 11756 8904 11762
rect 8852 11698 8904 11704
rect 8864 11014 8892 11698
rect 8956 11286 8984 13484
rect 9036 13466 9088 13472
rect 9310 13424 9366 13433
rect 9310 13359 9366 13368
rect 9494 13424 9550 13433
rect 9494 13359 9550 13368
rect 9036 12912 9088 12918
rect 9034 12880 9036 12889
rect 9088 12880 9090 12889
rect 9034 12815 9090 12824
rect 9220 12096 9272 12102
rect 9220 12038 9272 12044
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 8944 11280 8996 11286
rect 8944 11222 8996 11228
rect 8944 11144 8996 11150
rect 8944 11086 8996 11092
rect 8852 11008 8904 11014
rect 8852 10950 8904 10956
rect 8666 10704 8722 10713
rect 8666 10639 8722 10648
rect 8760 10668 8812 10674
rect 8760 10610 8812 10616
rect 8772 10266 8800 10610
rect 8864 10606 8892 10950
rect 8852 10600 8904 10606
rect 8852 10542 8904 10548
rect 8956 10305 8984 11086
rect 8942 10296 8998 10305
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8852 10260 8904 10266
rect 8942 10231 8998 10240
rect 8852 10202 8904 10208
rect 8864 10146 8892 10202
rect 8864 10118 8984 10146
rect 8758 10024 8814 10033
rect 8668 9988 8720 9994
rect 8758 9959 8814 9968
rect 8668 9930 8720 9936
rect 8680 9722 8708 9930
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 8574 9072 8630 9081
rect 8574 9007 8630 9016
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8298 8528 8354 8537
rect 8298 8463 8354 8472
rect 8588 8129 8616 8910
rect 8680 8838 8708 9522
rect 8772 8974 8800 9959
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8574 8120 8630 8129
rect 8574 8055 8630 8064
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8206 7712 8262 7721
rect 8206 7647 8262 7656
rect 8220 7154 8248 7647
rect 8220 7126 8294 7154
rect 8266 7002 8294 7126
rect 8254 6996 8306 7002
rect 8254 6938 8306 6944
rect 8404 6934 8432 7890
rect 8484 7200 8536 7206
rect 8484 7142 8536 7148
rect 8067 6888 8156 6916
rect 8392 6928 8444 6934
rect 8067 6882 8095 6888
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 8036 6854 8095 6882
rect 8392 6870 8444 6876
rect 8496 6866 8524 7142
rect 8484 6860 8536 6866
rect 7944 6730 7972 6802
rect 7932 6724 7984 6730
rect 7932 6666 7984 6672
rect 8036 6361 8064 6854
rect 8484 6802 8536 6808
rect 8680 6798 8708 8774
rect 8668 6792 8720 6798
rect 8668 6734 8720 6740
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8022 6352 8078 6361
rect 8022 6287 8078 6296
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7622 6012 7930 6032
rect 7622 6010 7628 6012
rect 7684 6010 7708 6012
rect 7764 6010 7788 6012
rect 7844 6010 7868 6012
rect 7924 6010 7930 6012
rect 7684 5958 7686 6010
rect 7866 5958 7868 6010
rect 7622 5956 7628 5958
rect 7684 5956 7708 5958
rect 7764 5956 7788 5958
rect 7844 5956 7868 5958
rect 7924 5956 7930 5958
rect 7622 5936 7930 5956
rect 8128 5778 8156 6598
rect 8404 6458 8432 6598
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8116 5772 8168 5778
rect 8116 5714 8168 5720
rect 8312 5710 8340 6054
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8116 5636 8168 5642
rect 8116 5578 8168 5584
rect 7378 5400 7434 5409
rect 7288 5364 7340 5370
rect 7208 5324 7288 5352
rect 7102 4856 7158 4865
rect 7102 4791 7158 4800
rect 6918 3023 6974 3032
rect 7012 3052 7064 3058
rect 6644 2916 6696 2922
rect 6644 2858 6696 2864
rect 6656 2689 6684 2858
rect 6642 2680 6698 2689
rect 6642 2615 6698 2624
rect 6642 2544 6698 2553
rect 6368 2508 6420 2514
rect 6642 2479 6698 2488
rect 6368 2450 6420 2456
rect 6656 2446 6684 2479
rect 6644 2440 6696 2446
rect 6644 2382 6696 2388
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 5920 734 6316 762
rect 6472 678 6500 2246
rect 6748 800 6776 3023
rect 6932 2825 6960 3023
rect 7012 2994 7064 3000
rect 6918 2816 6974 2825
rect 7116 2774 7144 4791
rect 7208 3233 7236 5324
rect 7378 5335 7434 5344
rect 7288 5306 7340 5312
rect 8128 5166 8156 5578
rect 7472 5160 7524 5166
rect 7472 5102 7524 5108
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 7380 5024 7432 5030
rect 7484 5001 7512 5102
rect 8024 5024 8076 5030
rect 7380 4966 7432 4972
rect 7470 4992 7526 5001
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7194 3224 7250 3233
rect 7194 3159 7196 3168
rect 7248 3159 7250 3168
rect 7196 3130 7248 3136
rect 7208 3099 7236 3130
rect 7196 2984 7248 2990
rect 7300 2972 7328 4422
rect 7392 3534 7420 4966
rect 8024 4966 8076 4972
rect 7470 4927 7526 4936
rect 7622 4924 7930 4944
rect 7622 4922 7628 4924
rect 7684 4922 7708 4924
rect 7764 4922 7788 4924
rect 7844 4922 7868 4924
rect 7924 4922 7930 4924
rect 7684 4870 7686 4922
rect 7866 4870 7868 4922
rect 7622 4868 7628 4870
rect 7684 4868 7708 4870
rect 7764 4868 7788 4870
rect 7844 4868 7868 4870
rect 7924 4868 7930 4870
rect 7622 4848 7930 4868
rect 8036 4826 8064 4966
rect 8024 4820 8076 4826
rect 8024 4762 8076 4768
rect 8024 4140 8076 4146
rect 8024 4082 8076 4088
rect 7622 3836 7930 3856
rect 7622 3834 7628 3836
rect 7684 3834 7708 3836
rect 7764 3834 7788 3836
rect 7844 3834 7868 3836
rect 7924 3834 7930 3836
rect 7684 3782 7686 3834
rect 7866 3782 7868 3834
rect 7622 3780 7628 3782
rect 7684 3780 7708 3782
rect 7764 3780 7788 3782
rect 7844 3780 7868 3782
rect 7924 3780 7930 3782
rect 7470 3768 7526 3777
rect 7622 3760 7930 3780
rect 7470 3703 7526 3712
rect 7484 3584 7512 3703
rect 7484 3556 7604 3584
rect 7380 3528 7432 3534
rect 7380 3470 7432 3476
rect 7576 3398 7604 3556
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7930 3360 7986 3369
rect 7930 3295 7986 3304
rect 7944 3058 7972 3295
rect 7932 3052 7984 3058
rect 7932 2994 7984 3000
rect 7380 2984 7432 2990
rect 7300 2944 7380 2972
rect 7196 2926 7248 2932
rect 7840 2984 7892 2990
rect 7380 2926 7432 2932
rect 7484 2944 7840 2972
rect 7208 2854 7236 2926
rect 7196 2848 7248 2854
rect 6918 2751 6974 2760
rect 7024 2746 7144 2774
rect 7194 2816 7196 2825
rect 7248 2816 7250 2825
rect 7194 2751 7250 2760
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 6840 1970 6868 2450
rect 7024 2310 7052 2746
rect 7102 2680 7158 2689
rect 7102 2615 7158 2624
rect 7116 2310 7144 2615
rect 7208 2582 7236 2751
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 7392 2514 7420 2926
rect 7380 2508 7432 2514
rect 7380 2450 7432 2456
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 7024 1698 7052 2246
rect 7012 1692 7064 1698
rect 7012 1634 7064 1640
rect 7116 1562 7144 2246
rect 7104 1556 7156 1562
rect 7484 1544 7512 2944
rect 7840 2926 7892 2932
rect 7622 2748 7930 2768
rect 7622 2746 7628 2748
rect 7684 2746 7708 2748
rect 7764 2746 7788 2748
rect 7844 2746 7868 2748
rect 7924 2746 7930 2748
rect 7684 2694 7686 2746
rect 7866 2694 7868 2746
rect 7622 2692 7628 2694
rect 7684 2692 7708 2694
rect 7764 2692 7788 2694
rect 7844 2692 7868 2694
rect 7924 2692 7930 2694
rect 7622 2672 7930 2692
rect 8036 2689 8064 4082
rect 8128 3602 8156 5102
rect 8312 4690 8340 5646
rect 8588 5370 8616 5782
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8680 5302 8708 6598
rect 8772 5817 8800 8774
rect 8864 7546 8892 8842
rect 8852 7540 8904 7546
rect 8852 7482 8904 7488
rect 8758 5808 8814 5817
rect 8758 5743 8814 5752
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8668 5296 8720 5302
rect 8668 5238 8720 5244
rect 8758 5264 8814 5273
rect 8496 5030 8524 5238
rect 8758 5199 8814 5208
rect 8484 5024 8536 5030
rect 8484 4966 8536 4972
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8208 4548 8260 4554
rect 8208 4490 8260 4496
rect 8220 4185 8248 4490
rect 8206 4176 8262 4185
rect 8312 4146 8340 4626
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8206 4111 8262 4120
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8206 3904 8262 3913
rect 8206 3839 8262 3848
rect 8220 3670 8248 3839
rect 8208 3664 8260 3670
rect 8208 3606 8260 3612
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8022 2680 8078 2689
rect 8022 2615 8078 2624
rect 8128 2514 8156 3538
rect 8220 3233 8248 3606
rect 8312 3602 8340 4082
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8206 3224 8262 3233
rect 8312 3194 8340 3538
rect 8206 3159 8262 3168
rect 8300 3188 8352 3194
rect 8300 3130 8352 3136
rect 8254 2916 8306 2922
rect 8254 2858 8306 2864
rect 8266 2774 8294 2858
rect 8220 2746 8294 2774
rect 8220 2582 8248 2746
rect 8208 2576 8260 2582
rect 8208 2518 8260 2524
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7944 1630 7972 2246
rect 8404 1766 8432 4422
rect 8496 4146 8524 4966
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8484 3732 8536 3738
rect 8484 3674 8536 3680
rect 8496 3398 8524 3674
rect 8484 3392 8536 3398
rect 8484 3334 8536 3340
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8496 2990 8524 3130
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 8496 2281 8524 2382
rect 8668 2304 8720 2310
rect 8482 2272 8538 2281
rect 8668 2246 8720 2252
rect 8482 2207 8538 2216
rect 8680 2106 8708 2246
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 8392 1760 8444 1766
rect 8392 1702 8444 1708
rect 7932 1624 7984 1630
rect 7932 1566 7984 1572
rect 7484 1516 7604 1544
rect 7104 1498 7156 1504
rect 7576 800 7604 1516
rect 8496 870 8616 898
rect 8496 800 8524 870
rect 6460 672 6512 678
rect 6460 614 6512 620
rect 6734 0 6790 800
rect 7562 0 7618 800
rect 8482 0 8538 800
rect 8588 762 8616 870
rect 8772 762 8800 5199
rect 8956 4622 8984 10118
rect 9048 5817 9076 11494
rect 9140 10674 9168 11766
rect 9128 10668 9180 10674
rect 9128 10610 9180 10616
rect 9126 10296 9182 10305
rect 9126 10231 9182 10240
rect 9140 6610 9168 10231
rect 9232 7993 9260 12038
rect 9324 11354 9352 13359
rect 9508 12986 9536 13359
rect 10232 13320 10284 13326
rect 10232 13262 10284 13268
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 9496 12980 9548 12986
rect 9496 12922 9548 12928
rect 9600 12918 9628 13087
rect 9846 13084 10154 13104
rect 9846 13082 9852 13084
rect 9908 13082 9932 13084
rect 9988 13082 10012 13084
rect 10068 13082 10092 13084
rect 10148 13082 10154 13084
rect 9908 13030 9910 13082
rect 10090 13030 10092 13082
rect 9846 13028 9852 13030
rect 9908 13028 9932 13030
rect 9988 13028 10012 13030
rect 10068 13028 10092 13030
rect 10148 13028 10154 13030
rect 9678 13016 9734 13025
rect 9846 13008 10154 13028
rect 9678 12951 9734 12960
rect 9588 12912 9640 12918
rect 9588 12854 9640 12860
rect 9404 12844 9456 12850
rect 9404 12786 9456 12792
rect 9416 12374 9444 12786
rect 9692 12442 9720 12951
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9770 12472 9826 12481
rect 9588 12436 9640 12442
rect 9588 12378 9640 12384
rect 9680 12436 9732 12442
rect 9732 12416 9770 12434
rect 9968 12434 9996 12718
rect 10138 12608 10194 12617
rect 10138 12543 10194 12552
rect 10152 12442 10180 12543
rect 10244 12442 10272 13262
rect 10336 12986 10364 15370
rect 10428 14278 10456 16510
rect 13910 16400 13966 17200
rect 15658 16960 15714 16969
rect 15658 16895 15714 16904
rect 13924 15502 13952 16400
rect 14832 15836 14884 15842
rect 14832 15778 14884 15784
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 10874 15192 10930 15201
rect 10508 15156 10560 15162
rect 10874 15127 10930 15136
rect 10508 15098 10560 15104
rect 10416 14272 10468 14278
rect 10416 14214 10468 14220
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10428 12986 10456 13466
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 9732 12407 9826 12416
rect 9732 12406 9812 12407
rect 9876 12406 9996 12434
rect 10140 12436 10192 12442
rect 9680 12378 9732 12384
rect 9404 12368 9456 12374
rect 9404 12310 9456 12316
rect 9600 12102 9628 12378
rect 9876 12322 9904 12406
rect 10140 12378 10192 12384
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 9784 12294 9904 12322
rect 10048 12368 10100 12374
rect 10336 12345 10364 12922
rect 10428 12374 10456 12922
rect 10416 12368 10468 12374
rect 10048 12310 10100 12316
rect 10322 12336 10378 12345
rect 9496 12096 9548 12102
rect 9496 12038 9548 12044
rect 9588 12096 9640 12102
rect 9588 12038 9640 12044
rect 9508 11914 9536 12038
rect 9784 11914 9812 12294
rect 10060 12152 10088 12310
rect 10416 12310 10468 12316
rect 10322 12271 10378 12280
rect 10520 12220 10548 15098
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 10612 14113 10640 14894
rect 10598 14104 10654 14113
rect 10598 14039 10654 14048
rect 10784 13864 10836 13870
rect 10784 13806 10836 13812
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10600 13184 10652 13190
rect 10704 13161 10732 13194
rect 10600 13126 10652 13132
rect 10690 13152 10746 13161
rect 10612 12782 10640 13126
rect 10690 13087 10746 13096
rect 10704 12986 10732 13087
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10692 12844 10744 12850
rect 10692 12786 10744 12792
rect 10600 12776 10652 12782
rect 10600 12718 10652 12724
rect 10600 12368 10652 12374
rect 10600 12310 10652 12316
rect 10244 12192 10548 12220
rect 10140 12164 10192 12170
rect 10060 12124 10140 12152
rect 10244 12152 10272 12192
rect 10192 12124 10272 12152
rect 10140 12106 10192 12112
rect 10324 12096 10376 12102
rect 10322 12064 10324 12073
rect 10416 12096 10468 12102
rect 10376 12064 10378 12073
rect 9846 11996 10154 12016
rect 10416 12038 10468 12044
rect 10322 11999 10378 12008
rect 9846 11994 9852 11996
rect 9908 11994 9932 11996
rect 9988 11994 10012 11996
rect 10068 11994 10092 11996
rect 10148 11994 10154 11996
rect 9908 11942 9910 11994
rect 10090 11942 10092 11994
rect 9846 11940 9852 11942
rect 9908 11940 9932 11942
rect 9988 11940 10012 11942
rect 10068 11940 10092 11942
rect 10148 11940 10154 11942
rect 9846 11920 10154 11940
rect 10428 11914 10456 12038
rect 9508 11886 9812 11914
rect 10244 11886 10456 11914
rect 9404 11552 9456 11558
rect 9404 11494 9456 11500
rect 9312 11348 9364 11354
rect 9312 11290 9364 11296
rect 9310 11112 9366 11121
rect 9310 11047 9366 11056
rect 9324 10062 9352 11047
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9324 9110 9352 9998
rect 9312 9104 9364 9110
rect 9312 9046 9364 9052
rect 9416 8974 9444 11494
rect 9692 11082 9720 11886
rect 10244 11762 10272 11886
rect 10416 11824 10468 11830
rect 10322 11792 10378 11801
rect 10232 11756 10284 11762
rect 10416 11766 10468 11772
rect 10322 11727 10378 11736
rect 10232 11698 10284 11704
rect 10232 11552 10284 11558
rect 10232 11494 10284 11500
rect 10244 11082 10272 11494
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 10232 11076 10284 11082
rect 10232 11018 10284 11024
rect 9846 10908 10154 10928
rect 9846 10906 9852 10908
rect 9908 10906 9932 10908
rect 9988 10906 10012 10908
rect 10068 10906 10092 10908
rect 10148 10906 10154 10908
rect 9908 10854 9910 10906
rect 10090 10854 10092 10906
rect 9846 10852 9852 10854
rect 9908 10852 9932 10854
rect 9988 10852 10012 10854
rect 10068 10852 10092 10854
rect 10148 10852 10154 10854
rect 9846 10832 10154 10852
rect 9496 10804 9548 10810
rect 9496 10746 9548 10752
rect 9508 10690 9536 10746
rect 9862 10704 9918 10713
rect 9508 10662 9812 10690
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9508 10266 9536 10542
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 9588 10260 9640 10266
rect 9588 10202 9640 10208
rect 9600 10130 9628 10202
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9508 9450 9536 9930
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9324 8566 9352 8910
rect 9312 8560 9364 8566
rect 9312 8502 9364 8508
rect 9508 8498 9536 9114
rect 9600 8537 9628 9862
rect 9784 9722 9812 10662
rect 9862 10639 9918 10648
rect 10140 10668 10192 10674
rect 9876 10062 9904 10639
rect 10140 10610 10192 10616
rect 10048 10464 10100 10470
rect 10152 10452 10180 10610
rect 10244 10606 10272 11018
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10152 10424 10272 10452
rect 10048 10406 10100 10412
rect 9864 10056 9916 10062
rect 9862 10024 9864 10033
rect 9916 10024 9918 10033
rect 9862 9959 9918 9968
rect 10060 9908 10088 10406
rect 10244 10198 10272 10424
rect 10232 10192 10284 10198
rect 10232 10134 10284 10140
rect 10244 10033 10272 10134
rect 10230 10024 10286 10033
rect 10230 9959 10286 9968
rect 10232 9920 10284 9926
rect 10060 9880 10232 9908
rect 10232 9862 10284 9868
rect 9846 9820 10154 9840
rect 9846 9818 9852 9820
rect 9908 9818 9932 9820
rect 9988 9818 10012 9820
rect 10068 9818 10092 9820
rect 10148 9818 10154 9820
rect 9908 9766 9910 9818
rect 10090 9766 10092 9818
rect 9846 9764 9852 9766
rect 9908 9764 9932 9766
rect 9988 9764 10012 9766
rect 10068 9764 10092 9766
rect 10148 9764 10154 9766
rect 9846 9744 10154 9764
rect 10230 9752 10286 9761
rect 9680 9716 9732 9722
rect 9680 9658 9732 9664
rect 9772 9716 9824 9722
rect 10230 9687 10286 9696
rect 9772 9658 9824 9664
rect 9692 9178 9720 9658
rect 10244 9586 10272 9687
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9772 9376 9824 9382
rect 9772 9318 9824 9324
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9678 9072 9734 9081
rect 9678 9007 9734 9016
rect 9586 8528 9642 8537
rect 9496 8492 9548 8498
rect 9692 8498 9720 9007
rect 9784 8838 9812 9318
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9846 8732 10154 8752
rect 9846 8730 9852 8732
rect 9908 8730 9932 8732
rect 9988 8730 10012 8732
rect 10068 8730 10092 8732
rect 10148 8730 10154 8732
rect 9908 8678 9910 8730
rect 10090 8678 10092 8730
rect 9846 8676 9852 8678
rect 9908 8676 9932 8678
rect 9988 8676 10012 8678
rect 10068 8676 10092 8678
rect 10148 8676 10154 8678
rect 9846 8656 10154 8676
rect 10244 8634 10272 9318
rect 10336 9081 10364 11727
rect 10428 11218 10456 11766
rect 10612 11665 10640 12310
rect 10704 12170 10732 12786
rect 10692 12164 10744 12170
rect 10692 12106 10744 12112
rect 10704 12073 10732 12106
rect 10690 12064 10746 12073
rect 10690 11999 10746 12008
rect 10598 11656 10654 11665
rect 10598 11591 10654 11600
rect 10692 11280 10744 11286
rect 10692 11222 10744 11228
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 10428 10441 10456 11154
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10508 10532 10560 10538
rect 10508 10474 10560 10480
rect 10414 10432 10470 10441
rect 10414 10367 10470 10376
rect 10520 10266 10548 10474
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10506 9752 10562 9761
rect 10416 9716 10468 9722
rect 10506 9687 10562 9696
rect 10416 9658 10468 9664
rect 10322 9072 10378 9081
rect 10322 9007 10378 9016
rect 10324 8968 10376 8974
rect 10324 8910 10376 8916
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 9586 8463 9642 8472
rect 9680 8492 9732 8498
rect 9496 8434 9548 8440
rect 9680 8434 9732 8440
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9404 8356 9456 8362
rect 9404 8298 9456 8304
rect 9218 7984 9274 7993
rect 9218 7919 9274 7928
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9232 6769 9260 7822
rect 9310 7304 9366 7313
rect 9310 7239 9366 7248
rect 9218 6760 9274 6769
rect 9218 6695 9274 6704
rect 9140 6582 9260 6610
rect 9128 6180 9180 6186
rect 9128 6122 9180 6128
rect 9034 5808 9090 5817
rect 9034 5743 9090 5752
rect 9036 5636 9088 5642
rect 9036 5578 9088 5584
rect 9048 5370 9076 5578
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9140 5166 9168 6122
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9036 5092 9088 5098
rect 9036 5034 9088 5040
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8864 882 8892 4422
rect 8944 4208 8996 4214
rect 8944 4150 8996 4156
rect 8956 2106 8984 4150
rect 9048 2446 9076 5034
rect 9128 4684 9180 4690
rect 9232 4672 9260 6582
rect 9324 5370 9352 7239
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9312 5228 9364 5234
rect 9312 5170 9364 5176
rect 9324 4690 9352 5170
rect 9180 4644 9260 4672
rect 9312 4684 9364 4690
rect 9128 4626 9180 4632
rect 9312 4626 9364 4632
rect 9312 4548 9364 4554
rect 9232 4508 9312 4536
rect 9232 4282 9260 4508
rect 9312 4490 9364 4496
rect 9310 4448 9366 4457
rect 9310 4383 9366 4392
rect 9220 4276 9272 4282
rect 9220 4218 9272 4224
rect 9324 4214 9352 4383
rect 9312 4208 9364 4214
rect 9312 4150 9364 4156
rect 9220 3936 9272 3942
rect 9220 3878 9272 3884
rect 9232 3466 9260 3878
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 9140 2650 9168 2790
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9232 2514 9260 3402
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9220 2508 9272 2514
rect 9220 2450 9272 2456
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8944 2100 8996 2106
rect 8944 2042 8996 2048
rect 9324 1442 9352 3334
rect 9416 3194 9444 8298
rect 9772 8288 9824 8294
rect 9692 8248 9772 8276
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 7546 9628 7754
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9692 7342 9720 8248
rect 9772 8230 9824 8236
rect 10152 7834 10180 8434
rect 10232 7948 10284 7954
rect 10336 7936 10364 8910
rect 10284 7908 10364 7936
rect 10232 7890 10284 7896
rect 10428 7886 10456 9658
rect 10416 7880 10468 7886
rect 10322 7848 10378 7857
rect 10152 7806 10272 7834
rect 9846 7644 10154 7664
rect 9846 7642 9852 7644
rect 9908 7642 9932 7644
rect 9988 7642 10012 7644
rect 10068 7642 10092 7644
rect 10148 7642 10154 7644
rect 9908 7590 9910 7642
rect 10090 7590 10092 7642
rect 9846 7588 9852 7590
rect 9908 7588 9932 7590
rect 9988 7588 10012 7590
rect 10068 7588 10092 7590
rect 10148 7588 10154 7590
rect 9846 7568 10154 7588
rect 9770 7440 9826 7449
rect 9770 7375 9826 7384
rect 9954 7440 10010 7449
rect 9954 7375 10010 7384
rect 9784 7342 9812 7375
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9772 7336 9824 7342
rect 9772 7278 9824 7284
rect 9692 6730 9720 7278
rect 9680 6724 9732 6730
rect 9680 6666 9732 6672
rect 9494 6488 9550 6497
rect 9494 6423 9550 6432
rect 9508 4282 9536 6423
rect 9692 6254 9720 6666
rect 9784 6458 9812 7278
rect 9968 7177 9996 7375
rect 9954 7168 10010 7177
rect 9954 7103 10010 7112
rect 9846 6556 10154 6576
rect 9846 6554 9852 6556
rect 9908 6554 9932 6556
rect 9988 6554 10012 6556
rect 10068 6554 10092 6556
rect 10148 6554 10154 6556
rect 9908 6502 9910 6554
rect 10090 6502 10092 6554
rect 9846 6500 9852 6502
rect 9908 6500 9932 6502
rect 9988 6500 10012 6502
rect 10068 6500 10092 6502
rect 10148 6500 10154 6502
rect 9846 6480 10154 6500
rect 9772 6452 9824 6458
rect 9772 6394 9824 6400
rect 10244 6254 10272 7806
rect 10416 7822 10468 7828
rect 10322 7783 10378 7792
rect 10336 6474 10364 7783
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 7002 10456 7346
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10336 6458 10456 6474
rect 10336 6452 10468 6458
rect 10336 6446 10416 6452
rect 10416 6394 10468 6400
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 10232 6248 10284 6254
rect 10428 6225 10456 6394
rect 10232 6190 10284 6196
rect 10414 6216 10470 6225
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9494 4176 9550 4185
rect 9494 4111 9550 4120
rect 9404 3188 9456 3194
rect 9404 3130 9456 3136
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 9416 2514 9444 2790
rect 9404 2508 9456 2514
rect 9404 2450 9456 2456
rect 9404 2372 9456 2378
rect 9404 2314 9456 2320
rect 9416 1834 9444 2314
rect 9404 1828 9456 1834
rect 9404 1770 9456 1776
rect 9508 1601 9536 4111
rect 9600 3126 9628 5578
rect 9692 5166 9720 6190
rect 9772 5568 9824 5574
rect 9772 5510 9824 5516
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9784 4826 9812 5510
rect 9846 5468 10154 5488
rect 9846 5466 9852 5468
rect 9908 5466 9932 5468
rect 9988 5466 10012 5468
rect 10068 5466 10092 5468
rect 10148 5466 10154 5468
rect 9908 5414 9910 5466
rect 10090 5414 10092 5466
rect 9846 5412 9852 5414
rect 9908 5412 9932 5414
rect 9988 5412 10012 5414
rect 10068 5412 10092 5414
rect 10148 5412 10154 5414
rect 9846 5392 10154 5412
rect 10140 5296 10192 5302
rect 10140 5238 10192 5244
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 9772 4820 9824 4826
rect 9772 4762 9824 4768
rect 9876 4690 9904 5170
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 10060 4604 10088 5102
rect 10152 4758 10180 5238
rect 10244 5137 10272 6190
rect 10414 6151 10470 6160
rect 10520 5710 10548 9687
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10508 5568 10560 5574
rect 10508 5510 10560 5516
rect 10520 5234 10548 5510
rect 10508 5228 10560 5234
rect 10508 5170 10560 5176
rect 10230 5128 10286 5137
rect 10230 5063 10286 5072
rect 10612 4758 10640 10950
rect 10704 10742 10732 11222
rect 10796 11121 10824 13806
rect 10888 13530 10916 15127
rect 11612 15088 11664 15094
rect 11612 15030 11664 15036
rect 11428 14884 11480 14890
rect 11428 14826 11480 14832
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 10876 13524 10928 13530
rect 10876 13466 10928 13472
rect 11060 13320 11112 13326
rect 11058 13288 11060 13297
rect 11112 13288 11114 13297
rect 10968 13252 11020 13258
rect 11164 13258 11192 13738
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11058 13223 11114 13232
rect 11152 13252 11204 13258
rect 10968 13194 11020 13200
rect 11152 13194 11204 13200
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 10876 12708 10928 12714
rect 10876 12650 10928 12656
rect 10782 11112 10838 11121
rect 10782 11047 10838 11056
rect 10784 11008 10836 11014
rect 10784 10950 10836 10956
rect 10796 10810 10824 10950
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 10692 10736 10744 10742
rect 10692 10678 10744 10684
rect 10692 10464 10744 10470
rect 10692 10406 10744 10412
rect 10704 10169 10732 10406
rect 10690 10160 10746 10169
rect 10690 10095 10746 10104
rect 10888 9704 10916 12650
rect 10980 12238 11008 13194
rect 11060 12300 11112 12306
rect 11060 12242 11112 12248
rect 10968 12232 11020 12238
rect 10968 12174 11020 12180
rect 10966 11928 11022 11937
rect 10966 11863 11022 11872
rect 10980 11257 11008 11863
rect 11072 11762 11100 12242
rect 11164 12102 11192 13194
rect 11256 12481 11284 13194
rect 11348 13025 11376 13670
rect 11440 13530 11468 14826
rect 11624 14550 11652 15030
rect 11886 14920 11942 14929
rect 11886 14855 11942 14864
rect 11794 14648 11850 14657
rect 11900 14618 11928 14855
rect 11992 14618 12020 15302
rect 12440 15292 12492 15298
rect 12440 15234 12492 15240
rect 12070 14716 12378 14736
rect 12070 14714 12076 14716
rect 12132 14714 12156 14716
rect 12212 14714 12236 14716
rect 12292 14714 12316 14716
rect 12372 14714 12378 14716
rect 12132 14662 12134 14714
rect 12314 14662 12316 14714
rect 12070 14660 12076 14662
rect 12132 14660 12156 14662
rect 12212 14660 12236 14662
rect 12292 14660 12316 14662
rect 12372 14660 12378 14662
rect 12070 14640 12378 14660
rect 12452 14618 12480 15234
rect 12624 15224 12676 15230
rect 12624 15166 12676 15172
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 11794 14583 11850 14592
rect 11888 14612 11940 14618
rect 11808 14550 11836 14583
rect 11888 14554 11940 14560
rect 11980 14612 12032 14618
rect 11980 14554 12032 14560
rect 12440 14612 12492 14618
rect 12440 14554 12492 14560
rect 11612 14544 11664 14550
rect 11612 14486 11664 14492
rect 11796 14544 11848 14550
rect 11796 14486 11848 14492
rect 11624 13734 11652 14486
rect 11716 14334 12112 14362
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11428 13524 11480 13530
rect 11428 13466 11480 13472
rect 11612 13524 11664 13530
rect 11612 13466 11664 13472
rect 11334 13016 11390 13025
rect 11440 12986 11468 13466
rect 11520 13388 11572 13394
rect 11520 13330 11572 13336
rect 11532 13297 11560 13330
rect 11518 13288 11574 13297
rect 11518 13223 11574 13232
rect 11334 12951 11390 12960
rect 11428 12980 11480 12986
rect 11428 12922 11480 12928
rect 11624 12889 11652 13466
rect 11610 12880 11666 12889
rect 11348 12838 11560 12866
rect 11348 12617 11376 12838
rect 11532 12782 11560 12838
rect 11610 12815 11666 12824
rect 11520 12776 11572 12782
rect 11426 12744 11482 12753
rect 11520 12718 11572 12724
rect 11426 12679 11482 12688
rect 11612 12708 11664 12714
rect 11334 12608 11390 12617
rect 11334 12543 11390 12552
rect 11242 12472 11298 12481
rect 11242 12407 11244 12416
rect 11296 12407 11298 12416
rect 11336 12436 11388 12442
rect 11244 12378 11296 12384
rect 11336 12378 11388 12384
rect 11244 12300 11296 12306
rect 11244 12242 11296 12248
rect 11256 12170 11284 12242
rect 11244 12164 11296 12170
rect 11244 12106 11296 12112
rect 11152 12096 11204 12102
rect 11152 12038 11204 12044
rect 11348 11914 11376 12378
rect 11164 11886 11376 11914
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10966 11248 11022 11257
rect 10966 11183 10968 11192
rect 11020 11183 11022 11192
rect 10968 11154 11020 11160
rect 11072 11082 11100 11698
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 11058 10976 11114 10985
rect 11058 10911 11114 10920
rect 10968 10600 11020 10606
rect 10968 10542 11020 10548
rect 10704 9676 10916 9704
rect 10704 9217 10732 9676
rect 10980 9636 11008 10542
rect 10782 9616 10838 9625
rect 10782 9551 10784 9560
rect 10836 9551 10838 9560
rect 10888 9608 11008 9636
rect 10784 9522 10836 9528
rect 10690 9208 10746 9217
rect 10690 9143 10746 9152
rect 10692 9104 10744 9110
rect 10692 9046 10744 9052
rect 10704 8498 10732 9046
rect 10888 8974 10916 9608
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10980 9042 11008 9454
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10968 8832 11020 8838
rect 10966 8800 10968 8809
rect 11020 8800 11022 8809
rect 10966 8735 11022 8744
rect 10784 8628 10836 8634
rect 10784 8570 10836 8576
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10704 6866 10732 8434
rect 10796 8022 10824 8570
rect 10784 8016 10836 8022
rect 10784 7958 10836 7964
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 10796 6730 10824 7958
rect 11072 7818 11100 10911
rect 11164 10606 11192 11886
rect 11336 11688 11388 11694
rect 11336 11630 11388 11636
rect 11242 11520 11298 11529
rect 11242 11455 11298 11464
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11150 10432 11206 10441
rect 11150 10367 11206 10376
rect 11060 7812 11112 7818
rect 11060 7754 11112 7760
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10690 6080 10746 6089
rect 10690 6015 10746 6024
rect 10140 4752 10192 4758
rect 10140 4694 10192 4700
rect 10324 4752 10376 4758
rect 10324 4694 10376 4700
rect 10600 4752 10652 4758
rect 10600 4694 10652 4700
rect 10232 4616 10284 4622
rect 10060 4576 10232 4604
rect 10232 4558 10284 4564
rect 9772 4548 9824 4554
rect 9864 4548 9916 4554
rect 9824 4508 9864 4536
rect 9772 4490 9824 4496
rect 9916 4508 9996 4536
rect 9864 4490 9916 4496
rect 9968 4468 9996 4508
rect 9968 4457 10272 4468
rect 9968 4448 10286 4457
rect 9968 4440 10230 4448
rect 9846 4380 10154 4400
rect 10230 4383 10286 4392
rect 9846 4378 9852 4380
rect 9908 4378 9932 4380
rect 9988 4378 10012 4380
rect 10068 4378 10092 4380
rect 10148 4378 10154 4380
rect 9908 4326 9910 4378
rect 10090 4326 10092 4378
rect 9846 4324 9852 4326
rect 9908 4324 9932 4326
rect 9988 4324 10012 4326
rect 10068 4324 10092 4326
rect 10148 4324 10154 4326
rect 9846 4304 10154 4324
rect 10230 4312 10286 4321
rect 9772 4276 9824 4282
rect 10230 4247 10232 4256
rect 9772 4218 9824 4224
rect 10284 4247 10286 4256
rect 10232 4218 10284 4224
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9588 3120 9640 3126
rect 9588 3062 9640 3068
rect 9692 2582 9720 3402
rect 9680 2576 9732 2582
rect 9680 2518 9732 2524
rect 9784 2446 9812 4218
rect 9956 4208 10008 4214
rect 10008 4168 10180 4196
rect 9956 4150 10008 4156
rect 10152 4162 10180 4168
rect 10152 4146 10272 4162
rect 10152 4140 10284 4146
rect 10152 4134 10232 4140
rect 10232 4082 10284 4088
rect 9956 4072 10008 4078
rect 9956 4014 10008 4020
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 9968 3942 9996 4014
rect 9956 3936 10008 3942
rect 9956 3878 10008 3884
rect 10152 3466 10180 4014
rect 10140 3460 10192 3466
rect 10140 3402 10192 3408
rect 10232 3460 10284 3466
rect 10232 3402 10284 3408
rect 9846 3292 10154 3312
rect 9846 3290 9852 3292
rect 9908 3290 9932 3292
rect 9988 3290 10012 3292
rect 10068 3290 10092 3292
rect 10148 3290 10154 3292
rect 9908 3238 9910 3290
rect 10090 3238 10092 3290
rect 9846 3236 9852 3238
rect 9908 3236 9932 3238
rect 9988 3236 10012 3238
rect 10068 3236 10092 3238
rect 10148 3236 10154 3238
rect 9846 3216 10154 3236
rect 10244 2774 10272 3402
rect 10336 3194 10364 4694
rect 10704 4690 10732 6015
rect 10888 5273 10916 7686
rect 11164 7528 11192 10367
rect 11256 9178 11284 11455
rect 11348 11218 11376 11630
rect 11336 11212 11388 11218
rect 11336 11154 11388 11160
rect 11348 10266 11376 11154
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 11336 10056 11388 10062
rect 11334 10024 11336 10033
rect 11388 10024 11390 10033
rect 11334 9959 11390 9968
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11242 9072 11298 9081
rect 11242 9007 11298 9016
rect 11256 8090 11284 9007
rect 11348 8430 11376 9959
rect 11336 8424 11388 8430
rect 11336 8366 11388 8372
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11256 7750 11284 8026
rect 11348 7954 11376 8366
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11336 7812 11388 7818
rect 11336 7754 11388 7760
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11348 7546 11376 7754
rect 11072 7500 11192 7528
rect 11336 7540 11388 7546
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6254 11008 6802
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 11072 6186 11100 7500
rect 11336 7482 11388 7488
rect 11440 7426 11468 12679
rect 11612 12650 11664 12656
rect 11520 12640 11572 12646
rect 11520 12582 11572 12588
rect 11532 11898 11560 12582
rect 11520 11892 11572 11898
rect 11520 11834 11572 11840
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11532 11150 11560 11630
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11532 10441 11560 10610
rect 11518 10432 11574 10441
rect 11518 10367 11574 10376
rect 11518 10296 11574 10305
rect 11518 10231 11574 10240
rect 11164 7398 11468 7426
rect 11060 6180 11112 6186
rect 11060 6122 11112 6128
rect 10874 5264 10930 5273
rect 10874 5199 10930 5208
rect 10968 5228 11020 5234
rect 10968 5170 11020 5176
rect 10416 4684 10468 4690
rect 10416 4626 10468 4632
rect 10692 4684 10744 4690
rect 10692 4626 10744 4632
rect 10428 3534 10456 4626
rect 10598 3904 10654 3913
rect 10598 3839 10654 3848
rect 10416 3528 10468 3534
rect 10416 3470 10468 3476
rect 10612 3346 10640 3839
rect 10704 3369 10732 4626
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10876 4480 10928 4486
rect 10876 4422 10928 4428
rect 10796 3738 10824 4422
rect 10888 4321 10916 4422
rect 10874 4312 10930 4321
rect 10874 4247 10930 4256
rect 10876 3936 10928 3942
rect 10876 3878 10928 3884
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10784 3392 10836 3398
rect 10520 3318 10640 3346
rect 10690 3360 10746 3369
rect 10324 3188 10376 3194
rect 10324 3130 10376 3136
rect 10520 3058 10548 3318
rect 10784 3334 10836 3340
rect 10690 3295 10746 3304
rect 10598 3224 10654 3233
rect 10598 3159 10654 3168
rect 10612 3126 10640 3159
rect 10600 3120 10652 3126
rect 10600 3062 10652 3068
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10508 3052 10560 3058
rect 10508 2994 10560 3000
rect 10506 2952 10562 2961
rect 10506 2887 10508 2896
rect 10560 2887 10562 2896
rect 10508 2858 10560 2864
rect 10244 2746 10364 2774
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 9846 2204 10154 2224
rect 9846 2202 9852 2204
rect 9908 2202 9932 2204
rect 9988 2202 10012 2204
rect 10068 2202 10092 2204
rect 10148 2202 10154 2204
rect 9908 2150 9910 2202
rect 10090 2150 10092 2202
rect 9846 2148 9852 2150
rect 9908 2148 9932 2150
rect 9988 2148 10012 2150
rect 10068 2148 10092 2150
rect 10148 2148 10154 2150
rect 9846 2128 10154 2148
rect 9494 1592 9550 1601
rect 9494 1527 9550 1536
rect 9324 1414 9444 1442
rect 8852 876 8904 882
rect 8852 818 8904 824
rect 9416 800 9444 1414
rect 10336 800 10364 2746
rect 10704 2650 10732 3062
rect 10796 3058 10824 3334
rect 10888 3194 10916 3878
rect 10980 3738 11008 5170
rect 11164 4162 11192 7398
rect 11244 7336 11296 7342
rect 11244 7278 11296 7284
rect 11256 6798 11284 7278
rect 11532 6798 11560 10231
rect 11624 10033 11652 12650
rect 11716 12374 11744 14334
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11794 14104 11850 14113
rect 11794 14039 11850 14048
rect 11808 12442 11836 14039
rect 11888 13728 11940 13734
rect 11886 13696 11888 13705
rect 11940 13696 11942 13705
rect 11886 13631 11942 13640
rect 11796 12436 11848 12442
rect 11900 12434 11928 13631
rect 11992 12850 12020 14214
rect 12084 13870 12112 14334
rect 12162 14104 12218 14113
rect 12162 14039 12218 14048
rect 12346 14104 12402 14113
rect 12346 14039 12402 14048
rect 12176 13938 12204 14039
rect 12360 14006 12388 14039
rect 12544 14006 12572 14826
rect 12636 14618 12664 15166
rect 12714 15056 12770 15065
rect 12898 15056 12954 15065
rect 12714 14991 12770 15000
rect 12808 15020 12860 15026
rect 12728 14657 12756 14991
rect 12898 14991 12954 15000
rect 12808 14962 12860 14968
rect 12714 14648 12770 14657
rect 12624 14612 12676 14618
rect 12820 14618 12848 14962
rect 12912 14958 12940 14991
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 12992 14816 13044 14822
rect 12898 14784 12954 14793
rect 12992 14758 13044 14764
rect 12898 14719 12954 14728
rect 12714 14583 12770 14592
rect 12808 14612 12860 14618
rect 12624 14554 12676 14560
rect 12728 14006 12756 14583
rect 12808 14554 12860 14560
rect 12912 14260 12940 14719
rect 13004 14618 13032 14758
rect 13188 14618 13216 14894
rect 12992 14612 13044 14618
rect 12992 14554 13044 14560
rect 13176 14612 13228 14618
rect 13176 14554 13228 14560
rect 13176 14476 13228 14482
rect 13176 14418 13228 14424
rect 12820 14232 12940 14260
rect 12820 14113 12848 14232
rect 12806 14104 12862 14113
rect 12806 14039 12862 14048
rect 12348 14000 12400 14006
rect 12348 13942 12400 13948
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12716 14000 12768 14006
rect 12716 13942 12768 13948
rect 13082 13968 13138 13977
rect 12164 13932 12216 13938
rect 13188 13938 13216 14418
rect 13082 13903 13084 13912
rect 12164 13874 12216 13880
rect 13136 13903 13138 13912
rect 13176 13932 13228 13938
rect 13084 13874 13136 13880
rect 13176 13874 13228 13880
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12806 13832 12862 13841
rect 12806 13767 12862 13776
rect 13082 13832 13138 13841
rect 13082 13767 13138 13776
rect 12714 13696 12770 13705
rect 12070 13628 12378 13648
rect 12714 13631 12770 13640
rect 12070 13626 12076 13628
rect 12132 13626 12156 13628
rect 12212 13626 12236 13628
rect 12292 13626 12316 13628
rect 12372 13626 12378 13628
rect 12132 13574 12134 13626
rect 12314 13574 12316 13626
rect 12070 13572 12076 13574
rect 12132 13572 12156 13574
rect 12212 13572 12236 13574
rect 12292 13572 12316 13574
rect 12372 13572 12378 13574
rect 12070 13552 12378 13572
rect 12622 13560 12678 13569
rect 12176 13484 12480 13512
rect 12622 13495 12678 13504
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12084 13326 12112 13398
rect 12072 13320 12124 13326
rect 12072 13262 12124 13268
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 13025 12112 13126
rect 12070 13016 12126 13025
rect 12070 12951 12126 12960
rect 12176 12918 12204 13484
rect 12254 13424 12310 13433
rect 12452 13410 12480 13484
rect 12452 13394 12572 13410
rect 12254 13359 12310 13368
rect 12348 13388 12400 13394
rect 12164 12912 12216 12918
rect 12164 12854 12216 12860
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 12164 12776 12216 12782
rect 12268 12764 12296 13359
rect 12452 13388 12584 13394
rect 12452 13382 12532 13388
rect 12348 13330 12400 13336
rect 12532 13330 12584 13336
rect 12360 12850 12388 13330
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12216 12736 12296 12764
rect 12164 12718 12216 12724
rect 12070 12540 12378 12560
rect 12070 12538 12076 12540
rect 12132 12538 12156 12540
rect 12212 12538 12236 12540
rect 12292 12538 12316 12540
rect 12372 12538 12378 12540
rect 12132 12486 12134 12538
rect 12314 12486 12316 12538
rect 12070 12484 12076 12486
rect 12132 12484 12156 12486
rect 12212 12484 12236 12486
rect 12292 12484 12316 12486
rect 12372 12484 12378 12486
rect 12070 12464 12378 12484
rect 11900 12406 12204 12434
rect 11796 12378 11848 12384
rect 11704 12368 11756 12374
rect 11702 12336 11704 12345
rect 11888 12368 11940 12374
rect 11756 12336 11758 12345
rect 11702 12271 11758 12280
rect 11886 12336 11888 12345
rect 11940 12336 11942 12345
rect 11886 12271 11942 12280
rect 11716 12245 11744 12271
rect 11796 12232 11848 12238
rect 11796 12174 11848 12180
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11716 10606 11744 12038
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11704 10464 11756 10470
rect 11704 10406 11756 10412
rect 11716 10062 11744 10406
rect 11704 10056 11756 10062
rect 11610 10024 11666 10033
rect 11704 9998 11756 10004
rect 11610 9959 11666 9968
rect 11610 9752 11666 9761
rect 11610 9687 11612 9696
rect 11664 9687 11666 9696
rect 11612 9658 11664 9664
rect 11702 9480 11758 9489
rect 11702 9415 11704 9424
rect 11756 9415 11758 9424
rect 11704 9386 11756 9392
rect 11612 9376 11664 9382
rect 11612 9318 11664 9324
rect 11244 6792 11296 6798
rect 11244 6734 11296 6740
rect 11520 6792 11572 6798
rect 11520 6734 11572 6740
rect 11256 5574 11284 6734
rect 11428 6656 11480 6662
rect 11334 6624 11390 6633
rect 11428 6598 11480 6604
rect 11334 6559 11390 6568
rect 11348 6458 11376 6559
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11336 5636 11388 5642
rect 11336 5578 11388 5584
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11256 5166 11284 5510
rect 11348 5302 11376 5578
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11244 5160 11296 5166
rect 11244 5102 11296 5108
rect 11072 4134 11192 4162
rect 10968 3732 11020 3738
rect 10968 3674 11020 3680
rect 10876 3188 10928 3194
rect 10876 3130 10928 3136
rect 10784 3052 10836 3058
rect 10784 2994 10836 3000
rect 10796 2774 10824 2994
rect 10968 2984 11020 2990
rect 10968 2926 11020 2932
rect 10796 2746 10916 2774
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10428 2446 10456 2586
rect 10508 2576 10560 2582
rect 10508 2518 10560 2524
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 10520 2310 10548 2518
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10888 2106 10916 2746
rect 10980 2582 11008 2926
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10876 2100 10928 2106
rect 10876 2042 10928 2048
rect 10980 1358 11008 2246
rect 10968 1352 11020 1358
rect 10968 1294 11020 1300
rect 11072 1222 11100 4134
rect 11152 4072 11204 4078
rect 11152 4014 11204 4020
rect 11164 3913 11192 4014
rect 11150 3904 11206 3913
rect 11150 3839 11206 3848
rect 11256 3534 11284 5102
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4690 11376 4966
rect 11336 4684 11388 4690
rect 11336 4626 11388 4632
rect 11348 4146 11376 4626
rect 11336 4140 11388 4146
rect 11336 4082 11388 4088
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 11164 2038 11192 2246
rect 11152 2032 11204 2038
rect 11152 1974 11204 1980
rect 11244 1488 11296 1494
rect 11244 1430 11296 1436
rect 11060 1216 11112 1222
rect 11060 1158 11112 1164
rect 11256 800 11284 1430
rect 11440 1290 11468 6598
rect 11624 5760 11652 9318
rect 11704 9172 11756 9178
rect 11704 9114 11756 9120
rect 11716 8294 11744 9114
rect 11808 8498 11836 12174
rect 12176 12102 12204 12406
rect 12452 12374 12480 13262
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12544 12714 12572 13194
rect 12636 13161 12664 13495
rect 12622 13152 12678 13161
rect 12622 13087 12678 13096
rect 12728 12986 12756 13631
rect 12820 13530 12848 13767
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 12716 12980 12768 12986
rect 12716 12922 12768 12928
rect 12714 12880 12770 12889
rect 12820 12850 12848 13466
rect 13096 13462 13124 13767
rect 13176 13728 13228 13734
rect 13176 13670 13228 13676
rect 13084 13456 13136 13462
rect 13084 13398 13136 13404
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 13025 12940 13262
rect 12898 13016 12954 13025
rect 12898 12951 12954 12960
rect 12714 12815 12770 12824
rect 12808 12844 12860 12850
rect 12532 12708 12584 12714
rect 12532 12650 12584 12656
rect 12728 12481 12756 12815
rect 13004 12832 13032 13330
rect 13188 12986 13216 13670
rect 13176 12980 13228 12986
rect 13176 12922 13228 12928
rect 13084 12844 13136 12850
rect 13004 12804 13084 12832
rect 12808 12786 12860 12792
rect 13084 12786 13136 12792
rect 13372 12782 13400 15438
rect 14004 14612 14056 14618
rect 14004 14554 14056 14560
rect 13910 14512 13966 14521
rect 13910 14447 13912 14456
rect 13964 14447 13966 14456
rect 13912 14418 13964 14424
rect 13820 14340 13872 14346
rect 13820 14282 13872 14288
rect 13832 14249 13860 14282
rect 13818 14240 13874 14249
rect 14016 14226 14044 14554
rect 14568 14414 14596 15642
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14556 14408 14608 14414
rect 14556 14350 14608 14356
rect 14096 14340 14148 14346
rect 14148 14300 14228 14328
rect 14096 14282 14148 14288
rect 14016 14198 14136 14226
rect 13818 14175 13874 14184
rect 14002 14104 14058 14113
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13912 14068 13964 14074
rect 14002 14039 14058 14048
rect 13912 14010 13964 14016
rect 13648 13938 13676 14010
rect 13636 13932 13688 13938
rect 13636 13874 13688 13880
rect 13636 13796 13688 13802
rect 13636 13738 13688 13744
rect 13544 13524 13596 13530
rect 13544 13466 13596 13472
rect 13556 13433 13584 13466
rect 13542 13424 13598 13433
rect 13542 13359 13598 13368
rect 13648 13326 13676 13738
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13452 13184 13504 13190
rect 13452 13126 13504 13132
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13464 12832 13492 13126
rect 13648 12889 13676 13126
rect 13634 12880 13690 12889
rect 13544 12844 13596 12850
rect 13464 12804 13544 12832
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 12992 12708 13044 12714
rect 12992 12650 13044 12656
rect 12714 12472 12770 12481
rect 12714 12407 12770 12416
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 11980 12096 12032 12102
rect 12164 12096 12216 12102
rect 11980 12038 12032 12044
rect 12162 12064 12164 12073
rect 12348 12096 12400 12102
rect 12216 12064 12218 12073
rect 11992 11937 12020 12038
rect 12348 12038 12400 12044
rect 12162 11999 12218 12008
rect 11978 11928 12034 11937
rect 11978 11863 11980 11872
rect 12032 11863 12034 11872
rect 11980 11834 12032 11840
rect 12360 11801 12388 12038
rect 12346 11792 12402 11801
rect 11980 11756 12032 11762
rect 12346 11727 12402 11736
rect 11980 11698 12032 11704
rect 11888 11552 11940 11558
rect 11888 11494 11940 11500
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11716 7478 11744 8026
rect 11808 7857 11836 8434
rect 11900 8401 11928 11494
rect 11886 8392 11942 8401
rect 11886 8327 11942 8336
rect 11888 8288 11940 8294
rect 11888 8230 11940 8236
rect 11794 7848 11850 7857
rect 11794 7783 11850 7792
rect 11704 7472 11756 7478
rect 11704 7414 11756 7420
rect 11796 7404 11848 7410
rect 11796 7346 11848 7352
rect 11704 6656 11756 6662
rect 11808 6644 11836 7346
rect 11756 6616 11836 6644
rect 11704 6598 11756 6604
rect 11716 6254 11744 6598
rect 11794 6488 11850 6497
rect 11794 6423 11796 6432
rect 11848 6423 11850 6432
rect 11796 6394 11848 6400
rect 11796 6316 11848 6322
rect 11796 6258 11848 6264
rect 11704 6248 11756 6254
rect 11704 6190 11756 6196
rect 11716 5914 11744 6190
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11624 5732 11744 5760
rect 11520 5024 11572 5030
rect 11520 4966 11572 4972
rect 11532 4758 11560 4966
rect 11520 4752 11572 4758
rect 11520 4694 11572 4700
rect 11520 4616 11572 4622
rect 11520 4558 11572 4564
rect 11610 4584 11666 4593
rect 11532 4214 11560 4558
rect 11610 4519 11666 4528
rect 11520 4208 11572 4214
rect 11520 4150 11572 4156
rect 11624 4146 11652 4519
rect 11612 4140 11664 4146
rect 11612 4082 11664 4088
rect 11520 4072 11572 4078
rect 11520 4014 11572 4020
rect 11532 3194 11560 4014
rect 11610 3768 11666 3777
rect 11610 3703 11666 3712
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11624 2922 11652 3703
rect 11716 3194 11744 5732
rect 11808 5642 11836 6258
rect 11796 5636 11848 5642
rect 11796 5578 11848 5584
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4554 11836 4966
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11900 4486 11928 8230
rect 11992 6474 12020 11698
rect 12070 11452 12378 11472
rect 12070 11450 12076 11452
rect 12132 11450 12156 11452
rect 12212 11450 12236 11452
rect 12292 11450 12316 11452
rect 12372 11450 12378 11452
rect 12132 11398 12134 11450
rect 12314 11398 12316 11450
rect 12070 11396 12076 11398
rect 12132 11396 12156 11398
rect 12212 11396 12236 11398
rect 12292 11396 12316 11398
rect 12372 11396 12378 11398
rect 12070 11376 12378 11396
rect 12254 11248 12310 11257
rect 12254 11183 12256 11192
rect 12308 11183 12310 11192
rect 12256 11154 12308 11160
rect 12452 11150 12480 12310
rect 13004 12306 13032 12650
rect 13268 12640 13320 12646
rect 13268 12582 13320 12588
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 12808 12232 12860 12238
rect 12530 12200 12586 12209
rect 12808 12174 12860 12180
rect 12900 12232 12952 12238
rect 12900 12174 12952 12180
rect 13176 12232 13228 12238
rect 13176 12174 13228 12180
rect 12530 12135 12586 12144
rect 12544 12102 12572 12135
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12820 11880 12848 12174
rect 12912 11914 12940 12174
rect 13084 12096 13136 12102
rect 13084 12038 13136 12044
rect 12912 11886 13032 11914
rect 12636 11852 12848 11880
rect 12532 11756 12584 11762
rect 12532 11698 12584 11704
rect 12440 11144 12492 11150
rect 12254 11112 12310 11121
rect 12440 11086 12492 11092
rect 12254 11047 12310 11056
rect 12164 11008 12216 11014
rect 12164 10950 12216 10956
rect 12176 10849 12204 10950
rect 12162 10840 12218 10849
rect 12162 10775 12218 10784
rect 12162 10568 12218 10577
rect 12268 10538 12296 11047
rect 12162 10503 12164 10512
rect 12216 10503 12218 10512
rect 12256 10532 12308 10538
rect 12164 10474 12216 10480
rect 12256 10474 12308 10480
rect 12070 10364 12378 10384
rect 12070 10362 12076 10364
rect 12132 10362 12156 10364
rect 12212 10362 12236 10364
rect 12292 10362 12316 10364
rect 12372 10362 12378 10364
rect 12132 10310 12134 10362
rect 12314 10310 12316 10362
rect 12070 10308 12076 10310
rect 12132 10308 12156 10310
rect 12212 10308 12236 10310
rect 12292 10308 12316 10310
rect 12372 10308 12378 10310
rect 12070 10288 12378 10308
rect 12348 9920 12400 9926
rect 12452 9897 12480 11086
rect 12348 9862 12400 9868
rect 12438 9888 12494 9897
rect 12360 9364 12388 9862
rect 12438 9823 12494 9832
rect 12440 9648 12492 9654
rect 12440 9590 12492 9596
rect 12452 9489 12480 9590
rect 12438 9480 12494 9489
rect 12438 9415 12494 9424
rect 12544 9382 12572 11698
rect 12636 11014 12664 11852
rect 12900 11824 12952 11830
rect 12806 11792 12862 11801
rect 12900 11766 12952 11772
rect 12806 11727 12862 11736
rect 12820 11626 12848 11727
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 12716 11552 12768 11558
rect 12716 11494 12768 11500
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12636 10690 12664 10950
rect 12728 10810 12756 11494
rect 12912 11393 12940 11766
rect 13004 11506 13032 11886
rect 13096 11801 13124 12038
rect 13188 11937 13216 12174
rect 13174 11928 13230 11937
rect 13174 11863 13230 11872
rect 13082 11792 13138 11801
rect 13082 11727 13138 11736
rect 13082 11656 13138 11665
rect 13082 11591 13084 11600
rect 13136 11591 13138 11600
rect 13084 11562 13136 11568
rect 13082 11520 13138 11529
rect 13004 11478 13082 11506
rect 13082 11455 13138 11464
rect 12898 11384 12954 11393
rect 12808 11348 12860 11354
rect 12898 11319 12954 11328
rect 12808 11290 12860 11296
rect 12716 10804 12768 10810
rect 12716 10746 12768 10752
rect 12636 10662 12756 10690
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12636 10305 12664 10406
rect 12622 10296 12678 10305
rect 12622 10231 12678 10240
rect 12624 9988 12676 9994
rect 12624 9930 12676 9936
rect 12636 9586 12664 9930
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 12532 9376 12584 9382
rect 12360 9336 12480 9364
rect 12070 9276 12378 9296
rect 12070 9274 12076 9276
rect 12132 9274 12156 9276
rect 12212 9274 12236 9276
rect 12292 9274 12316 9276
rect 12372 9274 12378 9276
rect 12132 9222 12134 9274
rect 12314 9222 12316 9274
rect 12070 9220 12076 9222
rect 12132 9220 12156 9222
rect 12212 9220 12236 9222
rect 12292 9220 12316 9222
rect 12372 9220 12378 9222
rect 12070 9200 12378 9220
rect 12452 9160 12480 9336
rect 12532 9318 12584 9324
rect 12360 9132 12480 9160
rect 12530 9208 12586 9217
rect 12530 9143 12586 9152
rect 12070 9072 12126 9081
rect 12070 9007 12126 9016
rect 12084 8974 12112 9007
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 8430 12112 8774
rect 12072 8424 12124 8430
rect 12072 8366 12124 8372
rect 12360 8344 12388 9132
rect 12438 8800 12494 8809
rect 12438 8735 12494 8744
rect 12452 8634 12480 8735
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12360 8316 12434 8344
rect 12070 8188 12378 8208
rect 12070 8186 12076 8188
rect 12132 8186 12156 8188
rect 12212 8186 12236 8188
rect 12292 8186 12316 8188
rect 12372 8186 12378 8188
rect 12132 8134 12134 8186
rect 12314 8134 12316 8186
rect 12070 8132 12076 8134
rect 12132 8132 12156 8134
rect 12212 8132 12236 8134
rect 12292 8132 12316 8134
rect 12372 8132 12378 8134
rect 12070 8112 12378 8132
rect 12406 7970 12434 8316
rect 12360 7942 12434 7970
rect 12360 7256 12388 7942
rect 12544 7562 12572 9143
rect 12636 9042 12664 9522
rect 12728 9058 12756 10662
rect 12820 9353 12848 11290
rect 13176 11280 13228 11286
rect 12990 11248 13046 11257
rect 13176 11222 13228 11228
rect 12990 11183 13046 11192
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12806 9344 12862 9353
rect 12806 9279 12862 9288
rect 12624 9036 12676 9042
rect 12728 9030 12848 9058
rect 12624 8978 12676 8984
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12624 8832 12676 8838
rect 12624 8774 12676 8780
rect 12636 8634 12664 8774
rect 12728 8634 12756 8910
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12716 7812 12768 7818
rect 12716 7754 12768 7760
rect 12544 7534 12664 7562
rect 12360 7228 12480 7256
rect 12070 7100 12378 7120
rect 12070 7098 12076 7100
rect 12132 7098 12156 7100
rect 12212 7098 12236 7100
rect 12292 7098 12316 7100
rect 12372 7098 12378 7100
rect 12132 7046 12134 7098
rect 12314 7046 12316 7098
rect 12070 7044 12076 7046
rect 12132 7044 12156 7046
rect 12212 7044 12236 7046
rect 12292 7044 12316 7046
rect 12372 7044 12378 7046
rect 12070 7024 12378 7044
rect 12452 6916 12480 7228
rect 12360 6888 12480 6916
rect 11992 6458 12204 6474
rect 11992 6452 12216 6458
rect 11992 6446 12164 6452
rect 12164 6394 12216 6400
rect 12072 6316 12124 6322
rect 12256 6316 12308 6322
rect 12124 6276 12256 6304
rect 12072 6258 12124 6264
rect 12256 6258 12308 6264
rect 12360 6202 12388 6888
rect 12360 6174 12480 6202
rect 12070 6012 12378 6032
rect 12070 6010 12076 6012
rect 12132 6010 12156 6012
rect 12212 6010 12236 6012
rect 12292 6010 12316 6012
rect 12372 6010 12378 6012
rect 12132 5958 12134 6010
rect 12314 5958 12316 6010
rect 12070 5956 12076 5958
rect 12132 5956 12156 5958
rect 12212 5956 12236 5958
rect 12292 5956 12316 5958
rect 12372 5956 12378 5958
rect 12070 5936 12378 5956
rect 12452 5794 12480 6174
rect 12360 5766 12480 5794
rect 12360 5137 12388 5766
rect 12636 5370 12664 7534
rect 12728 7410 12756 7754
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12728 5370 12756 7346
rect 12820 7002 12848 9030
rect 12912 7546 12940 11086
rect 13004 11082 13032 11183
rect 13084 11144 13136 11150
rect 13084 11086 13136 11092
rect 12992 11076 13044 11082
rect 12992 11018 13044 11024
rect 12992 10804 13044 10810
rect 12992 10746 13044 10752
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 12820 6186 12848 6394
rect 12912 6254 12940 7482
rect 13004 7041 13032 10746
rect 13096 8650 13124 11086
rect 13188 10554 13216 11222
rect 13280 10674 13308 12582
rect 13358 12336 13414 12345
rect 13358 12271 13414 12280
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13372 10606 13400 12271
rect 13464 11150 13492 12804
rect 13634 12815 13690 12824
rect 13544 12786 13596 12792
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 12481 13676 12582
rect 13634 12472 13690 12481
rect 13634 12407 13690 12416
rect 13740 12374 13768 14010
rect 13818 13832 13874 13841
rect 13818 13767 13874 13776
rect 13832 13462 13860 13767
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 13820 12980 13872 12986
rect 13820 12922 13872 12928
rect 13728 12368 13780 12374
rect 13832 12345 13860 12922
rect 13728 12310 13780 12316
rect 13818 12336 13874 12345
rect 13818 12271 13874 12280
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13634 12064 13690 12073
rect 13634 11999 13690 12008
rect 13648 11762 13676 11999
rect 13740 11812 13768 12174
rect 13820 12096 13872 12102
rect 13818 12064 13820 12073
rect 13872 12064 13874 12073
rect 13818 11999 13874 12008
rect 13740 11784 13860 11812
rect 13636 11756 13688 11762
rect 13688 11716 13768 11744
rect 13636 11698 13688 11704
rect 13636 11552 13688 11558
rect 13740 11529 13768 11716
rect 13832 11665 13860 11784
rect 13818 11656 13874 11665
rect 13818 11591 13874 11600
rect 13820 11552 13872 11558
rect 13636 11494 13688 11500
rect 13726 11520 13782 11529
rect 13648 11354 13676 11494
rect 13820 11494 13872 11500
rect 13726 11455 13782 11464
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13452 11144 13504 11150
rect 13832 11098 13860 11494
rect 13452 11086 13504 11092
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13648 11070 13860 11098
rect 13360 10600 13412 10606
rect 13188 10526 13308 10554
rect 13360 10542 13412 10548
rect 13176 10464 13228 10470
rect 13176 10406 13228 10412
rect 13188 8838 13216 10406
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13096 8622 13216 8650
rect 13084 8424 13136 8430
rect 13084 8366 13136 8372
rect 12990 7032 13046 7041
rect 12990 6967 13046 6976
rect 13096 6662 13124 8366
rect 13188 7410 13216 8622
rect 13280 8294 13308 10526
rect 13360 9512 13412 9518
rect 13360 9454 13412 9460
rect 13372 9178 13400 9454
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13464 9042 13492 9318
rect 13452 9036 13504 9042
rect 13452 8978 13504 8984
rect 13360 8900 13412 8906
rect 13360 8842 13412 8848
rect 13268 8288 13320 8294
rect 13268 8230 13320 8236
rect 13176 7404 13228 7410
rect 13176 7346 13228 7352
rect 13176 6996 13228 7002
rect 13176 6938 13228 6944
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13082 6488 13138 6497
rect 13082 6423 13084 6432
rect 13136 6423 13138 6432
rect 13084 6394 13136 6400
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12808 6180 12860 6186
rect 12808 6122 12860 6128
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 11978 5128 12034 5137
rect 11978 5063 12034 5072
rect 12346 5128 12402 5137
rect 12346 5063 12402 5072
rect 11992 4826 12020 5063
rect 12070 4924 12378 4944
rect 12070 4922 12076 4924
rect 12132 4922 12156 4924
rect 12212 4922 12236 4924
rect 12292 4922 12316 4924
rect 12372 4922 12378 4924
rect 12132 4870 12134 4922
rect 12314 4870 12316 4922
rect 12070 4868 12076 4870
rect 12132 4868 12156 4870
rect 12212 4868 12236 4870
rect 12292 4868 12316 4870
rect 12372 4868 12378 4870
rect 12070 4848 12378 4868
rect 11980 4820 12032 4826
rect 11980 4762 12032 4768
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 12348 4480 12400 4486
rect 12348 4422 12400 4428
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 11888 4208 11940 4214
rect 11888 4150 11940 4156
rect 11978 4176 12034 4185
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11808 3738 11836 3878
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 11704 3188 11756 3194
rect 11704 3130 11756 3136
rect 11612 2916 11664 2922
rect 11612 2858 11664 2864
rect 11900 2009 11928 4150
rect 11978 4111 12034 4120
rect 11992 2446 12020 4111
rect 12360 4026 12388 4422
rect 12544 4282 12572 4422
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12636 4146 12664 5306
rect 12900 4208 12952 4214
rect 13004 4196 13032 6326
rect 13188 6254 13216 6938
rect 13266 6896 13322 6905
rect 13372 6866 13400 8842
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13266 6831 13322 6840
rect 13360 6860 13412 6866
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13084 5296 13136 5302
rect 13084 5238 13136 5244
rect 13096 5030 13124 5238
rect 13084 5024 13136 5030
rect 13084 4966 13136 4972
rect 12952 4168 13032 4196
rect 12900 4150 12952 4156
rect 12624 4140 12676 4146
rect 12624 4082 12676 4088
rect 13084 4072 13136 4078
rect 12360 3998 12572 4026
rect 13084 4014 13136 4020
rect 12070 3836 12378 3856
rect 12070 3834 12076 3836
rect 12132 3834 12156 3836
rect 12212 3834 12236 3836
rect 12292 3834 12316 3836
rect 12372 3834 12378 3836
rect 12132 3782 12134 3834
rect 12314 3782 12316 3834
rect 12070 3780 12076 3782
rect 12132 3780 12156 3782
rect 12212 3780 12236 3782
rect 12292 3780 12316 3782
rect 12372 3780 12378 3782
rect 12070 3760 12378 3780
rect 12164 3664 12216 3670
rect 12084 3612 12164 3618
rect 12084 3606 12216 3612
rect 12084 3590 12204 3606
rect 12084 3369 12112 3590
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12070 3360 12126 3369
rect 12070 3295 12126 3304
rect 12070 3088 12126 3097
rect 12070 3023 12126 3032
rect 12084 2990 12112 3023
rect 12176 2990 12204 3470
rect 12544 3058 12572 3998
rect 12808 4004 12860 4010
rect 12808 3946 12860 3952
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12636 3534 12664 3567
rect 12624 3528 12676 3534
rect 12624 3470 12676 3476
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12072 2984 12124 2990
rect 12072 2926 12124 2932
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 12070 2748 12378 2768
rect 12070 2746 12076 2748
rect 12132 2746 12156 2748
rect 12212 2746 12236 2748
rect 12292 2746 12316 2748
rect 12372 2746 12378 2748
rect 12132 2694 12134 2746
rect 12314 2694 12316 2746
rect 12070 2692 12076 2694
rect 12132 2692 12156 2694
rect 12212 2692 12236 2694
rect 12292 2692 12316 2694
rect 12372 2692 12378 2694
rect 12070 2672 12378 2692
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 11980 2440 12032 2446
rect 11980 2382 12032 2388
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11886 2000 11942 2009
rect 11886 1935 11942 1944
rect 11992 1358 12020 2246
rect 12084 1766 12112 2450
rect 12256 2440 12308 2446
rect 12256 2382 12308 2388
rect 12072 1760 12124 1766
rect 12072 1702 12124 1708
rect 12164 1760 12216 1766
rect 12164 1702 12216 1708
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 11428 1284 11480 1290
rect 11428 1226 11480 1232
rect 12176 800 12204 1702
rect 12268 1630 12296 2382
rect 12348 2372 12400 2378
rect 12348 2314 12400 2320
rect 12360 1970 12388 2314
rect 12544 2038 12572 2994
rect 12624 2304 12676 2310
rect 12624 2246 12676 2252
rect 12716 2304 12768 2310
rect 12716 2246 12768 2252
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 12348 1964 12400 1970
rect 12348 1906 12400 1912
rect 12256 1624 12308 1630
rect 12256 1566 12308 1572
rect 12544 1465 12572 1974
rect 12636 1698 12664 2246
rect 12624 1692 12676 1698
rect 12624 1634 12676 1640
rect 12728 1630 12756 2246
rect 12716 1624 12768 1630
rect 12716 1566 12768 1572
rect 12820 1494 12848 3946
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 12912 3670 12940 3878
rect 13096 3738 13124 4014
rect 13084 3732 13136 3738
rect 13084 3674 13136 3680
rect 12900 3664 12952 3670
rect 12900 3606 12952 3612
rect 13174 3632 13230 3641
rect 13174 3567 13230 3576
rect 13188 3398 13216 3567
rect 13280 3482 13308 6831
rect 13360 6802 13412 6808
rect 13372 6662 13400 6802
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13464 6474 13492 8774
rect 13556 7886 13584 11018
rect 13544 7880 13596 7886
rect 13544 7822 13596 7828
rect 13372 6446 13492 6474
rect 13372 4593 13400 6446
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13464 5710 13492 6258
rect 13452 5704 13504 5710
rect 13452 5646 13504 5652
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13556 4690 13584 5170
rect 13544 4684 13596 4690
rect 13544 4626 13596 4632
rect 13358 4584 13414 4593
rect 13358 4519 13414 4528
rect 13360 4480 13412 4486
rect 13360 4422 13412 4428
rect 13372 3738 13400 4422
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13464 3505 13492 4082
rect 13556 4078 13584 4626
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 13450 3496 13506 3505
rect 13280 3454 13400 3482
rect 13372 3398 13400 3454
rect 13450 3431 13506 3440
rect 13176 3392 13228 3398
rect 13176 3334 13228 3340
rect 13360 3392 13412 3398
rect 13360 3334 13412 3340
rect 13544 3392 13596 3398
rect 13544 3334 13596 3340
rect 13556 3233 13584 3334
rect 13542 3224 13598 3233
rect 13542 3159 13598 3168
rect 12900 2848 12952 2854
rect 12900 2790 12952 2796
rect 13268 2848 13320 2854
rect 13268 2790 13320 2796
rect 12912 2378 12940 2790
rect 12900 2372 12952 2378
rect 12900 2314 12952 2320
rect 12808 1488 12860 1494
rect 12530 1456 12586 1465
rect 13280 1442 13308 2790
rect 12808 1430 12860 1436
rect 12530 1391 12586 1400
rect 13096 1414 13308 1442
rect 13096 800 13124 1414
rect 13648 1358 13676 11070
rect 13818 10840 13874 10849
rect 13818 10775 13874 10784
rect 13832 10554 13860 10775
rect 13740 10526 13860 10554
rect 13740 10146 13768 10526
rect 13740 10118 13860 10146
rect 13728 9920 13780 9926
rect 13728 9862 13780 9868
rect 13740 9450 13768 9862
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 8974 13768 9386
rect 13832 9110 13860 10118
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13924 9058 13952 14010
rect 14016 13920 14044 14039
rect 14108 13988 14136 14198
rect 14200 14056 14228 14300
rect 14294 14172 14602 14192
rect 14294 14170 14300 14172
rect 14356 14170 14380 14172
rect 14436 14170 14460 14172
rect 14516 14170 14540 14172
rect 14596 14170 14602 14172
rect 14356 14118 14358 14170
rect 14538 14118 14540 14170
rect 14294 14116 14300 14118
rect 14356 14116 14380 14118
rect 14436 14116 14460 14118
rect 14516 14116 14540 14118
rect 14596 14116 14602 14118
rect 14294 14096 14602 14116
rect 14200 14028 14320 14056
rect 14108 13960 14228 13988
rect 14016 13892 14136 13920
rect 14004 13184 14056 13190
rect 14004 13126 14056 13132
rect 14016 11830 14044 13126
rect 14108 12986 14136 13892
rect 14200 13326 14228 13960
rect 14292 13394 14320 14028
rect 14660 13988 14688 15574
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 14113 14780 14214
rect 14738 14104 14794 14113
rect 14844 14074 14872 15778
rect 15476 15292 15528 15298
rect 15476 15234 15528 15240
rect 15488 15094 15516 15234
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15476 15088 15528 15094
rect 15476 15030 15528 15036
rect 15028 14906 15056 15030
rect 15028 14878 15240 14906
rect 15106 14648 15162 14657
rect 15106 14583 15162 14592
rect 15120 14550 15148 14583
rect 15016 14544 15068 14550
rect 14922 14512 14978 14521
rect 15016 14486 15068 14492
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 14922 14447 14978 14456
rect 14936 14074 14964 14447
rect 15028 14414 15056 14486
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15212 14346 15240 14878
rect 15108 14340 15160 14346
rect 15108 14282 15160 14288
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14738 14039 14794 14048
rect 14832 14068 14884 14074
rect 14832 14010 14884 14016
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 14660 13960 14780 13988
rect 14648 13864 14700 13870
rect 14370 13832 14426 13841
rect 14648 13806 14700 13812
rect 14370 13767 14372 13776
rect 14424 13767 14426 13776
rect 14372 13738 14424 13744
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14568 13569 14596 13670
rect 14554 13560 14610 13569
rect 14554 13495 14610 13504
rect 14370 13424 14426 13433
rect 14280 13388 14332 13394
rect 14370 13359 14426 13368
rect 14280 13330 14332 13336
rect 14188 13320 14240 13326
rect 14188 13262 14240 13268
rect 14188 13184 14240 13190
rect 14384 13172 14412 13359
rect 14240 13144 14412 13172
rect 14188 13126 14240 13132
rect 14294 13084 14602 13104
rect 14294 13082 14300 13084
rect 14356 13082 14380 13084
rect 14436 13082 14460 13084
rect 14516 13082 14540 13084
rect 14596 13082 14602 13084
rect 14356 13030 14358 13082
rect 14538 13030 14540 13082
rect 14294 13028 14300 13030
rect 14356 13028 14380 13030
rect 14436 13028 14460 13030
rect 14516 13028 14540 13030
rect 14596 13028 14602 13030
rect 14294 13008 14602 13028
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14094 12880 14150 12889
rect 14094 12815 14096 12824
rect 14148 12815 14150 12824
rect 14556 12844 14608 12850
rect 14096 12786 14148 12792
rect 14556 12786 14608 12792
rect 14278 12744 14334 12753
rect 14188 12708 14240 12714
rect 14278 12679 14280 12688
rect 14188 12650 14240 12656
rect 14332 12679 14334 12688
rect 14462 12744 14518 12753
rect 14462 12679 14518 12688
rect 14280 12650 14332 12656
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 11824 14056 11830
rect 14004 11766 14056 11772
rect 14108 11746 14136 12582
rect 14200 12345 14228 12650
rect 14476 12442 14504 12679
rect 14568 12481 14596 12786
rect 14554 12472 14610 12481
rect 14464 12436 14516 12442
rect 14554 12407 14610 12416
rect 14464 12378 14516 12384
rect 14186 12336 14242 12345
rect 14186 12271 14242 12280
rect 14188 12232 14240 12238
rect 14188 12174 14240 12180
rect 14096 11740 14148 11746
rect 14096 11682 14148 11688
rect 14002 11656 14058 11665
rect 14002 11591 14058 11600
rect 14016 11354 14044 11591
rect 14094 11384 14150 11393
rect 14004 11348 14056 11354
rect 14094 11319 14150 11328
rect 14004 11290 14056 11296
rect 14004 11076 14056 11082
rect 14004 11018 14056 11024
rect 14016 9178 14044 11018
rect 14108 10606 14136 11319
rect 14200 10810 14228 12174
rect 14294 11996 14602 12016
rect 14294 11994 14300 11996
rect 14356 11994 14380 11996
rect 14436 11994 14460 11996
rect 14516 11994 14540 11996
rect 14596 11994 14602 11996
rect 14356 11942 14358 11994
rect 14538 11942 14540 11994
rect 14294 11940 14300 11942
rect 14356 11940 14380 11942
rect 14436 11940 14460 11942
rect 14516 11940 14540 11942
rect 14596 11940 14602 11942
rect 14294 11920 14602 11940
rect 14556 11824 14608 11830
rect 14556 11766 14608 11772
rect 14372 11552 14424 11558
rect 14372 11494 14424 11500
rect 14384 11393 14412 11494
rect 14370 11384 14426 11393
rect 14370 11319 14426 11328
rect 14568 11082 14596 11766
rect 14660 11762 14688 13806
rect 14752 12850 14780 13960
rect 15028 13818 15056 14214
rect 15120 14006 15148 14282
rect 15304 14278 15332 15030
rect 15672 14958 15700 16895
rect 16302 16552 16358 16561
rect 16302 16487 16358 16496
rect 15842 15056 15898 15065
rect 15842 14991 15898 15000
rect 16026 15056 16082 15065
rect 16316 15026 16344 16487
rect 17866 16400 17922 17200
rect 17682 16144 17738 16153
rect 17682 16079 17738 16088
rect 17590 15736 17646 15745
rect 17590 15671 17646 15680
rect 17604 15162 17632 15671
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 16026 14991 16082 15000
rect 16304 15020 16356 15026
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15672 14414 15700 14894
rect 15856 14414 15884 14991
rect 16040 14822 16068 14991
rect 16304 14962 16356 14968
rect 16028 14816 16080 14822
rect 16028 14758 16080 14764
rect 16210 14784 16266 14793
rect 16040 14414 16068 14758
rect 16210 14719 16266 14728
rect 15660 14408 15712 14414
rect 15474 14376 15530 14385
rect 15660 14350 15712 14356
rect 15844 14408 15896 14414
rect 15844 14350 15896 14356
rect 16028 14408 16080 14414
rect 16028 14350 16080 14356
rect 15474 14311 15530 14320
rect 15292 14272 15344 14278
rect 15292 14214 15344 14220
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15382 13968 15438 13977
rect 15292 13932 15344 13938
rect 15382 13903 15384 13912
rect 15292 13874 15344 13880
rect 15436 13903 15438 13912
rect 15384 13874 15436 13880
rect 15304 13841 15332 13874
rect 15290 13832 15346 13841
rect 15028 13790 15240 13818
rect 14924 13728 14976 13734
rect 15108 13728 15160 13734
rect 14976 13688 15056 13716
rect 14924 13670 14976 13676
rect 14922 13560 14978 13569
rect 14922 13495 14978 13504
rect 14936 13462 14964 13495
rect 14924 13456 14976 13462
rect 14830 13424 14886 13433
rect 14924 13398 14976 13404
rect 14830 13359 14886 13368
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14844 12424 14872 13359
rect 14924 13252 14976 13258
rect 14924 13194 14976 13200
rect 14936 13161 14964 13194
rect 14922 13152 14978 13161
rect 14922 13087 14978 13096
rect 15028 12866 15056 13688
rect 15108 13670 15160 13676
rect 15120 13297 15148 13670
rect 15212 13512 15240 13790
rect 15290 13767 15346 13776
rect 15212 13484 15332 13512
rect 15200 13388 15252 13394
rect 15200 13330 15252 13336
rect 15106 13288 15162 13297
rect 15106 13223 15162 13232
rect 14936 12838 15056 12866
rect 14936 12442 14964 12838
rect 15212 12730 15240 13330
rect 15120 12702 15240 12730
rect 14752 12396 14872 12424
rect 14924 12436 14976 12442
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14556 11076 14608 11082
rect 14556 11018 14608 11024
rect 14294 10908 14602 10928
rect 14294 10906 14300 10908
rect 14356 10906 14380 10908
rect 14436 10906 14460 10908
rect 14516 10906 14540 10908
rect 14596 10906 14602 10908
rect 14356 10854 14358 10906
rect 14538 10854 14540 10906
rect 14294 10852 14300 10854
rect 14356 10852 14380 10854
rect 14436 10852 14460 10854
rect 14516 10852 14540 10854
rect 14596 10852 14602 10854
rect 14294 10832 14602 10852
rect 14188 10804 14240 10810
rect 14188 10746 14240 10752
rect 14660 10742 14688 11494
rect 14648 10736 14700 10742
rect 14648 10678 14700 10684
rect 14096 10600 14148 10606
rect 14096 10542 14148 10548
rect 14370 10432 14426 10441
rect 14370 10367 14426 10376
rect 14096 10124 14148 10130
rect 14096 10066 14148 10072
rect 14108 9722 14136 10066
rect 14384 10062 14412 10367
rect 14554 10296 14610 10305
rect 14752 10266 14780 12396
rect 14924 12378 14976 12384
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14844 11121 14872 12242
rect 15120 12186 15148 12702
rect 15200 12640 15252 12646
rect 15198 12608 15200 12617
rect 15252 12608 15254 12617
rect 15198 12543 15254 12552
rect 15120 12158 15240 12186
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15106 12064 15162 12073
rect 14936 11898 14964 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 14830 11112 14886 11121
rect 14830 11047 14886 11056
rect 14832 10464 14884 10470
rect 14936 10418 14964 11698
rect 15028 11354 15056 12038
rect 15106 11999 15162 12008
rect 15120 11830 15148 11999
rect 15108 11824 15160 11830
rect 15108 11766 15160 11772
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14884 10412 14964 10418
rect 14832 10406 14964 10412
rect 14844 10390 14964 10406
rect 14554 10231 14610 10240
rect 14740 10260 14792 10266
rect 14372 10056 14424 10062
rect 14372 9998 14424 10004
rect 14568 9908 14596 10231
rect 14740 10202 14792 10208
rect 14936 10198 14964 10390
rect 14924 10192 14976 10198
rect 14646 10160 14702 10169
rect 14702 10118 14780 10146
rect 14924 10134 14976 10140
rect 14646 10095 14702 10104
rect 14568 9880 14688 9908
rect 14752 9897 14780 10118
rect 14832 9920 14884 9926
rect 14294 9820 14602 9840
rect 14294 9818 14300 9820
rect 14356 9818 14380 9820
rect 14436 9818 14460 9820
rect 14516 9818 14540 9820
rect 14596 9818 14602 9820
rect 14356 9766 14358 9818
rect 14538 9766 14540 9818
rect 14294 9764 14300 9766
rect 14356 9764 14380 9766
rect 14436 9764 14460 9766
rect 14516 9764 14540 9766
rect 14596 9764 14602 9766
rect 14294 9744 14602 9764
rect 14096 9716 14148 9722
rect 14096 9658 14148 9664
rect 14108 9178 14136 9658
rect 14188 9648 14240 9654
rect 14188 9590 14240 9596
rect 14004 9172 14056 9178
rect 14004 9114 14056 9120
rect 14096 9172 14148 9178
rect 14096 9114 14148 9120
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13728 8628 13780 8634
rect 13832 8616 13860 9046
rect 13924 9030 14044 9058
rect 13912 8628 13964 8634
rect 13832 8588 13912 8616
rect 13728 8570 13780 8576
rect 13912 8570 13964 8576
rect 13740 8514 13768 8570
rect 13740 8486 13860 8514
rect 13832 8090 13860 8486
rect 13912 8424 13964 8430
rect 13912 8366 13964 8372
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13818 7984 13874 7993
rect 13818 7919 13874 7928
rect 13832 7750 13860 7919
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13740 7274 13768 7686
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 6866 13768 7210
rect 13832 6882 13860 7686
rect 13924 7546 13952 8366
rect 14016 7886 14044 9030
rect 14108 8430 14136 9114
rect 14200 8974 14228 9590
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14200 7886 14228 8910
rect 14294 8732 14602 8752
rect 14294 8730 14300 8732
rect 14356 8730 14380 8732
rect 14436 8730 14460 8732
rect 14516 8730 14540 8732
rect 14596 8730 14602 8732
rect 14356 8678 14358 8730
rect 14538 8678 14540 8730
rect 14294 8676 14300 8678
rect 14356 8676 14380 8678
rect 14436 8676 14460 8678
rect 14516 8676 14540 8678
rect 14596 8676 14602 8678
rect 14294 8656 14602 8676
rect 14556 8288 14608 8294
rect 14556 8230 14608 8236
rect 14568 7886 14596 8230
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14556 7880 14608 7886
rect 14556 7822 14608 7828
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 14004 7200 14056 7206
rect 14004 7142 14056 7148
rect 14016 7002 14044 7142
rect 14004 6996 14056 7002
rect 14004 6938 14056 6944
rect 13728 6860 13780 6866
rect 13832 6854 13952 6882
rect 13728 6802 13780 6808
rect 13820 6724 13872 6730
rect 13820 6666 13872 6672
rect 13728 6316 13780 6322
rect 13728 6258 13780 6264
rect 13740 6066 13768 6258
rect 13832 6254 13860 6666
rect 13820 6248 13872 6254
rect 13820 6190 13872 6196
rect 13924 6066 13952 6854
rect 14002 6624 14058 6633
rect 14002 6559 14058 6568
rect 14016 6390 14044 6559
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 14002 6216 14058 6225
rect 14002 6151 14058 6160
rect 13740 6038 13952 6066
rect 13832 5234 13860 6038
rect 14016 5930 14044 6151
rect 13924 5902 14044 5930
rect 13924 5710 13952 5902
rect 13912 5704 13964 5710
rect 13912 5646 13964 5652
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13726 4448 13782 4457
rect 13726 4383 13782 4392
rect 13740 4146 13768 4383
rect 13832 4282 13860 4558
rect 13924 4486 13952 5646
rect 14002 5536 14058 5545
rect 14002 5471 14058 5480
rect 14016 5370 14044 5471
rect 14004 5364 14056 5370
rect 14004 5306 14056 5312
rect 13912 4480 13964 4486
rect 13912 4422 13964 4428
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13924 4185 13952 4422
rect 14016 4282 14044 5306
rect 14108 4298 14136 7686
rect 14200 7206 14228 7822
rect 14294 7644 14602 7664
rect 14294 7642 14300 7644
rect 14356 7642 14380 7644
rect 14436 7642 14460 7644
rect 14516 7642 14540 7644
rect 14596 7642 14602 7644
rect 14356 7590 14358 7642
rect 14538 7590 14540 7642
rect 14294 7588 14300 7590
rect 14356 7588 14380 7590
rect 14436 7588 14460 7590
rect 14516 7588 14540 7590
rect 14596 7588 14602 7590
rect 14294 7568 14602 7588
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14294 6556 14602 6576
rect 14294 6554 14300 6556
rect 14356 6554 14380 6556
rect 14436 6554 14460 6556
rect 14516 6554 14540 6556
rect 14596 6554 14602 6556
rect 14356 6502 14358 6554
rect 14538 6502 14540 6554
rect 14294 6500 14300 6502
rect 14356 6500 14380 6502
rect 14436 6500 14460 6502
rect 14516 6500 14540 6502
rect 14596 6500 14602 6502
rect 14294 6480 14602 6500
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14568 5778 14596 6054
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14660 5681 14688 9880
rect 14738 9888 14794 9897
rect 14832 9862 14884 9868
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14738 9823 14794 9832
rect 14844 9722 14872 9862
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14936 9586 14964 9862
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14752 9382 14780 9454
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14922 8392 14978 8401
rect 14922 8327 14978 8336
rect 14740 7744 14792 7750
rect 14740 7686 14792 7692
rect 14646 5672 14702 5681
rect 14646 5607 14702 5616
rect 14294 5468 14602 5488
rect 14294 5466 14300 5468
rect 14356 5466 14380 5468
rect 14436 5466 14460 5468
rect 14516 5466 14540 5468
rect 14596 5466 14602 5468
rect 14356 5414 14358 5466
rect 14538 5414 14540 5466
rect 14294 5412 14300 5414
rect 14356 5412 14380 5414
rect 14436 5412 14460 5414
rect 14516 5412 14540 5414
rect 14596 5412 14602 5414
rect 14294 5392 14602 5412
rect 14646 5264 14702 5273
rect 14646 5199 14702 5208
rect 14294 4380 14602 4400
rect 14294 4378 14300 4380
rect 14356 4378 14380 4380
rect 14436 4378 14460 4380
rect 14516 4378 14540 4380
rect 14596 4378 14602 4380
rect 14356 4326 14358 4378
rect 14538 4326 14540 4378
rect 14294 4324 14300 4326
rect 14356 4324 14380 4326
rect 14436 4324 14460 4326
rect 14516 4324 14540 4326
rect 14596 4324 14602 4326
rect 14294 4304 14602 4324
rect 14004 4276 14056 4282
rect 14108 4270 14228 4298
rect 14004 4218 14056 4224
rect 14096 4208 14148 4214
rect 13910 4176 13966 4185
rect 13728 4140 13780 4146
rect 14096 4150 14148 4156
rect 13910 4111 13966 4120
rect 13728 4082 13780 4088
rect 14004 4072 14056 4078
rect 13818 4040 13874 4049
rect 14004 4014 14056 4020
rect 13818 3975 13820 3984
rect 13872 3975 13874 3984
rect 13820 3946 13872 3952
rect 13728 3460 13780 3466
rect 13728 3402 13780 3408
rect 13740 2990 13768 3402
rect 13820 3188 13872 3194
rect 13820 3130 13872 3136
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 13832 1442 13860 3130
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13924 2650 13952 2994
rect 14016 2961 14044 4014
rect 14108 3194 14136 4150
rect 14200 3194 14228 4270
rect 14462 3768 14518 3777
rect 14660 3738 14688 5199
rect 14752 4706 14780 7686
rect 14832 6724 14884 6730
rect 14832 6666 14884 6672
rect 14844 6254 14872 6666
rect 14832 6248 14884 6254
rect 14832 6190 14884 6196
rect 14844 5914 14872 6190
rect 14832 5908 14884 5914
rect 14832 5850 14884 5856
rect 14844 5574 14872 5850
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14752 4678 14872 4706
rect 14740 4548 14792 4554
rect 14740 4490 14792 4496
rect 14752 4078 14780 4490
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14462 3703 14518 3712
rect 14648 3732 14700 3738
rect 14476 3534 14504 3703
rect 14648 3674 14700 3680
rect 14752 3602 14780 4014
rect 14740 3596 14792 3602
rect 14660 3556 14740 3584
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14294 3292 14602 3312
rect 14294 3290 14300 3292
rect 14356 3290 14380 3292
rect 14436 3290 14460 3292
rect 14516 3290 14540 3292
rect 14596 3290 14602 3292
rect 14356 3238 14358 3290
rect 14538 3238 14540 3290
rect 14294 3236 14300 3238
rect 14356 3236 14380 3238
rect 14436 3236 14460 3238
rect 14516 3236 14540 3238
rect 14596 3236 14602 3238
rect 14294 3216 14602 3236
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14462 3088 14518 3097
rect 14462 3023 14464 3032
rect 14516 3023 14518 3032
rect 14464 2994 14516 3000
rect 14660 2990 14688 3556
rect 14740 3538 14792 3544
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14372 2984 14424 2990
rect 14002 2952 14058 2961
rect 14372 2926 14424 2932
rect 14648 2984 14700 2990
rect 14648 2926 14700 2932
rect 14002 2887 14058 2896
rect 14384 2650 14412 2926
rect 14660 2854 14688 2926
rect 14648 2848 14700 2854
rect 14648 2790 14700 2796
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14372 2644 14424 2650
rect 14372 2586 14424 2592
rect 14200 2496 14228 2586
rect 14752 2582 14780 3062
rect 14844 2938 14872 4678
rect 14936 3058 14964 8327
rect 15028 6633 15056 11018
rect 15108 10600 15160 10606
rect 15108 10542 15160 10548
rect 15120 7342 15148 10542
rect 15212 9994 15240 12158
rect 15304 12102 15332 13484
rect 15488 13410 15516 14311
rect 15856 14249 15884 14350
rect 15842 14240 15898 14249
rect 15842 14175 15898 14184
rect 15660 14068 15712 14074
rect 15712 14028 15792 14056
rect 15660 14010 15712 14016
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15396 13382 15516 13410
rect 15568 13456 15620 13462
rect 15568 13398 15620 13404
rect 15396 13326 15424 13382
rect 15384 13320 15436 13326
rect 15384 13262 15436 13268
rect 15476 13320 15528 13326
rect 15580 13297 15608 13398
rect 15476 13262 15528 13268
rect 15566 13288 15622 13297
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 13025 15424 13126
rect 15382 13016 15438 13025
rect 15382 12951 15438 12960
rect 15488 12850 15516 13262
rect 15566 13223 15622 13232
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15304 11529 15332 11834
rect 15290 11520 15346 11529
rect 15290 11455 15346 11464
rect 15396 11014 15424 12650
rect 15580 11642 15608 13126
rect 15672 12850 15700 13466
rect 15764 13190 15792 14028
rect 15844 13932 15896 13938
rect 15844 13874 15896 13880
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 15856 13433 15884 13874
rect 16026 13832 16082 13841
rect 16026 13767 16082 13776
rect 15842 13424 15898 13433
rect 15842 13359 15898 13368
rect 15752 13184 15804 13190
rect 15752 13126 15804 13132
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 15660 12844 15712 12850
rect 15660 12786 15712 12792
rect 15672 11937 15700 12786
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15658 11928 15714 11937
rect 15658 11863 15714 11872
rect 15764 11830 15792 12038
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15580 11614 15792 11642
rect 15568 11552 15620 11558
rect 15474 11520 15530 11529
rect 15568 11494 15620 11500
rect 15660 11552 15712 11558
rect 15660 11494 15712 11500
rect 15474 11455 15530 11464
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15200 9988 15252 9994
rect 15200 9930 15252 9936
rect 15384 9988 15436 9994
rect 15384 9930 15436 9936
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 8945 15332 9658
rect 15396 9217 15424 9930
rect 15382 9208 15438 9217
rect 15382 9143 15438 9152
rect 15290 8936 15346 8945
rect 15200 8900 15252 8906
rect 15290 8871 15346 8880
rect 15200 8842 15252 8848
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15212 7274 15240 8842
rect 15488 8650 15516 11455
rect 15580 9654 15608 11494
rect 15672 11082 15700 11494
rect 15660 11076 15712 11082
rect 15660 11018 15712 11024
rect 15658 10976 15714 10985
rect 15658 10911 15714 10920
rect 15672 9994 15700 10911
rect 15660 9988 15712 9994
rect 15660 9930 15712 9936
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15658 9344 15714 9353
rect 15658 9279 15714 9288
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15396 8622 15516 8650
rect 15304 8498 15332 8570
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15396 7426 15424 8622
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 15488 7546 15516 8502
rect 15476 7540 15528 7546
rect 15476 7482 15528 7488
rect 15396 7410 15516 7426
rect 15396 7404 15528 7410
rect 15396 7398 15476 7404
rect 15292 7336 15344 7342
rect 15396 7313 15424 7398
rect 15476 7346 15528 7352
rect 15292 7278 15344 7284
rect 15382 7304 15438 7313
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15304 7177 15332 7278
rect 15382 7239 15438 7248
rect 15290 7168 15346 7177
rect 15290 7103 15346 7112
rect 15106 7032 15162 7041
rect 15106 6967 15162 6976
rect 15200 6996 15252 7002
rect 15014 6624 15070 6633
rect 15014 6559 15070 6568
rect 15016 6452 15068 6458
rect 15016 6394 15068 6400
rect 15028 6361 15056 6394
rect 15014 6352 15070 6361
rect 15014 6287 15070 6296
rect 15014 5944 15070 5953
rect 15014 5879 15070 5888
rect 15028 5642 15056 5879
rect 15016 5636 15068 5642
rect 15016 5578 15068 5584
rect 15028 5302 15056 5578
rect 15016 5296 15068 5302
rect 15016 5238 15068 5244
rect 15120 4826 15148 6967
rect 15200 6938 15252 6944
rect 15212 6390 15240 6938
rect 15384 6792 15436 6798
rect 15384 6734 15436 6740
rect 15292 6656 15344 6662
rect 15292 6598 15344 6604
rect 15200 6384 15252 6390
rect 15200 6326 15252 6332
rect 15198 5808 15254 5817
rect 15198 5743 15254 5752
rect 15108 4820 15160 4826
rect 15108 4762 15160 4768
rect 15014 4720 15070 4729
rect 15014 4655 15070 4664
rect 15028 3942 15056 4655
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15120 4049 15148 4082
rect 15106 4040 15162 4049
rect 15106 3975 15162 3984
rect 15016 3936 15068 3942
rect 15016 3878 15068 3884
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 15028 2990 15056 3878
rect 15212 3534 15240 5743
rect 15304 5574 15332 6598
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15396 5030 15424 6734
rect 15580 6730 15608 8842
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15476 6384 15528 6390
rect 15672 6361 15700 9279
rect 15764 8378 15792 11614
rect 15856 11529 15884 12922
rect 16040 12850 16068 13767
rect 16132 13530 16160 13874
rect 16224 13530 16252 14719
rect 16316 14414 16344 14962
rect 17314 14920 17370 14929
rect 16396 14884 16448 14890
rect 17314 14855 17370 14864
rect 16396 14826 16448 14832
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16408 14249 16436 14826
rect 16518 14716 16826 14736
rect 16518 14714 16524 14716
rect 16580 14714 16604 14716
rect 16660 14714 16684 14716
rect 16740 14714 16764 14716
rect 16820 14714 16826 14716
rect 16580 14662 16582 14714
rect 16762 14662 16764 14714
rect 16518 14660 16524 14662
rect 16580 14660 16604 14662
rect 16660 14660 16684 14662
rect 16740 14660 16764 14662
rect 16820 14660 16826 14662
rect 16518 14640 16826 14660
rect 16946 14648 17002 14657
rect 16946 14583 17002 14592
rect 16960 14482 16988 14583
rect 17328 14482 17356 14855
rect 17604 14482 17632 15098
rect 17696 15094 17724 16079
rect 17684 15088 17736 15094
rect 17684 15030 17736 15036
rect 16948 14476 17000 14482
rect 16948 14418 17000 14424
rect 17316 14476 17368 14482
rect 17316 14418 17368 14424
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17408 14340 17460 14346
rect 17408 14282 17460 14288
rect 16394 14240 16450 14249
rect 16394 14175 16450 14184
rect 16408 13870 16436 14175
rect 16396 13864 16448 13870
rect 16396 13806 16448 13812
rect 17132 13864 17184 13870
rect 17132 13806 17184 13812
rect 17040 13728 17092 13734
rect 17040 13670 17092 13676
rect 16518 13628 16826 13648
rect 16518 13626 16524 13628
rect 16580 13626 16604 13628
rect 16660 13626 16684 13628
rect 16740 13626 16764 13628
rect 16820 13626 16826 13628
rect 16580 13574 16582 13626
rect 16762 13574 16764 13626
rect 16518 13572 16524 13574
rect 16580 13572 16604 13574
rect 16660 13572 16684 13574
rect 16740 13572 16764 13574
rect 16820 13572 16826 13574
rect 16302 13560 16358 13569
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 16212 13524 16264 13530
rect 16518 13552 16826 13572
rect 16358 13504 16528 13512
rect 16302 13495 16528 13504
rect 16316 13484 16528 13495
rect 16212 13466 16264 13472
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16210 12744 16266 12753
rect 16210 12679 16212 12688
rect 16264 12679 16266 12688
rect 16212 12650 16264 12656
rect 16408 12646 16436 13194
rect 16500 13161 16528 13484
rect 16856 13388 16908 13394
rect 16856 13330 16908 13336
rect 16486 13152 16542 13161
rect 16486 13087 16542 13096
rect 16500 12850 16528 13087
rect 16488 12844 16540 12850
rect 16488 12786 16540 12792
rect 16396 12640 16448 12646
rect 16396 12582 16448 12588
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 15936 12096 15988 12102
rect 15936 12038 15988 12044
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 15842 11520 15898 11529
rect 15842 11455 15898 11464
rect 15844 11348 15896 11354
rect 15844 11290 15896 11296
rect 15856 10130 15884 11290
rect 15844 10124 15896 10130
rect 15844 10066 15896 10072
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8498 15884 8910
rect 15948 8498 15976 12038
rect 16132 11898 16160 12038
rect 16224 11898 16252 12106
rect 16120 11892 16172 11898
rect 16120 11834 16172 11840
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 16040 10266 16068 11494
rect 16028 10260 16080 10266
rect 16028 10202 16080 10208
rect 16040 10130 16068 10202
rect 16028 10124 16080 10130
rect 16028 10066 16080 10072
rect 16132 9450 16160 11630
rect 16224 11234 16252 11834
rect 16304 11756 16356 11762
rect 16304 11698 16356 11704
rect 16316 11354 16344 11698
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16224 11206 16344 11234
rect 16212 11144 16264 11150
rect 16212 11086 16264 11092
rect 16224 10606 16252 11086
rect 16316 10713 16344 11206
rect 16408 10742 16436 12582
rect 16518 12540 16826 12560
rect 16518 12538 16524 12540
rect 16580 12538 16604 12540
rect 16660 12538 16684 12540
rect 16740 12538 16764 12540
rect 16820 12538 16826 12540
rect 16580 12486 16582 12538
rect 16762 12486 16764 12538
rect 16518 12484 16524 12486
rect 16580 12484 16604 12486
rect 16660 12484 16684 12486
rect 16740 12484 16764 12486
rect 16820 12484 16826 12486
rect 16518 12464 16826 12484
rect 16518 11452 16826 11472
rect 16518 11450 16524 11452
rect 16580 11450 16604 11452
rect 16660 11450 16684 11452
rect 16740 11450 16764 11452
rect 16820 11450 16826 11452
rect 16580 11398 16582 11450
rect 16762 11398 16764 11450
rect 16518 11396 16524 11398
rect 16580 11396 16604 11398
rect 16660 11396 16684 11398
rect 16740 11396 16764 11398
rect 16820 11396 16826 11398
rect 16518 11376 16826 11396
rect 16868 10742 16896 13330
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16960 12073 16988 12378
rect 16946 12064 17002 12073
rect 16946 11999 17002 12008
rect 16396 10736 16448 10742
rect 16302 10704 16358 10713
rect 16396 10678 16448 10684
rect 16856 10736 16908 10742
rect 16856 10678 16908 10684
rect 16302 10639 16358 10648
rect 16212 10600 16264 10606
rect 16212 10542 16264 10548
rect 16304 10600 16356 10606
rect 16304 10542 16356 10548
rect 16856 10600 16908 10606
rect 16856 10542 16908 10548
rect 16120 9444 16172 9450
rect 16120 9386 16172 9392
rect 16132 9042 16160 9386
rect 16120 9036 16172 9042
rect 16120 8978 16172 8984
rect 16224 8974 16252 10542
rect 16316 10062 16344 10542
rect 16518 10364 16826 10384
rect 16518 10362 16524 10364
rect 16580 10362 16604 10364
rect 16660 10362 16684 10364
rect 16740 10362 16764 10364
rect 16820 10362 16826 10364
rect 16580 10310 16582 10362
rect 16762 10310 16764 10362
rect 16518 10308 16524 10310
rect 16580 10308 16604 10310
rect 16660 10308 16684 10310
rect 16740 10308 16764 10310
rect 16820 10308 16826 10310
rect 16518 10288 16826 10308
rect 16394 10160 16450 10169
rect 16394 10095 16450 10104
rect 16304 10056 16356 10062
rect 16304 9998 16356 10004
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16304 8900 16356 8906
rect 16304 8842 16356 8848
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 15844 8492 15896 8498
rect 15844 8434 15896 8440
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 15764 8350 15884 8378
rect 15476 6326 15528 6332
rect 15658 6352 15714 6361
rect 15488 6254 15516 6326
rect 15658 6287 15714 6296
rect 15752 6316 15804 6322
rect 15752 6258 15804 6264
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15488 5778 15516 6190
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5846 15608 6054
rect 15568 5840 15620 5846
rect 15568 5782 15620 5788
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 15764 5574 15792 6258
rect 15856 6089 15884 8350
rect 15934 7576 15990 7585
rect 15934 7511 15990 7520
rect 15948 7002 15976 7511
rect 15936 6996 15988 7002
rect 15936 6938 15988 6944
rect 16040 6338 16068 8570
rect 16316 8498 16344 8842
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16120 8356 16172 8362
rect 16120 8298 16172 8304
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16132 6916 16160 8298
rect 16224 7954 16252 8298
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16210 7848 16266 7857
rect 16210 7783 16266 7792
rect 16224 7478 16252 7783
rect 16316 7585 16344 8230
rect 16302 7576 16358 7585
rect 16302 7511 16358 7520
rect 16212 7472 16264 7478
rect 16212 7414 16264 7420
rect 16302 7168 16358 7177
rect 16302 7103 16358 7112
rect 16132 6888 16252 6916
rect 15948 6310 16068 6338
rect 15842 6080 15898 6089
rect 15842 6015 15898 6024
rect 15948 5930 15976 6310
rect 16120 6248 16172 6254
rect 16026 6216 16082 6225
rect 16120 6190 16172 6196
rect 16026 6151 16082 6160
rect 15856 5902 15976 5930
rect 15752 5568 15804 5574
rect 15752 5510 15804 5516
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4622 15424 4966
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15292 4480 15344 4486
rect 15292 4422 15344 4428
rect 15304 3670 15332 4422
rect 15396 4214 15424 4558
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15384 4208 15436 4214
rect 15384 4150 15436 4156
rect 15384 4004 15436 4010
rect 15384 3946 15436 3952
rect 15292 3664 15344 3670
rect 15292 3606 15344 3612
rect 15396 3602 15424 3946
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15384 3596 15436 3602
rect 15384 3538 15436 3544
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15304 3058 15332 3334
rect 15382 3224 15438 3233
rect 15382 3159 15384 3168
rect 15436 3159 15438 3168
rect 15384 3130 15436 3136
rect 15292 3052 15344 3058
rect 15292 2994 15344 3000
rect 15016 2984 15068 2990
rect 14844 2910 14964 2938
rect 15488 2961 15516 3674
rect 15580 3194 15608 4422
rect 15660 3596 15712 3602
rect 15660 3538 15712 3544
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15016 2926 15068 2932
rect 15474 2952 15530 2961
rect 14936 2854 14964 2910
rect 15474 2887 15530 2896
rect 14924 2848 14976 2854
rect 14830 2816 14886 2825
rect 14924 2790 14976 2796
rect 14830 2751 14886 2760
rect 14740 2576 14792 2582
rect 14740 2518 14792 2524
rect 14372 2508 14424 2514
rect 14200 2468 14372 2496
rect 14372 2450 14424 2456
rect 14294 2204 14602 2224
rect 14294 2202 14300 2204
rect 14356 2202 14380 2204
rect 14436 2202 14460 2204
rect 14516 2202 14540 2204
rect 14596 2202 14602 2204
rect 14356 2150 14358 2202
rect 14538 2150 14540 2202
rect 14294 2148 14300 2150
rect 14356 2148 14380 2150
rect 14436 2148 14460 2150
rect 14516 2148 14540 2150
rect 14596 2148 14602 2150
rect 14294 2128 14602 2148
rect 13832 1414 13952 1442
rect 13636 1352 13688 1358
rect 13636 1294 13688 1300
rect 13924 800 13952 1414
rect 14844 800 14872 2751
rect 15672 2446 15700 3538
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 15660 2440 15712 2446
rect 15660 2382 15712 2388
rect 14936 2106 14964 2382
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 15764 1698 15792 3334
rect 15856 3058 15884 5902
rect 15936 5840 15988 5846
rect 15936 5782 15988 5788
rect 15948 4622 15976 5782
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 15948 1737 15976 3334
rect 16040 3126 16068 6151
rect 16132 5914 16160 6190
rect 16120 5908 16172 5914
rect 16120 5850 16172 5856
rect 16120 5704 16172 5710
rect 16120 5646 16172 5652
rect 16132 3466 16160 5646
rect 16224 5545 16252 6888
rect 16210 5536 16266 5545
rect 16210 5471 16266 5480
rect 16316 5114 16344 7103
rect 16408 6916 16436 10095
rect 16488 9920 16540 9926
rect 16488 9862 16540 9868
rect 16500 9654 16528 9862
rect 16762 9752 16818 9761
rect 16762 9687 16818 9696
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16776 9586 16804 9687
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16518 9276 16826 9296
rect 16518 9274 16524 9276
rect 16580 9274 16604 9276
rect 16660 9274 16684 9276
rect 16740 9274 16764 9276
rect 16820 9274 16826 9276
rect 16580 9222 16582 9274
rect 16762 9222 16764 9274
rect 16518 9220 16524 9222
rect 16580 9220 16604 9222
rect 16660 9220 16684 9222
rect 16740 9220 16764 9222
rect 16820 9220 16826 9222
rect 16518 9200 16826 9220
rect 16868 8566 16896 10542
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16960 10062 16988 10406
rect 17052 10266 17080 13670
rect 17144 12434 17172 13806
rect 17144 12406 17356 12434
rect 17222 12200 17278 12209
rect 17222 12135 17224 12144
rect 17276 12135 17278 12144
rect 17224 12106 17276 12112
rect 17132 11552 17184 11558
rect 17132 11494 17184 11500
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17040 9648 17092 9654
rect 17038 9616 17040 9625
rect 17092 9616 17094 9625
rect 17038 9551 17094 9560
rect 17144 8974 17172 11494
rect 17236 10849 17264 12106
rect 17328 10985 17356 12406
rect 17314 10976 17370 10985
rect 17314 10911 17370 10920
rect 17222 10840 17278 10849
rect 17222 10775 17278 10784
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 17236 9722 17264 10134
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17132 8968 17184 8974
rect 17132 8910 17184 8916
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17144 8634 17172 8774
rect 17132 8628 17184 8634
rect 17132 8570 17184 8576
rect 16856 8560 16908 8566
rect 16856 8502 16908 8508
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16518 8188 16826 8208
rect 16518 8186 16524 8188
rect 16580 8186 16604 8188
rect 16660 8186 16684 8188
rect 16740 8186 16764 8188
rect 16820 8186 16826 8188
rect 16580 8134 16582 8186
rect 16762 8134 16764 8186
rect 16518 8132 16524 8134
rect 16580 8132 16604 8134
rect 16660 8132 16684 8134
rect 16740 8132 16764 8134
rect 16820 8132 16826 8134
rect 16518 8112 16826 8132
rect 17052 7857 17080 8434
rect 17236 8430 17264 8774
rect 17328 8634 17356 10610
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17236 7954 17264 8366
rect 17316 8084 17368 8090
rect 17316 8026 17368 8032
rect 17224 7948 17276 7954
rect 17224 7890 17276 7896
rect 17038 7848 17094 7857
rect 16948 7812 17000 7818
rect 17038 7783 17094 7792
rect 16948 7754 17000 7760
rect 16672 7744 16724 7750
rect 16672 7686 16724 7692
rect 16856 7744 16908 7750
rect 16856 7686 16908 7692
rect 16684 7478 16712 7686
rect 16672 7472 16724 7478
rect 16672 7414 16724 7420
rect 16670 7304 16726 7313
rect 16670 7239 16672 7248
rect 16724 7239 16726 7248
rect 16672 7210 16724 7216
rect 16518 7100 16826 7120
rect 16518 7098 16524 7100
rect 16580 7098 16604 7100
rect 16660 7098 16684 7100
rect 16740 7098 16764 7100
rect 16820 7098 16826 7100
rect 16580 7046 16582 7098
rect 16762 7046 16764 7098
rect 16518 7044 16524 7046
rect 16580 7044 16604 7046
rect 16660 7044 16684 7046
rect 16740 7044 16764 7046
rect 16820 7044 16826 7046
rect 16518 7024 16826 7044
rect 16408 6888 16528 6916
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16224 5086 16344 5114
rect 16224 4486 16252 5086
rect 16304 5024 16356 5030
rect 16304 4966 16356 4972
rect 16316 4690 16344 4966
rect 16304 4684 16356 4690
rect 16304 4626 16356 4632
rect 16212 4480 16264 4486
rect 16212 4422 16264 4428
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16118 3224 16174 3233
rect 16118 3159 16174 3168
rect 16028 3120 16080 3126
rect 16028 3062 16080 3068
rect 16132 3058 16160 3159
rect 16224 3097 16252 4422
rect 16316 4146 16344 4626
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 16408 4010 16436 6666
rect 16500 6662 16528 6888
rect 16672 6792 16724 6798
rect 16868 6769 16896 7686
rect 16960 7546 16988 7754
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 17236 6934 17264 7890
rect 17328 7342 17356 8026
rect 17316 7336 17368 7342
rect 17316 7278 17368 7284
rect 17224 6928 17276 6934
rect 17130 6896 17186 6905
rect 17224 6870 17276 6876
rect 17130 6831 17186 6840
rect 17144 6798 17172 6831
rect 17132 6792 17184 6798
rect 16672 6734 16724 6740
rect 16854 6760 16910 6769
rect 16488 6656 16540 6662
rect 16488 6598 16540 6604
rect 16684 6254 16712 6734
rect 17132 6734 17184 6740
rect 16854 6695 16910 6704
rect 16856 6656 16908 6662
rect 16856 6598 16908 6604
rect 17040 6656 17092 6662
rect 17040 6598 17092 6604
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16518 6012 16826 6032
rect 16518 6010 16524 6012
rect 16580 6010 16604 6012
rect 16660 6010 16684 6012
rect 16740 6010 16764 6012
rect 16820 6010 16826 6012
rect 16580 5958 16582 6010
rect 16762 5958 16764 6010
rect 16518 5956 16524 5958
rect 16580 5956 16604 5958
rect 16660 5956 16684 5958
rect 16740 5956 16764 5958
rect 16820 5956 16826 5958
rect 16518 5936 16826 5956
rect 16762 5808 16818 5817
rect 16762 5743 16818 5752
rect 16776 5234 16804 5743
rect 16868 5574 16896 6598
rect 17052 6390 17080 6598
rect 17040 6384 17092 6390
rect 16946 6352 17002 6361
rect 17040 6326 17092 6332
rect 16946 6287 17002 6296
rect 16960 5953 16988 6287
rect 16946 5944 17002 5953
rect 16946 5879 17002 5888
rect 16856 5568 16908 5574
rect 16856 5510 16908 5516
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16518 4924 16826 4944
rect 16518 4922 16524 4924
rect 16580 4922 16604 4924
rect 16660 4922 16684 4924
rect 16740 4922 16764 4924
rect 16820 4922 16826 4924
rect 16580 4870 16582 4922
rect 16762 4870 16764 4922
rect 16518 4868 16524 4870
rect 16580 4868 16604 4870
rect 16660 4868 16684 4870
rect 16740 4868 16764 4870
rect 16820 4868 16826 4870
rect 16518 4848 16826 4868
rect 16396 4004 16448 4010
rect 16396 3946 16448 3952
rect 16518 3836 16826 3856
rect 16518 3834 16524 3836
rect 16580 3834 16604 3836
rect 16660 3834 16684 3836
rect 16740 3834 16764 3836
rect 16820 3834 16826 3836
rect 16580 3782 16582 3834
rect 16762 3782 16764 3834
rect 16518 3780 16524 3782
rect 16580 3780 16604 3782
rect 16660 3780 16684 3782
rect 16740 3780 16764 3782
rect 16820 3780 16826 3782
rect 16518 3760 16826 3780
rect 16670 3632 16726 3641
rect 16868 3618 16896 5510
rect 17040 5296 17092 5302
rect 17040 5238 17092 5244
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16670 3567 16726 3576
rect 16776 3590 16896 3618
rect 16488 3460 16540 3466
rect 16488 3402 16540 3408
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 16408 3194 16436 3334
rect 16500 3194 16528 3402
rect 16396 3188 16448 3194
rect 16396 3130 16448 3136
rect 16488 3188 16540 3194
rect 16488 3130 16540 3136
rect 16210 3088 16266 3097
rect 16120 3052 16172 3058
rect 16684 3058 16712 3567
rect 16776 3058 16804 3590
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16210 3023 16266 3032
rect 16672 3052 16724 3058
rect 16120 2994 16172 3000
rect 16672 2994 16724 3000
rect 16764 3052 16816 3058
rect 16764 2994 16816 3000
rect 16518 2748 16826 2768
rect 16518 2746 16524 2748
rect 16580 2746 16604 2748
rect 16660 2746 16684 2748
rect 16740 2746 16764 2748
rect 16820 2746 16826 2748
rect 16580 2694 16582 2746
rect 16762 2694 16764 2746
rect 16518 2692 16524 2694
rect 16580 2692 16604 2694
rect 16660 2692 16684 2694
rect 16740 2692 16764 2694
rect 16820 2692 16826 2694
rect 16518 2672 16826 2692
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16408 2038 16436 2246
rect 16396 2032 16448 2038
rect 16396 1974 16448 1980
rect 16684 1834 16712 2382
rect 16672 1828 16724 1834
rect 16672 1770 16724 1776
rect 15934 1728 15990 1737
rect 15752 1692 15804 1698
rect 15934 1663 15990 1672
rect 15752 1634 15804 1640
rect 16868 1442 16896 3402
rect 16684 1414 16896 1442
rect 15200 1352 15252 1358
rect 15200 1294 15252 1300
rect 15934 1320 15990 1329
rect 8588 734 8800 762
rect 9402 0 9458 800
rect 10322 0 10378 800
rect 11242 0 11298 800
rect 12162 0 12218 800
rect 13082 0 13138 800
rect 13910 0 13966 800
rect 14830 0 14886 800
rect 15212 241 15240 1294
rect 15934 1255 15936 1264
rect 15988 1255 15990 1264
rect 15936 1226 15988 1232
rect 15844 1216 15896 1222
rect 15844 1158 15896 1164
rect 15672 870 15792 898
rect 15198 232 15254 241
rect 15198 167 15254 176
rect 15672 66 15700 870
rect 15764 800 15792 870
rect 15660 60 15712 66
rect 15660 2 15712 8
rect 15750 0 15806 800
rect 15856 513 15884 1158
rect 16684 800 16712 1414
rect 16960 921 16988 4966
rect 17052 4690 17080 5238
rect 17132 5024 17184 5030
rect 17132 4966 17184 4972
rect 17040 4684 17092 4690
rect 17040 4626 17092 4632
rect 17038 4176 17094 4185
rect 17038 4111 17094 4120
rect 17052 3126 17080 4111
rect 17144 3534 17172 4966
rect 17328 4146 17356 7278
rect 17420 5710 17448 14282
rect 17592 14272 17644 14278
rect 17592 14214 17644 14220
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17512 10538 17540 12174
rect 17604 11132 17632 14214
rect 17696 13870 17724 15030
rect 17880 14618 17908 16400
rect 17960 15564 18012 15570
rect 17960 15506 18012 15512
rect 17868 14612 17920 14618
rect 17868 14554 17920 14560
rect 17684 13864 17736 13870
rect 17684 13806 17736 13812
rect 17868 13388 17920 13394
rect 17868 13330 17920 13336
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17682 12744 17738 12753
rect 17682 12679 17738 12688
rect 17696 12345 17724 12679
rect 17682 12336 17738 12345
rect 17682 12271 17684 12280
rect 17736 12271 17738 12280
rect 17684 12242 17736 12248
rect 17684 11688 17736 11694
rect 17788 11665 17816 13194
rect 17880 12345 17908 13330
rect 17866 12336 17922 12345
rect 17972 12306 18000 15506
rect 18510 15464 18566 15473
rect 18510 15399 18566 15408
rect 19892 15428 19944 15434
rect 18524 15366 18552 15399
rect 19892 15370 19944 15376
rect 18512 15360 18564 15366
rect 18512 15302 18564 15308
rect 18234 15192 18290 15201
rect 18234 15127 18290 15136
rect 18248 14414 18276 15127
rect 18524 14482 18552 15302
rect 18512 14476 18564 14482
rect 18512 14418 18564 14424
rect 18236 14408 18288 14414
rect 18236 14350 18288 14356
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19432 14068 19484 14074
rect 19432 14010 19484 14016
rect 19064 13932 19116 13938
rect 19064 13874 19116 13880
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 18064 12306 18092 13262
rect 18510 13016 18566 13025
rect 18510 12951 18566 12960
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18144 12708 18196 12714
rect 18144 12650 18196 12656
rect 17866 12271 17922 12280
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18052 12300 18104 12306
rect 18052 12242 18104 12248
rect 18052 12164 18104 12170
rect 18052 12106 18104 12112
rect 17960 11688 18012 11694
rect 17684 11630 17736 11636
rect 17774 11656 17830 11665
rect 17696 11257 17724 11630
rect 17960 11630 18012 11636
rect 17774 11591 17830 11600
rect 17972 11393 18000 11630
rect 17958 11384 18014 11393
rect 17958 11319 18014 11328
rect 17682 11248 17738 11257
rect 17682 11183 17738 11192
rect 17604 11104 17908 11132
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17592 10736 17644 10742
rect 17592 10678 17644 10684
rect 17500 10532 17552 10538
rect 17500 10474 17552 10480
rect 17512 10169 17540 10474
rect 17498 10160 17554 10169
rect 17498 10095 17554 10104
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17512 9722 17540 9930
rect 17500 9716 17552 9722
rect 17500 9658 17552 9664
rect 17500 7880 17552 7886
rect 17500 7822 17552 7828
rect 17604 7834 17632 10678
rect 17696 10538 17724 10950
rect 17684 10532 17736 10538
rect 17684 10474 17736 10480
rect 17696 9450 17724 10474
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17788 9722 17816 9862
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17880 9602 17908 11104
rect 17960 11008 18012 11014
rect 17960 10950 18012 10956
rect 17972 10606 18000 10950
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 17972 10130 18000 10542
rect 17960 10124 18012 10130
rect 17960 10066 18012 10072
rect 17958 9888 18014 9897
rect 17958 9823 18014 9832
rect 17788 9574 17908 9602
rect 17684 9444 17736 9450
rect 17684 9386 17736 9392
rect 17512 7342 17540 7822
rect 17604 7806 17724 7834
rect 17592 7744 17644 7750
rect 17592 7686 17644 7692
rect 17604 7546 17632 7686
rect 17592 7540 17644 7546
rect 17592 7482 17644 7488
rect 17500 7336 17552 7342
rect 17500 7278 17552 7284
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17408 5704 17460 5710
rect 17408 5646 17460 5652
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17316 4140 17368 4146
rect 17316 4082 17368 4088
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17236 3670 17264 4014
rect 17420 3738 17448 4422
rect 17408 3732 17460 3738
rect 17408 3674 17460 3680
rect 17224 3664 17276 3670
rect 17224 3606 17276 3612
rect 17132 3528 17184 3534
rect 17224 3528 17276 3534
rect 17132 3470 17184 3476
rect 17222 3496 17224 3505
rect 17276 3496 17278 3505
rect 17222 3431 17278 3440
rect 17040 3120 17092 3126
rect 17040 3062 17092 3068
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 17316 2304 17368 2310
rect 17316 2246 17368 2252
rect 17328 1601 17356 2246
rect 17420 1902 17448 2382
rect 17408 1896 17460 1902
rect 17408 1838 17460 1844
rect 17512 1737 17540 6598
rect 17696 6202 17724 7806
rect 17788 6866 17816 9574
rect 17868 9444 17920 9450
rect 17868 9386 17920 9392
rect 17880 8362 17908 9386
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 17972 7886 18000 9823
rect 18064 8922 18092 12106
rect 18156 10810 18184 12650
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18144 10668 18196 10674
rect 18144 10610 18196 10616
rect 18156 9178 18184 10610
rect 18248 10062 18276 12718
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11762 18368 12038
rect 18328 11756 18380 11762
rect 18328 11698 18380 11704
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18340 9994 18368 11698
rect 18432 10198 18460 12242
rect 18524 10538 18552 12951
rect 18616 11801 18644 13806
rect 18972 12436 19024 12442
rect 18972 12378 19024 12384
rect 18880 12368 18932 12374
rect 18880 12310 18932 12316
rect 18602 11792 18658 11801
rect 18602 11727 18658 11736
rect 18512 10532 18564 10538
rect 18512 10474 18564 10480
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18510 10024 18566 10033
rect 18328 9988 18380 9994
rect 18510 9959 18566 9968
rect 18328 9930 18380 9936
rect 18236 9648 18288 9654
rect 18236 9590 18288 9596
rect 18248 9353 18276 9590
rect 18234 9344 18290 9353
rect 18234 9279 18290 9288
rect 18340 9194 18368 9930
rect 18420 9920 18472 9926
rect 18420 9862 18472 9868
rect 18432 9353 18460 9862
rect 18524 9761 18552 9959
rect 18510 9752 18566 9761
rect 18510 9687 18566 9696
rect 18418 9344 18474 9353
rect 18418 9279 18474 9288
rect 18144 9172 18196 9178
rect 18340 9166 18460 9194
rect 18196 9132 18276 9160
rect 18144 9114 18196 9120
rect 18064 8894 18184 8922
rect 18052 8832 18104 8838
rect 18052 8774 18104 8780
rect 18064 8537 18092 8774
rect 18050 8528 18106 8537
rect 18050 8463 18106 8472
rect 18050 8392 18106 8401
rect 18050 8327 18106 8336
rect 17960 7880 18012 7886
rect 17960 7822 18012 7828
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17972 7449 18000 7686
rect 17958 7440 18014 7449
rect 17868 7404 17920 7410
rect 17958 7375 17960 7384
rect 17868 7346 17920 7352
rect 18012 7375 18014 7384
rect 17960 7346 18012 7352
rect 17880 7002 17908 7346
rect 17972 7315 18000 7346
rect 18064 7256 18092 8327
rect 17972 7228 18092 7256
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17776 6860 17828 6866
rect 17776 6802 17828 6808
rect 17776 6384 17828 6390
rect 17776 6326 17828 6332
rect 17604 6174 17724 6202
rect 17604 5642 17632 6174
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17696 5778 17724 6054
rect 17684 5772 17736 5778
rect 17684 5714 17736 5720
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17696 5302 17724 5714
rect 17684 5296 17736 5302
rect 17684 5238 17736 5244
rect 17592 5160 17644 5166
rect 17592 5102 17644 5108
rect 17604 4282 17632 5102
rect 17592 4276 17644 4282
rect 17592 4218 17644 4224
rect 17788 4078 17816 6326
rect 17972 4826 18000 7228
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17868 4480 17920 4486
rect 17868 4422 17920 4428
rect 17776 4072 17828 4078
rect 17590 4040 17646 4049
rect 17776 4014 17828 4020
rect 17590 3975 17646 3984
rect 17604 3398 17632 3975
rect 17684 3936 17736 3942
rect 17684 3878 17736 3884
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17696 2774 17724 3878
rect 17788 3602 17816 4014
rect 17880 3738 17908 4422
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17788 2990 17816 3538
rect 17972 3194 18000 4490
rect 18064 4282 18092 5510
rect 18052 4276 18104 4282
rect 18052 4218 18104 4224
rect 18064 3534 18092 4218
rect 18156 3942 18184 8894
rect 18248 8498 18276 9132
rect 18328 8968 18380 8974
rect 18328 8910 18380 8916
rect 18340 8634 18368 8910
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18326 8120 18382 8129
rect 18326 8055 18382 8064
rect 18236 7200 18288 7206
rect 18236 7142 18288 7148
rect 18248 5234 18276 7142
rect 18340 6458 18368 8055
rect 18328 6452 18380 6458
rect 18328 6394 18380 6400
rect 18432 6338 18460 9166
rect 18524 8974 18552 9687
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18616 8566 18644 11727
rect 18694 11520 18750 11529
rect 18694 11455 18750 11464
rect 18708 9042 18736 11455
rect 18788 10668 18840 10674
rect 18788 10610 18840 10616
rect 18696 9036 18748 9042
rect 18696 8978 18748 8984
rect 18694 8936 18750 8945
rect 18694 8871 18750 8880
rect 18604 8560 18656 8566
rect 18604 8502 18656 8508
rect 18510 7848 18566 7857
rect 18510 7783 18566 7792
rect 18340 6310 18460 6338
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18236 5024 18288 5030
rect 18236 4966 18288 4972
rect 18248 4146 18276 4966
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18144 3936 18196 3942
rect 18144 3878 18196 3884
rect 18052 3528 18104 3534
rect 18052 3470 18104 3476
rect 18340 3466 18368 6310
rect 18420 5568 18472 5574
rect 18420 5510 18472 5516
rect 18432 4729 18460 5510
rect 18524 4826 18552 7783
rect 18602 7440 18658 7449
rect 18602 7375 18658 7384
rect 18512 4820 18564 4826
rect 18512 4762 18564 4768
rect 18418 4720 18474 4729
rect 18418 4655 18474 4664
rect 18420 4548 18472 4554
rect 18420 4490 18472 4496
rect 18328 3460 18380 3466
rect 18328 3402 18380 3408
rect 17960 3188 18012 3194
rect 17960 3130 18012 3136
rect 18328 3188 18380 3194
rect 18328 3130 18380 3136
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17972 2854 18000 2926
rect 17960 2848 18012 2854
rect 17960 2790 18012 2796
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17604 2746 17724 2774
rect 17498 1728 17554 1737
rect 17498 1663 17554 1672
rect 17314 1592 17370 1601
rect 17314 1527 17370 1536
rect 16946 912 17002 921
rect 16946 847 17002 856
rect 17604 800 17632 2746
rect 18052 2576 18104 2582
rect 18050 2544 18052 2553
rect 18104 2544 18106 2553
rect 18050 2479 18106 2488
rect 17960 2440 18012 2446
rect 18248 2417 18276 2790
rect 17960 2382 18012 2388
rect 18234 2408 18290 2417
rect 17972 1873 18000 2382
rect 18234 2343 18290 2352
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 17958 1864 18014 1873
rect 17958 1799 18014 1808
rect 18156 1766 18184 2246
rect 18340 2145 18368 3130
rect 18432 3126 18460 4490
rect 18616 4010 18644 7375
rect 18708 5370 18736 8871
rect 18800 7750 18828 10610
rect 18788 7744 18840 7750
rect 18788 7686 18840 7692
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18800 5250 18828 7686
rect 18708 5222 18828 5250
rect 18708 4214 18736 5222
rect 18696 4208 18748 4214
rect 18696 4150 18748 4156
rect 18604 4004 18656 4010
rect 18604 3946 18656 3952
rect 18420 3120 18472 3126
rect 18420 3062 18472 3068
rect 18512 2984 18564 2990
rect 18512 2926 18564 2932
rect 18326 2136 18382 2145
rect 18326 2071 18382 2080
rect 18144 1760 18196 1766
rect 18144 1702 18196 1708
rect 18524 800 18552 2926
rect 18708 1970 18736 4150
rect 18892 3641 18920 12310
rect 18984 9586 19012 12378
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18984 6798 19012 9522
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18972 6384 19024 6390
rect 18972 6326 19024 6332
rect 18984 3738 19012 6326
rect 19076 5710 19104 13874
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19064 5704 19116 5710
rect 19064 5646 19116 5652
rect 18972 3732 19024 3738
rect 18972 3674 19024 3680
rect 19168 3670 19196 13126
rect 19248 11824 19300 11830
rect 19248 11766 19300 11772
rect 19156 3664 19208 3670
rect 18878 3632 18934 3641
rect 19156 3606 19208 3612
rect 18878 3567 18934 3576
rect 19260 2774 19288 11766
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19352 3194 19380 8978
rect 19444 7886 19472 14010
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19536 4078 19564 9590
rect 19628 6186 19656 14350
rect 19708 10532 19760 10538
rect 19708 10474 19760 10480
rect 19720 6322 19748 10474
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19616 6180 19668 6186
rect 19616 6122 19668 6128
rect 19628 4554 19656 6122
rect 19616 4548 19668 4554
rect 19616 4490 19668 4496
rect 19524 4072 19576 4078
rect 19524 4014 19576 4020
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19904 3058 19932 15370
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19432 2916 19484 2922
rect 19432 2858 19484 2864
rect 18800 2746 19288 2774
rect 18800 2417 18828 2746
rect 18786 2408 18842 2417
rect 18786 2343 18842 2352
rect 18696 1964 18748 1970
rect 18696 1906 18748 1912
rect 19444 800 19472 2858
rect 15842 504 15898 513
rect 15842 439 15898 448
rect 16670 0 16726 800
rect 17590 0 17646 800
rect 18510 0 18566 800
rect 19430 0 19486 800
<< via2 >>
rect 3790 16904 3846 16960
rect 2134 15952 2190 16008
rect 1490 14864 1546 14920
rect 1122 12960 1178 13016
rect 938 12552 994 12608
rect 846 7894 902 7950
rect 1030 12416 1086 12472
rect 1122 7384 1178 7440
rect 938 6704 994 6760
rect 1122 6160 1178 6216
rect 1122 4664 1178 4720
rect 1030 3304 1086 3360
rect 1950 14476 2006 14512
rect 1950 14456 1952 14476
rect 1952 14456 2004 14476
rect 2004 14456 2006 14476
rect 2226 14184 2282 14240
rect 1858 13368 1914 13424
rect 1674 12144 1730 12200
rect 1490 9968 1546 10024
rect 1306 9424 1362 9480
rect 1398 8744 1454 8800
rect 2410 13912 2466 13968
rect 2410 13232 2466 13288
rect 2134 11736 2190 11792
rect 1950 11192 2006 11248
rect 1950 9968 2006 10024
rect 1950 9580 2006 9616
rect 1950 9560 1952 9580
rect 1952 9560 2004 9580
rect 2004 9560 2006 9580
rect 1858 9288 1914 9344
rect 1674 9036 1730 9072
rect 1674 9016 1676 9036
rect 1676 9016 1728 9036
rect 1728 9016 1730 9036
rect 1858 8744 1914 8800
rect 1674 5636 1730 5672
rect 1674 5616 1676 5636
rect 1676 5616 1728 5636
rect 1728 5616 1730 5636
rect 1766 5344 1822 5400
rect 1490 5072 1546 5128
rect 1398 4528 1454 4584
rect 1398 2896 1454 2952
rect 2226 10648 2282 10704
rect 2226 10512 2282 10568
rect 2226 9696 2282 9752
rect 1950 6704 2006 6760
rect 2226 8472 2282 8528
rect 4066 16632 4122 16688
rect 3882 15272 3938 15328
rect 2778 15000 2834 15056
rect 3180 14714 3236 14716
rect 3260 14714 3316 14716
rect 3340 14714 3396 14716
rect 3420 14714 3476 14716
rect 3180 14662 3226 14714
rect 3226 14662 3236 14714
rect 3260 14662 3290 14714
rect 3290 14662 3302 14714
rect 3302 14662 3316 14714
rect 3340 14662 3354 14714
rect 3354 14662 3366 14714
rect 3366 14662 3396 14714
rect 3420 14662 3430 14714
rect 3430 14662 3476 14714
rect 3180 14660 3236 14662
rect 3260 14660 3316 14662
rect 3340 14660 3396 14662
rect 3420 14660 3476 14662
rect 2962 14612 3018 14648
rect 2962 14592 2964 14612
rect 2964 14592 3016 14612
rect 3016 14592 3018 14612
rect 4342 16224 4398 16280
rect 2778 14320 2834 14376
rect 3054 14048 3110 14104
rect 3238 13932 3294 13968
rect 4618 15544 4674 15600
rect 4986 15000 5042 15056
rect 3238 13912 3240 13932
rect 3240 13912 3292 13932
rect 3292 13912 3294 13932
rect 4066 13776 4122 13832
rect 3180 13626 3236 13628
rect 3260 13626 3316 13628
rect 3340 13626 3396 13628
rect 3420 13626 3476 13628
rect 3180 13574 3226 13626
rect 3226 13574 3236 13626
rect 3260 13574 3290 13626
rect 3290 13574 3302 13626
rect 3302 13574 3316 13626
rect 3340 13574 3354 13626
rect 3354 13574 3366 13626
rect 3366 13574 3396 13626
rect 3420 13574 3430 13626
rect 3430 13574 3476 13626
rect 3180 13572 3236 13574
rect 3260 13572 3316 13574
rect 3340 13572 3396 13574
rect 3420 13572 3476 13574
rect 3606 13504 3662 13560
rect 3790 13368 3846 13424
rect 4066 13368 4122 13424
rect 3422 13268 3424 13288
rect 3424 13268 3476 13288
rect 3476 13268 3478 13288
rect 3422 13232 3478 13268
rect 3238 12960 3294 13016
rect 2778 12824 2834 12880
rect 3054 12844 3110 12880
rect 3054 12824 3056 12844
rect 3056 12824 3108 12844
rect 3108 12824 3110 12844
rect 2870 12688 2926 12744
rect 2962 12416 3018 12472
rect 2502 12280 2558 12336
rect 2778 12008 2834 12064
rect 2870 11600 2926 11656
rect 3180 12538 3236 12540
rect 3260 12538 3316 12540
rect 3340 12538 3396 12540
rect 3420 12538 3476 12540
rect 3180 12486 3226 12538
rect 3226 12486 3236 12538
rect 3260 12486 3290 12538
rect 3290 12486 3302 12538
rect 3302 12486 3316 12538
rect 3340 12486 3354 12538
rect 3354 12486 3366 12538
rect 3366 12486 3396 12538
rect 3420 12486 3430 12538
rect 3430 12486 3476 12538
rect 3180 12484 3236 12486
rect 3260 12484 3316 12486
rect 3340 12484 3396 12486
rect 3420 12484 3476 12486
rect 3422 12300 3478 12336
rect 3422 12280 3424 12300
rect 3424 12280 3476 12300
rect 3476 12280 3478 12300
rect 2962 11328 3018 11384
rect 2962 10920 3018 10976
rect 3180 11450 3236 11452
rect 3260 11450 3316 11452
rect 3340 11450 3396 11452
rect 3420 11450 3476 11452
rect 3180 11398 3226 11450
rect 3226 11398 3236 11450
rect 3260 11398 3290 11450
rect 3290 11398 3302 11450
rect 3302 11398 3316 11450
rect 3340 11398 3354 11450
rect 3354 11398 3366 11450
rect 3366 11398 3396 11450
rect 3420 11398 3430 11450
rect 3430 11398 3476 11450
rect 3180 11396 3236 11398
rect 3260 11396 3316 11398
rect 3340 11396 3396 11398
rect 3420 11396 3476 11398
rect 2778 10412 2780 10432
rect 2780 10412 2832 10432
rect 2832 10412 2834 10432
rect 2778 10376 2834 10412
rect 2502 8880 2558 8936
rect 2594 8200 2650 8256
rect 2778 8200 2834 8256
rect 3180 10362 3236 10364
rect 3260 10362 3316 10364
rect 3340 10362 3396 10364
rect 3420 10362 3476 10364
rect 3180 10310 3226 10362
rect 3226 10310 3236 10362
rect 3260 10310 3290 10362
rect 3290 10310 3302 10362
rect 3302 10310 3316 10362
rect 3340 10310 3354 10362
rect 3354 10310 3366 10362
rect 3366 10310 3396 10362
rect 3420 10310 3430 10362
rect 3430 10310 3476 10362
rect 3180 10308 3236 10310
rect 3260 10308 3316 10310
rect 3340 10308 3396 10310
rect 3420 10308 3476 10310
rect 2962 8472 3018 8528
rect 3790 12824 3846 12880
rect 3606 12552 3662 12608
rect 3790 12552 3846 12608
rect 3790 12416 3846 12472
rect 3606 10376 3662 10432
rect 3606 10240 3662 10296
rect 3790 10648 3846 10704
rect 4342 13096 4398 13152
rect 4250 12960 4306 13016
rect 4250 12844 4306 12880
rect 4250 12824 4252 12844
rect 4252 12824 4304 12844
rect 4304 12824 4306 12844
rect 3974 12044 3976 12064
rect 3976 12044 4028 12064
rect 4028 12044 4030 12064
rect 3974 12008 4030 12044
rect 3180 9274 3236 9276
rect 3260 9274 3316 9276
rect 3340 9274 3396 9276
rect 3420 9274 3476 9276
rect 3180 9222 3226 9274
rect 3226 9222 3236 9274
rect 3260 9222 3290 9274
rect 3290 9222 3302 9274
rect 3302 9222 3316 9274
rect 3340 9222 3354 9274
rect 3354 9222 3366 9274
rect 3366 9222 3396 9274
rect 3420 9222 3430 9274
rect 3430 9222 3476 9274
rect 3180 9220 3236 9222
rect 3260 9220 3316 9222
rect 3340 9220 3396 9222
rect 3420 9220 3476 9222
rect 3146 8880 3202 8936
rect 3238 8508 3240 8528
rect 3240 8508 3292 8528
rect 3292 8508 3294 8528
rect 3238 8472 3294 8508
rect 3882 9696 3938 9752
rect 3698 9016 3754 9072
rect 3698 8880 3754 8936
rect 4342 11872 4398 11928
rect 4250 11056 4306 11112
rect 4066 10784 4122 10840
rect 4710 13776 4766 13832
rect 5078 14184 5134 14240
rect 4986 14068 5042 14104
rect 4986 14048 4988 14068
rect 4988 14048 5040 14068
rect 5040 14048 5042 14068
rect 4894 13640 4950 13696
rect 4710 12960 4766 13016
rect 4158 9968 4214 10024
rect 3974 9016 4030 9072
rect 3180 8186 3236 8188
rect 3260 8186 3316 8188
rect 3340 8186 3396 8188
rect 3420 8186 3476 8188
rect 3180 8134 3226 8186
rect 3226 8134 3236 8186
rect 3260 8134 3290 8186
rect 3290 8134 3302 8186
rect 3302 8134 3316 8186
rect 3340 8134 3354 8186
rect 3354 8134 3366 8186
rect 3366 8134 3396 8186
rect 3420 8134 3430 8186
rect 3430 8134 3476 8186
rect 3180 8132 3236 8134
rect 3260 8132 3316 8134
rect 3340 8132 3396 8134
rect 3420 8132 3476 8134
rect 3974 8336 4030 8392
rect 3882 8254 3884 8256
rect 3884 8254 3936 8256
rect 3936 8254 3938 8256
rect 3606 8064 3662 8120
rect 3882 8200 3938 8254
rect 3238 7948 3294 7984
rect 3238 7928 3240 7948
rect 3240 7928 3292 7948
rect 3292 7928 3294 7948
rect 1950 5208 2006 5264
rect 2042 3576 2098 3632
rect 1766 2896 1822 2952
rect 1766 2624 1822 2680
rect 1490 176 1546 232
rect 2686 7520 2742 7576
rect 3330 7792 3386 7848
rect 2778 6976 2834 7032
rect 2686 5480 2742 5536
rect 2410 4800 2466 4856
rect 2318 4684 2374 4720
rect 2318 4664 2320 4684
rect 2320 4664 2372 4684
rect 2372 4664 2374 4684
rect 2502 4664 2558 4720
rect 2962 6024 3018 6080
rect 2962 5888 3018 5944
rect 3606 7656 3662 7712
rect 3180 7098 3236 7100
rect 3260 7098 3316 7100
rect 3340 7098 3396 7100
rect 3420 7098 3476 7100
rect 3180 7046 3226 7098
rect 3226 7046 3236 7098
rect 3260 7046 3290 7098
rect 3290 7046 3302 7098
rect 3302 7046 3316 7098
rect 3340 7046 3354 7098
rect 3354 7046 3366 7098
rect 3366 7046 3396 7098
rect 3420 7046 3430 7098
rect 3430 7046 3476 7098
rect 3180 7044 3236 7046
rect 3260 7044 3316 7046
rect 3340 7044 3396 7046
rect 3420 7044 3476 7046
rect 3422 6860 3478 6896
rect 3422 6840 3424 6860
rect 3424 6840 3476 6860
rect 3476 6840 3478 6860
rect 3146 6316 3202 6352
rect 3146 6296 3148 6316
rect 3148 6296 3200 6316
rect 3200 6296 3202 6316
rect 3180 6010 3236 6012
rect 3260 6010 3316 6012
rect 3340 6010 3396 6012
rect 3420 6010 3476 6012
rect 3180 5958 3226 6010
rect 3226 5958 3236 6010
rect 3260 5958 3290 6010
rect 3290 5958 3302 6010
rect 3302 5958 3316 6010
rect 3340 5958 3354 6010
rect 3354 5958 3366 6010
rect 3366 5958 3396 6010
rect 3420 5958 3430 6010
rect 3430 5958 3476 6010
rect 3180 5956 3236 5958
rect 3260 5956 3316 5958
rect 3340 5956 3396 5958
rect 3420 5956 3476 5958
rect 2962 5072 3018 5128
rect 3180 4922 3236 4924
rect 3260 4922 3316 4924
rect 3340 4922 3396 4924
rect 3420 4922 3476 4924
rect 3180 4870 3226 4922
rect 3226 4870 3236 4922
rect 3260 4870 3290 4922
rect 3290 4870 3302 4922
rect 3302 4870 3316 4922
rect 3340 4870 3354 4922
rect 3354 4870 3366 4922
rect 3366 4870 3396 4922
rect 3420 4870 3430 4922
rect 3430 4870 3476 4922
rect 3180 4868 3236 4870
rect 3260 4868 3316 4870
rect 3340 4868 3396 4870
rect 3420 4868 3476 4870
rect 3422 4684 3478 4720
rect 3422 4664 3424 4684
rect 3424 4664 3476 4684
rect 3476 4664 3478 4684
rect 2962 2760 3018 2816
rect 3238 4256 3294 4312
rect 3180 3834 3236 3836
rect 3260 3834 3316 3836
rect 3340 3834 3396 3836
rect 3420 3834 3476 3836
rect 3180 3782 3226 3834
rect 3226 3782 3236 3834
rect 3260 3782 3290 3834
rect 3290 3782 3302 3834
rect 3302 3782 3316 3834
rect 3340 3782 3354 3834
rect 3354 3782 3366 3834
rect 3366 3782 3396 3834
rect 3420 3782 3430 3834
rect 3430 3782 3476 3834
rect 3180 3780 3236 3782
rect 3260 3780 3316 3782
rect 3340 3780 3396 3782
rect 3420 3780 3476 3782
rect 3698 7248 3754 7304
rect 4158 8200 4214 8256
rect 4526 8780 4528 8800
rect 4528 8780 4580 8800
rect 4580 8780 4582 8800
rect 4526 8744 4582 8780
rect 4250 8064 4306 8120
rect 4066 7656 4122 7712
rect 4342 7656 4398 7712
rect 3790 7112 3846 7168
rect 3790 6568 3846 6624
rect 3790 3984 3846 4040
rect 3514 3440 3570 3496
rect 3180 2746 3236 2748
rect 3260 2746 3316 2748
rect 3340 2746 3396 2748
rect 3420 2746 3476 2748
rect 3180 2694 3226 2746
rect 3226 2694 3236 2746
rect 3260 2694 3290 2746
rect 3290 2694 3302 2746
rect 3302 2694 3316 2746
rect 3340 2694 3354 2746
rect 3354 2694 3366 2746
rect 3366 2694 3396 2746
rect 3420 2694 3430 2746
rect 3430 2694 3476 2746
rect 3180 2692 3236 2694
rect 3260 2692 3316 2694
rect 3340 2692 3396 2694
rect 3420 2692 3476 2694
rect 3422 1944 3478 2000
rect 3698 3032 3754 3088
rect 4526 7812 4582 7848
rect 4526 7792 4528 7812
rect 4528 7792 4580 7812
rect 4580 7792 4582 7812
rect 4618 7520 4674 7576
rect 4618 7284 4620 7304
rect 4620 7284 4672 7304
rect 4672 7284 4674 7304
rect 4618 7248 4674 7284
rect 4618 6976 4674 7032
rect 4618 6876 4620 6896
rect 4620 6876 4672 6896
rect 4672 6876 4674 6896
rect 4618 6840 4674 6876
rect 4434 6432 4490 6488
rect 4342 6160 4398 6216
rect 4250 4528 4306 4584
rect 4066 4392 4122 4448
rect 4250 3712 4306 3768
rect 3790 2760 3846 2816
rect 3882 2644 3938 2680
rect 3882 2624 3884 2644
rect 3884 2624 3936 2644
rect 3936 2624 3938 2644
rect 4894 12824 4950 12880
rect 5722 14864 5778 14920
rect 5354 14592 5410 14648
rect 5722 14320 5778 14376
rect 5404 14170 5460 14172
rect 5484 14170 5540 14172
rect 5564 14170 5620 14172
rect 5644 14170 5700 14172
rect 5404 14118 5450 14170
rect 5450 14118 5460 14170
rect 5484 14118 5514 14170
rect 5514 14118 5526 14170
rect 5526 14118 5540 14170
rect 5564 14118 5578 14170
rect 5578 14118 5590 14170
rect 5590 14118 5620 14170
rect 5644 14118 5654 14170
rect 5654 14118 5700 14170
rect 5404 14116 5460 14118
rect 5484 14116 5540 14118
rect 5564 14116 5620 14118
rect 5644 14116 5700 14118
rect 5814 14068 5870 14104
rect 5814 14048 5816 14068
rect 5816 14048 5868 14068
rect 5868 14048 5870 14068
rect 5262 13640 5318 13696
rect 5446 13640 5502 13696
rect 5354 13368 5410 13424
rect 5170 12708 5226 12744
rect 5170 12688 5172 12708
rect 5172 12688 5224 12708
rect 5224 12688 5226 12708
rect 5404 13082 5460 13084
rect 5484 13082 5540 13084
rect 5564 13082 5620 13084
rect 5644 13082 5700 13084
rect 5404 13030 5450 13082
rect 5450 13030 5460 13082
rect 5484 13030 5514 13082
rect 5514 13030 5526 13082
rect 5526 13030 5540 13082
rect 5564 13030 5578 13082
rect 5578 13030 5590 13082
rect 5590 13030 5620 13082
rect 5644 13030 5654 13082
rect 5654 13030 5700 13082
rect 5404 13028 5460 13030
rect 5484 13028 5540 13030
rect 5564 13028 5620 13030
rect 5644 13028 5700 13030
rect 6274 14320 6330 14376
rect 6090 13368 6146 13424
rect 6182 12824 6238 12880
rect 7102 14592 7158 14648
rect 6826 14184 6882 14240
rect 6918 13948 6920 13968
rect 6920 13948 6972 13968
rect 6972 13948 6974 13968
rect 6918 13912 6974 13948
rect 6550 13252 6606 13288
rect 6550 13232 6552 13252
rect 6552 13232 6604 13252
rect 6604 13232 6606 13252
rect 6090 12688 6146 12744
rect 5630 12280 5686 12336
rect 5998 12552 6054 12608
rect 6182 12552 6238 12608
rect 6182 12416 6238 12472
rect 5354 12144 5410 12200
rect 5078 11600 5134 11656
rect 4986 10920 5042 10976
rect 5078 9324 5080 9344
rect 5080 9324 5132 9344
rect 5132 9324 5134 9344
rect 5078 9288 5134 9324
rect 5078 6704 5134 6760
rect 4710 5480 4766 5536
rect 4434 4528 4490 4584
rect 4986 6160 5042 6216
rect 4894 6024 4950 6080
rect 5998 12164 6054 12200
rect 5998 12144 6000 12164
rect 6000 12144 6052 12164
rect 6052 12144 6054 12164
rect 5404 11994 5460 11996
rect 5484 11994 5540 11996
rect 5564 11994 5620 11996
rect 5644 11994 5700 11996
rect 5404 11942 5450 11994
rect 5450 11942 5460 11994
rect 5484 11942 5514 11994
rect 5514 11942 5526 11994
rect 5526 11942 5540 11994
rect 5564 11942 5578 11994
rect 5578 11942 5590 11994
rect 5590 11942 5620 11994
rect 5644 11942 5654 11994
rect 5654 11942 5700 11994
rect 5404 11940 5460 11942
rect 5484 11940 5540 11942
rect 5564 11940 5620 11942
rect 5644 11940 5700 11942
rect 5354 11464 5410 11520
rect 5722 11328 5778 11384
rect 5404 10906 5460 10908
rect 5484 10906 5540 10908
rect 5564 10906 5620 10908
rect 5644 10906 5700 10908
rect 5404 10854 5450 10906
rect 5450 10854 5460 10906
rect 5484 10854 5514 10906
rect 5514 10854 5526 10906
rect 5526 10854 5540 10906
rect 5564 10854 5578 10906
rect 5578 10854 5590 10906
rect 5590 10854 5620 10906
rect 5644 10854 5654 10906
rect 5654 10854 5700 10906
rect 5404 10852 5460 10854
rect 5484 10852 5540 10854
rect 5564 10852 5620 10854
rect 5644 10852 5700 10854
rect 5404 9818 5460 9820
rect 5484 9818 5540 9820
rect 5564 9818 5620 9820
rect 5644 9818 5700 9820
rect 5404 9766 5450 9818
rect 5450 9766 5460 9818
rect 5484 9766 5514 9818
rect 5514 9766 5526 9818
rect 5526 9766 5540 9818
rect 5564 9766 5578 9818
rect 5578 9766 5590 9818
rect 5590 9766 5620 9818
rect 5644 9766 5654 9818
rect 5654 9766 5700 9818
rect 5404 9764 5460 9766
rect 5484 9764 5540 9766
rect 5564 9764 5620 9766
rect 5644 9764 5700 9766
rect 5906 12008 5962 12064
rect 5906 11772 5908 11792
rect 5908 11772 5960 11792
rect 5960 11772 5962 11792
rect 5906 11736 5962 11772
rect 5906 10784 5962 10840
rect 5404 8730 5460 8732
rect 5484 8730 5540 8732
rect 5564 8730 5620 8732
rect 5644 8730 5700 8732
rect 5404 8678 5450 8730
rect 5450 8678 5460 8730
rect 5484 8678 5514 8730
rect 5514 8678 5526 8730
rect 5526 8678 5540 8730
rect 5564 8678 5578 8730
rect 5578 8678 5590 8730
rect 5590 8678 5620 8730
rect 5644 8678 5654 8730
rect 5654 8678 5700 8730
rect 5404 8676 5460 8678
rect 5484 8676 5540 8678
rect 5564 8676 5620 8678
rect 5644 8676 5700 8678
rect 5262 8608 5318 8664
rect 5262 8336 5318 8392
rect 5262 7792 5318 7848
rect 5404 7642 5460 7644
rect 5484 7642 5540 7644
rect 5564 7642 5620 7644
rect 5644 7642 5700 7644
rect 5404 7590 5450 7642
rect 5450 7590 5460 7642
rect 5484 7590 5514 7642
rect 5514 7590 5526 7642
rect 5526 7590 5540 7642
rect 5564 7590 5578 7642
rect 5578 7590 5590 7642
rect 5590 7590 5620 7642
rect 5644 7590 5654 7642
rect 5654 7590 5700 7642
rect 5404 7588 5460 7590
rect 5484 7588 5540 7590
rect 5564 7588 5620 7590
rect 5644 7588 5700 7590
rect 5446 7112 5502 7168
rect 5630 7112 5686 7168
rect 5262 6976 5318 7032
rect 5404 6554 5460 6556
rect 5484 6554 5540 6556
rect 5564 6554 5620 6556
rect 5644 6554 5700 6556
rect 5404 6502 5450 6554
rect 5450 6502 5460 6554
rect 5484 6502 5514 6554
rect 5514 6502 5526 6554
rect 5526 6502 5540 6554
rect 5564 6502 5578 6554
rect 5578 6502 5590 6554
rect 5590 6502 5620 6554
rect 5644 6502 5654 6554
rect 5654 6502 5700 6554
rect 5404 6500 5460 6502
rect 5484 6500 5540 6502
rect 5564 6500 5620 6502
rect 5644 6500 5700 6502
rect 5078 5616 5134 5672
rect 4710 3848 4766 3904
rect 4342 2624 4398 2680
rect 5170 4664 5226 4720
rect 5078 4120 5134 4176
rect 6090 11192 6146 11248
rect 5998 7520 6054 7576
rect 5404 5466 5460 5468
rect 5484 5466 5540 5468
rect 5564 5466 5620 5468
rect 5644 5466 5700 5468
rect 5404 5414 5450 5466
rect 5450 5414 5460 5466
rect 5484 5414 5514 5466
rect 5514 5414 5526 5466
rect 5526 5414 5540 5466
rect 5564 5414 5578 5466
rect 5578 5414 5590 5466
rect 5590 5414 5620 5466
rect 5644 5414 5654 5466
rect 5654 5414 5700 5466
rect 5404 5412 5460 5414
rect 5484 5412 5540 5414
rect 5564 5412 5620 5414
rect 5644 5412 5700 5414
rect 5814 5344 5870 5400
rect 6274 9560 6330 9616
rect 7628 14714 7684 14716
rect 7708 14714 7764 14716
rect 7788 14714 7844 14716
rect 7868 14714 7924 14716
rect 7628 14662 7674 14714
rect 7674 14662 7684 14714
rect 7708 14662 7738 14714
rect 7738 14662 7750 14714
rect 7750 14662 7764 14714
rect 7788 14662 7802 14714
rect 7802 14662 7814 14714
rect 7814 14662 7844 14714
rect 7868 14662 7878 14714
rect 7878 14662 7924 14714
rect 7628 14660 7684 14662
rect 7708 14660 7764 14662
rect 7788 14660 7844 14662
rect 7868 14660 7924 14662
rect 8298 14048 8354 14104
rect 7378 13640 7434 13696
rect 7628 13626 7684 13628
rect 7708 13626 7764 13628
rect 7788 13626 7844 13628
rect 7868 13626 7924 13628
rect 7628 13574 7674 13626
rect 7674 13574 7684 13626
rect 7708 13574 7738 13626
rect 7738 13574 7750 13626
rect 7750 13574 7764 13626
rect 7788 13574 7802 13626
rect 7802 13574 7814 13626
rect 7814 13574 7844 13626
rect 7868 13574 7878 13626
rect 7878 13574 7924 13626
rect 7628 13572 7684 13574
rect 7708 13572 7764 13574
rect 7788 13572 7844 13574
rect 7868 13572 7924 13574
rect 8114 13776 8170 13832
rect 7194 13388 7250 13424
rect 7194 13368 7196 13388
rect 7196 13368 7248 13388
rect 7248 13368 7250 13388
rect 7010 13232 7066 13288
rect 8114 13232 8170 13288
rect 7746 13132 7748 13152
rect 7748 13132 7800 13152
rect 7800 13132 7802 13152
rect 7010 12960 7066 13016
rect 6918 12552 6974 12608
rect 6826 12416 6882 12472
rect 7010 12416 7066 12472
rect 6550 12280 6606 12336
rect 6550 11056 6606 11112
rect 6642 10784 6698 10840
rect 6550 10240 6606 10296
rect 6458 9560 6514 9616
rect 7746 13096 7802 13132
rect 7628 12538 7684 12540
rect 7708 12538 7764 12540
rect 7788 12538 7844 12540
rect 7868 12538 7924 12540
rect 7628 12486 7674 12538
rect 7674 12486 7684 12538
rect 7708 12486 7738 12538
rect 7738 12486 7750 12538
rect 7750 12486 7764 12538
rect 7788 12486 7802 12538
rect 7802 12486 7814 12538
rect 7814 12486 7844 12538
rect 7868 12486 7878 12538
rect 7878 12486 7924 12538
rect 7628 12484 7684 12486
rect 7708 12484 7764 12486
rect 7788 12484 7844 12486
rect 7868 12484 7924 12486
rect 7378 12280 7434 12336
rect 7562 12280 7618 12336
rect 6918 10104 6974 10160
rect 6826 9832 6882 9888
rect 6274 6876 6276 6896
rect 6276 6876 6328 6896
rect 6328 6876 6330 6896
rect 6274 6840 6330 6876
rect 6918 9696 6974 9752
rect 6642 7656 6698 7712
rect 7286 12008 7342 12064
rect 7286 11736 7342 11792
rect 8758 15000 8814 15056
rect 8114 12552 8170 12608
rect 8114 11872 8170 11928
rect 8022 11772 8024 11792
rect 8024 11772 8076 11792
rect 8076 11772 8078 11792
rect 8022 11736 8078 11772
rect 7628 11450 7684 11452
rect 7708 11450 7764 11452
rect 7788 11450 7844 11452
rect 7868 11450 7924 11452
rect 7628 11398 7674 11450
rect 7674 11398 7684 11450
rect 7708 11398 7738 11450
rect 7738 11398 7750 11450
rect 7750 11398 7764 11450
rect 7788 11398 7802 11450
rect 7802 11398 7814 11450
rect 7814 11398 7844 11450
rect 7868 11398 7878 11450
rect 7878 11398 7924 11450
rect 7628 11396 7684 11398
rect 7708 11396 7764 11398
rect 7788 11396 7844 11398
rect 7868 11396 7924 11398
rect 7378 10376 7434 10432
rect 7286 10240 7342 10296
rect 7194 10104 7250 10160
rect 7628 10362 7684 10364
rect 7708 10362 7764 10364
rect 7788 10362 7844 10364
rect 7868 10362 7924 10364
rect 7628 10310 7674 10362
rect 7674 10310 7684 10362
rect 7708 10310 7738 10362
rect 7738 10310 7750 10362
rect 7750 10310 7764 10362
rect 7788 10310 7802 10362
rect 7802 10310 7814 10362
rect 7814 10310 7844 10362
rect 7868 10310 7878 10362
rect 7878 10310 7924 10362
rect 7628 10308 7684 10310
rect 7708 10308 7764 10310
rect 7788 10308 7844 10310
rect 7868 10308 7924 10310
rect 8114 10784 8170 10840
rect 7378 9424 7434 9480
rect 7654 9832 7710 9888
rect 7746 9696 7802 9752
rect 7930 9696 7986 9752
rect 7562 9424 7618 9480
rect 7286 8608 7342 8664
rect 6826 6296 6882 6352
rect 5998 5072 6054 5128
rect 5404 4378 5460 4380
rect 5484 4378 5540 4380
rect 5564 4378 5620 4380
rect 5644 4378 5700 4380
rect 5404 4326 5450 4378
rect 5450 4326 5460 4378
rect 5484 4326 5514 4378
rect 5514 4326 5526 4378
rect 5526 4326 5540 4378
rect 5564 4326 5578 4378
rect 5578 4326 5590 4378
rect 5590 4326 5620 4378
rect 5644 4326 5654 4378
rect 5654 4326 5700 4378
rect 5404 4324 5460 4326
rect 5484 4324 5540 4326
rect 5564 4324 5620 4326
rect 5644 4324 5700 4326
rect 5170 3984 5226 4040
rect 4894 2216 4950 2272
rect 4066 1808 4122 1864
rect 4066 1400 4122 1456
rect 4066 1128 4122 1184
rect 5262 3712 5318 3768
rect 5404 3290 5460 3292
rect 5484 3290 5540 3292
rect 5564 3290 5620 3292
rect 5644 3290 5700 3292
rect 5404 3238 5450 3290
rect 5450 3238 5460 3290
rect 5484 3238 5514 3290
rect 5514 3238 5526 3290
rect 5526 3238 5540 3290
rect 5564 3238 5578 3290
rect 5578 3238 5590 3290
rect 5590 3238 5620 3290
rect 5644 3238 5654 3290
rect 5654 3238 5700 3290
rect 5404 3236 5460 3238
rect 5484 3236 5540 3238
rect 5564 3236 5620 3238
rect 5644 3236 5700 3238
rect 5814 3168 5870 3224
rect 5404 2202 5460 2204
rect 5484 2202 5540 2204
rect 5564 2202 5620 2204
rect 5644 2202 5700 2204
rect 5404 2150 5450 2202
rect 5450 2150 5460 2202
rect 5484 2150 5514 2202
rect 5514 2150 5526 2202
rect 5526 2150 5540 2202
rect 5564 2150 5578 2202
rect 5578 2150 5590 2202
rect 5590 2150 5620 2202
rect 5644 2150 5654 2202
rect 5654 2150 5700 2202
rect 5404 2148 5460 2150
rect 5484 2148 5540 2150
rect 5564 2148 5620 2150
rect 5644 2148 5700 2150
rect 5262 2080 5318 2136
rect 5262 1672 5318 1728
rect 6458 5108 6460 5128
rect 6460 5108 6512 5128
rect 6512 5108 6514 5128
rect 6458 5072 6514 5108
rect 6182 4392 6238 4448
rect 6274 3440 6330 3496
rect 6182 2524 6184 2544
rect 6184 2524 6236 2544
rect 6236 2524 6238 2544
rect 6182 2488 6238 2524
rect 5814 1400 5870 1456
rect 3422 720 3478 776
rect 3698 448 3754 504
rect 6642 3304 6698 3360
rect 6826 3848 6882 3904
rect 6918 3440 6974 3496
rect 6734 3032 6790 3088
rect 6918 3032 6974 3088
rect 7470 9288 7526 9344
rect 7628 9274 7684 9276
rect 7708 9274 7764 9276
rect 7788 9274 7844 9276
rect 7868 9274 7924 9276
rect 7628 9222 7674 9274
rect 7674 9222 7684 9274
rect 7708 9222 7738 9274
rect 7738 9222 7750 9274
rect 7750 9222 7764 9274
rect 7788 9222 7802 9274
rect 7802 9222 7814 9274
rect 7814 9222 7844 9274
rect 7868 9222 7878 9274
rect 7878 9222 7924 9274
rect 7628 9220 7684 9222
rect 7708 9220 7764 9222
rect 7788 9220 7844 9222
rect 7868 9220 7924 9222
rect 7746 8880 7802 8936
rect 8114 8880 8170 8936
rect 7470 8744 7526 8800
rect 7562 8608 7618 8664
rect 8114 8744 8170 8800
rect 7470 8200 7526 8256
rect 7628 8186 7684 8188
rect 7708 8186 7764 8188
rect 7788 8186 7844 8188
rect 7868 8186 7924 8188
rect 7628 8134 7674 8186
rect 7674 8134 7684 8186
rect 7708 8134 7738 8186
rect 7738 8134 7750 8186
rect 7750 8134 7764 8186
rect 7788 8134 7802 8186
rect 7802 8134 7814 8186
rect 7814 8134 7844 8186
rect 7868 8134 7878 8186
rect 7878 8134 7924 8186
rect 7628 8132 7684 8134
rect 7708 8132 7764 8134
rect 7788 8132 7844 8134
rect 7868 8132 7924 8134
rect 7930 7520 7986 7576
rect 7628 7098 7684 7100
rect 7708 7098 7764 7100
rect 7788 7098 7844 7100
rect 7868 7098 7924 7100
rect 7628 7046 7674 7098
rect 7674 7046 7684 7098
rect 7708 7046 7738 7098
rect 7738 7046 7750 7098
rect 7750 7046 7764 7098
rect 7788 7046 7802 7098
rect 7802 7046 7814 7098
rect 7814 7046 7844 7098
rect 7868 7046 7878 7098
rect 7878 7046 7924 7098
rect 7628 7044 7684 7046
rect 7708 7044 7764 7046
rect 7788 7044 7844 7046
rect 7868 7044 7924 7046
rect 7562 6432 7618 6488
rect 9402 14592 9458 14648
rect 10230 14184 10286 14240
rect 9852 14170 9908 14172
rect 9932 14170 9988 14172
rect 10012 14170 10068 14172
rect 10092 14170 10148 14172
rect 9852 14118 9898 14170
rect 9898 14118 9908 14170
rect 9932 14118 9962 14170
rect 9962 14118 9974 14170
rect 9974 14118 9988 14170
rect 10012 14118 10026 14170
rect 10026 14118 10038 14170
rect 10038 14118 10068 14170
rect 10092 14118 10102 14170
rect 10102 14118 10148 14170
rect 9852 14116 9908 14118
rect 9932 14116 9988 14118
rect 10012 14116 10068 14118
rect 10092 14116 10148 14118
rect 9402 13640 9458 13696
rect 8850 12844 8906 12880
rect 8850 12824 8852 12844
rect 8852 12824 8904 12844
rect 8904 12824 8906 12844
rect 8390 10956 8392 10976
rect 8392 10956 8444 10976
rect 8444 10956 8446 10976
rect 8390 10920 8446 10956
rect 8390 10512 8446 10568
rect 9310 13368 9366 13424
rect 9494 13368 9550 13424
rect 9034 12860 9036 12880
rect 9036 12860 9088 12880
rect 9088 12860 9090 12880
rect 9034 12824 9090 12860
rect 8666 10648 8722 10704
rect 8942 10240 8998 10296
rect 8758 9968 8814 10024
rect 8574 9016 8630 9072
rect 8298 8472 8354 8528
rect 8574 8064 8630 8120
rect 8206 7656 8262 7712
rect 8022 6296 8078 6352
rect 7628 6010 7684 6012
rect 7708 6010 7764 6012
rect 7788 6010 7844 6012
rect 7868 6010 7924 6012
rect 7628 5958 7674 6010
rect 7674 5958 7684 6010
rect 7708 5958 7738 6010
rect 7738 5958 7750 6010
rect 7750 5958 7764 6010
rect 7788 5958 7802 6010
rect 7802 5958 7814 6010
rect 7814 5958 7844 6010
rect 7868 5958 7878 6010
rect 7878 5958 7924 6010
rect 7628 5956 7684 5958
rect 7708 5956 7764 5958
rect 7788 5956 7844 5958
rect 7868 5956 7924 5958
rect 7102 4800 7158 4856
rect 6642 2624 6698 2680
rect 6642 2488 6698 2544
rect 6918 2760 6974 2816
rect 7378 5344 7434 5400
rect 7194 3188 7250 3224
rect 7194 3168 7196 3188
rect 7196 3168 7248 3188
rect 7248 3168 7250 3188
rect 7470 4936 7526 4992
rect 7628 4922 7684 4924
rect 7708 4922 7764 4924
rect 7788 4922 7844 4924
rect 7868 4922 7924 4924
rect 7628 4870 7674 4922
rect 7674 4870 7684 4922
rect 7708 4870 7738 4922
rect 7738 4870 7750 4922
rect 7750 4870 7764 4922
rect 7788 4870 7802 4922
rect 7802 4870 7814 4922
rect 7814 4870 7844 4922
rect 7868 4870 7878 4922
rect 7878 4870 7924 4922
rect 7628 4868 7684 4870
rect 7708 4868 7764 4870
rect 7788 4868 7844 4870
rect 7868 4868 7924 4870
rect 7628 3834 7684 3836
rect 7708 3834 7764 3836
rect 7788 3834 7844 3836
rect 7868 3834 7924 3836
rect 7628 3782 7674 3834
rect 7674 3782 7684 3834
rect 7708 3782 7738 3834
rect 7738 3782 7750 3834
rect 7750 3782 7764 3834
rect 7788 3782 7802 3834
rect 7802 3782 7814 3834
rect 7814 3782 7844 3834
rect 7868 3782 7878 3834
rect 7878 3782 7924 3834
rect 7628 3780 7684 3782
rect 7708 3780 7764 3782
rect 7788 3780 7844 3782
rect 7868 3780 7924 3782
rect 7470 3712 7526 3768
rect 7930 3304 7986 3360
rect 7194 2796 7196 2816
rect 7196 2796 7248 2816
rect 7248 2796 7250 2816
rect 7194 2760 7250 2796
rect 7102 2624 7158 2680
rect 7628 2746 7684 2748
rect 7708 2746 7764 2748
rect 7788 2746 7844 2748
rect 7868 2746 7924 2748
rect 7628 2694 7674 2746
rect 7674 2694 7684 2746
rect 7708 2694 7738 2746
rect 7738 2694 7750 2746
rect 7750 2694 7764 2746
rect 7788 2694 7802 2746
rect 7802 2694 7814 2746
rect 7814 2694 7844 2746
rect 7868 2694 7878 2746
rect 7878 2694 7924 2746
rect 7628 2692 7684 2694
rect 7708 2692 7764 2694
rect 7788 2692 7844 2694
rect 7868 2692 7924 2694
rect 8758 5752 8814 5808
rect 8758 5208 8814 5264
rect 8206 4120 8262 4176
rect 8206 3848 8262 3904
rect 8022 2624 8078 2680
rect 8206 3168 8262 3224
rect 8482 2216 8538 2272
rect 9126 10240 9182 10296
rect 9586 13096 9642 13152
rect 9852 13082 9908 13084
rect 9932 13082 9988 13084
rect 10012 13082 10068 13084
rect 10092 13082 10148 13084
rect 9852 13030 9898 13082
rect 9898 13030 9908 13082
rect 9932 13030 9962 13082
rect 9962 13030 9974 13082
rect 9974 13030 9988 13082
rect 10012 13030 10026 13082
rect 10026 13030 10038 13082
rect 10038 13030 10068 13082
rect 10092 13030 10102 13082
rect 10102 13030 10148 13082
rect 9852 13028 9908 13030
rect 9932 13028 9988 13030
rect 10012 13028 10068 13030
rect 10092 13028 10148 13030
rect 9678 12960 9734 13016
rect 9770 12416 9826 12472
rect 10138 12552 10194 12608
rect 15658 16904 15714 16960
rect 10874 15136 10930 15192
rect 10322 12280 10378 12336
rect 10598 14048 10654 14104
rect 10690 13096 10746 13152
rect 10322 12044 10324 12064
rect 10324 12044 10376 12064
rect 10376 12044 10378 12064
rect 10322 12008 10378 12044
rect 9852 11994 9908 11996
rect 9932 11994 9988 11996
rect 10012 11994 10068 11996
rect 10092 11994 10148 11996
rect 9852 11942 9898 11994
rect 9898 11942 9908 11994
rect 9932 11942 9962 11994
rect 9962 11942 9974 11994
rect 9974 11942 9988 11994
rect 10012 11942 10026 11994
rect 10026 11942 10038 11994
rect 10038 11942 10068 11994
rect 10092 11942 10102 11994
rect 10102 11942 10148 11994
rect 9852 11940 9908 11942
rect 9932 11940 9988 11942
rect 10012 11940 10068 11942
rect 10092 11940 10148 11942
rect 9310 11056 9366 11112
rect 10322 11736 10378 11792
rect 9852 10906 9908 10908
rect 9932 10906 9988 10908
rect 10012 10906 10068 10908
rect 10092 10906 10148 10908
rect 9852 10854 9898 10906
rect 9898 10854 9908 10906
rect 9932 10854 9962 10906
rect 9962 10854 9974 10906
rect 9974 10854 9988 10906
rect 10012 10854 10026 10906
rect 10026 10854 10038 10906
rect 10038 10854 10068 10906
rect 10092 10854 10102 10906
rect 10102 10854 10148 10906
rect 9852 10852 9908 10854
rect 9932 10852 9988 10854
rect 10012 10852 10068 10854
rect 10092 10852 10148 10854
rect 9862 10648 9918 10704
rect 9862 10004 9864 10024
rect 9864 10004 9916 10024
rect 9916 10004 9918 10024
rect 9862 9968 9918 10004
rect 10230 9968 10286 10024
rect 9852 9818 9908 9820
rect 9932 9818 9988 9820
rect 10012 9818 10068 9820
rect 10092 9818 10148 9820
rect 9852 9766 9898 9818
rect 9898 9766 9908 9818
rect 9932 9766 9962 9818
rect 9962 9766 9974 9818
rect 9974 9766 9988 9818
rect 10012 9766 10026 9818
rect 10026 9766 10038 9818
rect 10038 9766 10068 9818
rect 10092 9766 10102 9818
rect 10102 9766 10148 9818
rect 9852 9764 9908 9766
rect 9932 9764 9988 9766
rect 10012 9764 10068 9766
rect 10092 9764 10148 9766
rect 10230 9696 10286 9752
rect 9678 9016 9734 9072
rect 9586 8472 9642 8528
rect 9852 8730 9908 8732
rect 9932 8730 9988 8732
rect 10012 8730 10068 8732
rect 10092 8730 10148 8732
rect 9852 8678 9898 8730
rect 9898 8678 9908 8730
rect 9932 8678 9962 8730
rect 9962 8678 9974 8730
rect 9974 8678 9988 8730
rect 10012 8678 10026 8730
rect 10026 8678 10038 8730
rect 10038 8678 10068 8730
rect 10092 8678 10102 8730
rect 10102 8678 10148 8730
rect 9852 8676 9908 8678
rect 9932 8676 9988 8678
rect 10012 8676 10068 8678
rect 10092 8676 10148 8678
rect 10690 12008 10746 12064
rect 10598 11600 10654 11656
rect 10414 10376 10470 10432
rect 10506 9696 10562 9752
rect 10322 9016 10378 9072
rect 9218 7928 9274 7984
rect 9310 7248 9366 7304
rect 9218 6704 9274 6760
rect 9034 5752 9090 5808
rect 9310 4392 9366 4448
rect 9852 7642 9908 7644
rect 9932 7642 9988 7644
rect 10012 7642 10068 7644
rect 10092 7642 10148 7644
rect 9852 7590 9898 7642
rect 9898 7590 9908 7642
rect 9932 7590 9962 7642
rect 9962 7590 9974 7642
rect 9974 7590 9988 7642
rect 10012 7590 10026 7642
rect 10026 7590 10038 7642
rect 10038 7590 10068 7642
rect 10092 7590 10102 7642
rect 10102 7590 10148 7642
rect 9852 7588 9908 7590
rect 9932 7588 9988 7590
rect 10012 7588 10068 7590
rect 10092 7588 10148 7590
rect 9770 7384 9826 7440
rect 9954 7384 10010 7440
rect 9494 6432 9550 6488
rect 9954 7112 10010 7168
rect 9852 6554 9908 6556
rect 9932 6554 9988 6556
rect 10012 6554 10068 6556
rect 10092 6554 10148 6556
rect 9852 6502 9898 6554
rect 9898 6502 9908 6554
rect 9932 6502 9962 6554
rect 9962 6502 9974 6554
rect 9974 6502 9988 6554
rect 10012 6502 10026 6554
rect 10026 6502 10038 6554
rect 10038 6502 10068 6554
rect 10092 6502 10102 6554
rect 10102 6502 10148 6554
rect 9852 6500 9908 6502
rect 9932 6500 9988 6502
rect 10012 6500 10068 6502
rect 10092 6500 10148 6502
rect 10322 7792 10378 7848
rect 9494 4120 9550 4176
rect 9852 5466 9908 5468
rect 9932 5466 9988 5468
rect 10012 5466 10068 5468
rect 10092 5466 10148 5468
rect 9852 5414 9898 5466
rect 9898 5414 9908 5466
rect 9932 5414 9962 5466
rect 9962 5414 9974 5466
rect 9974 5414 9988 5466
rect 10012 5414 10026 5466
rect 10026 5414 10038 5466
rect 10038 5414 10068 5466
rect 10092 5414 10102 5466
rect 10102 5414 10148 5466
rect 9852 5412 9908 5414
rect 9932 5412 9988 5414
rect 10012 5412 10068 5414
rect 10092 5412 10148 5414
rect 10414 6160 10470 6216
rect 10230 5072 10286 5128
rect 11058 13268 11060 13288
rect 11060 13268 11112 13288
rect 11112 13268 11114 13288
rect 11058 13232 11114 13268
rect 10782 11056 10838 11112
rect 10690 10104 10746 10160
rect 10966 11872 11022 11928
rect 11886 14864 11942 14920
rect 11794 14592 11850 14648
rect 12076 14714 12132 14716
rect 12156 14714 12212 14716
rect 12236 14714 12292 14716
rect 12316 14714 12372 14716
rect 12076 14662 12122 14714
rect 12122 14662 12132 14714
rect 12156 14662 12186 14714
rect 12186 14662 12198 14714
rect 12198 14662 12212 14714
rect 12236 14662 12250 14714
rect 12250 14662 12262 14714
rect 12262 14662 12292 14714
rect 12316 14662 12326 14714
rect 12326 14662 12372 14714
rect 12076 14660 12132 14662
rect 12156 14660 12212 14662
rect 12236 14660 12292 14662
rect 12316 14660 12372 14662
rect 11334 12960 11390 13016
rect 11518 13232 11574 13288
rect 11610 12824 11666 12880
rect 11426 12688 11482 12744
rect 11334 12552 11390 12608
rect 11242 12436 11298 12472
rect 11242 12416 11244 12436
rect 11244 12416 11296 12436
rect 11296 12416 11298 12436
rect 10966 11212 11022 11248
rect 10966 11192 10968 11212
rect 10968 11192 11020 11212
rect 11020 11192 11022 11212
rect 11058 10920 11114 10976
rect 10782 9580 10838 9616
rect 10782 9560 10784 9580
rect 10784 9560 10836 9580
rect 10836 9560 10838 9580
rect 10690 9152 10746 9208
rect 10966 8780 10968 8800
rect 10968 8780 11020 8800
rect 11020 8780 11022 8800
rect 10966 8744 11022 8780
rect 11242 11464 11298 11520
rect 11150 10376 11206 10432
rect 10690 6024 10746 6080
rect 10230 4392 10286 4448
rect 9852 4378 9908 4380
rect 9932 4378 9988 4380
rect 10012 4378 10068 4380
rect 10092 4378 10148 4380
rect 9852 4326 9898 4378
rect 9898 4326 9908 4378
rect 9932 4326 9962 4378
rect 9962 4326 9974 4378
rect 9974 4326 9988 4378
rect 10012 4326 10026 4378
rect 10026 4326 10038 4378
rect 10038 4326 10068 4378
rect 10092 4326 10102 4378
rect 10102 4326 10148 4378
rect 9852 4324 9908 4326
rect 9932 4324 9988 4326
rect 10012 4324 10068 4326
rect 10092 4324 10148 4326
rect 10230 4276 10286 4312
rect 10230 4256 10232 4276
rect 10232 4256 10284 4276
rect 10284 4256 10286 4276
rect 9852 3290 9908 3292
rect 9932 3290 9988 3292
rect 10012 3290 10068 3292
rect 10092 3290 10148 3292
rect 9852 3238 9898 3290
rect 9898 3238 9908 3290
rect 9932 3238 9962 3290
rect 9962 3238 9974 3290
rect 9974 3238 9988 3290
rect 10012 3238 10026 3290
rect 10026 3238 10038 3290
rect 10038 3238 10068 3290
rect 10092 3238 10102 3290
rect 10102 3238 10148 3290
rect 9852 3236 9908 3238
rect 9932 3236 9988 3238
rect 10012 3236 10068 3238
rect 10092 3236 10148 3238
rect 11334 10004 11336 10024
rect 11336 10004 11388 10024
rect 11388 10004 11390 10024
rect 11334 9968 11390 10004
rect 11242 9016 11298 9072
rect 11518 10376 11574 10432
rect 11518 10240 11574 10296
rect 10874 5208 10930 5264
rect 10598 3848 10654 3904
rect 10874 4256 10930 4312
rect 10690 3304 10746 3360
rect 10598 3168 10654 3224
rect 10506 2916 10562 2952
rect 10506 2896 10508 2916
rect 10508 2896 10560 2916
rect 10560 2896 10562 2916
rect 9852 2202 9908 2204
rect 9932 2202 9988 2204
rect 10012 2202 10068 2204
rect 10092 2202 10148 2204
rect 9852 2150 9898 2202
rect 9898 2150 9908 2202
rect 9932 2150 9962 2202
rect 9962 2150 9974 2202
rect 9974 2150 9988 2202
rect 10012 2150 10026 2202
rect 10026 2150 10038 2202
rect 10038 2150 10068 2202
rect 10092 2150 10102 2202
rect 10102 2150 10148 2202
rect 9852 2148 9908 2150
rect 9932 2148 9988 2150
rect 10012 2148 10068 2150
rect 10092 2148 10148 2150
rect 9494 1536 9550 1592
rect 11794 14048 11850 14104
rect 11886 13676 11888 13696
rect 11888 13676 11940 13696
rect 11940 13676 11942 13696
rect 11886 13640 11942 13676
rect 12162 14048 12218 14104
rect 12346 14048 12402 14104
rect 12714 15000 12770 15056
rect 12898 15000 12954 15056
rect 12714 14592 12770 14648
rect 12898 14728 12954 14784
rect 12806 14048 12862 14104
rect 13082 13932 13138 13968
rect 13082 13912 13084 13932
rect 13084 13912 13136 13932
rect 13136 13912 13138 13932
rect 12806 13776 12862 13832
rect 13082 13776 13138 13832
rect 12714 13640 12770 13696
rect 12076 13626 12132 13628
rect 12156 13626 12212 13628
rect 12236 13626 12292 13628
rect 12316 13626 12372 13628
rect 12076 13574 12122 13626
rect 12122 13574 12132 13626
rect 12156 13574 12186 13626
rect 12186 13574 12198 13626
rect 12198 13574 12212 13626
rect 12236 13574 12250 13626
rect 12250 13574 12262 13626
rect 12262 13574 12292 13626
rect 12316 13574 12326 13626
rect 12326 13574 12372 13626
rect 12076 13572 12132 13574
rect 12156 13572 12212 13574
rect 12236 13572 12292 13574
rect 12316 13572 12372 13574
rect 12622 13504 12678 13560
rect 12070 12960 12126 13016
rect 12254 13368 12310 13424
rect 12076 12538 12132 12540
rect 12156 12538 12212 12540
rect 12236 12538 12292 12540
rect 12316 12538 12372 12540
rect 12076 12486 12122 12538
rect 12122 12486 12132 12538
rect 12156 12486 12186 12538
rect 12186 12486 12198 12538
rect 12198 12486 12212 12538
rect 12236 12486 12250 12538
rect 12250 12486 12262 12538
rect 12262 12486 12292 12538
rect 12316 12486 12326 12538
rect 12326 12486 12372 12538
rect 12076 12484 12132 12486
rect 12156 12484 12212 12486
rect 12236 12484 12292 12486
rect 12316 12484 12372 12486
rect 11702 12316 11704 12336
rect 11704 12316 11756 12336
rect 11756 12316 11758 12336
rect 11702 12280 11758 12316
rect 11886 12316 11888 12336
rect 11888 12316 11940 12336
rect 11940 12316 11942 12336
rect 11886 12280 11942 12316
rect 11610 9968 11666 10024
rect 11610 9716 11666 9752
rect 11610 9696 11612 9716
rect 11612 9696 11664 9716
rect 11664 9696 11666 9716
rect 11702 9444 11758 9480
rect 11702 9424 11704 9444
rect 11704 9424 11756 9444
rect 11756 9424 11758 9444
rect 11334 6568 11390 6624
rect 11150 3848 11206 3904
rect 12622 13096 12678 13152
rect 12714 12824 12770 12880
rect 12898 12960 12954 13016
rect 13910 14476 13966 14512
rect 13910 14456 13912 14476
rect 13912 14456 13964 14476
rect 13964 14456 13966 14476
rect 13818 14184 13874 14240
rect 14002 14048 14058 14104
rect 13542 13368 13598 13424
rect 12714 12416 12770 12472
rect 12162 12044 12164 12064
rect 12164 12044 12216 12064
rect 12216 12044 12218 12064
rect 12162 12008 12218 12044
rect 11978 11892 12034 11928
rect 11978 11872 11980 11892
rect 11980 11872 12032 11892
rect 12032 11872 12034 11892
rect 12346 11736 12402 11792
rect 11886 8336 11942 8392
rect 11794 7792 11850 7848
rect 11794 6452 11850 6488
rect 11794 6432 11796 6452
rect 11796 6432 11848 6452
rect 11848 6432 11850 6452
rect 11610 4528 11666 4584
rect 11610 3712 11666 3768
rect 12076 11450 12132 11452
rect 12156 11450 12212 11452
rect 12236 11450 12292 11452
rect 12316 11450 12372 11452
rect 12076 11398 12122 11450
rect 12122 11398 12132 11450
rect 12156 11398 12186 11450
rect 12186 11398 12198 11450
rect 12198 11398 12212 11450
rect 12236 11398 12250 11450
rect 12250 11398 12262 11450
rect 12262 11398 12292 11450
rect 12316 11398 12326 11450
rect 12326 11398 12372 11450
rect 12076 11396 12132 11398
rect 12156 11396 12212 11398
rect 12236 11396 12292 11398
rect 12316 11396 12372 11398
rect 12254 11212 12310 11248
rect 12254 11192 12256 11212
rect 12256 11192 12308 11212
rect 12308 11192 12310 11212
rect 12530 12144 12586 12200
rect 12254 11056 12310 11112
rect 12162 10784 12218 10840
rect 12162 10532 12218 10568
rect 12162 10512 12164 10532
rect 12164 10512 12216 10532
rect 12216 10512 12218 10532
rect 12076 10362 12132 10364
rect 12156 10362 12212 10364
rect 12236 10362 12292 10364
rect 12316 10362 12372 10364
rect 12076 10310 12122 10362
rect 12122 10310 12132 10362
rect 12156 10310 12186 10362
rect 12186 10310 12198 10362
rect 12198 10310 12212 10362
rect 12236 10310 12250 10362
rect 12250 10310 12262 10362
rect 12262 10310 12292 10362
rect 12316 10310 12326 10362
rect 12326 10310 12372 10362
rect 12076 10308 12132 10310
rect 12156 10308 12212 10310
rect 12236 10308 12292 10310
rect 12316 10308 12372 10310
rect 12438 9832 12494 9888
rect 12438 9424 12494 9480
rect 12806 11736 12862 11792
rect 13174 11872 13230 11928
rect 13082 11736 13138 11792
rect 13082 11620 13138 11656
rect 13082 11600 13084 11620
rect 13084 11600 13136 11620
rect 13136 11600 13138 11620
rect 13082 11464 13138 11520
rect 12898 11328 12954 11384
rect 12622 10240 12678 10296
rect 12076 9274 12132 9276
rect 12156 9274 12212 9276
rect 12236 9274 12292 9276
rect 12316 9274 12372 9276
rect 12076 9222 12122 9274
rect 12122 9222 12132 9274
rect 12156 9222 12186 9274
rect 12186 9222 12198 9274
rect 12198 9222 12212 9274
rect 12236 9222 12250 9274
rect 12250 9222 12262 9274
rect 12262 9222 12292 9274
rect 12316 9222 12326 9274
rect 12326 9222 12372 9274
rect 12076 9220 12132 9222
rect 12156 9220 12212 9222
rect 12236 9220 12292 9222
rect 12316 9220 12372 9222
rect 12530 9152 12586 9208
rect 12070 9016 12126 9072
rect 12438 8744 12494 8800
rect 12076 8186 12132 8188
rect 12156 8186 12212 8188
rect 12236 8186 12292 8188
rect 12316 8186 12372 8188
rect 12076 8134 12122 8186
rect 12122 8134 12132 8186
rect 12156 8134 12186 8186
rect 12186 8134 12198 8186
rect 12198 8134 12212 8186
rect 12236 8134 12250 8186
rect 12250 8134 12262 8186
rect 12262 8134 12292 8186
rect 12316 8134 12326 8186
rect 12326 8134 12372 8186
rect 12076 8132 12132 8134
rect 12156 8132 12212 8134
rect 12236 8132 12292 8134
rect 12316 8132 12372 8134
rect 12990 11192 13046 11248
rect 12806 9288 12862 9344
rect 12076 7098 12132 7100
rect 12156 7098 12212 7100
rect 12236 7098 12292 7100
rect 12316 7098 12372 7100
rect 12076 7046 12122 7098
rect 12122 7046 12132 7098
rect 12156 7046 12186 7098
rect 12186 7046 12198 7098
rect 12198 7046 12212 7098
rect 12236 7046 12250 7098
rect 12250 7046 12262 7098
rect 12262 7046 12292 7098
rect 12316 7046 12326 7098
rect 12326 7046 12372 7098
rect 12076 7044 12132 7046
rect 12156 7044 12212 7046
rect 12236 7044 12292 7046
rect 12316 7044 12372 7046
rect 12076 6010 12132 6012
rect 12156 6010 12212 6012
rect 12236 6010 12292 6012
rect 12316 6010 12372 6012
rect 12076 5958 12122 6010
rect 12122 5958 12132 6010
rect 12156 5958 12186 6010
rect 12186 5958 12198 6010
rect 12198 5958 12212 6010
rect 12236 5958 12250 6010
rect 12250 5958 12262 6010
rect 12262 5958 12292 6010
rect 12316 5958 12326 6010
rect 12326 5958 12372 6010
rect 12076 5956 12132 5958
rect 12156 5956 12212 5958
rect 12236 5956 12292 5958
rect 12316 5956 12372 5958
rect 13358 12280 13414 12336
rect 13634 12824 13690 12880
rect 13634 12416 13690 12472
rect 13818 13776 13874 13832
rect 13818 12280 13874 12336
rect 13634 12008 13690 12064
rect 13818 12044 13820 12064
rect 13820 12044 13872 12064
rect 13872 12044 13874 12064
rect 13818 12008 13874 12044
rect 13818 11600 13874 11656
rect 13726 11464 13782 11520
rect 12990 6976 13046 7032
rect 13082 6452 13138 6488
rect 13082 6432 13084 6452
rect 13084 6432 13136 6452
rect 13136 6432 13138 6452
rect 11978 5072 12034 5128
rect 12346 5072 12402 5128
rect 12076 4922 12132 4924
rect 12156 4922 12212 4924
rect 12236 4922 12292 4924
rect 12316 4922 12372 4924
rect 12076 4870 12122 4922
rect 12122 4870 12132 4922
rect 12156 4870 12186 4922
rect 12186 4870 12198 4922
rect 12198 4870 12212 4922
rect 12236 4870 12250 4922
rect 12250 4870 12262 4922
rect 12262 4870 12292 4922
rect 12316 4870 12326 4922
rect 12326 4870 12372 4922
rect 12076 4868 12132 4870
rect 12156 4868 12212 4870
rect 12236 4868 12292 4870
rect 12316 4868 12372 4870
rect 11978 4120 12034 4176
rect 13266 6840 13322 6896
rect 12076 3834 12132 3836
rect 12156 3834 12212 3836
rect 12236 3834 12292 3836
rect 12316 3834 12372 3836
rect 12076 3782 12122 3834
rect 12122 3782 12132 3834
rect 12156 3782 12186 3834
rect 12186 3782 12198 3834
rect 12198 3782 12212 3834
rect 12236 3782 12250 3834
rect 12250 3782 12262 3834
rect 12262 3782 12292 3834
rect 12316 3782 12326 3834
rect 12326 3782 12372 3834
rect 12076 3780 12132 3782
rect 12156 3780 12212 3782
rect 12236 3780 12292 3782
rect 12316 3780 12372 3782
rect 12070 3304 12126 3360
rect 12070 3032 12126 3088
rect 12622 3576 12678 3632
rect 12076 2746 12132 2748
rect 12156 2746 12212 2748
rect 12236 2746 12292 2748
rect 12316 2746 12372 2748
rect 12076 2694 12122 2746
rect 12122 2694 12132 2746
rect 12156 2694 12186 2746
rect 12186 2694 12198 2746
rect 12198 2694 12212 2746
rect 12236 2694 12250 2746
rect 12250 2694 12262 2746
rect 12262 2694 12292 2746
rect 12316 2694 12326 2746
rect 12326 2694 12372 2746
rect 12076 2692 12132 2694
rect 12156 2692 12212 2694
rect 12236 2692 12292 2694
rect 12316 2692 12372 2694
rect 11886 1944 11942 2000
rect 13174 3576 13230 3632
rect 13358 4528 13414 4584
rect 13450 3440 13506 3496
rect 13542 3168 13598 3224
rect 12530 1400 12586 1456
rect 13818 10784 13874 10840
rect 14300 14170 14356 14172
rect 14380 14170 14436 14172
rect 14460 14170 14516 14172
rect 14540 14170 14596 14172
rect 14300 14118 14346 14170
rect 14346 14118 14356 14170
rect 14380 14118 14410 14170
rect 14410 14118 14422 14170
rect 14422 14118 14436 14170
rect 14460 14118 14474 14170
rect 14474 14118 14486 14170
rect 14486 14118 14516 14170
rect 14540 14118 14550 14170
rect 14550 14118 14596 14170
rect 14300 14116 14356 14118
rect 14380 14116 14436 14118
rect 14460 14116 14516 14118
rect 14540 14116 14596 14118
rect 14738 14048 14794 14104
rect 15106 14592 15162 14648
rect 14922 14456 14978 14512
rect 14370 13796 14426 13832
rect 14370 13776 14372 13796
rect 14372 13776 14424 13796
rect 14424 13776 14426 13796
rect 14554 13504 14610 13560
rect 14370 13368 14426 13424
rect 14300 13082 14356 13084
rect 14380 13082 14436 13084
rect 14460 13082 14516 13084
rect 14540 13082 14596 13084
rect 14300 13030 14346 13082
rect 14346 13030 14356 13082
rect 14380 13030 14410 13082
rect 14410 13030 14422 13082
rect 14422 13030 14436 13082
rect 14460 13030 14474 13082
rect 14474 13030 14486 13082
rect 14486 13030 14516 13082
rect 14540 13030 14550 13082
rect 14550 13030 14596 13082
rect 14300 13028 14356 13030
rect 14380 13028 14436 13030
rect 14460 13028 14516 13030
rect 14540 13028 14596 13030
rect 14094 12844 14150 12880
rect 14094 12824 14096 12844
rect 14096 12824 14148 12844
rect 14148 12824 14150 12844
rect 14278 12708 14334 12744
rect 14278 12688 14280 12708
rect 14280 12688 14332 12708
rect 14332 12688 14334 12708
rect 14462 12688 14518 12744
rect 14554 12416 14610 12472
rect 14186 12280 14242 12336
rect 14002 11600 14058 11656
rect 14094 11328 14150 11384
rect 14300 11994 14356 11996
rect 14380 11994 14436 11996
rect 14460 11994 14516 11996
rect 14540 11994 14596 11996
rect 14300 11942 14346 11994
rect 14346 11942 14356 11994
rect 14380 11942 14410 11994
rect 14410 11942 14422 11994
rect 14422 11942 14436 11994
rect 14460 11942 14474 11994
rect 14474 11942 14486 11994
rect 14486 11942 14516 11994
rect 14540 11942 14550 11994
rect 14550 11942 14596 11994
rect 14300 11940 14356 11942
rect 14380 11940 14436 11942
rect 14460 11940 14516 11942
rect 14540 11940 14596 11942
rect 14370 11328 14426 11384
rect 16302 16496 16358 16552
rect 15842 15000 15898 15056
rect 16026 15000 16082 15056
rect 17682 16088 17738 16144
rect 17590 15680 17646 15736
rect 16210 14728 16266 14784
rect 15474 14320 15530 14376
rect 15382 13932 15438 13968
rect 15382 13912 15384 13932
rect 15384 13912 15436 13932
rect 15436 13912 15438 13932
rect 14922 13504 14978 13560
rect 14830 13368 14886 13424
rect 14922 13096 14978 13152
rect 15290 13776 15346 13832
rect 15106 13232 15162 13288
rect 14300 10906 14356 10908
rect 14380 10906 14436 10908
rect 14460 10906 14516 10908
rect 14540 10906 14596 10908
rect 14300 10854 14346 10906
rect 14346 10854 14356 10906
rect 14380 10854 14410 10906
rect 14410 10854 14422 10906
rect 14422 10854 14436 10906
rect 14460 10854 14474 10906
rect 14474 10854 14486 10906
rect 14486 10854 14516 10906
rect 14540 10854 14550 10906
rect 14550 10854 14596 10906
rect 14300 10852 14356 10854
rect 14380 10852 14436 10854
rect 14460 10852 14516 10854
rect 14540 10852 14596 10854
rect 14370 10376 14426 10432
rect 14554 10240 14610 10296
rect 15198 12588 15200 12608
rect 15200 12588 15252 12608
rect 15252 12588 15254 12608
rect 15198 12552 15254 12588
rect 14830 11056 14886 11112
rect 15106 12008 15162 12064
rect 14646 10104 14702 10160
rect 14300 9818 14356 9820
rect 14380 9818 14436 9820
rect 14460 9818 14516 9820
rect 14540 9818 14596 9820
rect 14300 9766 14346 9818
rect 14346 9766 14356 9818
rect 14380 9766 14410 9818
rect 14410 9766 14422 9818
rect 14422 9766 14436 9818
rect 14460 9766 14474 9818
rect 14474 9766 14486 9818
rect 14486 9766 14516 9818
rect 14540 9766 14550 9818
rect 14550 9766 14596 9818
rect 14300 9764 14356 9766
rect 14380 9764 14436 9766
rect 14460 9764 14516 9766
rect 14540 9764 14596 9766
rect 13818 7928 13874 7984
rect 14300 8730 14356 8732
rect 14380 8730 14436 8732
rect 14460 8730 14516 8732
rect 14540 8730 14596 8732
rect 14300 8678 14346 8730
rect 14346 8678 14356 8730
rect 14380 8678 14410 8730
rect 14410 8678 14422 8730
rect 14422 8678 14436 8730
rect 14460 8678 14474 8730
rect 14474 8678 14486 8730
rect 14486 8678 14516 8730
rect 14540 8678 14550 8730
rect 14550 8678 14596 8730
rect 14300 8676 14356 8678
rect 14380 8676 14436 8678
rect 14460 8676 14516 8678
rect 14540 8676 14596 8678
rect 14002 6568 14058 6624
rect 14002 6160 14058 6216
rect 13726 4392 13782 4448
rect 14002 5480 14058 5536
rect 14300 7642 14356 7644
rect 14380 7642 14436 7644
rect 14460 7642 14516 7644
rect 14540 7642 14596 7644
rect 14300 7590 14346 7642
rect 14346 7590 14356 7642
rect 14380 7590 14410 7642
rect 14410 7590 14422 7642
rect 14422 7590 14436 7642
rect 14460 7590 14474 7642
rect 14474 7590 14486 7642
rect 14486 7590 14516 7642
rect 14540 7590 14550 7642
rect 14550 7590 14596 7642
rect 14300 7588 14356 7590
rect 14380 7588 14436 7590
rect 14460 7588 14516 7590
rect 14540 7588 14596 7590
rect 14300 6554 14356 6556
rect 14380 6554 14436 6556
rect 14460 6554 14516 6556
rect 14540 6554 14596 6556
rect 14300 6502 14346 6554
rect 14346 6502 14356 6554
rect 14380 6502 14410 6554
rect 14410 6502 14422 6554
rect 14422 6502 14436 6554
rect 14460 6502 14474 6554
rect 14474 6502 14486 6554
rect 14486 6502 14516 6554
rect 14540 6502 14550 6554
rect 14550 6502 14596 6554
rect 14300 6500 14356 6502
rect 14380 6500 14436 6502
rect 14460 6500 14516 6502
rect 14540 6500 14596 6502
rect 14738 9832 14794 9888
rect 14922 8336 14978 8392
rect 14646 5616 14702 5672
rect 14300 5466 14356 5468
rect 14380 5466 14436 5468
rect 14460 5466 14516 5468
rect 14540 5466 14596 5468
rect 14300 5414 14346 5466
rect 14346 5414 14356 5466
rect 14380 5414 14410 5466
rect 14410 5414 14422 5466
rect 14422 5414 14436 5466
rect 14460 5414 14474 5466
rect 14474 5414 14486 5466
rect 14486 5414 14516 5466
rect 14540 5414 14550 5466
rect 14550 5414 14596 5466
rect 14300 5412 14356 5414
rect 14380 5412 14436 5414
rect 14460 5412 14516 5414
rect 14540 5412 14596 5414
rect 14646 5208 14702 5264
rect 14300 4378 14356 4380
rect 14380 4378 14436 4380
rect 14460 4378 14516 4380
rect 14540 4378 14596 4380
rect 14300 4326 14346 4378
rect 14346 4326 14356 4378
rect 14380 4326 14410 4378
rect 14410 4326 14422 4378
rect 14422 4326 14436 4378
rect 14460 4326 14474 4378
rect 14474 4326 14486 4378
rect 14486 4326 14516 4378
rect 14540 4326 14550 4378
rect 14550 4326 14596 4378
rect 14300 4324 14356 4326
rect 14380 4324 14436 4326
rect 14460 4324 14516 4326
rect 14540 4324 14596 4326
rect 13910 4120 13966 4176
rect 13818 4004 13874 4040
rect 13818 3984 13820 4004
rect 13820 3984 13872 4004
rect 13872 3984 13874 4004
rect 14462 3712 14518 3768
rect 14300 3290 14356 3292
rect 14380 3290 14436 3292
rect 14460 3290 14516 3292
rect 14540 3290 14596 3292
rect 14300 3238 14346 3290
rect 14346 3238 14356 3290
rect 14380 3238 14410 3290
rect 14410 3238 14422 3290
rect 14422 3238 14436 3290
rect 14460 3238 14474 3290
rect 14474 3238 14486 3290
rect 14486 3238 14516 3290
rect 14540 3238 14550 3290
rect 14550 3238 14596 3290
rect 14300 3236 14356 3238
rect 14380 3236 14436 3238
rect 14460 3236 14516 3238
rect 14540 3236 14596 3238
rect 14462 3052 14518 3088
rect 14462 3032 14464 3052
rect 14464 3032 14516 3052
rect 14516 3032 14518 3052
rect 14002 2896 14058 2952
rect 15842 14184 15898 14240
rect 15382 12960 15438 13016
rect 15566 13232 15622 13288
rect 15290 11464 15346 11520
rect 16026 13776 16082 13832
rect 15842 13368 15898 13424
rect 15658 11872 15714 11928
rect 15474 11464 15530 11520
rect 15382 9152 15438 9208
rect 15290 8880 15346 8936
rect 15658 10920 15714 10976
rect 15658 9288 15714 9344
rect 15382 7248 15438 7304
rect 15290 7112 15346 7168
rect 15106 6976 15162 7032
rect 15014 6568 15070 6624
rect 15014 6296 15070 6352
rect 15014 5888 15070 5944
rect 15198 5752 15254 5808
rect 15014 4664 15070 4720
rect 15106 3984 15162 4040
rect 17314 14864 17370 14920
rect 16524 14714 16580 14716
rect 16604 14714 16660 14716
rect 16684 14714 16740 14716
rect 16764 14714 16820 14716
rect 16524 14662 16570 14714
rect 16570 14662 16580 14714
rect 16604 14662 16634 14714
rect 16634 14662 16646 14714
rect 16646 14662 16660 14714
rect 16684 14662 16698 14714
rect 16698 14662 16710 14714
rect 16710 14662 16740 14714
rect 16764 14662 16774 14714
rect 16774 14662 16820 14714
rect 16524 14660 16580 14662
rect 16604 14660 16660 14662
rect 16684 14660 16740 14662
rect 16764 14660 16820 14662
rect 16946 14592 17002 14648
rect 16394 14184 16450 14240
rect 16524 13626 16580 13628
rect 16604 13626 16660 13628
rect 16684 13626 16740 13628
rect 16764 13626 16820 13628
rect 16524 13574 16570 13626
rect 16570 13574 16580 13626
rect 16604 13574 16634 13626
rect 16634 13574 16646 13626
rect 16646 13574 16660 13626
rect 16684 13574 16698 13626
rect 16698 13574 16710 13626
rect 16710 13574 16740 13626
rect 16764 13574 16774 13626
rect 16774 13574 16820 13626
rect 16524 13572 16580 13574
rect 16604 13572 16660 13574
rect 16684 13572 16740 13574
rect 16764 13572 16820 13574
rect 16302 13504 16358 13560
rect 16210 12708 16266 12744
rect 16210 12688 16212 12708
rect 16212 12688 16264 12708
rect 16264 12688 16266 12708
rect 16486 13096 16542 13152
rect 15842 11464 15898 11520
rect 16524 12538 16580 12540
rect 16604 12538 16660 12540
rect 16684 12538 16740 12540
rect 16764 12538 16820 12540
rect 16524 12486 16570 12538
rect 16570 12486 16580 12538
rect 16604 12486 16634 12538
rect 16634 12486 16646 12538
rect 16646 12486 16660 12538
rect 16684 12486 16698 12538
rect 16698 12486 16710 12538
rect 16710 12486 16740 12538
rect 16764 12486 16774 12538
rect 16774 12486 16820 12538
rect 16524 12484 16580 12486
rect 16604 12484 16660 12486
rect 16684 12484 16740 12486
rect 16764 12484 16820 12486
rect 16524 11450 16580 11452
rect 16604 11450 16660 11452
rect 16684 11450 16740 11452
rect 16764 11450 16820 11452
rect 16524 11398 16570 11450
rect 16570 11398 16580 11450
rect 16604 11398 16634 11450
rect 16634 11398 16646 11450
rect 16646 11398 16660 11450
rect 16684 11398 16698 11450
rect 16698 11398 16710 11450
rect 16710 11398 16740 11450
rect 16764 11398 16774 11450
rect 16774 11398 16820 11450
rect 16524 11396 16580 11398
rect 16604 11396 16660 11398
rect 16684 11396 16740 11398
rect 16764 11396 16820 11398
rect 16946 12008 17002 12064
rect 16302 10648 16358 10704
rect 16524 10362 16580 10364
rect 16604 10362 16660 10364
rect 16684 10362 16740 10364
rect 16764 10362 16820 10364
rect 16524 10310 16570 10362
rect 16570 10310 16580 10362
rect 16604 10310 16634 10362
rect 16634 10310 16646 10362
rect 16646 10310 16660 10362
rect 16684 10310 16698 10362
rect 16698 10310 16710 10362
rect 16710 10310 16740 10362
rect 16764 10310 16774 10362
rect 16774 10310 16820 10362
rect 16524 10308 16580 10310
rect 16604 10308 16660 10310
rect 16684 10308 16740 10310
rect 16764 10308 16820 10310
rect 16394 10104 16450 10160
rect 15658 6296 15714 6352
rect 15934 7520 15990 7576
rect 16210 7792 16266 7848
rect 16302 7520 16358 7576
rect 16302 7112 16358 7168
rect 15842 6024 15898 6080
rect 16026 6160 16082 6216
rect 15382 3188 15438 3224
rect 15382 3168 15384 3188
rect 15384 3168 15436 3188
rect 15436 3168 15438 3188
rect 15474 2896 15530 2952
rect 14830 2760 14886 2816
rect 14300 2202 14356 2204
rect 14380 2202 14436 2204
rect 14460 2202 14516 2204
rect 14540 2202 14596 2204
rect 14300 2150 14346 2202
rect 14346 2150 14356 2202
rect 14380 2150 14410 2202
rect 14410 2150 14422 2202
rect 14422 2150 14436 2202
rect 14460 2150 14474 2202
rect 14474 2150 14486 2202
rect 14486 2150 14516 2202
rect 14540 2150 14550 2202
rect 14550 2150 14596 2202
rect 14300 2148 14356 2150
rect 14380 2148 14436 2150
rect 14460 2148 14516 2150
rect 14540 2148 14596 2150
rect 16210 5480 16266 5536
rect 16762 9696 16818 9752
rect 16524 9274 16580 9276
rect 16604 9274 16660 9276
rect 16684 9274 16740 9276
rect 16764 9274 16820 9276
rect 16524 9222 16570 9274
rect 16570 9222 16580 9274
rect 16604 9222 16634 9274
rect 16634 9222 16646 9274
rect 16646 9222 16660 9274
rect 16684 9222 16698 9274
rect 16698 9222 16710 9274
rect 16710 9222 16740 9274
rect 16764 9222 16774 9274
rect 16774 9222 16820 9274
rect 16524 9220 16580 9222
rect 16604 9220 16660 9222
rect 16684 9220 16740 9222
rect 16764 9220 16820 9222
rect 17222 12164 17278 12200
rect 17222 12144 17224 12164
rect 17224 12144 17276 12164
rect 17276 12144 17278 12164
rect 17038 9596 17040 9616
rect 17040 9596 17092 9616
rect 17092 9596 17094 9616
rect 17038 9560 17094 9596
rect 17314 10920 17370 10976
rect 17222 10784 17278 10840
rect 16524 8186 16580 8188
rect 16604 8186 16660 8188
rect 16684 8186 16740 8188
rect 16764 8186 16820 8188
rect 16524 8134 16570 8186
rect 16570 8134 16580 8186
rect 16604 8134 16634 8186
rect 16634 8134 16646 8186
rect 16646 8134 16660 8186
rect 16684 8134 16698 8186
rect 16698 8134 16710 8186
rect 16710 8134 16740 8186
rect 16764 8134 16774 8186
rect 16774 8134 16820 8186
rect 16524 8132 16580 8134
rect 16604 8132 16660 8134
rect 16684 8132 16740 8134
rect 16764 8132 16820 8134
rect 17038 7792 17094 7848
rect 16670 7268 16726 7304
rect 16670 7248 16672 7268
rect 16672 7248 16724 7268
rect 16724 7248 16726 7268
rect 16524 7098 16580 7100
rect 16604 7098 16660 7100
rect 16684 7098 16740 7100
rect 16764 7098 16820 7100
rect 16524 7046 16570 7098
rect 16570 7046 16580 7098
rect 16604 7046 16634 7098
rect 16634 7046 16646 7098
rect 16646 7046 16660 7098
rect 16684 7046 16698 7098
rect 16698 7046 16710 7098
rect 16710 7046 16740 7098
rect 16764 7046 16774 7098
rect 16774 7046 16820 7098
rect 16524 7044 16580 7046
rect 16604 7044 16660 7046
rect 16684 7044 16740 7046
rect 16764 7044 16820 7046
rect 16118 3168 16174 3224
rect 17130 6840 17186 6896
rect 16854 6704 16910 6760
rect 16524 6010 16580 6012
rect 16604 6010 16660 6012
rect 16684 6010 16740 6012
rect 16764 6010 16820 6012
rect 16524 5958 16570 6010
rect 16570 5958 16580 6010
rect 16604 5958 16634 6010
rect 16634 5958 16646 6010
rect 16646 5958 16660 6010
rect 16684 5958 16698 6010
rect 16698 5958 16710 6010
rect 16710 5958 16740 6010
rect 16764 5958 16774 6010
rect 16774 5958 16820 6010
rect 16524 5956 16580 5958
rect 16604 5956 16660 5958
rect 16684 5956 16740 5958
rect 16764 5956 16820 5958
rect 16762 5752 16818 5808
rect 16946 6296 17002 6352
rect 16946 5888 17002 5944
rect 16524 4922 16580 4924
rect 16604 4922 16660 4924
rect 16684 4922 16740 4924
rect 16764 4922 16820 4924
rect 16524 4870 16570 4922
rect 16570 4870 16580 4922
rect 16604 4870 16634 4922
rect 16634 4870 16646 4922
rect 16646 4870 16660 4922
rect 16684 4870 16698 4922
rect 16698 4870 16710 4922
rect 16710 4870 16740 4922
rect 16764 4870 16774 4922
rect 16774 4870 16820 4922
rect 16524 4868 16580 4870
rect 16604 4868 16660 4870
rect 16684 4868 16740 4870
rect 16764 4868 16820 4870
rect 16524 3834 16580 3836
rect 16604 3834 16660 3836
rect 16684 3834 16740 3836
rect 16764 3834 16820 3836
rect 16524 3782 16570 3834
rect 16570 3782 16580 3834
rect 16604 3782 16634 3834
rect 16634 3782 16646 3834
rect 16646 3782 16660 3834
rect 16684 3782 16698 3834
rect 16698 3782 16710 3834
rect 16710 3782 16740 3834
rect 16764 3782 16774 3834
rect 16774 3782 16820 3834
rect 16524 3780 16580 3782
rect 16604 3780 16660 3782
rect 16684 3780 16740 3782
rect 16764 3780 16820 3782
rect 16670 3576 16726 3632
rect 16210 3032 16266 3088
rect 16524 2746 16580 2748
rect 16604 2746 16660 2748
rect 16684 2746 16740 2748
rect 16764 2746 16820 2748
rect 16524 2694 16570 2746
rect 16570 2694 16580 2746
rect 16604 2694 16634 2746
rect 16634 2694 16646 2746
rect 16646 2694 16660 2746
rect 16684 2694 16698 2746
rect 16698 2694 16710 2746
rect 16710 2694 16740 2746
rect 16764 2694 16774 2746
rect 16774 2694 16820 2746
rect 16524 2692 16580 2694
rect 16604 2692 16660 2694
rect 16684 2692 16740 2694
rect 16764 2692 16820 2694
rect 15934 1672 15990 1728
rect 15934 1284 15990 1320
rect 15934 1264 15936 1284
rect 15936 1264 15988 1284
rect 15988 1264 15990 1284
rect 15198 176 15254 232
rect 17038 4120 17094 4176
rect 17682 12688 17738 12744
rect 17682 12300 17738 12336
rect 17682 12280 17684 12300
rect 17684 12280 17736 12300
rect 17736 12280 17738 12300
rect 17866 12280 17922 12336
rect 18510 15408 18566 15464
rect 18234 15136 18290 15192
rect 18510 12960 18566 13016
rect 17774 11600 17830 11656
rect 17958 11328 18014 11384
rect 17682 11192 17738 11248
rect 17498 10104 17554 10160
rect 17958 9832 18014 9888
rect 17222 3476 17224 3496
rect 17224 3476 17276 3496
rect 17276 3476 17278 3496
rect 17222 3440 17278 3476
rect 18602 11736 18658 11792
rect 18510 9968 18566 10024
rect 18234 9288 18290 9344
rect 18510 9696 18566 9752
rect 18418 9288 18474 9344
rect 18050 8472 18106 8528
rect 18050 8336 18106 8392
rect 17958 7404 18014 7440
rect 17958 7384 17960 7404
rect 17960 7384 18012 7404
rect 18012 7384 18014 7404
rect 17590 3984 17646 4040
rect 18326 8064 18382 8120
rect 18694 11464 18750 11520
rect 18694 8880 18750 8936
rect 18510 7792 18566 7848
rect 18602 7384 18658 7440
rect 18418 4664 18474 4720
rect 17498 1672 17554 1728
rect 17314 1536 17370 1592
rect 16946 856 17002 912
rect 18050 2524 18052 2544
rect 18052 2524 18104 2544
rect 18104 2524 18106 2544
rect 18050 2488 18106 2524
rect 18234 2352 18290 2408
rect 17958 1808 18014 1864
rect 18326 2080 18382 2136
rect 18878 3576 18934 3632
rect 18786 2352 18842 2408
rect 15842 448 15898 504
<< metal3 >>
rect 0 16962 800 16992
rect 3785 16962 3851 16965
rect 0 16960 3851 16962
rect 0 16904 3790 16960
rect 3846 16904 3851 16960
rect 0 16902 3851 16904
rect 0 16872 800 16902
rect 3785 16899 3851 16902
rect 15653 16962 15719 16965
rect 19200 16962 20000 16992
rect 15653 16960 20000 16962
rect 15653 16904 15658 16960
rect 15714 16904 20000 16960
rect 15653 16902 20000 16904
rect 15653 16899 15719 16902
rect 19200 16872 20000 16902
rect 0 16690 800 16720
rect 4061 16690 4127 16693
rect 0 16688 4127 16690
rect 0 16632 4066 16688
rect 4122 16632 4127 16688
rect 0 16630 4127 16632
rect 0 16600 800 16630
rect 4061 16627 4127 16630
rect 16297 16554 16363 16557
rect 19200 16554 20000 16584
rect 16297 16552 20000 16554
rect 16297 16496 16302 16552
rect 16358 16496 20000 16552
rect 16297 16494 20000 16496
rect 16297 16491 16363 16494
rect 19200 16464 20000 16494
rect 0 16282 800 16312
rect 4337 16282 4403 16285
rect 0 16280 4403 16282
rect 0 16224 4342 16280
rect 4398 16224 4403 16280
rect 0 16222 4403 16224
rect 0 16192 800 16222
rect 4337 16219 4403 16222
rect 17677 16146 17743 16149
rect 19200 16146 20000 16176
rect 17677 16144 20000 16146
rect 17677 16088 17682 16144
rect 17738 16088 20000 16144
rect 17677 16086 20000 16088
rect 17677 16083 17743 16086
rect 19200 16056 20000 16086
rect 0 16010 800 16040
rect 2129 16010 2195 16013
rect 0 16008 2195 16010
rect 0 15952 2134 16008
rect 2190 15952 2195 16008
rect 0 15950 2195 15952
rect 0 15920 800 15950
rect 2129 15947 2195 15950
rect 974 15812 980 15876
rect 1044 15874 1050 15876
rect 12750 15874 12756 15876
rect 1044 15814 12756 15874
rect 1044 15812 1050 15814
rect 12750 15812 12756 15814
rect 12820 15812 12826 15876
rect 1158 15676 1164 15740
rect 1228 15738 1234 15740
rect 9438 15738 9444 15740
rect 1228 15678 9444 15738
rect 1228 15676 1234 15678
rect 9438 15676 9444 15678
rect 9508 15676 9514 15740
rect 17585 15738 17651 15741
rect 19200 15738 20000 15768
rect 17585 15736 20000 15738
rect 17585 15680 17590 15736
rect 17646 15680 20000 15736
rect 17585 15678 20000 15680
rect 17585 15675 17651 15678
rect 19200 15648 20000 15678
rect 0 15602 800 15632
rect 4613 15602 4679 15605
rect 0 15600 4679 15602
rect 0 15544 4618 15600
rect 4674 15544 4679 15600
rect 0 15542 4679 15544
rect 0 15512 800 15542
rect 4613 15539 4679 15542
rect 2630 15404 2636 15468
rect 2700 15466 2706 15468
rect 12566 15466 12572 15468
rect 2700 15406 12572 15466
rect 2700 15404 2706 15406
rect 12566 15404 12572 15406
rect 12636 15404 12642 15468
rect 18505 15466 18571 15469
rect 19200 15466 20000 15496
rect 18505 15464 20000 15466
rect 18505 15408 18510 15464
rect 18566 15408 20000 15464
rect 18505 15406 20000 15408
rect 18505 15403 18571 15406
rect 19200 15376 20000 15406
rect 0 15330 800 15360
rect 3877 15330 3943 15333
rect 0 15328 3943 15330
rect 0 15272 3882 15328
rect 3938 15272 3943 15328
rect 0 15270 3943 15272
rect 0 15240 800 15270
rect 3877 15267 3943 15270
rect 10869 15194 10935 15197
rect 18229 15194 18295 15197
rect 10869 15192 18295 15194
rect 10869 15136 10874 15192
rect 10930 15136 18234 15192
rect 18290 15136 18295 15192
rect 10869 15134 18295 15136
rect 10869 15131 10935 15134
rect 18229 15131 18295 15134
rect 0 15058 800 15088
rect 2773 15058 2839 15061
rect 0 15056 2839 15058
rect 0 15000 2778 15056
rect 2834 15000 2839 15056
rect 0 14998 2839 15000
rect 0 14968 800 14998
rect 2773 14995 2839 14998
rect 4981 15058 5047 15061
rect 8753 15058 8819 15061
rect 10910 15058 10916 15060
rect 4981 15056 10916 15058
rect 4981 15000 4986 15056
rect 5042 15000 8758 15056
rect 8814 15000 10916 15056
rect 4981 14998 10916 15000
rect 4981 14995 5047 14998
rect 8753 14995 8819 14998
rect 10910 14996 10916 14998
rect 10980 15058 10986 15060
rect 12709 15058 12775 15061
rect 10980 15056 12775 15058
rect 10980 15000 12714 15056
rect 12770 15000 12775 15056
rect 10980 14998 12775 15000
rect 10980 14996 10986 14998
rect 12709 14995 12775 14998
rect 12893 15058 12959 15061
rect 15837 15058 15903 15061
rect 12893 15056 15903 15058
rect 12893 15000 12898 15056
rect 12954 15000 15842 15056
rect 15898 15000 15903 15056
rect 12893 14998 15903 15000
rect 12893 14995 12959 14998
rect 15837 14995 15903 14998
rect 16021 15058 16087 15061
rect 19200 15058 20000 15088
rect 16021 15056 20000 15058
rect 16021 15000 16026 15056
rect 16082 15000 20000 15056
rect 16021 14998 20000 15000
rect 16021 14995 16087 14998
rect 19200 14968 20000 14998
rect 1485 14922 1551 14925
rect 5717 14922 5783 14925
rect 1485 14920 5783 14922
rect 1485 14864 1490 14920
rect 1546 14864 5722 14920
rect 5778 14864 5783 14920
rect 1485 14862 5783 14864
rect 1485 14859 1551 14862
rect 5717 14859 5783 14862
rect 11881 14922 11947 14925
rect 16062 14922 16068 14924
rect 11881 14920 16068 14922
rect 11881 14864 11886 14920
rect 11942 14864 16068 14920
rect 11881 14862 16068 14864
rect 11881 14859 11947 14862
rect 16062 14860 16068 14862
rect 16132 14922 16138 14924
rect 17309 14922 17375 14925
rect 16132 14920 17375 14922
rect 16132 14864 17314 14920
rect 17370 14864 17375 14920
rect 16132 14862 17375 14864
rect 16132 14860 16138 14862
rect 17309 14859 17375 14862
rect 12893 14786 12959 14789
rect 16205 14786 16271 14789
rect 12893 14784 16271 14786
rect 12893 14728 12898 14784
rect 12954 14728 16210 14784
rect 16266 14728 16271 14784
rect 12893 14726 16271 14728
rect 12893 14723 12959 14726
rect 16205 14723 16271 14726
rect 3168 14720 3488 14721
rect 0 14650 800 14680
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 14655 3488 14656
rect 7616 14720 7936 14721
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 14655 7936 14656
rect 12064 14720 12384 14721
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 14655 12384 14656
rect 16512 14720 16832 14721
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16512 14655 16832 14656
rect 2957 14650 3023 14653
rect 0 14648 3023 14650
rect 0 14592 2962 14648
rect 3018 14592 3023 14648
rect 0 14590 3023 14592
rect 0 14560 800 14590
rect 2957 14587 3023 14590
rect 4470 14588 4476 14652
rect 4540 14650 4546 14652
rect 5349 14650 5415 14653
rect 7097 14650 7163 14653
rect 4540 14648 7163 14650
rect 4540 14592 5354 14648
rect 5410 14592 7102 14648
rect 7158 14592 7163 14648
rect 4540 14590 7163 14592
rect 4540 14588 4546 14590
rect 5349 14587 5415 14590
rect 7097 14587 7163 14590
rect 9397 14650 9463 14653
rect 10726 14650 10732 14652
rect 9397 14648 10732 14650
rect 9397 14592 9402 14648
rect 9458 14592 10732 14648
rect 9397 14590 10732 14592
rect 9397 14587 9463 14590
rect 10726 14588 10732 14590
rect 10796 14650 10802 14652
rect 11789 14650 11855 14653
rect 10796 14648 11855 14650
rect 10796 14592 11794 14648
rect 11850 14592 11855 14648
rect 10796 14590 11855 14592
rect 10796 14588 10802 14590
rect 11789 14587 11855 14590
rect 12709 14650 12775 14653
rect 15101 14650 15167 14653
rect 12709 14648 15167 14650
rect 12709 14592 12714 14648
rect 12770 14592 15106 14648
rect 15162 14592 15167 14648
rect 12709 14590 15167 14592
rect 12709 14587 12775 14590
rect 15101 14587 15167 14590
rect 16941 14650 17007 14653
rect 19200 14650 20000 14680
rect 16941 14648 20000 14650
rect 16941 14592 16946 14648
rect 17002 14592 20000 14648
rect 16941 14590 20000 14592
rect 16941 14587 17007 14590
rect 19200 14560 20000 14590
rect 1945 14514 2011 14517
rect 13905 14514 13971 14517
rect 14917 14514 14983 14517
rect 1945 14512 13784 14514
rect 1945 14456 1950 14512
rect 2006 14456 13784 14512
rect 1945 14454 13784 14456
rect 1945 14451 2011 14454
rect 0 14378 800 14408
rect 2773 14378 2839 14381
rect 0 14376 2839 14378
rect 0 14320 2778 14376
rect 2834 14320 2839 14376
rect 0 14318 2839 14320
rect 0 14288 800 14318
rect 2773 14315 2839 14318
rect 5717 14378 5783 14381
rect 6269 14378 6335 14381
rect 10358 14378 10364 14380
rect 5717 14376 6194 14378
rect 5717 14320 5722 14376
rect 5778 14320 6194 14376
rect 5717 14318 6194 14320
rect 5717 14315 5783 14318
rect 2221 14242 2287 14245
rect 5073 14242 5139 14245
rect 2221 14240 5139 14242
rect 2221 14184 2226 14240
rect 2282 14184 5078 14240
rect 5134 14184 5139 14240
rect 2221 14182 5139 14184
rect 6134 14242 6194 14318
rect 6269 14376 10364 14378
rect 6269 14320 6274 14376
rect 6330 14320 10364 14376
rect 6269 14318 10364 14320
rect 6269 14315 6335 14318
rect 10358 14316 10364 14318
rect 10428 14316 10434 14380
rect 13724 14378 13784 14454
rect 13905 14512 14983 14514
rect 13905 14456 13910 14512
rect 13966 14456 14922 14512
rect 14978 14456 14983 14512
rect 13905 14454 14983 14456
rect 13905 14451 13971 14454
rect 14917 14451 14983 14454
rect 15469 14378 15535 14381
rect 13724 14376 15535 14378
rect 13724 14320 15474 14376
rect 15530 14320 15535 14376
rect 13724 14318 15535 14320
rect 15469 14315 15535 14318
rect 6821 14242 6887 14245
rect 6134 14240 6887 14242
rect 6134 14184 6826 14240
rect 6882 14184 6887 14240
rect 6134 14182 6887 14184
rect 2221 14179 2287 14182
rect 5073 14179 5139 14182
rect 6821 14179 6887 14182
rect 10225 14242 10291 14245
rect 13813 14242 13879 14245
rect 10225 14240 13879 14242
rect 10225 14184 10230 14240
rect 10286 14184 13818 14240
rect 13874 14184 13879 14240
rect 10225 14182 13879 14184
rect 10225 14179 10291 14182
rect 13813 14179 13879 14182
rect 15837 14242 15903 14245
rect 16246 14242 16252 14244
rect 15837 14240 16252 14242
rect 15837 14184 15842 14240
rect 15898 14184 16252 14240
rect 15837 14182 16252 14184
rect 15837 14179 15903 14182
rect 16246 14180 16252 14182
rect 16316 14180 16322 14244
rect 16389 14242 16455 14245
rect 19200 14242 20000 14272
rect 16389 14240 20000 14242
rect 16389 14184 16394 14240
rect 16450 14184 20000 14240
rect 16389 14182 20000 14184
rect 16389 14179 16455 14182
rect 5392 14176 5712 14177
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5392 14111 5712 14112
rect 9840 14176 10160 14177
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9840 14111 10160 14112
rect 14288 14176 14608 14177
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 19200 14152 20000 14182
rect 14288 14111 14608 14112
rect 3049 14106 3115 14109
rect 4981 14106 5047 14109
rect 3049 14104 5047 14106
rect 3049 14048 3054 14104
rect 3110 14048 4986 14104
rect 5042 14048 5047 14104
rect 3049 14046 5047 14048
rect 3049 14043 3115 14046
rect 4981 14043 5047 14046
rect 5809 14106 5875 14109
rect 8293 14106 8359 14109
rect 10593 14108 10659 14109
rect 5809 14104 8359 14106
rect 5809 14048 5814 14104
rect 5870 14048 8298 14104
rect 8354 14048 8359 14104
rect 5809 14046 8359 14048
rect 5809 14043 5875 14046
rect 8293 14043 8359 14046
rect 10542 14044 10548 14108
rect 10612 14106 10659 14108
rect 11789 14106 11855 14109
rect 12157 14106 12223 14109
rect 10612 14104 10704 14106
rect 10654 14048 10704 14104
rect 10612 14046 10704 14048
rect 11789 14104 12223 14106
rect 11789 14048 11794 14104
rect 11850 14048 12162 14104
rect 12218 14048 12223 14104
rect 11789 14046 12223 14048
rect 10612 14044 10659 14046
rect 10593 14043 10659 14044
rect 11789 14043 11855 14046
rect 12157 14043 12223 14046
rect 12341 14106 12407 14109
rect 12801 14106 12867 14109
rect 13997 14106 14063 14109
rect 12341 14104 12867 14106
rect 12341 14048 12346 14104
rect 12402 14048 12806 14104
rect 12862 14048 12867 14104
rect 12341 14046 12867 14048
rect 12341 14043 12407 14046
rect 12801 14043 12867 14046
rect 12942 14104 14063 14106
rect 12942 14048 14002 14104
rect 14058 14048 14063 14104
rect 12942 14046 14063 14048
rect 0 13970 800 14000
rect 2405 13970 2471 13973
rect 3233 13970 3299 13973
rect 6913 13970 6979 13973
rect 12942 13970 13002 14046
rect 13997 14043 14063 14046
rect 14733 14106 14799 14109
rect 17350 14106 17356 14108
rect 14733 14104 17356 14106
rect 14733 14048 14738 14104
rect 14794 14048 17356 14104
rect 14733 14046 17356 14048
rect 14733 14043 14799 14046
rect 17350 14044 17356 14046
rect 17420 14044 17426 14108
rect 0 13968 2471 13970
rect 0 13912 2410 13968
rect 2466 13912 2471 13968
rect 0 13910 2471 13912
rect 0 13880 800 13910
rect 2405 13907 2471 13910
rect 2730 13968 6979 13970
rect 2730 13912 3238 13968
rect 3294 13912 6918 13968
rect 6974 13912 6979 13968
rect 2730 13910 6979 13912
rect 0 13698 800 13728
rect 2730 13698 2790 13910
rect 3233 13907 3299 13910
rect 6913 13907 6979 13910
rect 7054 13910 13002 13970
rect 13077 13970 13143 13973
rect 15377 13970 15443 13973
rect 13077 13968 15443 13970
rect 13077 13912 13082 13968
rect 13138 13912 15382 13968
rect 15438 13912 15443 13968
rect 13077 13910 15443 13912
rect 4061 13834 4127 13837
rect 4705 13834 4771 13837
rect 7054 13834 7114 13910
rect 13077 13907 13143 13910
rect 15377 13907 15443 13910
rect 4061 13832 7114 13834
rect 4061 13776 4066 13832
rect 4122 13776 4710 13832
rect 4766 13776 7114 13832
rect 4061 13774 7114 13776
rect 8109 13834 8175 13837
rect 12801 13834 12867 13837
rect 8109 13832 12867 13834
rect 8109 13776 8114 13832
rect 8170 13776 12806 13832
rect 12862 13776 12867 13832
rect 8109 13774 12867 13776
rect 4061 13771 4127 13774
rect 4705 13771 4771 13774
rect 8109 13771 8175 13774
rect 12801 13771 12867 13774
rect 13077 13834 13143 13837
rect 13813 13834 13879 13837
rect 13077 13832 13879 13834
rect 13077 13776 13082 13832
rect 13138 13776 13818 13832
rect 13874 13776 13879 13832
rect 13077 13774 13879 13776
rect 13077 13771 13143 13774
rect 13813 13771 13879 13774
rect 14038 13772 14044 13836
rect 14108 13834 14114 13836
rect 14365 13834 14431 13837
rect 14108 13832 14431 13834
rect 14108 13776 14370 13832
rect 14426 13776 14431 13832
rect 14108 13774 14431 13776
rect 14108 13772 14114 13774
rect 14365 13771 14431 13774
rect 15285 13834 15351 13837
rect 15510 13834 15516 13836
rect 15285 13832 15516 13834
rect 15285 13776 15290 13832
rect 15346 13776 15516 13832
rect 15285 13774 15516 13776
rect 15285 13771 15351 13774
rect 15510 13772 15516 13774
rect 15580 13772 15586 13836
rect 16021 13834 16087 13837
rect 19200 13834 20000 13864
rect 16021 13832 20000 13834
rect 16021 13776 16026 13832
rect 16082 13776 20000 13832
rect 16021 13774 20000 13776
rect 16021 13771 16087 13774
rect 0 13638 2790 13698
rect 0 13608 800 13638
rect 3550 13636 3556 13700
rect 3620 13698 3626 13700
rect 4889 13698 4955 13701
rect 3620 13696 4955 13698
rect 3620 13640 4894 13696
rect 4950 13640 4955 13696
rect 3620 13638 4955 13640
rect 3620 13636 3626 13638
rect 4889 13635 4955 13638
rect 5022 13636 5028 13700
rect 5092 13698 5098 13700
rect 5257 13698 5323 13701
rect 5092 13696 5323 13698
rect 5092 13640 5262 13696
rect 5318 13640 5323 13696
rect 5092 13638 5323 13640
rect 5092 13636 5098 13638
rect 5257 13635 5323 13638
rect 5441 13698 5507 13701
rect 7373 13698 7439 13701
rect 5441 13696 7439 13698
rect 5441 13640 5446 13696
rect 5502 13640 7378 13696
rect 7434 13640 7439 13696
rect 5441 13638 7439 13640
rect 5441 13635 5507 13638
rect 7373 13635 7439 13638
rect 9397 13698 9463 13701
rect 11881 13698 11947 13701
rect 9397 13696 11947 13698
rect 9397 13640 9402 13696
rect 9458 13640 11886 13696
rect 11942 13640 11947 13696
rect 9397 13638 11947 13640
rect 9397 13635 9463 13638
rect 11881 13635 11947 13638
rect 12709 13698 12775 13701
rect 16024 13698 16084 13771
rect 19200 13744 20000 13774
rect 12709 13696 16084 13698
rect 12709 13640 12714 13696
rect 12770 13640 16084 13696
rect 12709 13638 16084 13640
rect 12709 13635 12775 13638
rect 3168 13632 3488 13633
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3168 13567 3488 13568
rect 7616 13632 7936 13633
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 7616 13567 7936 13568
rect 12064 13632 12384 13633
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 12064 13567 12384 13568
rect 16512 13632 16832 13633
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 13567 16832 13568
rect 3601 13562 3667 13565
rect 12617 13562 12683 13565
rect 14549 13562 14615 13565
rect 14774 13562 14780 13564
rect 3601 13560 7528 13562
rect 3601 13504 3606 13560
rect 3662 13504 7528 13560
rect 3601 13502 7528 13504
rect 3601 13499 3667 13502
rect 1853 13426 1919 13429
rect 3785 13426 3851 13429
rect 1853 13424 3851 13426
rect 1853 13368 1858 13424
rect 1914 13368 3790 13424
rect 3846 13368 3851 13424
rect 1853 13366 3851 13368
rect 1853 13363 1919 13366
rect 3785 13363 3851 13366
rect 4061 13426 4127 13429
rect 5349 13426 5415 13429
rect 4061 13424 5415 13426
rect 4061 13368 4066 13424
rect 4122 13368 5354 13424
rect 5410 13368 5415 13424
rect 4061 13366 5415 13368
rect 4061 13363 4127 13366
rect 5349 13363 5415 13366
rect 6085 13426 6151 13429
rect 7189 13426 7255 13429
rect 6085 13424 7255 13426
rect 6085 13368 6090 13424
rect 6146 13368 7194 13424
rect 7250 13368 7255 13424
rect 6085 13366 7255 13368
rect 7468 13426 7528 13502
rect 12617 13560 14780 13562
rect 12617 13504 12622 13560
rect 12678 13504 14554 13560
rect 14610 13504 14780 13560
rect 12617 13502 14780 13504
rect 12617 13499 12683 13502
rect 14549 13499 14615 13502
rect 14774 13500 14780 13502
rect 14844 13500 14850 13564
rect 14917 13562 14983 13565
rect 16297 13562 16363 13565
rect 19200 13562 20000 13592
rect 14917 13560 16363 13562
rect 14917 13504 14922 13560
rect 14978 13504 16302 13560
rect 16358 13504 16363 13560
rect 14917 13502 16363 13504
rect 14917 13499 14983 13502
rect 16297 13499 16363 13502
rect 16944 13502 20000 13562
rect 9305 13426 9371 13429
rect 9489 13428 9555 13429
rect 7468 13424 9371 13426
rect 7468 13368 9310 13424
rect 9366 13368 9371 13424
rect 7468 13366 9371 13368
rect 6085 13363 6151 13366
rect 7189 13363 7255 13366
rect 9305 13363 9371 13366
rect 9438 13364 9444 13428
rect 9508 13426 9555 13428
rect 12249 13426 12315 13429
rect 13537 13426 13603 13429
rect 9508 13424 12082 13426
rect 9550 13368 12082 13424
rect 9508 13366 12082 13368
rect 9508 13364 9555 13366
rect 9489 13363 9555 13364
rect 0 13290 800 13320
rect 2405 13290 2471 13293
rect 0 13288 2471 13290
rect 0 13232 2410 13288
rect 2466 13232 2471 13288
rect 0 13230 2471 13232
rect 0 13200 800 13230
rect 2405 13227 2471 13230
rect 3417 13290 3483 13293
rect 3550 13290 3556 13292
rect 3417 13288 3556 13290
rect 3417 13232 3422 13288
rect 3478 13232 3556 13288
rect 3417 13230 3556 13232
rect 3417 13227 3483 13230
rect 3550 13228 3556 13230
rect 3620 13228 3626 13292
rect 3918 13228 3924 13292
rect 3988 13290 3994 13292
rect 6545 13290 6611 13293
rect 3988 13288 6611 13290
rect 3988 13232 6550 13288
rect 6606 13232 6611 13288
rect 3988 13230 6611 13232
rect 3988 13228 3994 13230
rect 6545 13227 6611 13230
rect 6678 13228 6684 13292
rect 6748 13290 6754 13292
rect 7005 13290 7071 13293
rect 8109 13290 8175 13293
rect 11053 13290 11119 13293
rect 6748 13288 11119 13290
rect 6748 13232 7010 13288
rect 7066 13232 8114 13288
rect 8170 13232 11058 13288
rect 11114 13232 11119 13288
rect 6748 13230 11119 13232
rect 6748 13228 6754 13230
rect 7005 13227 7071 13230
rect 8109 13227 8175 13230
rect 11053 13227 11119 13230
rect 11513 13290 11579 13293
rect 11646 13290 11652 13292
rect 11513 13288 11652 13290
rect 11513 13232 11518 13288
rect 11574 13232 11652 13288
rect 11513 13230 11652 13232
rect 11513 13227 11579 13230
rect 11646 13228 11652 13230
rect 11716 13228 11722 13292
rect 12022 13290 12082 13366
rect 12249 13424 13603 13426
rect 12249 13368 12254 13424
rect 12310 13368 13542 13424
rect 13598 13368 13603 13424
rect 12249 13366 13603 13368
rect 12249 13363 12315 13366
rect 13537 13363 13603 13366
rect 14365 13426 14431 13429
rect 14825 13426 14891 13429
rect 14365 13424 14891 13426
rect 14365 13368 14370 13424
rect 14426 13368 14830 13424
rect 14886 13368 14891 13424
rect 14365 13366 14891 13368
rect 14365 13363 14431 13366
rect 14825 13363 14891 13366
rect 15837 13426 15903 13429
rect 16944 13426 17004 13502
rect 19200 13472 20000 13502
rect 15837 13424 17004 13426
rect 15837 13368 15842 13424
rect 15898 13368 17004 13424
rect 15837 13366 17004 13368
rect 15837 13363 15903 13366
rect 15101 13290 15167 13293
rect 12022 13288 15167 13290
rect 12022 13232 15106 13288
rect 15162 13232 15167 13288
rect 12022 13230 15167 13232
rect 15101 13227 15167 13230
rect 15561 13290 15627 13293
rect 15694 13290 15700 13292
rect 15561 13288 15700 13290
rect 15561 13232 15566 13288
rect 15622 13232 15700 13288
rect 15561 13230 15700 13232
rect 15561 13227 15627 13230
rect 15694 13228 15700 13230
rect 15764 13228 15770 13292
rect 2446 13092 2452 13156
rect 2516 13154 2522 13156
rect 4337 13154 4403 13157
rect 7741 13154 7807 13157
rect 9581 13154 9647 13157
rect 2516 13152 4403 13154
rect 2516 13096 4342 13152
rect 4398 13096 4403 13152
rect 2516 13094 4403 13096
rect 2516 13092 2522 13094
rect 4337 13091 4403 13094
rect 5950 13152 9647 13154
rect 5950 13096 7746 13152
rect 7802 13096 9586 13152
rect 9642 13096 9647 13152
rect 5950 13094 9647 13096
rect 5392 13088 5712 13089
rect 0 13018 800 13048
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5392 13023 5712 13024
rect 1117 13018 1183 13021
rect 0 13016 1183 13018
rect 0 12960 1122 13016
rect 1178 12960 1183 13016
rect 0 12958 1183 12960
rect 0 12928 800 12958
rect 1117 12955 1183 12958
rect 3233 13018 3299 13021
rect 4245 13018 4311 13021
rect 4705 13018 4771 13021
rect 3233 13016 3986 13018
rect 3233 12960 3238 13016
rect 3294 12960 3986 13016
rect 3233 12958 3986 12960
rect 3233 12955 3299 12958
rect 1342 12820 1348 12884
rect 1412 12882 1418 12884
rect 2773 12882 2839 12885
rect 3049 12884 3115 12885
rect 1412 12880 2839 12882
rect 1412 12824 2778 12880
rect 2834 12824 2839 12880
rect 1412 12822 2839 12824
rect 1412 12820 1418 12822
rect 2773 12819 2839 12822
rect 2998 12820 3004 12884
rect 3068 12882 3115 12884
rect 3785 12882 3851 12885
rect 3068 12880 3851 12882
rect 3110 12824 3790 12880
rect 3846 12824 3851 12880
rect 3068 12822 3851 12824
rect 3926 12882 3986 12958
rect 4245 13016 4771 13018
rect 4245 12960 4250 13016
rect 4306 12960 4710 13016
rect 4766 12960 4771 13016
rect 4245 12958 4771 12960
rect 4245 12955 4311 12958
rect 4705 12955 4771 12958
rect 4245 12882 4311 12885
rect 4889 12884 4955 12885
rect 4838 12882 4844 12884
rect 3926 12880 4311 12882
rect 3926 12824 4250 12880
rect 4306 12824 4311 12880
rect 3926 12822 4311 12824
rect 4798 12822 4844 12882
rect 4908 12880 4955 12884
rect 4950 12824 4955 12880
rect 3068 12820 3115 12822
rect 3049 12819 3115 12820
rect 3785 12819 3851 12822
rect 4245 12819 4311 12822
rect 4838 12820 4844 12822
rect 4908 12820 4955 12824
rect 5206 12820 5212 12884
rect 5276 12882 5282 12884
rect 5950 12882 6010 13094
rect 7741 13091 7807 13094
rect 9581 13091 9647 13094
rect 10685 13154 10751 13157
rect 12617 13154 12683 13157
rect 10685 13152 12683 13154
rect 10685 13096 10690 13152
rect 10746 13096 12622 13152
rect 12678 13096 12683 13152
rect 10685 13094 12683 13096
rect 10685 13091 10751 13094
rect 12617 13091 12683 13094
rect 14917 13154 14983 13157
rect 15326 13154 15332 13156
rect 14917 13152 15332 13154
rect 14917 13096 14922 13152
rect 14978 13096 15332 13152
rect 14917 13094 15332 13096
rect 14917 13091 14983 13094
rect 15326 13092 15332 13094
rect 15396 13092 15402 13156
rect 16481 13154 16547 13157
rect 19200 13154 20000 13184
rect 16481 13152 20000 13154
rect 16481 13096 16486 13152
rect 16542 13096 20000 13152
rect 16481 13094 20000 13096
rect 16481 13091 16547 13094
rect 9840 13088 10160 13089
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 9840 13023 10160 13024
rect 14288 13088 14608 13089
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 19200 13064 20000 13094
rect 14288 13023 14608 13024
rect 7005 13018 7071 13021
rect 9673 13018 9739 13021
rect 7005 13016 9739 13018
rect 7005 12960 7010 13016
rect 7066 12960 9678 13016
rect 9734 12960 9739 13016
rect 7005 12958 9739 12960
rect 7005 12955 7071 12958
rect 9673 12955 9739 12958
rect 11329 13018 11395 13021
rect 12065 13018 12131 13021
rect 12893 13018 12959 13021
rect 13302 13018 13308 13020
rect 11329 13016 12266 13018
rect 11329 12960 11334 13016
rect 11390 12960 12070 13016
rect 12126 12960 12266 13016
rect 11329 12958 12266 12960
rect 11329 12955 11395 12958
rect 12065 12955 12131 12958
rect 5276 12822 6010 12882
rect 6177 12882 6243 12885
rect 8845 12882 8911 12885
rect 6177 12880 8911 12882
rect 6177 12824 6182 12880
rect 6238 12824 8850 12880
rect 8906 12824 8911 12880
rect 6177 12822 8911 12824
rect 5276 12820 5282 12822
rect 4889 12819 4955 12820
rect 6177 12819 6243 12822
rect 8845 12819 8911 12822
rect 9029 12882 9095 12885
rect 11605 12882 11671 12885
rect 9029 12880 11671 12882
rect 9029 12824 9034 12880
rect 9090 12824 11610 12880
rect 11666 12824 11671 12880
rect 9029 12822 11671 12824
rect 12206 12882 12266 12958
rect 12893 13016 13308 13018
rect 12893 12960 12898 13016
rect 12954 12960 13308 13016
rect 12893 12958 13308 12960
rect 12893 12955 12959 12958
rect 13302 12956 13308 12958
rect 13372 12956 13378 13020
rect 15377 13018 15443 13021
rect 18505 13018 18571 13021
rect 15377 13016 18571 13018
rect 15377 12960 15382 13016
rect 15438 12960 18510 13016
rect 18566 12960 18571 13016
rect 15377 12958 18571 12960
rect 15377 12955 15443 12958
rect 18505 12955 18571 12958
rect 12709 12882 12775 12885
rect 13629 12884 13695 12885
rect 12206 12880 12775 12882
rect 12206 12824 12714 12880
rect 12770 12824 12775 12880
rect 12206 12822 12775 12824
rect 9029 12819 9095 12822
rect 11605 12819 11671 12822
rect 12709 12819 12775 12822
rect 12934 12820 12940 12884
rect 13004 12882 13010 12884
rect 13486 12882 13492 12884
rect 13004 12822 13492 12882
rect 13004 12820 13010 12822
rect 13486 12820 13492 12822
rect 13556 12820 13562 12884
rect 13629 12880 13676 12884
rect 13740 12882 13746 12884
rect 14089 12882 14155 12885
rect 16982 12882 16988 12884
rect 13629 12824 13634 12880
rect 13629 12820 13676 12824
rect 13740 12822 13786 12882
rect 14089 12880 16988 12882
rect 14089 12824 14094 12880
rect 14150 12824 16988 12880
rect 14089 12822 16988 12824
rect 13740 12820 13746 12822
rect 13629 12819 13695 12820
rect 14089 12819 14155 12822
rect 16982 12820 16988 12822
rect 17052 12820 17058 12884
rect 0 12746 800 12776
rect 2865 12746 2931 12749
rect 5165 12746 5231 12749
rect 0 12744 2931 12746
rect 0 12688 2870 12744
rect 2926 12688 2931 12744
rect 0 12686 2931 12688
rect 0 12656 800 12686
rect 2865 12683 2931 12686
rect 3006 12744 5231 12746
rect 3006 12688 5170 12744
rect 5226 12688 5231 12744
rect 3006 12686 5231 12688
rect 933 12610 999 12613
rect 3006 12610 3066 12686
rect 5165 12683 5231 12686
rect 6085 12746 6151 12749
rect 8886 12746 8892 12748
rect 6085 12744 8892 12746
rect 6085 12688 6090 12744
rect 6146 12688 8892 12744
rect 6085 12686 8892 12688
rect 6085 12683 6151 12686
rect 8886 12684 8892 12686
rect 8956 12684 8962 12748
rect 11421 12746 11487 12749
rect 14273 12746 14339 12749
rect 11421 12744 14339 12746
rect 11421 12688 11426 12744
rect 11482 12688 14278 12744
rect 14334 12688 14339 12744
rect 11421 12686 14339 12688
rect 11421 12683 11487 12686
rect 14273 12683 14339 12686
rect 14457 12746 14523 12749
rect 16205 12746 16271 12749
rect 14457 12744 16271 12746
rect 14457 12688 14462 12744
rect 14518 12688 16210 12744
rect 16266 12688 16271 12744
rect 14457 12686 16271 12688
rect 14457 12683 14523 12686
rect 16205 12683 16271 12686
rect 17677 12746 17743 12749
rect 19200 12746 20000 12776
rect 17677 12744 20000 12746
rect 17677 12688 17682 12744
rect 17738 12688 20000 12744
rect 17677 12686 20000 12688
rect 17677 12683 17743 12686
rect 19200 12656 20000 12686
rect 933 12608 3066 12610
rect 933 12552 938 12608
rect 994 12552 3066 12608
rect 933 12550 3066 12552
rect 3601 12608 3667 12613
rect 3601 12552 3606 12608
rect 3662 12552 3667 12608
rect 933 12547 999 12550
rect 3601 12547 3667 12552
rect 3785 12610 3851 12613
rect 5993 12610 6059 12613
rect 3785 12608 6059 12610
rect 3785 12552 3790 12608
rect 3846 12552 5998 12608
rect 6054 12552 6059 12608
rect 3785 12550 6059 12552
rect 3785 12547 3851 12550
rect 5993 12547 6059 12550
rect 6177 12610 6243 12613
rect 6310 12610 6316 12612
rect 6177 12608 6316 12610
rect 6177 12552 6182 12608
rect 6238 12552 6316 12608
rect 6177 12550 6316 12552
rect 6177 12547 6243 12550
rect 6310 12548 6316 12550
rect 6380 12548 6386 12612
rect 6494 12548 6500 12612
rect 6564 12610 6570 12612
rect 6913 12610 6979 12613
rect 8109 12612 8175 12613
rect 8109 12610 8156 12612
rect 6564 12608 6979 12610
rect 6564 12552 6918 12608
rect 6974 12552 6979 12608
rect 6564 12550 6979 12552
rect 8064 12608 8156 12610
rect 8064 12552 8114 12608
rect 8064 12550 8156 12552
rect 6564 12548 6570 12550
rect 6913 12547 6979 12550
rect 8109 12548 8156 12550
rect 8220 12548 8226 12612
rect 10133 12610 10199 12613
rect 10542 12610 10548 12612
rect 10133 12608 10548 12610
rect 10133 12552 10138 12608
rect 10194 12552 10548 12608
rect 10133 12550 10548 12552
rect 8109 12547 8175 12548
rect 10133 12547 10199 12550
rect 10542 12548 10548 12550
rect 10612 12548 10618 12612
rect 11329 12610 11395 12613
rect 11462 12610 11468 12612
rect 11329 12608 11468 12610
rect 11329 12552 11334 12608
rect 11390 12552 11468 12608
rect 11329 12550 11468 12552
rect 11329 12547 11395 12550
rect 11462 12548 11468 12550
rect 11532 12548 11538 12612
rect 15193 12610 15259 12613
rect 15878 12610 15884 12612
rect 13310 12608 15884 12610
rect 13310 12552 15198 12608
rect 15254 12552 15884 12608
rect 13310 12550 15884 12552
rect 3168 12544 3488 12545
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 12479 3488 12480
rect 1025 12474 1091 12477
rect 2957 12474 3023 12477
rect 1025 12472 3023 12474
rect 1025 12416 1030 12472
rect 1086 12416 2962 12472
rect 3018 12416 3023 12472
rect 1025 12414 3023 12416
rect 3604 12474 3664 12547
rect 7616 12544 7936 12545
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7616 12479 7936 12480
rect 12064 12544 12384 12545
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 12064 12479 12384 12480
rect 3785 12474 3851 12477
rect 3604 12472 3851 12474
rect 3604 12416 3790 12472
rect 3846 12416 3851 12472
rect 3604 12414 3851 12416
rect 1025 12411 1091 12414
rect 2957 12411 3023 12414
rect 3785 12411 3851 12414
rect 4102 12412 4108 12476
rect 4172 12474 4178 12476
rect 6177 12474 6243 12477
rect 6821 12474 6887 12477
rect 4172 12414 6056 12474
rect 4172 12412 4178 12414
rect 0 12338 800 12368
rect 2497 12338 2563 12341
rect 0 12336 2563 12338
rect 0 12280 2502 12336
rect 2558 12280 2563 12336
rect 0 12278 2563 12280
rect 0 12248 800 12278
rect 2497 12275 2563 12278
rect 3417 12338 3483 12341
rect 5625 12338 5691 12341
rect 3417 12336 5691 12338
rect 3417 12280 3422 12336
rect 3478 12280 5630 12336
rect 5686 12280 5691 12336
rect 3417 12278 5691 12280
rect 5996 12338 6056 12414
rect 6177 12472 6887 12474
rect 6177 12416 6182 12472
rect 6238 12416 6826 12472
rect 6882 12416 6887 12472
rect 6177 12414 6887 12416
rect 6177 12411 6243 12414
rect 6821 12411 6887 12414
rect 7005 12476 7071 12477
rect 7005 12472 7052 12476
rect 7116 12474 7122 12476
rect 9765 12474 9831 12477
rect 7005 12416 7010 12472
rect 7005 12412 7052 12416
rect 7116 12414 7162 12474
rect 9765 12472 10610 12474
rect 9765 12416 9770 12472
rect 9826 12416 10610 12472
rect 9765 12414 10610 12416
rect 7116 12412 7122 12414
rect 7005 12411 7071 12412
rect 9765 12411 9831 12414
rect 6545 12338 6611 12341
rect 5996 12336 6611 12338
rect 5996 12280 6550 12336
rect 6606 12280 6611 12336
rect 5996 12278 6611 12280
rect 3417 12275 3483 12278
rect 5625 12275 5691 12278
rect 6545 12275 6611 12278
rect 7230 12276 7236 12340
rect 7300 12338 7306 12340
rect 7373 12338 7439 12341
rect 7300 12336 7439 12338
rect 7300 12280 7378 12336
rect 7434 12280 7439 12336
rect 7300 12278 7439 12280
rect 7300 12276 7306 12278
rect 7373 12275 7439 12278
rect 7557 12338 7623 12341
rect 10317 12338 10383 12341
rect 7557 12336 10383 12338
rect 7557 12280 7562 12336
rect 7618 12280 10322 12336
rect 10378 12280 10383 12336
rect 7557 12278 10383 12280
rect 10550 12338 10610 12414
rect 11094 12412 11100 12476
rect 11164 12474 11170 12476
rect 11237 12474 11303 12477
rect 11164 12472 11303 12474
rect 11164 12416 11242 12472
rect 11298 12416 11303 12472
rect 11164 12414 11303 12416
rect 11164 12412 11170 12414
rect 11237 12411 11303 12414
rect 12709 12474 12775 12477
rect 13310 12474 13370 12550
rect 15193 12547 15259 12550
rect 15878 12548 15884 12550
rect 15948 12548 15954 12612
rect 16512 12544 16832 12545
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 12479 16832 12480
rect 12709 12472 13370 12474
rect 12709 12416 12714 12472
rect 12770 12416 13370 12472
rect 12709 12414 13370 12416
rect 12709 12411 12775 12414
rect 13486 12412 13492 12476
rect 13556 12474 13562 12476
rect 13629 12474 13695 12477
rect 13556 12472 13695 12474
rect 13556 12416 13634 12472
rect 13690 12416 13695 12472
rect 13556 12414 13695 12416
rect 13556 12412 13562 12414
rect 13629 12411 13695 12414
rect 14549 12474 14615 12477
rect 14774 12474 14780 12476
rect 14549 12472 14780 12474
rect 14549 12416 14554 12472
rect 14610 12416 14780 12472
rect 14549 12414 14780 12416
rect 14549 12411 14615 12414
rect 14774 12412 14780 12414
rect 14844 12412 14850 12476
rect 11697 12338 11763 12341
rect 10550 12336 11763 12338
rect 10550 12280 11702 12336
rect 11758 12280 11763 12336
rect 10550 12278 11763 12280
rect 7557 12275 7623 12278
rect 10317 12275 10383 12278
rect 11697 12275 11763 12278
rect 11881 12338 11947 12341
rect 13353 12338 13419 12341
rect 13813 12338 13879 12341
rect 11881 12336 12772 12338
rect 11881 12280 11886 12336
rect 11942 12280 12772 12336
rect 11881 12278 12772 12280
rect 11881 12275 11947 12278
rect 1669 12202 1735 12205
rect 5349 12202 5415 12205
rect 1669 12200 5415 12202
rect 1669 12144 1674 12200
rect 1730 12144 5354 12200
rect 5410 12144 5415 12200
rect 1669 12142 5415 12144
rect 1669 12139 1735 12142
rect 5349 12139 5415 12142
rect 5993 12202 6059 12205
rect 12525 12202 12591 12205
rect 5993 12200 12591 12202
rect 5993 12144 5998 12200
rect 6054 12144 12530 12200
rect 12586 12144 12591 12200
rect 5993 12142 12591 12144
rect 12712 12202 12772 12278
rect 13353 12336 13879 12338
rect 13353 12280 13358 12336
rect 13414 12280 13818 12336
rect 13874 12280 13879 12336
rect 13353 12278 13879 12280
rect 13353 12275 13419 12278
rect 13813 12275 13879 12278
rect 14181 12338 14247 12341
rect 17677 12338 17743 12341
rect 14181 12336 17743 12338
rect 14181 12280 14186 12336
rect 14242 12280 17682 12336
rect 17738 12280 17743 12336
rect 14181 12278 17743 12280
rect 14181 12275 14247 12278
rect 17677 12275 17743 12278
rect 17861 12338 17927 12341
rect 19200 12338 20000 12368
rect 17861 12336 20000 12338
rect 17861 12280 17866 12336
rect 17922 12280 20000 12336
rect 17861 12278 20000 12280
rect 17861 12275 17927 12278
rect 19200 12248 20000 12278
rect 17217 12202 17283 12205
rect 12712 12200 17283 12202
rect 12712 12144 17222 12200
rect 17278 12144 17283 12200
rect 12712 12142 17283 12144
rect 5993 12139 6059 12142
rect 12525 12139 12591 12142
rect 17217 12139 17283 12142
rect 0 12066 800 12096
rect 2773 12066 2839 12069
rect 0 12064 2839 12066
rect 0 12008 2778 12064
rect 2834 12008 2839 12064
rect 0 12006 2839 12008
rect 0 11976 800 12006
rect 2773 12003 2839 12006
rect 3969 12066 4035 12069
rect 4102 12066 4108 12068
rect 3969 12064 4108 12066
rect 3969 12008 3974 12064
rect 4030 12008 4108 12064
rect 3969 12006 4108 12008
rect 3969 12003 4035 12006
rect 4102 12004 4108 12006
rect 4172 12004 4178 12068
rect 5901 12066 5967 12069
rect 7281 12066 7347 12069
rect 8150 12066 8156 12068
rect 5901 12064 8156 12066
rect 5901 12008 5906 12064
rect 5962 12008 7286 12064
rect 7342 12008 8156 12064
rect 5901 12006 8156 12008
rect 5901 12003 5967 12006
rect 7281 12003 7347 12006
rect 8150 12004 8156 12006
rect 8220 12004 8226 12068
rect 10317 12064 10383 12069
rect 10317 12008 10322 12064
rect 10378 12008 10383 12064
rect 10317 12003 10383 12008
rect 10685 12066 10751 12069
rect 11278 12066 11284 12068
rect 10685 12064 11284 12066
rect 10685 12008 10690 12064
rect 10746 12008 11284 12064
rect 10685 12006 11284 12008
rect 10685 12003 10751 12006
rect 11278 12004 11284 12006
rect 11348 12004 11354 12068
rect 12157 12066 12223 12069
rect 13629 12066 13695 12069
rect 13813 12068 13879 12069
rect 13813 12066 13860 12068
rect 12157 12064 13695 12066
rect 12157 12008 12162 12064
rect 12218 12008 13634 12064
rect 13690 12008 13695 12064
rect 12157 12006 13695 12008
rect 13768 12064 13860 12066
rect 13768 12008 13818 12064
rect 13768 12006 13860 12008
rect 12157 12003 12223 12006
rect 13629 12003 13695 12006
rect 13813 12004 13860 12006
rect 13924 12004 13930 12068
rect 15101 12066 15167 12069
rect 16941 12066 17007 12069
rect 15101 12064 17007 12066
rect 15101 12008 15106 12064
rect 15162 12008 16946 12064
rect 17002 12008 17007 12064
rect 15101 12006 17007 12008
rect 13813 12003 13879 12004
rect 15101 12003 15167 12006
rect 16941 12003 17007 12006
rect 5392 12000 5712 12001
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 11935 5712 11936
rect 9840 12000 10160 12001
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9840 11935 10160 11936
rect 2262 11868 2268 11932
rect 2332 11930 2338 11932
rect 4337 11930 4403 11933
rect 2332 11928 4403 11930
rect 2332 11872 4342 11928
rect 4398 11872 4403 11928
rect 2332 11870 4403 11872
rect 2332 11868 2338 11870
rect 4337 11867 4403 11870
rect 7414 11868 7420 11932
rect 7484 11930 7490 11932
rect 8109 11930 8175 11933
rect 7484 11928 8175 11930
rect 7484 11872 8114 11928
rect 8170 11872 8175 11928
rect 7484 11870 8175 11872
rect 10320 11930 10380 12003
rect 14288 12000 14608 12001
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 11935 14608 11936
rect 10961 11930 11027 11933
rect 10320 11928 11027 11930
rect 10320 11872 10966 11928
rect 11022 11872 11027 11928
rect 10320 11870 11027 11872
rect 7484 11868 7490 11870
rect 8109 11867 8175 11870
rect 10961 11867 11027 11870
rect 11973 11930 12039 11933
rect 13169 11930 13235 11933
rect 13486 11930 13492 11932
rect 11973 11928 13492 11930
rect 11973 11872 11978 11928
rect 12034 11872 13174 11928
rect 13230 11872 13492 11928
rect 11973 11870 13492 11872
rect 11973 11867 12039 11870
rect 13169 11867 13235 11870
rect 13486 11868 13492 11870
rect 13556 11868 13562 11932
rect 15653 11930 15719 11933
rect 19200 11930 20000 11960
rect 15653 11928 20000 11930
rect 15653 11872 15658 11928
rect 15714 11872 20000 11928
rect 15653 11870 20000 11872
rect 15653 11867 15719 11870
rect 19200 11840 20000 11870
rect 2129 11794 2195 11797
rect 5901 11794 5967 11797
rect 2129 11792 5967 11794
rect 2129 11736 2134 11792
rect 2190 11736 5906 11792
rect 5962 11736 5967 11792
rect 2129 11734 5967 11736
rect 2129 11731 2195 11734
rect 5901 11731 5967 11734
rect 6862 11732 6868 11796
rect 6932 11794 6938 11796
rect 7281 11794 7347 11797
rect 6932 11792 7347 11794
rect 6932 11736 7286 11792
rect 7342 11736 7347 11792
rect 6932 11734 7347 11736
rect 6932 11732 6938 11734
rect 7281 11731 7347 11734
rect 8017 11794 8083 11797
rect 9622 11794 9628 11796
rect 8017 11792 9628 11794
rect 8017 11736 8022 11792
rect 8078 11736 9628 11792
rect 8017 11734 9628 11736
rect 8017 11731 8083 11734
rect 9622 11732 9628 11734
rect 9692 11732 9698 11796
rect 10317 11794 10383 11797
rect 10726 11794 10732 11796
rect 10317 11792 10732 11794
rect 10317 11736 10322 11792
rect 10378 11736 10732 11792
rect 10317 11734 10732 11736
rect 10317 11731 10383 11734
rect 10726 11732 10732 11734
rect 10796 11732 10802 11796
rect 11830 11732 11836 11796
rect 11900 11794 11906 11796
rect 12341 11794 12407 11797
rect 11900 11792 12407 11794
rect 11900 11736 12346 11792
rect 12402 11736 12407 11792
rect 11900 11734 12407 11736
rect 11900 11732 11906 11734
rect 12341 11731 12407 11734
rect 12566 11732 12572 11796
rect 12636 11794 12642 11796
rect 12801 11794 12867 11797
rect 12636 11792 12867 11794
rect 12636 11736 12806 11792
rect 12862 11736 12867 11792
rect 12636 11734 12867 11736
rect 12636 11732 12642 11734
rect 12801 11731 12867 11734
rect 13077 11794 13143 11797
rect 15142 11794 15148 11796
rect 13077 11792 15148 11794
rect 13077 11736 13082 11792
rect 13138 11736 15148 11792
rect 13077 11734 15148 11736
rect 13077 11731 13143 11734
rect 15142 11732 15148 11734
rect 15212 11732 15218 11796
rect 18597 11794 18663 11797
rect 15288 11792 18663 11794
rect 15288 11736 18602 11792
rect 18658 11736 18663 11792
rect 15288 11734 18663 11736
rect 0 11658 800 11688
rect 2865 11658 2931 11661
rect 0 11656 2931 11658
rect 0 11600 2870 11656
rect 2926 11600 2931 11656
rect 0 11598 2931 11600
rect 0 11568 800 11598
rect 2865 11595 2931 11598
rect 5073 11658 5139 11661
rect 6126 11658 6132 11660
rect 5073 11656 6132 11658
rect 5073 11600 5078 11656
rect 5134 11600 6132 11656
rect 5073 11598 6132 11600
rect 5073 11595 5139 11598
rect 6126 11596 6132 11598
rect 6196 11596 6202 11660
rect 10593 11658 10659 11661
rect 13077 11658 13143 11661
rect 13813 11658 13879 11661
rect 6318 11656 10659 11658
rect 6318 11600 10598 11656
rect 10654 11600 10659 11656
rect 6318 11598 10659 11600
rect 5349 11522 5415 11525
rect 6318 11522 6378 11598
rect 10593 11595 10659 11598
rect 10734 11656 13143 11658
rect 10734 11600 13082 11656
rect 13138 11600 13143 11656
rect 10734 11598 13143 11600
rect 5349 11520 6378 11522
rect 5349 11464 5354 11520
rect 5410 11464 6378 11520
rect 5349 11462 6378 11464
rect 5349 11459 5415 11462
rect 10542 11460 10548 11524
rect 10612 11522 10618 11524
rect 10734 11522 10794 11598
rect 13077 11595 13143 11598
rect 13494 11656 13879 11658
rect 13494 11600 13818 11656
rect 13874 11600 13879 11656
rect 13494 11598 13879 11600
rect 10612 11462 10794 11522
rect 10612 11460 10618 11462
rect 10910 11460 10916 11524
rect 10980 11522 10986 11524
rect 11237 11522 11303 11525
rect 10980 11520 11303 11522
rect 10980 11464 11242 11520
rect 11298 11464 11303 11520
rect 10980 11462 11303 11464
rect 10980 11460 10986 11462
rect 11237 11459 11303 11462
rect 12750 11460 12756 11524
rect 12820 11522 12826 11524
rect 13077 11522 13143 11525
rect 12820 11520 13143 11522
rect 12820 11464 13082 11520
rect 13138 11464 13143 11520
rect 12820 11462 13143 11464
rect 12820 11460 12826 11462
rect 13077 11459 13143 11462
rect 3168 11456 3488 11457
rect 0 11386 800 11416
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 11391 3488 11392
rect 7616 11456 7936 11457
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 11391 7936 11392
rect 12064 11456 12384 11457
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 11391 12384 11392
rect 2957 11386 3023 11389
rect 0 11384 3023 11386
rect 0 11328 2962 11384
rect 3018 11328 3023 11384
rect 0 11326 3023 11328
rect 0 11296 800 11326
rect 2957 11323 3023 11326
rect 5717 11386 5783 11389
rect 12893 11386 12959 11389
rect 13118 11386 13124 11388
rect 5717 11384 7482 11386
rect 5717 11328 5722 11384
rect 5778 11328 7482 11384
rect 5717 11326 7482 11328
rect 5717 11323 5783 11326
rect 1945 11250 2011 11253
rect 1945 11248 5826 11250
rect 1945 11192 1950 11248
rect 2006 11192 5826 11248
rect 1945 11190 5826 11192
rect 1945 11187 2011 11190
rect 2078 11052 2084 11116
rect 2148 11114 2154 11116
rect 4245 11114 4311 11117
rect 2148 11112 4311 11114
rect 2148 11056 4250 11112
rect 4306 11056 4311 11112
rect 2148 11054 4311 11056
rect 5766 11114 5826 11190
rect 5942 11188 5948 11252
rect 6012 11250 6018 11252
rect 6085 11250 6151 11253
rect 6012 11248 6151 11250
rect 6012 11192 6090 11248
rect 6146 11192 6151 11248
rect 6012 11190 6151 11192
rect 7422 11250 7482 11326
rect 12893 11384 13124 11386
rect 12893 11328 12898 11384
rect 12954 11328 13124 11384
rect 12893 11326 13124 11328
rect 12893 11323 12959 11326
rect 13118 11324 13124 11326
rect 13188 11324 13194 11388
rect 13494 11386 13554 11598
rect 13813 11595 13879 11598
rect 13997 11658 14063 11661
rect 15288 11658 15348 11734
rect 18597 11731 18663 11734
rect 17769 11658 17835 11661
rect 19200 11658 20000 11688
rect 13997 11656 15348 11658
rect 13997 11600 14002 11656
rect 14058 11600 15348 11656
rect 13997 11598 15348 11600
rect 16254 11598 17648 11658
rect 13997 11595 14063 11598
rect 13721 11522 13787 11525
rect 14958 11522 14964 11524
rect 13721 11520 14964 11522
rect 13721 11464 13726 11520
rect 13782 11464 14964 11520
rect 13721 11462 14964 11464
rect 13721 11459 13787 11462
rect 14958 11460 14964 11462
rect 15028 11522 15034 11524
rect 15285 11522 15351 11525
rect 15028 11520 15351 11522
rect 15028 11464 15290 11520
rect 15346 11464 15351 11520
rect 15028 11462 15351 11464
rect 15028 11460 15034 11462
rect 15285 11459 15351 11462
rect 15469 11522 15535 11525
rect 15837 11522 15903 11525
rect 15469 11520 15903 11522
rect 15469 11464 15474 11520
rect 15530 11464 15842 11520
rect 15898 11464 15903 11520
rect 15469 11462 15903 11464
rect 15469 11459 15535 11462
rect 15837 11459 15903 11462
rect 14089 11386 14155 11389
rect 13494 11384 14155 11386
rect 13494 11328 14094 11384
rect 14150 11328 14155 11384
rect 13494 11326 14155 11328
rect 14089 11323 14155 11326
rect 14365 11386 14431 11389
rect 16254 11386 16314 11598
rect 17588 11522 17648 11598
rect 17769 11656 20000 11658
rect 17769 11600 17774 11656
rect 17830 11600 20000 11656
rect 17769 11598 20000 11600
rect 17769 11595 17835 11598
rect 19200 11568 20000 11598
rect 18689 11522 18755 11525
rect 17588 11520 18755 11522
rect 17588 11464 18694 11520
rect 18750 11464 18755 11520
rect 17588 11462 18755 11464
rect 18689 11459 18755 11462
rect 16512 11456 16832 11457
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 11391 16832 11392
rect 17953 11386 18019 11389
rect 14365 11384 16314 11386
rect 14365 11328 14370 11384
rect 14426 11328 16314 11384
rect 14365 11326 16314 11328
rect 16944 11384 18019 11386
rect 16944 11328 17958 11384
rect 18014 11328 18019 11384
rect 16944 11326 18019 11328
rect 14365 11323 14431 11326
rect 9438 11250 9444 11252
rect 7422 11190 9444 11250
rect 6012 11188 6018 11190
rect 6085 11187 6151 11190
rect 9438 11188 9444 11190
rect 9508 11188 9514 11252
rect 10961 11250 11027 11253
rect 12249 11250 12315 11253
rect 10961 11248 12315 11250
rect 10961 11192 10966 11248
rect 11022 11192 12254 11248
rect 12310 11192 12315 11248
rect 10961 11190 12315 11192
rect 10961 11187 11027 11190
rect 12249 11187 12315 11190
rect 12985 11250 13051 11253
rect 16944 11250 17004 11326
rect 17953 11323 18019 11326
rect 12985 11248 17004 11250
rect 12985 11192 12990 11248
rect 13046 11192 17004 11248
rect 12985 11190 17004 11192
rect 17677 11250 17743 11253
rect 19200 11250 20000 11280
rect 17677 11248 20000 11250
rect 17677 11192 17682 11248
rect 17738 11192 20000 11248
rect 17677 11190 20000 11192
rect 12985 11187 13051 11190
rect 17677 11187 17743 11190
rect 19200 11160 20000 11190
rect 6545 11114 6611 11117
rect 8518 11114 8524 11116
rect 5766 11054 6378 11114
rect 2148 11052 2154 11054
rect 4245 11051 4311 11054
rect 0 10978 800 11008
rect 2957 10978 3023 10981
rect 4981 10978 5047 10981
rect 0 10976 5047 10978
rect 0 10920 2962 10976
rect 3018 10920 4986 10976
rect 5042 10920 5047 10976
rect 0 10918 5047 10920
rect 6318 10978 6378 11054
rect 6545 11112 8524 11114
rect 6545 11056 6550 11112
rect 6606 11056 8524 11112
rect 6545 11054 8524 11056
rect 6545 11051 6611 11054
rect 8518 11052 8524 11054
rect 8588 11052 8594 11116
rect 9305 11114 9371 11117
rect 10777 11114 10843 11117
rect 8664 11112 10843 11114
rect 8664 11056 9310 11112
rect 9366 11056 10782 11112
rect 10838 11056 10843 11112
rect 8664 11054 10843 11056
rect 8385 10978 8451 10981
rect 8664 10978 8724 11054
rect 9305 11051 9371 11054
rect 10777 11051 10843 11054
rect 11646 11052 11652 11116
rect 11716 11114 11722 11116
rect 12249 11114 12315 11117
rect 14825 11114 14891 11117
rect 11716 11112 12315 11114
rect 11716 11056 12254 11112
rect 12310 11056 12315 11112
rect 11716 11054 12315 11056
rect 11716 11052 11722 11054
rect 12249 11051 12315 11054
rect 12390 11112 14891 11114
rect 12390 11056 14830 11112
rect 14886 11056 14891 11112
rect 12390 11054 14891 11056
rect 6318 10976 8724 10978
rect 6318 10920 8390 10976
rect 8446 10920 8724 10976
rect 6318 10918 8724 10920
rect 11053 10978 11119 10981
rect 12390 10978 12450 11054
rect 14825 11051 14891 11054
rect 11053 10976 12450 10978
rect 11053 10920 11058 10976
rect 11114 10920 12450 10976
rect 11053 10918 12450 10920
rect 15653 10978 15719 10981
rect 17309 10978 17375 10981
rect 15653 10976 17375 10978
rect 15653 10920 15658 10976
rect 15714 10920 17314 10976
rect 17370 10920 17375 10976
rect 15653 10918 17375 10920
rect 0 10888 800 10918
rect 2957 10915 3023 10918
rect 4981 10915 5047 10918
rect 8385 10915 8451 10918
rect 11053 10915 11119 10918
rect 15653 10915 15719 10918
rect 17309 10915 17375 10918
rect 5392 10912 5712 10913
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 10847 5712 10848
rect 9840 10912 10160 10913
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 10847 10160 10848
rect 14288 10912 14608 10913
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 10847 14608 10848
rect 2630 10780 2636 10844
rect 2700 10842 2706 10844
rect 4061 10842 4127 10845
rect 2700 10840 4127 10842
rect 2700 10784 4066 10840
rect 4122 10784 4127 10840
rect 2700 10782 4127 10784
rect 2700 10780 2706 10782
rect 4061 10779 4127 10782
rect 5901 10842 5967 10845
rect 6637 10842 6703 10845
rect 8109 10842 8175 10845
rect 5901 10840 8175 10842
rect 5901 10784 5906 10840
rect 5962 10784 6642 10840
rect 6698 10784 8114 10840
rect 8170 10784 8175 10840
rect 5901 10782 8175 10784
rect 5901 10779 5967 10782
rect 6637 10779 6703 10782
rect 8109 10779 8175 10782
rect 12157 10842 12223 10845
rect 13813 10842 13879 10845
rect 12157 10840 13879 10842
rect 12157 10784 12162 10840
rect 12218 10784 13818 10840
rect 13874 10784 13879 10840
rect 12157 10782 13879 10784
rect 12157 10779 12223 10782
rect 13813 10779 13879 10782
rect 17217 10842 17283 10845
rect 19200 10842 20000 10872
rect 17217 10840 20000 10842
rect 17217 10784 17222 10840
rect 17278 10784 20000 10840
rect 17217 10782 20000 10784
rect 17217 10779 17283 10782
rect 19200 10752 20000 10782
rect 0 10706 800 10736
rect 2221 10706 2287 10709
rect 0 10704 2287 10706
rect 0 10648 2226 10704
rect 2282 10648 2287 10704
rect 0 10646 2287 10648
rect 0 10616 800 10646
rect 2221 10643 2287 10646
rect 2814 10644 2820 10708
rect 2884 10706 2890 10708
rect 3550 10706 3556 10708
rect 2884 10646 3556 10706
rect 2884 10644 2890 10646
rect 3550 10644 3556 10646
rect 3620 10644 3626 10708
rect 3785 10706 3851 10709
rect 8661 10706 8727 10709
rect 3785 10704 8727 10706
rect 3785 10648 3790 10704
rect 3846 10648 8666 10704
rect 8722 10648 8727 10704
rect 3785 10646 8727 10648
rect 3785 10643 3851 10646
rect 8661 10643 8727 10646
rect 9857 10706 9923 10709
rect 16297 10706 16363 10709
rect 9857 10704 16363 10706
rect 9857 10648 9862 10704
rect 9918 10648 16302 10704
rect 16358 10648 16363 10704
rect 9857 10646 16363 10648
rect 9857 10643 9923 10646
rect 16297 10643 16363 10646
rect 2221 10570 2287 10573
rect 7230 10570 7236 10572
rect 2221 10568 7236 10570
rect 2221 10512 2226 10568
rect 2282 10512 7236 10568
rect 2221 10510 7236 10512
rect 2221 10507 2287 10510
rect 7230 10508 7236 10510
rect 7300 10508 7306 10572
rect 8385 10570 8451 10573
rect 11094 10570 11100 10572
rect 8385 10568 11100 10570
rect 8385 10512 8390 10568
rect 8446 10512 11100 10568
rect 8385 10510 11100 10512
rect 8385 10507 8451 10510
rect 11094 10508 11100 10510
rect 11164 10508 11170 10572
rect 11646 10508 11652 10572
rect 11716 10570 11722 10572
rect 12157 10570 12223 10573
rect 11716 10568 12223 10570
rect 11716 10512 12162 10568
rect 12218 10512 12223 10568
rect 11716 10510 12223 10512
rect 11716 10508 11722 10510
rect 12157 10507 12223 10510
rect 13302 10508 13308 10572
rect 13372 10570 13378 10572
rect 13372 10510 17004 10570
rect 13372 10508 13378 10510
rect 0 10434 800 10464
rect 2773 10434 2839 10437
rect 0 10432 2839 10434
rect 0 10376 2778 10432
rect 2834 10376 2839 10432
rect 0 10374 2839 10376
rect 0 10344 800 10374
rect 2773 10371 2839 10374
rect 3601 10434 3667 10437
rect 7373 10434 7439 10437
rect 3601 10432 7439 10434
rect 3601 10376 3606 10432
rect 3662 10376 7378 10432
rect 7434 10376 7439 10432
rect 3601 10374 7439 10376
rect 3601 10371 3667 10374
rect 7373 10371 7439 10374
rect 10409 10434 10475 10437
rect 11145 10434 11211 10437
rect 11513 10434 11579 10437
rect 10409 10432 10978 10434
rect 10409 10376 10414 10432
rect 10470 10376 10978 10432
rect 10409 10374 10978 10376
rect 10409 10371 10475 10374
rect 3168 10368 3488 10369
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 10303 3488 10304
rect 7616 10368 7936 10369
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7616 10303 7936 10304
rect 3601 10298 3667 10301
rect 6545 10298 6611 10301
rect 3601 10296 6611 10298
rect 3601 10240 3606 10296
rect 3662 10240 6550 10296
rect 6606 10240 6611 10296
rect 3601 10238 6611 10240
rect 3601 10235 3667 10238
rect 6545 10235 6611 10238
rect 7281 10298 7347 10301
rect 7414 10298 7420 10300
rect 7281 10296 7420 10298
rect 7281 10240 7286 10296
rect 7342 10240 7420 10296
rect 7281 10238 7420 10240
rect 7281 10235 7347 10238
rect 7414 10236 7420 10238
rect 7484 10236 7490 10300
rect 8937 10298 9003 10301
rect 9121 10298 9187 10301
rect 8937 10296 9187 10298
rect 8937 10240 8942 10296
rect 8998 10240 9126 10296
rect 9182 10240 9187 10296
rect 8937 10238 9187 10240
rect 8937 10235 9003 10238
rect 9121 10235 9187 10238
rect 606 10134 612 10198
rect 676 10196 682 10198
rect 676 10162 996 10196
rect 6913 10162 6979 10165
rect 676 10160 6979 10162
rect 676 10136 6918 10160
rect 676 10134 682 10136
rect 936 10104 6918 10136
rect 6974 10104 6979 10160
rect 936 10102 6979 10104
rect 6913 10099 6979 10102
rect 7189 10162 7255 10165
rect 10685 10162 10751 10165
rect 7189 10160 10751 10162
rect 7189 10104 7194 10160
rect 7250 10104 10690 10160
rect 10746 10104 10751 10160
rect 7189 10102 10751 10104
rect 7189 10099 7255 10102
rect 10685 10099 10751 10102
rect 0 10026 800 10056
rect 1485 10026 1551 10029
rect 1945 10026 2011 10029
rect 0 10024 2011 10026
rect 0 9968 1490 10024
rect 1546 9968 1950 10024
rect 2006 9968 2011 10024
rect 0 9966 2011 9968
rect 0 9936 800 9966
rect 1485 9963 1551 9966
rect 1945 9963 2011 9966
rect 4153 10026 4219 10029
rect 8753 10026 8819 10029
rect 9857 10026 9923 10029
rect 4153 10024 8819 10026
rect 4153 9968 4158 10024
rect 4214 9968 8758 10024
rect 8814 9968 8819 10024
rect 4153 9966 8819 9968
rect 4153 9963 4219 9966
rect 8753 9963 8819 9966
rect 9630 10024 9923 10026
rect 9630 9968 9862 10024
rect 9918 9968 9923 10024
rect 9630 9966 9923 9968
rect 6678 9828 6684 9892
rect 6748 9890 6754 9892
rect 6821 9890 6887 9893
rect 6748 9888 6887 9890
rect 6748 9832 6826 9888
rect 6882 9832 6887 9888
rect 6748 9830 6887 9832
rect 6748 9828 6754 9830
rect 6821 9827 6887 9830
rect 7414 9828 7420 9892
rect 7484 9890 7490 9892
rect 7649 9890 7715 9893
rect 9630 9890 9690 9966
rect 9857 9963 9923 9966
rect 10225 10026 10291 10029
rect 10918 10026 10978 10374
rect 11145 10432 11579 10434
rect 11145 10376 11150 10432
rect 11206 10376 11518 10432
rect 11574 10376 11579 10432
rect 11145 10374 11579 10376
rect 11145 10371 11211 10374
rect 11513 10371 11579 10374
rect 14365 10434 14431 10437
rect 16062 10434 16068 10436
rect 14365 10432 16068 10434
rect 14365 10376 14370 10432
rect 14426 10376 16068 10432
rect 14365 10374 16068 10376
rect 14365 10371 14431 10374
rect 16062 10372 16068 10374
rect 16132 10372 16138 10436
rect 16944 10434 17004 10510
rect 19200 10434 20000 10464
rect 16944 10374 20000 10434
rect 12064 10368 12384 10369
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 12064 10303 12384 10304
rect 16512 10368 16832 10369
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 19200 10344 20000 10374
rect 16512 10303 16832 10304
rect 11513 10300 11579 10301
rect 11462 10236 11468 10300
rect 11532 10298 11579 10300
rect 12617 10298 12683 10301
rect 14549 10298 14615 10301
rect 11532 10296 11624 10298
rect 11574 10240 11624 10296
rect 11532 10238 11624 10240
rect 12617 10296 14615 10298
rect 12617 10240 12622 10296
rect 12678 10240 14554 10296
rect 14610 10240 14615 10296
rect 12617 10238 14615 10240
rect 11532 10236 11579 10238
rect 11513 10235 11579 10236
rect 12617 10235 12683 10238
rect 14549 10235 14615 10238
rect 11278 10100 11284 10164
rect 11348 10162 11354 10164
rect 14641 10162 14707 10165
rect 11348 10160 14707 10162
rect 11348 10104 14646 10160
rect 14702 10104 14707 10160
rect 11348 10102 14707 10104
rect 11348 10100 11354 10102
rect 14641 10099 14707 10102
rect 15326 10100 15332 10164
rect 15396 10162 15402 10164
rect 16389 10162 16455 10165
rect 15396 10160 16455 10162
rect 15396 10104 16394 10160
rect 16450 10104 16455 10160
rect 15396 10102 16455 10104
rect 15396 10100 15402 10102
rect 16389 10099 16455 10102
rect 17493 10162 17559 10165
rect 17493 10160 18706 10162
rect 17493 10104 17498 10160
rect 17554 10104 18706 10160
rect 17493 10102 18706 10104
rect 17493 10099 17559 10102
rect 11329 10026 11395 10029
rect 10225 10024 10426 10026
rect 10225 9968 10230 10024
rect 10286 9968 10426 10024
rect 10225 9966 10426 9968
rect 10918 10024 11395 10026
rect 10918 9968 11334 10024
rect 11390 9968 11395 10024
rect 10918 9966 11395 9968
rect 10225 9963 10291 9966
rect 7484 9828 7528 9890
rect 5392 9824 5712 9825
rect 0 9754 800 9784
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 9759 5712 9760
rect 2221 9754 2287 9757
rect 0 9752 2287 9754
rect 0 9696 2226 9752
rect 2282 9696 2287 9752
rect 0 9694 2287 9696
rect 0 9664 800 9694
rect 2221 9691 2287 9694
rect 3877 9754 3943 9757
rect 4286 9754 4292 9756
rect 3877 9752 4292 9754
rect 3877 9696 3882 9752
rect 3938 9696 4292 9752
rect 3877 9694 4292 9696
rect 3877 9691 3943 9694
rect 4286 9692 4292 9694
rect 4356 9692 4362 9756
rect 6494 9754 6500 9756
rect 5996 9694 6500 9754
rect 1945 9618 2011 9621
rect 5996 9618 6056 9694
rect 6494 9692 6500 9694
rect 6564 9754 6570 9756
rect 6913 9754 6979 9757
rect 6564 9752 6979 9754
rect 6564 9696 6918 9752
rect 6974 9696 6979 9752
rect 6564 9694 6979 9696
rect 7468 9754 7528 9828
rect 7649 9888 9690 9890
rect 7649 9832 7654 9888
rect 7710 9832 9690 9888
rect 7649 9830 9690 9832
rect 7649 9827 7715 9830
rect 9840 9824 10160 9825
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 9759 10160 9760
rect 7741 9754 7807 9757
rect 7468 9752 7807 9754
rect 7468 9696 7746 9752
rect 7802 9696 7807 9752
rect 7468 9694 7807 9696
rect 6564 9692 6570 9694
rect 6913 9691 6979 9694
rect 7741 9691 7807 9694
rect 7925 9754 7991 9757
rect 8150 9754 8156 9756
rect 7925 9752 8156 9754
rect 7925 9696 7930 9752
rect 7986 9696 8156 9752
rect 7925 9694 8156 9696
rect 7925 9691 7991 9694
rect 8150 9692 8156 9694
rect 8220 9692 8226 9756
rect 10225 9754 10291 9757
rect 10366 9754 10426 9966
rect 11329 9963 11395 9966
rect 11605 10026 11671 10029
rect 18505 10026 18571 10029
rect 11605 10024 18571 10026
rect 11605 9968 11610 10024
rect 11666 9968 18510 10024
rect 18566 9968 18571 10024
rect 11605 9966 18571 9968
rect 18646 10026 18706 10102
rect 19200 10026 20000 10056
rect 18646 9966 20000 10026
rect 11605 9963 11671 9966
rect 18505 9963 18571 9966
rect 19200 9936 20000 9966
rect 11646 9828 11652 9892
rect 11716 9890 11722 9892
rect 12433 9890 12499 9893
rect 11716 9888 12499 9890
rect 11716 9832 12438 9888
rect 12494 9832 12499 9888
rect 11716 9830 12499 9832
rect 11716 9828 11722 9830
rect 12433 9827 12499 9830
rect 14733 9890 14799 9893
rect 17953 9890 18019 9893
rect 14733 9888 18019 9890
rect 14733 9832 14738 9888
rect 14794 9832 17958 9888
rect 18014 9832 18019 9888
rect 14733 9830 18019 9832
rect 14733 9827 14799 9830
rect 17953 9827 18019 9830
rect 14288 9824 14608 9825
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14288 9759 14608 9760
rect 10225 9752 10426 9754
rect 10225 9696 10230 9752
rect 10286 9696 10426 9752
rect 10225 9694 10426 9696
rect 10501 9754 10567 9757
rect 11462 9754 11468 9756
rect 10501 9752 11468 9754
rect 10501 9696 10506 9752
rect 10562 9696 11468 9752
rect 10501 9694 11468 9696
rect 10225 9691 10291 9694
rect 10501 9691 10567 9694
rect 11462 9692 11468 9694
rect 11532 9692 11538 9756
rect 11605 9754 11671 9757
rect 11830 9754 11836 9756
rect 11605 9752 11836 9754
rect 11605 9696 11610 9752
rect 11666 9696 11836 9752
rect 11605 9694 11836 9696
rect 11605 9691 11671 9694
rect 11830 9692 11836 9694
rect 11900 9692 11906 9756
rect 16062 9692 16068 9756
rect 16132 9754 16138 9756
rect 16757 9754 16823 9757
rect 16132 9752 16823 9754
rect 16132 9696 16762 9752
rect 16818 9696 16823 9752
rect 16132 9694 16823 9696
rect 16132 9692 16138 9694
rect 16757 9691 16823 9694
rect 18505 9754 18571 9757
rect 19200 9754 20000 9784
rect 18505 9752 20000 9754
rect 18505 9696 18510 9752
rect 18566 9696 20000 9752
rect 18505 9694 20000 9696
rect 18505 9691 18571 9694
rect 19200 9664 20000 9694
rect 1945 9616 6056 9618
rect 1945 9560 1950 9616
rect 2006 9560 6056 9616
rect 1945 9558 6056 9560
rect 1945 9555 2011 9558
rect 6126 9556 6132 9620
rect 6196 9618 6202 9620
rect 6269 9618 6335 9621
rect 6196 9616 6335 9618
rect 6196 9560 6274 9616
rect 6330 9560 6335 9616
rect 6196 9558 6335 9560
rect 6196 9556 6202 9558
rect 6269 9555 6335 9558
rect 6453 9618 6519 9621
rect 10777 9618 10843 9621
rect 17033 9618 17099 9621
rect 6453 9616 17099 9618
rect 6453 9560 6458 9616
rect 6514 9560 10782 9616
rect 10838 9560 17038 9616
rect 17094 9560 17099 9616
rect 6453 9558 17099 9560
rect 6453 9555 6519 9558
rect 10777 9555 10843 9558
rect 17033 9555 17099 9558
rect 1301 9482 1367 9485
rect 7373 9482 7439 9485
rect 1301 9480 7439 9482
rect 1301 9424 1306 9480
rect 1362 9424 7378 9480
rect 7434 9424 7439 9480
rect 1301 9422 7439 9424
rect 1301 9419 1367 9422
rect 7373 9419 7439 9422
rect 7557 9482 7623 9485
rect 11697 9482 11763 9485
rect 7557 9480 11763 9482
rect 7557 9424 7562 9480
rect 7618 9424 11702 9480
rect 11758 9424 11763 9480
rect 7557 9422 11763 9424
rect 7557 9419 7623 9422
rect 11697 9419 11763 9422
rect 12433 9482 12499 9485
rect 14038 9482 14044 9484
rect 12433 9480 14044 9482
rect 12433 9424 12438 9480
rect 12494 9424 14044 9480
rect 12433 9422 14044 9424
rect 12433 9419 12499 9422
rect 14038 9420 14044 9422
rect 14108 9420 14114 9484
rect 0 9346 800 9376
rect 1853 9346 1919 9349
rect 0 9344 1919 9346
rect 0 9288 1858 9344
rect 1914 9288 1919 9344
rect 0 9286 1919 9288
rect 0 9256 800 9286
rect 1853 9283 1919 9286
rect 4102 9284 4108 9348
rect 4172 9346 4178 9348
rect 5073 9346 5139 9349
rect 7465 9346 7531 9349
rect 4172 9344 7531 9346
rect 4172 9288 5078 9344
rect 5134 9288 7470 9344
rect 7526 9288 7531 9344
rect 4172 9286 7531 9288
rect 4172 9284 4178 9286
rect 5073 9283 5139 9286
rect 7465 9283 7531 9286
rect 12801 9346 12867 9349
rect 15653 9346 15719 9349
rect 12801 9344 15719 9346
rect 12801 9288 12806 9344
rect 12862 9288 15658 9344
rect 15714 9288 15719 9344
rect 12801 9286 15719 9288
rect 12801 9283 12867 9286
rect 15653 9283 15719 9286
rect 18229 9344 18295 9349
rect 18229 9288 18234 9344
rect 18290 9288 18295 9344
rect 18229 9283 18295 9288
rect 18413 9346 18479 9349
rect 19200 9346 20000 9376
rect 18413 9344 20000 9346
rect 18413 9288 18418 9344
rect 18474 9288 20000 9344
rect 18413 9286 20000 9288
rect 18413 9283 18479 9286
rect 3168 9280 3488 9281
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 9215 3488 9216
rect 7616 9280 7936 9281
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7616 9215 7936 9216
rect 12064 9280 12384 9281
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 12064 9215 12384 9216
rect 16512 9280 16832 9281
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 9215 16832 9216
rect 10685 9212 10751 9213
rect 7046 9210 7052 9212
rect 3558 9150 7052 9210
rect 0 9074 800 9104
rect 1669 9074 1735 9077
rect 3558 9074 3618 9150
rect 7046 9148 7052 9150
rect 7116 9148 7122 9212
rect 10685 9210 10732 9212
rect 10640 9208 10732 9210
rect 10640 9152 10690 9208
rect 10640 9150 10732 9152
rect 10685 9148 10732 9150
rect 10796 9148 10802 9212
rect 12525 9210 12591 9213
rect 15377 9210 15443 9213
rect 12525 9208 15443 9210
rect 12525 9152 12530 9208
rect 12586 9152 15382 9208
rect 15438 9152 15443 9208
rect 12525 9150 15443 9152
rect 10685 9147 10751 9148
rect 12525 9147 12591 9150
rect 15377 9147 15443 9150
rect 0 9014 1594 9074
rect 0 8984 800 9014
rect 1534 8938 1594 9014
rect 1669 9072 3618 9074
rect 1669 9016 1674 9072
rect 1730 9016 3618 9072
rect 1669 9014 3618 9016
rect 3693 9076 3759 9077
rect 3693 9072 3740 9076
rect 3804 9074 3810 9076
rect 3969 9074 4035 9077
rect 8569 9074 8635 9077
rect 3693 9016 3698 9072
rect 1669 9011 1735 9014
rect 3693 9012 3740 9016
rect 3804 9014 3850 9074
rect 3969 9072 8635 9074
rect 3969 9016 3974 9072
rect 4030 9016 8574 9072
rect 8630 9016 8635 9072
rect 3969 9014 8635 9016
rect 3804 9012 3810 9014
rect 3693 9011 3759 9012
rect 3969 9011 4035 9014
rect 8569 9011 8635 9014
rect 9673 9074 9739 9077
rect 10317 9074 10383 9077
rect 9673 9072 10383 9074
rect 9673 9016 9678 9072
rect 9734 9016 10322 9072
rect 10378 9016 10383 9072
rect 9673 9014 10383 9016
rect 9673 9011 9739 9014
rect 10317 9011 10383 9014
rect 11237 9074 11303 9077
rect 12065 9074 12131 9077
rect 12934 9074 12940 9076
rect 11237 9072 12940 9074
rect 11237 9016 11242 9072
rect 11298 9016 12070 9072
rect 12126 9016 12940 9072
rect 11237 9014 12940 9016
rect 11237 9011 11303 9014
rect 12065 9011 12131 9014
rect 12934 9012 12940 9014
rect 13004 9012 13010 9076
rect 13486 9012 13492 9076
rect 13556 9074 13562 9076
rect 18232 9074 18292 9283
rect 19200 9256 20000 9286
rect 13556 9014 18292 9074
rect 13556 9012 13562 9014
rect 2497 8938 2563 8941
rect 1534 8936 2563 8938
rect 1534 8880 2502 8936
rect 2558 8880 2563 8936
rect 1534 8878 2563 8880
rect 2497 8875 2563 8878
rect 2814 8876 2820 8940
rect 2884 8938 2890 8940
rect 3141 8938 3207 8941
rect 2884 8936 3207 8938
rect 2884 8880 3146 8936
rect 3202 8880 3207 8936
rect 2884 8878 3207 8880
rect 2884 8876 2890 8878
rect 3141 8875 3207 8878
rect 3693 8938 3759 8941
rect 6862 8938 6868 8940
rect 3693 8936 6868 8938
rect 3693 8880 3698 8936
rect 3754 8880 6868 8936
rect 3693 8878 6868 8880
rect 3693 8875 3759 8878
rect 6862 8876 6868 8878
rect 6932 8876 6938 8940
rect 7414 8876 7420 8940
rect 7484 8938 7490 8940
rect 7741 8938 7807 8941
rect 7484 8936 7807 8938
rect 7484 8880 7746 8936
rect 7802 8880 7807 8936
rect 7484 8878 7807 8880
rect 7484 8876 7490 8878
rect 7741 8875 7807 8878
rect 8109 8938 8175 8941
rect 13486 8938 13492 8940
rect 8109 8936 13492 8938
rect 8109 8880 8114 8936
rect 8170 8880 13492 8936
rect 8109 8878 13492 8880
rect 8109 8875 8175 8878
rect 13486 8876 13492 8878
rect 13556 8876 13562 8940
rect 15285 8938 15351 8941
rect 13678 8936 15351 8938
rect 13678 8880 15290 8936
rect 15346 8880 15351 8936
rect 13678 8878 15351 8880
rect 0 8802 800 8832
rect 1393 8802 1459 8805
rect 0 8800 1459 8802
rect 0 8744 1398 8800
rect 1454 8744 1459 8800
rect 0 8742 1459 8744
rect 0 8712 800 8742
rect 1393 8739 1459 8742
rect 1853 8802 1919 8805
rect 4521 8802 4587 8805
rect 1853 8800 4587 8802
rect 1853 8744 1858 8800
rect 1914 8744 4526 8800
rect 4582 8744 4587 8800
rect 1853 8742 4587 8744
rect 1853 8739 1919 8742
rect 4521 8739 4587 8742
rect 7465 8802 7531 8805
rect 8109 8802 8175 8805
rect 7465 8800 8175 8802
rect 7465 8744 7470 8800
rect 7526 8744 8114 8800
rect 8170 8744 8175 8800
rect 7465 8742 8175 8744
rect 7465 8739 7531 8742
rect 8109 8739 8175 8742
rect 10961 8802 11027 8805
rect 12433 8802 12499 8805
rect 13678 8802 13738 8878
rect 15285 8875 15351 8878
rect 18689 8938 18755 8941
rect 19200 8938 20000 8968
rect 18689 8936 20000 8938
rect 18689 8880 18694 8936
rect 18750 8880 20000 8936
rect 18689 8878 20000 8880
rect 18689 8875 18755 8878
rect 19200 8848 20000 8878
rect 10961 8800 13738 8802
rect 10961 8744 10966 8800
rect 11022 8744 12438 8800
rect 12494 8744 13738 8800
rect 10961 8742 13738 8744
rect 10961 8739 11027 8742
rect 12433 8739 12499 8742
rect 5392 8736 5712 8737
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5392 8671 5712 8672
rect 9840 8736 10160 8737
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 8671 10160 8672
rect 14288 8736 14608 8737
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14288 8671 14608 8672
rect 5257 8668 5323 8669
rect 5206 8666 5212 8668
rect 2730 8606 5212 8666
rect 5276 8664 5323 8668
rect 5318 8608 5323 8664
rect 2221 8530 2287 8533
rect 2730 8530 2790 8606
rect 5206 8604 5212 8606
rect 5276 8604 5323 8608
rect 5257 8603 5323 8604
rect 7281 8666 7347 8669
rect 7557 8666 7623 8669
rect 7281 8664 7623 8666
rect 7281 8608 7286 8664
rect 7342 8608 7562 8664
rect 7618 8608 7623 8664
rect 7281 8606 7623 8608
rect 7281 8603 7347 8606
rect 7557 8603 7623 8606
rect 2221 8528 2790 8530
rect 2221 8472 2226 8528
rect 2282 8472 2790 8528
rect 2221 8470 2790 8472
rect 2957 8528 3023 8533
rect 2957 8472 2962 8528
rect 3018 8472 3023 8528
rect 2221 8467 2287 8470
rect 2957 8467 3023 8472
rect 3233 8530 3299 8533
rect 8293 8530 8359 8533
rect 3233 8528 8359 8530
rect 3233 8472 3238 8528
rect 3294 8472 8298 8528
rect 8354 8472 8359 8528
rect 3233 8470 8359 8472
rect 3233 8467 3299 8470
rect 8293 8467 8359 8470
rect 9581 8530 9647 8533
rect 18045 8530 18111 8533
rect 19200 8530 20000 8560
rect 9581 8528 17418 8530
rect 9581 8472 9586 8528
rect 9642 8472 17418 8528
rect 9581 8470 17418 8472
rect 9581 8467 9647 8470
rect 0 8394 800 8424
rect 2960 8394 3020 8467
rect 3969 8396 4035 8397
rect 3734 8394 3740 8396
rect 0 8334 3020 8394
rect 0 8304 800 8334
rect 3696 8332 3740 8394
rect 3804 8332 3810 8396
rect 3918 8332 3924 8396
rect 3988 8394 4035 8396
rect 5257 8394 5323 8397
rect 11881 8396 11947 8397
rect 8150 8394 8156 8396
rect 3988 8392 4080 8394
rect 4030 8336 4080 8392
rect 3988 8334 4080 8336
rect 5257 8392 8156 8394
rect 5257 8336 5262 8392
rect 5318 8336 8156 8392
rect 5257 8334 8156 8336
rect 3988 8332 4035 8334
rect 2589 8260 2655 8261
rect 2773 8260 2839 8261
rect 3696 8260 3756 8332
rect 3969 8331 4035 8332
rect 5257 8331 5323 8334
rect 8150 8332 8156 8334
rect 8220 8332 8226 8396
rect 11830 8394 11836 8396
rect 11790 8334 11836 8394
rect 11900 8392 11947 8396
rect 11942 8336 11947 8392
rect 11830 8332 11836 8334
rect 11900 8332 11947 8336
rect 13670 8332 13676 8396
rect 13740 8394 13746 8396
rect 14917 8394 14983 8397
rect 13740 8392 14983 8394
rect 13740 8336 14922 8392
rect 14978 8336 14983 8392
rect 13740 8334 14983 8336
rect 13740 8332 13746 8334
rect 11881 8331 11947 8332
rect 14917 8331 14983 8334
rect 15694 8332 15700 8396
rect 15764 8394 15770 8396
rect 17166 8394 17172 8396
rect 15764 8334 17172 8394
rect 15764 8332 15770 8334
rect 17166 8332 17172 8334
rect 17236 8332 17242 8396
rect 17358 8394 17418 8470
rect 18045 8528 20000 8530
rect 18045 8472 18050 8528
rect 18106 8472 20000 8528
rect 18045 8470 20000 8472
rect 18045 8467 18111 8470
rect 19200 8440 20000 8470
rect 18045 8394 18111 8397
rect 17358 8392 18111 8394
rect 17358 8336 18050 8392
rect 18106 8336 18111 8392
rect 17358 8334 18111 8336
rect 18045 8331 18111 8334
rect 2589 8258 2636 8260
rect 2544 8256 2636 8258
rect 2544 8200 2594 8256
rect 2544 8198 2636 8200
rect 2589 8196 2636 8198
rect 2700 8196 2706 8260
rect 2773 8256 2820 8260
rect 2884 8258 2890 8260
rect 2773 8200 2778 8256
rect 2773 8196 2820 8200
rect 2884 8198 2930 8258
rect 3696 8198 3740 8260
rect 2884 8196 2890 8198
rect 3734 8196 3740 8198
rect 3804 8196 3810 8260
rect 3877 8258 3943 8261
rect 4153 8258 4219 8261
rect 7465 8260 7531 8261
rect 7414 8258 7420 8260
rect 3877 8256 4219 8258
rect 3877 8200 3882 8256
rect 3938 8200 4158 8256
rect 4214 8200 4219 8256
rect 3877 8198 4219 8200
rect 7374 8198 7420 8258
rect 7484 8256 7531 8260
rect 7526 8200 7531 8256
rect 2589 8195 2655 8196
rect 2773 8195 2839 8196
rect 3877 8195 3943 8198
rect 4153 8195 4219 8198
rect 7414 8196 7420 8198
rect 7484 8196 7531 8200
rect 7465 8195 7531 8196
rect 3168 8192 3488 8193
rect 0 8122 800 8152
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 8127 3488 8128
rect 7616 8192 7936 8193
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 8127 7936 8128
rect 12064 8192 12384 8193
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 8127 12384 8128
rect 16512 8192 16832 8193
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 8127 16832 8128
rect 3601 8124 3667 8125
rect 0 8062 1594 8122
rect 0 8032 800 8062
rect 841 7952 907 7955
rect 798 7950 907 7952
rect 798 7894 846 7950
rect 902 7894 907 7950
rect 798 7889 907 7894
rect 798 7744 858 7889
rect 1534 7850 1594 8062
rect 3550 8060 3556 8124
rect 3620 8122 3667 8124
rect 3620 8120 3712 8122
rect 3662 8064 3712 8120
rect 3620 8062 3712 8064
rect 3620 8060 3667 8062
rect 3918 8060 3924 8124
rect 3988 8122 3994 8124
rect 4245 8122 4311 8125
rect 3988 8120 4311 8122
rect 3988 8064 4250 8120
rect 4306 8064 4311 8120
rect 3988 8062 4311 8064
rect 3988 8060 3994 8062
rect 3601 8059 3667 8060
rect 4245 8059 4311 8062
rect 8569 8122 8635 8125
rect 18321 8122 18387 8125
rect 19200 8122 20000 8152
rect 8569 8120 9506 8122
rect 8569 8064 8574 8120
rect 8630 8064 9506 8120
rect 8569 8062 9506 8064
rect 8569 8059 8635 8062
rect 3233 7986 3299 7989
rect 9213 7986 9279 7989
rect 2638 7984 9279 7986
rect 2638 7928 3238 7984
rect 3294 7928 9218 7984
rect 9274 7928 9279 7984
rect 2638 7926 9279 7928
rect 9446 7986 9506 8062
rect 18321 8120 20000 8122
rect 18321 8064 18326 8120
rect 18382 8064 20000 8120
rect 18321 8062 20000 8064
rect 18321 8059 18387 8062
rect 19200 8032 20000 8062
rect 13813 7986 13879 7989
rect 9446 7984 13879 7986
rect 9446 7928 13818 7984
rect 13874 7928 13879 7984
rect 9446 7926 13879 7928
rect 2638 7850 2698 7926
rect 3233 7923 3299 7926
rect 9213 7923 9279 7926
rect 13813 7923 13879 7926
rect 1534 7790 2698 7850
rect 3325 7850 3391 7853
rect 4521 7850 4587 7853
rect 3325 7848 4587 7850
rect 3325 7792 3330 7848
rect 3386 7792 4526 7848
rect 4582 7792 4587 7848
rect 3325 7790 4587 7792
rect 3325 7787 3391 7790
rect 4521 7787 4587 7790
rect 5022 7788 5028 7852
rect 5092 7850 5098 7852
rect 5257 7850 5323 7853
rect 10317 7850 10383 7853
rect 5092 7848 10383 7850
rect 5092 7792 5262 7848
rect 5318 7792 10322 7848
rect 10378 7792 10383 7848
rect 5092 7790 10383 7792
rect 5092 7788 5098 7790
rect 5257 7787 5323 7790
rect 10317 7787 10383 7790
rect 11789 7850 11855 7853
rect 14038 7850 14044 7852
rect 11789 7848 14044 7850
rect 11789 7792 11794 7848
rect 11850 7792 14044 7848
rect 11789 7790 14044 7792
rect 11789 7787 11855 7790
rect 14038 7788 14044 7790
rect 14108 7850 14114 7852
rect 16205 7850 16271 7853
rect 17033 7850 17099 7853
rect 14108 7848 17099 7850
rect 14108 7792 16210 7848
rect 16266 7792 17038 7848
rect 17094 7792 17099 7848
rect 14108 7790 17099 7792
rect 14108 7788 14114 7790
rect 16205 7787 16271 7790
rect 17033 7787 17099 7790
rect 18505 7850 18571 7853
rect 19200 7850 20000 7880
rect 18505 7848 20000 7850
rect 18505 7792 18510 7848
rect 18566 7792 20000 7848
rect 18505 7790 20000 7792
rect 18505 7787 18571 7790
rect 19200 7760 20000 7790
rect 0 7654 858 7744
rect 3601 7714 3667 7717
rect 4061 7714 4127 7717
rect 982 7712 4127 7714
rect 982 7656 3606 7712
rect 3662 7656 4066 7712
rect 4122 7656 4127 7712
rect 982 7654 4127 7656
rect 0 7624 800 7654
rect 0 7442 800 7472
rect 982 7442 1042 7654
rect 3601 7651 3667 7654
rect 4061 7651 4127 7654
rect 4337 7714 4403 7717
rect 4470 7714 4476 7716
rect 4337 7712 4476 7714
rect 4337 7656 4342 7712
rect 4398 7656 4476 7712
rect 4337 7654 4476 7656
rect 4337 7651 4403 7654
rect 4470 7652 4476 7654
rect 4540 7652 4546 7716
rect 6637 7714 6703 7717
rect 8201 7714 8267 7717
rect 6637 7712 8267 7714
rect 6637 7656 6642 7712
rect 6698 7656 8206 7712
rect 8262 7656 8267 7712
rect 6637 7654 8267 7656
rect 6637 7651 6703 7654
rect 8201 7651 8267 7654
rect 2681 7578 2747 7581
rect 4102 7578 4108 7580
rect 2681 7576 4108 7578
rect 2681 7520 2686 7576
rect 2742 7520 4108 7576
rect 2681 7518 4108 7520
rect 2681 7515 2747 7518
rect 4102 7516 4108 7518
rect 4172 7578 4178 7580
rect 4340 7578 4400 7651
rect 5392 7648 5712 7649
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 5392 7583 5712 7584
rect 9840 7648 10160 7649
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9840 7583 10160 7584
rect 14288 7648 14608 7649
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 7583 14608 7584
rect 4613 7580 4679 7581
rect 4613 7578 4660 7580
rect 4172 7518 4400 7578
rect 4568 7576 4660 7578
rect 4568 7520 4618 7576
rect 4568 7518 4660 7520
rect 4172 7516 4178 7518
rect 4613 7516 4660 7518
rect 4724 7516 4730 7580
rect 5993 7578 6059 7581
rect 7925 7578 7991 7581
rect 15929 7580 15995 7581
rect 5993 7576 7991 7578
rect 5993 7520 5998 7576
rect 6054 7520 7930 7576
rect 7986 7520 7991 7576
rect 5993 7518 7991 7520
rect 4613 7515 4679 7516
rect 5993 7515 6059 7518
rect 7925 7515 7991 7518
rect 15878 7516 15884 7580
rect 15948 7578 15995 7580
rect 16297 7578 16363 7581
rect 15948 7576 16040 7578
rect 15990 7520 16040 7576
rect 15948 7518 16040 7520
rect 16297 7576 18154 7578
rect 16297 7520 16302 7576
rect 16358 7520 18154 7576
rect 16297 7518 18154 7520
rect 15948 7516 15995 7518
rect 15929 7515 15995 7516
rect 16297 7515 16363 7518
rect 0 7382 1042 7442
rect 1117 7442 1183 7445
rect 9765 7442 9831 7445
rect 1117 7440 9831 7442
rect 1117 7384 1122 7440
rect 1178 7384 9770 7440
rect 9826 7384 9831 7440
rect 1117 7382 9831 7384
rect 0 7352 800 7382
rect 1117 7379 1183 7382
rect 9765 7379 9831 7382
rect 9949 7442 10015 7445
rect 17953 7442 18019 7445
rect 9949 7440 18019 7442
rect 9949 7384 9954 7440
rect 10010 7384 17958 7440
rect 18014 7384 18019 7440
rect 9949 7382 18019 7384
rect 9949 7379 10015 7382
rect 17953 7379 18019 7382
rect 3693 7308 3759 7309
rect 3693 7306 3740 7308
rect 3648 7304 3740 7306
rect 3648 7248 3698 7304
rect 3648 7246 3740 7248
rect 3693 7244 3740 7246
rect 3804 7244 3810 7308
rect 4613 7306 4679 7309
rect 9305 7306 9371 7309
rect 4613 7304 9506 7306
rect 4613 7248 4618 7304
rect 4674 7248 9310 7304
rect 9366 7248 9506 7304
rect 4613 7246 9506 7248
rect 3693 7243 3759 7244
rect 4613 7243 4679 7246
rect 9305 7243 9371 7246
rect 3785 7172 3851 7173
rect 3734 7108 3740 7172
rect 3804 7170 3851 7172
rect 3804 7168 3896 7170
rect 3846 7112 3896 7168
rect 3804 7110 3896 7112
rect 3804 7108 3851 7110
rect 4470 7108 4476 7172
rect 4540 7170 4546 7172
rect 5441 7170 5507 7173
rect 4540 7168 5507 7170
rect 4540 7112 5446 7168
rect 5502 7112 5507 7168
rect 4540 7110 5507 7112
rect 4540 7108 4546 7110
rect 3785 7107 3851 7108
rect 5441 7107 5507 7110
rect 5625 7170 5691 7173
rect 6126 7170 6132 7172
rect 5625 7168 6132 7170
rect 5625 7112 5630 7168
rect 5686 7112 6132 7168
rect 5625 7110 6132 7112
rect 5625 7107 5691 7110
rect 6126 7108 6132 7110
rect 6196 7108 6202 7172
rect 9446 7170 9506 7246
rect 9622 7244 9628 7308
rect 9692 7306 9698 7308
rect 15377 7306 15443 7309
rect 9692 7304 15443 7306
rect 9692 7248 15382 7304
rect 15438 7248 15443 7304
rect 9692 7246 15443 7248
rect 9692 7244 9698 7246
rect 15377 7243 15443 7246
rect 16665 7306 16731 7309
rect 16982 7306 16988 7308
rect 16665 7304 16988 7306
rect 16665 7248 16670 7304
rect 16726 7248 16988 7304
rect 16665 7246 16988 7248
rect 16665 7243 16731 7246
rect 16982 7244 16988 7246
rect 17052 7244 17058 7308
rect 9949 7170 10015 7173
rect 9446 7168 10015 7170
rect 9446 7112 9954 7168
rect 10010 7112 10015 7168
rect 9446 7110 10015 7112
rect 9949 7107 10015 7110
rect 15285 7170 15351 7173
rect 15878 7170 15884 7172
rect 15285 7168 15884 7170
rect 15285 7112 15290 7168
rect 15346 7112 15884 7168
rect 15285 7110 15884 7112
rect 15285 7107 15351 7110
rect 15878 7108 15884 7110
rect 15948 7170 15954 7172
rect 16297 7170 16363 7173
rect 15948 7168 16363 7170
rect 15948 7112 16302 7168
rect 16358 7112 16363 7168
rect 15948 7110 16363 7112
rect 15948 7108 15954 7110
rect 16297 7107 16363 7110
rect 3168 7104 3488 7105
rect 0 7034 800 7064
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3168 7039 3488 7040
rect 7616 7104 7936 7105
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 7039 7936 7040
rect 12064 7104 12384 7105
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 7039 12384 7040
rect 16512 7104 16832 7105
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 7039 16832 7040
rect 2773 7034 2839 7037
rect 4613 7034 4679 7037
rect 0 7032 2839 7034
rect 0 6976 2778 7032
rect 2834 6976 2839 7032
rect 0 6974 2839 6976
rect 0 6944 800 6974
rect 2773 6971 2839 6974
rect 4110 7032 4679 7034
rect 4110 6976 4618 7032
rect 4674 6976 4679 7032
rect 4110 6974 4679 6976
rect 2998 6836 3004 6900
rect 3068 6898 3074 6900
rect 3417 6898 3483 6901
rect 4110 6898 4170 6974
rect 4613 6971 4679 6974
rect 5257 7034 5323 7037
rect 11278 7034 11284 7036
rect 5257 7032 6516 7034
rect 5257 6976 5262 7032
rect 5318 6976 6516 7032
rect 5257 6974 6516 6976
rect 5257 6971 5323 6974
rect 3068 6896 4170 6898
rect 3068 6840 3422 6896
rect 3478 6840 4170 6896
rect 3068 6838 4170 6840
rect 3068 6836 3074 6838
rect 3417 6835 3483 6838
rect 4470 6836 4476 6900
rect 4540 6898 4546 6900
rect 4613 6898 4679 6901
rect 4540 6896 4679 6898
rect 4540 6840 4618 6896
rect 4674 6840 4679 6896
rect 4540 6838 4679 6840
rect 4540 6836 4546 6838
rect 4613 6835 4679 6838
rect 4838 6836 4844 6900
rect 4908 6898 4914 6900
rect 6269 6898 6335 6901
rect 4908 6896 6335 6898
rect 4908 6840 6274 6896
rect 6330 6840 6335 6896
rect 4908 6838 6335 6840
rect 6456 6898 6516 6974
rect 8250 6974 11284 7034
rect 8250 6898 8310 6974
rect 11278 6972 11284 6974
rect 11348 6972 11354 7036
rect 12985 7034 13051 7037
rect 12985 7032 13508 7034
rect 12985 6976 12990 7032
rect 13046 6976 13508 7032
rect 12985 6974 13508 6976
rect 12985 6971 13051 6974
rect 6456 6838 8310 6898
rect 4908 6836 4914 6838
rect 6269 6835 6335 6838
rect 13118 6836 13124 6900
rect 13188 6898 13194 6900
rect 13261 6898 13327 6901
rect 13188 6896 13327 6898
rect 13188 6840 13266 6896
rect 13322 6840 13327 6896
rect 13188 6838 13327 6840
rect 13448 6898 13508 6974
rect 14774 6972 14780 7036
rect 14844 7034 14850 7036
rect 15101 7034 15167 7037
rect 14844 7032 15167 7034
rect 14844 6976 15106 7032
rect 15162 6976 15167 7032
rect 14844 6974 15167 6976
rect 18094 7034 18154 7518
rect 18597 7442 18663 7445
rect 19200 7442 20000 7472
rect 18597 7440 20000 7442
rect 18597 7384 18602 7440
rect 18658 7384 20000 7440
rect 18597 7382 20000 7384
rect 18597 7379 18663 7382
rect 19200 7352 20000 7382
rect 19200 7034 20000 7064
rect 18094 6974 20000 7034
rect 14844 6972 14850 6974
rect 15101 6971 15167 6974
rect 19200 6944 20000 6974
rect 15694 6898 15700 6900
rect 13448 6838 15700 6898
rect 13188 6836 13194 6838
rect 13261 6835 13327 6838
rect 15694 6836 15700 6838
rect 15764 6836 15770 6900
rect 17125 6898 17191 6901
rect 17350 6898 17356 6900
rect 17125 6896 17356 6898
rect 17125 6840 17130 6896
rect 17186 6840 17356 6896
rect 17125 6838 17356 6840
rect 17125 6835 17191 6838
rect 17350 6836 17356 6838
rect 17420 6836 17426 6900
rect 0 6762 800 6792
rect 933 6762 999 6765
rect 0 6760 999 6762
rect 0 6704 938 6760
rect 994 6704 999 6760
rect 0 6702 999 6704
rect 0 6672 800 6702
rect 933 6699 999 6702
rect 1945 6762 2011 6765
rect 5073 6762 5139 6765
rect 7046 6762 7052 6764
rect 1945 6760 4906 6762
rect 1945 6704 1950 6760
rect 2006 6704 4906 6760
rect 1945 6702 4906 6704
rect 1945 6699 2011 6702
rect 3550 6564 3556 6628
rect 3620 6626 3626 6628
rect 3785 6626 3851 6629
rect 3620 6624 3851 6626
rect 3620 6568 3790 6624
rect 3846 6568 3851 6624
rect 3620 6566 3851 6568
rect 3620 6564 3626 6566
rect 3785 6563 3851 6566
rect 0 6490 800 6520
rect 4429 6490 4495 6493
rect 0 6488 4495 6490
rect 0 6432 4434 6488
rect 4490 6432 4495 6488
rect 0 6430 4495 6432
rect 0 6400 800 6430
rect 4429 6427 4495 6430
rect 3141 6354 3207 6357
rect 3550 6354 3556 6356
rect 3141 6352 3556 6354
rect 3141 6296 3146 6352
rect 3202 6296 3556 6352
rect 3141 6294 3556 6296
rect 3141 6291 3207 6294
rect 3550 6292 3556 6294
rect 3620 6292 3626 6356
rect 4846 6354 4906 6702
rect 5073 6760 7052 6762
rect 5073 6704 5078 6760
rect 5134 6704 7052 6760
rect 5073 6702 7052 6704
rect 5073 6699 5139 6702
rect 7046 6700 7052 6702
rect 7116 6762 7122 6764
rect 9213 6762 9279 6765
rect 16849 6762 16915 6765
rect 7116 6760 9279 6762
rect 7116 6704 9218 6760
rect 9274 6704 9279 6760
rect 7116 6702 9279 6704
rect 7116 6700 7122 6702
rect 9213 6699 9279 6702
rect 9630 6760 16915 6762
rect 9630 6704 16854 6760
rect 16910 6704 16915 6760
rect 9630 6702 16915 6704
rect 5392 6560 5712 6561
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 5392 6495 5712 6496
rect 7230 6428 7236 6492
rect 7300 6490 7306 6492
rect 7557 6490 7623 6493
rect 9489 6490 9555 6493
rect 9630 6490 9690 6702
rect 16849 6699 16915 6702
rect 11329 6626 11395 6629
rect 13997 6626 14063 6629
rect 11329 6624 14063 6626
rect 11329 6568 11334 6624
rect 11390 6568 14002 6624
rect 14058 6568 14063 6624
rect 11329 6566 14063 6568
rect 11329 6563 11395 6566
rect 13997 6563 14063 6566
rect 15009 6626 15075 6629
rect 19200 6626 20000 6656
rect 15009 6624 20000 6626
rect 15009 6568 15014 6624
rect 15070 6568 20000 6624
rect 15009 6566 20000 6568
rect 15009 6563 15075 6566
rect 9840 6560 10160 6561
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 6495 10160 6496
rect 14288 6560 14608 6561
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 19200 6536 20000 6566
rect 14288 6495 14608 6496
rect 7300 6488 9690 6490
rect 7300 6432 7562 6488
rect 7618 6432 9494 6488
rect 9550 6432 9690 6488
rect 7300 6430 9690 6432
rect 11789 6490 11855 6493
rect 13077 6490 13143 6493
rect 11789 6488 13143 6490
rect 11789 6432 11794 6488
rect 11850 6432 13082 6488
rect 13138 6432 13143 6488
rect 11789 6430 13143 6432
rect 7300 6428 7306 6430
rect 7557 6427 7623 6430
rect 9489 6427 9555 6430
rect 11789 6427 11855 6430
rect 13077 6427 13143 6430
rect 6821 6354 6887 6357
rect 8017 6354 8083 6357
rect 15009 6354 15075 6357
rect 4846 6294 6194 6354
rect 1117 6218 1183 6221
rect 3918 6218 3924 6220
rect 1117 6216 3924 6218
rect 1117 6160 1122 6216
rect 1178 6160 3924 6216
rect 1117 6158 3924 6160
rect 1117 6155 1183 6158
rect 3918 6156 3924 6158
rect 3988 6156 3994 6220
rect 4337 6218 4403 6221
rect 4981 6218 5047 6221
rect 6134 6220 6194 6294
rect 6821 6352 15075 6354
rect 6821 6296 6826 6352
rect 6882 6296 8022 6352
rect 8078 6296 15014 6352
rect 15070 6296 15075 6352
rect 6821 6294 15075 6296
rect 6821 6291 6887 6294
rect 8017 6291 8083 6294
rect 15009 6291 15075 6294
rect 15653 6354 15719 6357
rect 16941 6354 17007 6357
rect 15653 6352 17007 6354
rect 15653 6296 15658 6352
rect 15714 6296 16946 6352
rect 17002 6296 17007 6352
rect 15653 6294 17007 6296
rect 15653 6291 15719 6294
rect 16941 6291 17007 6294
rect 4337 6216 5047 6218
rect 4337 6160 4342 6216
rect 4398 6160 4986 6216
rect 5042 6160 5047 6216
rect 4337 6158 5047 6160
rect 4337 6155 4403 6158
rect 4981 6155 5047 6158
rect 6126 6156 6132 6220
rect 6196 6218 6202 6220
rect 10409 6218 10475 6221
rect 13997 6218 14063 6221
rect 6196 6158 8080 6218
rect 6196 6156 6202 6158
rect 0 6082 800 6112
rect 2957 6082 3023 6085
rect 0 6080 3023 6082
rect 0 6024 2962 6080
rect 3018 6024 3023 6080
rect 0 6022 3023 6024
rect 0 5992 800 6022
rect 2957 6019 3023 6022
rect 4654 6020 4660 6084
rect 4724 6082 4730 6084
rect 4889 6082 4955 6085
rect 4724 6080 4955 6082
rect 4724 6024 4894 6080
rect 4950 6024 4955 6080
rect 4724 6022 4955 6024
rect 8020 6082 8080 6158
rect 10409 6216 14063 6218
rect 10409 6160 10414 6216
rect 10470 6160 14002 6216
rect 14058 6160 14063 6216
rect 10409 6158 14063 6160
rect 10409 6155 10475 6158
rect 13997 6155 14063 6158
rect 16021 6218 16087 6221
rect 19200 6218 20000 6248
rect 16021 6216 20000 6218
rect 16021 6160 16026 6216
rect 16082 6160 20000 6216
rect 16021 6158 20000 6160
rect 16021 6155 16087 6158
rect 19200 6128 20000 6158
rect 10685 6082 10751 6085
rect 8020 6080 10751 6082
rect 8020 6024 10690 6080
rect 10746 6024 10751 6080
rect 8020 6022 10751 6024
rect 4724 6020 4730 6022
rect 4889 6019 4955 6022
rect 10685 6019 10751 6022
rect 15837 6082 15903 6085
rect 15837 6080 15946 6082
rect 15837 6024 15842 6080
rect 15898 6024 15946 6080
rect 15837 6019 15946 6024
rect 3168 6016 3488 6017
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 3168 5951 3488 5952
rect 7616 6016 7936 6017
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 5951 7936 5952
rect 12064 6016 12384 6017
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 5951 12384 5952
rect 2814 5884 2820 5948
rect 2884 5946 2890 5948
rect 2957 5946 3023 5949
rect 15009 5948 15075 5949
rect 2884 5944 3023 5946
rect 2884 5888 2962 5944
rect 3018 5888 3023 5944
rect 2884 5886 3023 5888
rect 2884 5884 2890 5886
rect 2957 5883 3023 5886
rect 14958 5884 14964 5948
rect 15028 5946 15075 5948
rect 15028 5944 15120 5946
rect 15070 5888 15120 5944
rect 15028 5886 15120 5888
rect 15028 5884 15075 5886
rect 15009 5883 15075 5884
rect 0 5810 800 5840
rect 8753 5810 8819 5813
rect 0 5808 8819 5810
rect 0 5752 8758 5808
rect 8814 5752 8819 5808
rect 0 5750 8819 5752
rect 0 5720 800 5750
rect 8753 5747 8819 5750
rect 9029 5810 9095 5813
rect 15193 5810 15259 5813
rect 9029 5808 15259 5810
rect 9029 5752 9034 5808
rect 9090 5752 15198 5808
rect 15254 5752 15259 5808
rect 9029 5750 15259 5752
rect 15886 5810 15946 6019
rect 16512 6016 16832 6017
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 5951 16832 5952
rect 16941 5946 17007 5949
rect 19200 5946 20000 5976
rect 16941 5944 20000 5946
rect 16941 5888 16946 5944
rect 17002 5888 20000 5944
rect 16941 5886 20000 5888
rect 16941 5883 17007 5886
rect 19200 5856 20000 5886
rect 16757 5810 16823 5813
rect 15886 5808 16823 5810
rect 15886 5752 16762 5808
rect 16818 5752 16823 5808
rect 15886 5750 16823 5752
rect 9029 5747 9095 5750
rect 15193 5747 15259 5750
rect 16757 5747 16823 5750
rect 1669 5674 1735 5677
rect 5073 5674 5139 5677
rect 1669 5672 5139 5674
rect 1669 5616 1674 5672
rect 1730 5616 5078 5672
rect 5134 5616 5139 5672
rect 1669 5614 5139 5616
rect 1669 5611 1735 5614
rect 5073 5611 5139 5614
rect 14641 5674 14707 5677
rect 14958 5674 14964 5676
rect 14641 5672 14964 5674
rect 14641 5616 14646 5672
rect 14702 5616 14964 5672
rect 14641 5614 14964 5616
rect 14641 5611 14707 5614
rect 14958 5612 14964 5614
rect 15028 5612 15034 5676
rect 2681 5538 2747 5541
rect 4705 5538 4771 5541
rect 13997 5538 14063 5541
rect 2681 5536 4771 5538
rect 2681 5480 2686 5536
rect 2742 5480 4710 5536
rect 4766 5480 4771 5536
rect 2681 5478 4771 5480
rect 2681 5475 2747 5478
rect 4705 5475 4771 5478
rect 10366 5536 14063 5538
rect 10366 5480 14002 5536
rect 14058 5480 14063 5536
rect 10366 5478 14063 5480
rect 5392 5472 5712 5473
rect 0 5402 800 5432
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 5407 5712 5408
rect 9840 5472 10160 5473
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 5407 10160 5408
rect 1761 5402 1827 5405
rect 0 5400 1827 5402
rect 0 5344 1766 5400
rect 1822 5344 1827 5400
rect 0 5342 1827 5344
rect 0 5312 800 5342
rect 1761 5339 1827 5342
rect 5809 5402 5875 5405
rect 5942 5402 5948 5404
rect 5809 5400 5948 5402
rect 5809 5344 5814 5400
rect 5870 5344 5948 5400
rect 5809 5342 5948 5344
rect 5809 5339 5875 5342
rect 5942 5340 5948 5342
rect 6012 5340 6018 5404
rect 7230 5340 7236 5404
rect 7300 5402 7306 5404
rect 7373 5402 7439 5405
rect 7300 5400 9690 5402
rect 7300 5344 7378 5400
rect 7434 5344 9690 5400
rect 7300 5342 9690 5344
rect 7300 5340 7306 5342
rect 7373 5339 7439 5342
rect 1945 5266 2011 5269
rect 8753 5266 8819 5269
rect 1945 5264 8819 5266
rect 1945 5208 1950 5264
rect 2006 5208 8758 5264
rect 8814 5208 8819 5264
rect 1945 5206 8819 5208
rect 9630 5266 9690 5342
rect 10366 5266 10426 5478
rect 13997 5475 14063 5478
rect 16205 5538 16271 5541
rect 19200 5538 20000 5568
rect 16205 5536 20000 5538
rect 16205 5480 16210 5536
rect 16266 5480 20000 5536
rect 16205 5478 20000 5480
rect 16205 5475 16271 5478
rect 14288 5472 14608 5473
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 19200 5448 20000 5478
rect 14288 5407 14608 5408
rect 9630 5206 10426 5266
rect 10869 5266 10935 5269
rect 14641 5266 14707 5269
rect 10869 5264 14707 5266
rect 10869 5208 10874 5264
rect 10930 5208 14646 5264
rect 14702 5208 14707 5264
rect 10869 5206 14707 5208
rect 1945 5203 2011 5206
rect 8753 5203 8819 5206
rect 10869 5203 10935 5206
rect 14641 5203 14707 5206
rect 0 5130 800 5160
rect 1485 5130 1551 5133
rect 0 5128 1551 5130
rect 0 5072 1490 5128
rect 1546 5072 1551 5128
rect 0 5070 1551 5072
rect 0 5040 800 5070
rect 1485 5067 1551 5070
rect 2957 5130 3023 5133
rect 5993 5130 6059 5133
rect 2957 5128 6059 5130
rect 2957 5072 2962 5128
rect 3018 5072 5998 5128
rect 6054 5072 6059 5128
rect 2957 5070 6059 5072
rect 2957 5067 3023 5070
rect 5993 5067 6059 5070
rect 6453 5130 6519 5133
rect 10225 5130 10291 5133
rect 6453 5128 10291 5130
rect 6453 5072 6458 5128
rect 6514 5072 10230 5128
rect 10286 5072 10291 5128
rect 6453 5070 10291 5072
rect 6453 5067 6519 5070
rect 10225 5067 10291 5070
rect 10358 5068 10364 5132
rect 10428 5130 10434 5132
rect 11973 5130 12039 5133
rect 10428 5128 12039 5130
rect 10428 5072 11978 5128
rect 12034 5072 12039 5128
rect 10428 5070 12039 5072
rect 10428 5068 10434 5070
rect 11973 5067 12039 5070
rect 12341 5130 12407 5133
rect 19200 5130 20000 5160
rect 12341 5128 20000 5130
rect 12341 5072 12346 5128
rect 12402 5072 20000 5128
rect 12341 5070 20000 5072
rect 12341 5067 12407 5070
rect 19200 5040 20000 5070
rect 4102 4932 4108 4996
rect 4172 4994 4178 4996
rect 7465 4994 7531 4997
rect 4172 4992 7531 4994
rect 4172 4936 7470 4992
rect 7526 4936 7531 4992
rect 4172 4934 7531 4936
rect 4172 4932 4178 4934
rect 7465 4931 7531 4934
rect 3168 4928 3488 4929
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 3168 4863 3488 4864
rect 7616 4928 7936 4929
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 4863 7936 4864
rect 12064 4928 12384 4929
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 4863 12384 4864
rect 16512 4928 16832 4929
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 4863 16832 4864
rect 2405 4860 2471 4861
rect 2405 4858 2452 4860
rect 2360 4856 2452 4858
rect 2360 4800 2410 4856
rect 2360 4798 2452 4800
rect 2405 4796 2452 4798
rect 2516 4796 2522 4860
rect 6862 4796 6868 4860
rect 6932 4858 6938 4860
rect 7097 4858 7163 4861
rect 6932 4856 7163 4858
rect 6932 4800 7102 4856
rect 7158 4800 7163 4856
rect 6932 4798 7163 4800
rect 6932 4796 6938 4798
rect 2405 4795 2471 4796
rect 7097 4795 7163 4798
rect 0 4722 800 4752
rect 1117 4722 1183 4725
rect 2313 4724 2379 4725
rect 0 4720 1183 4722
rect 0 4664 1122 4720
rect 1178 4664 1183 4720
rect 0 4662 1183 4664
rect 0 4632 800 4662
rect 1117 4659 1183 4662
rect 2262 4660 2268 4724
rect 2332 4722 2379 4724
rect 2497 4722 2563 4725
rect 2630 4722 2636 4724
rect 2332 4720 2424 4722
rect 2374 4664 2424 4720
rect 2332 4662 2424 4664
rect 2497 4720 2636 4722
rect 2497 4664 2502 4720
rect 2558 4664 2636 4720
rect 2497 4662 2636 4664
rect 2332 4660 2379 4662
rect 2313 4659 2379 4660
rect 2497 4659 2563 4662
rect 2630 4660 2636 4662
rect 2700 4722 2706 4724
rect 3417 4722 3483 4725
rect 2700 4720 3483 4722
rect 2700 4664 3422 4720
rect 3478 4664 3483 4720
rect 2700 4662 3483 4664
rect 2700 4660 2706 4662
rect 3417 4659 3483 4662
rect 5165 4722 5231 4725
rect 15009 4722 15075 4725
rect 5165 4720 15075 4722
rect 5165 4664 5170 4720
rect 5226 4664 15014 4720
rect 15070 4664 15075 4720
rect 5165 4662 15075 4664
rect 5165 4659 5231 4662
rect 15009 4659 15075 4662
rect 18413 4722 18479 4725
rect 19200 4722 20000 4752
rect 18413 4720 20000 4722
rect 18413 4664 18418 4720
rect 18474 4664 20000 4720
rect 18413 4662 20000 4664
rect 18413 4659 18479 4662
rect 19200 4632 20000 4662
rect 1393 4586 1459 4589
rect 4245 4586 4311 4589
rect 1393 4584 4311 4586
rect 1393 4528 1398 4584
rect 1454 4528 4250 4584
rect 4306 4528 4311 4584
rect 1393 4526 4311 4528
rect 1393 4523 1459 4526
rect 4245 4523 4311 4526
rect 4429 4586 4495 4589
rect 11605 4586 11671 4589
rect 4429 4584 11671 4586
rect 4429 4528 4434 4584
rect 4490 4528 11610 4584
rect 11666 4528 11671 4584
rect 4429 4526 11671 4528
rect 4429 4523 4495 4526
rect 11605 4523 11671 4526
rect 13353 4586 13419 4589
rect 13353 4584 15256 4586
rect 13353 4528 13358 4584
rect 13414 4528 15256 4584
rect 13353 4526 15256 4528
rect 13353 4523 13419 4526
rect 0 4450 800 4480
rect 4061 4450 4127 4453
rect 0 4448 4127 4450
rect 0 4392 4066 4448
rect 4122 4392 4127 4448
rect 0 4390 4127 4392
rect 0 4360 800 4390
rect 4061 4387 4127 4390
rect 6177 4450 6243 4453
rect 9305 4450 9371 4453
rect 6177 4448 9371 4450
rect 6177 4392 6182 4448
rect 6238 4392 9310 4448
rect 9366 4392 9371 4448
rect 6177 4390 9371 4392
rect 6177 4387 6243 4390
rect 9305 4387 9371 4390
rect 10225 4450 10291 4453
rect 10726 4450 10732 4452
rect 10225 4448 10732 4450
rect 10225 4392 10230 4448
rect 10286 4392 10732 4448
rect 10225 4390 10732 4392
rect 10225 4387 10291 4390
rect 10726 4388 10732 4390
rect 10796 4450 10802 4452
rect 13721 4450 13787 4453
rect 10796 4448 13787 4450
rect 10796 4392 13726 4448
rect 13782 4392 13787 4448
rect 10796 4390 13787 4392
rect 10796 4388 10802 4390
rect 13721 4387 13787 4390
rect 5392 4384 5712 4385
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 4319 5712 4320
rect 9840 4384 10160 4385
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9840 4319 10160 4320
rect 14288 4384 14608 4385
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14288 4319 14608 4320
rect 3233 4314 3299 4317
rect 10225 4314 10291 4317
rect 10869 4314 10935 4317
rect 3233 4312 5274 4314
rect 3233 4256 3238 4312
rect 3294 4256 5274 4312
rect 3233 4254 5274 4256
rect 3233 4251 3299 4254
rect 0 4178 800 4208
rect 5073 4178 5139 4181
rect 0 4176 5139 4178
rect 0 4120 5078 4176
rect 5134 4120 5139 4176
rect 0 4118 5139 4120
rect 5214 4178 5274 4254
rect 8020 4254 9690 4314
rect 8020 4178 8080 4254
rect 5214 4118 8080 4178
rect 8201 4178 8267 4181
rect 9489 4178 9555 4181
rect 8201 4176 9555 4178
rect 8201 4120 8206 4176
rect 8262 4120 9494 4176
rect 9550 4120 9555 4176
rect 8201 4118 9555 4120
rect 9630 4178 9690 4254
rect 10225 4312 10935 4314
rect 10225 4256 10230 4312
rect 10286 4256 10874 4312
rect 10930 4256 10935 4312
rect 10225 4254 10935 4256
rect 15196 4314 15256 4526
rect 19200 4314 20000 4344
rect 15196 4254 20000 4314
rect 10225 4251 10291 4254
rect 10869 4251 10935 4254
rect 19200 4224 20000 4254
rect 11646 4178 11652 4180
rect 9630 4118 11652 4178
rect 0 4088 800 4118
rect 5073 4115 5139 4118
rect 8201 4115 8267 4118
rect 9489 4115 9555 4118
rect 11646 4116 11652 4118
rect 11716 4178 11722 4180
rect 11973 4178 12039 4181
rect 11716 4176 12039 4178
rect 11716 4120 11978 4176
rect 12034 4120 12039 4176
rect 11716 4118 12039 4120
rect 11716 4116 11722 4118
rect 11973 4115 12039 4118
rect 13905 4178 13971 4181
rect 17033 4178 17099 4181
rect 13905 4176 17099 4178
rect 13905 4120 13910 4176
rect 13966 4120 17038 4176
rect 17094 4120 17099 4176
rect 13905 4118 17099 4120
rect 13905 4115 13971 4118
rect 17033 4115 17099 4118
rect 3785 4044 3851 4045
rect 3734 4042 3740 4044
rect 3694 3982 3740 4042
rect 3804 4040 3851 4044
rect 3846 3984 3851 4040
rect 3734 3980 3740 3982
rect 3804 3980 3851 3984
rect 3785 3979 3851 3980
rect 5165 4042 5231 4045
rect 13813 4042 13879 4045
rect 15101 4044 15167 4045
rect 15101 4042 15148 4044
rect 5165 4040 13879 4042
rect 5165 3984 5170 4040
rect 5226 3984 13818 4040
rect 13874 3984 13879 4040
rect 5165 3982 13879 3984
rect 15056 4040 15148 4042
rect 15056 3984 15106 4040
rect 15056 3982 15148 3984
rect 5165 3979 5231 3982
rect 13813 3979 13879 3982
rect 15101 3980 15148 3982
rect 15212 3980 15218 4044
rect 17585 4042 17651 4045
rect 19200 4042 20000 4072
rect 17585 4040 20000 4042
rect 17585 3984 17590 4040
rect 17646 3984 20000 4040
rect 17585 3982 20000 3984
rect 15101 3979 15167 3980
rect 17585 3979 17651 3982
rect 19200 3952 20000 3982
rect 2078 3906 2084 3908
rect 798 3846 2084 3906
rect 798 3800 858 3846
rect 2078 3844 2084 3846
rect 2148 3844 2154 3908
rect 4705 3906 4771 3909
rect 6821 3906 6887 3909
rect 4705 3904 6887 3906
rect 4705 3848 4710 3904
rect 4766 3848 6826 3904
rect 6882 3848 6887 3904
rect 4705 3846 6887 3848
rect 4705 3843 4771 3846
rect 6821 3843 6887 3846
rect 8201 3906 8267 3909
rect 9622 3906 9628 3908
rect 8201 3904 9628 3906
rect 8201 3848 8206 3904
rect 8262 3848 9628 3904
rect 8201 3846 9628 3848
rect 8201 3843 8267 3846
rect 9622 3844 9628 3846
rect 9692 3844 9698 3908
rect 10593 3906 10659 3909
rect 11145 3906 11211 3909
rect 10593 3904 11211 3906
rect 10593 3848 10598 3904
rect 10654 3848 11150 3904
rect 11206 3848 11211 3904
rect 10593 3846 11211 3848
rect 10593 3843 10659 3846
rect 11145 3843 11211 3846
rect 13854 3844 13860 3908
rect 13924 3906 13930 3908
rect 14774 3906 14780 3908
rect 13924 3846 14780 3906
rect 13924 3844 13930 3846
rect 14774 3844 14780 3846
rect 14844 3844 14850 3908
rect 0 3710 858 3800
rect 3168 3840 3488 3841
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 3168 3775 3488 3776
rect 7616 3840 7936 3841
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7616 3775 7936 3776
rect 12064 3840 12384 3841
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 3775 12384 3776
rect 16512 3840 16832 3841
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16512 3775 16832 3776
rect 4245 3770 4311 3773
rect 5257 3770 5323 3773
rect 4245 3768 5323 3770
rect 4245 3712 4250 3768
rect 4306 3712 5262 3768
rect 5318 3712 5323 3768
rect 4245 3710 5323 3712
rect 0 3680 800 3710
rect 4245 3707 4311 3710
rect 5257 3707 5323 3710
rect 7230 3708 7236 3772
rect 7300 3770 7306 3772
rect 7465 3770 7531 3773
rect 7300 3768 7531 3770
rect 7300 3712 7470 3768
rect 7526 3712 7531 3768
rect 7300 3710 7531 3712
rect 7300 3708 7306 3710
rect 7465 3707 7531 3710
rect 9438 3708 9444 3772
rect 9508 3770 9514 3772
rect 11605 3770 11671 3773
rect 9508 3768 11671 3770
rect 9508 3712 11610 3768
rect 11666 3712 11671 3768
rect 9508 3710 11671 3712
rect 9508 3708 9514 3710
rect 11605 3707 11671 3710
rect 14038 3708 14044 3772
rect 14108 3770 14114 3772
rect 14457 3770 14523 3773
rect 14108 3768 14523 3770
rect 14108 3712 14462 3768
rect 14518 3712 14523 3768
rect 14108 3710 14523 3712
rect 14108 3708 14114 3710
rect 14457 3707 14523 3710
rect 2037 3634 2103 3637
rect 12617 3634 12683 3637
rect 2037 3632 12683 3634
rect 2037 3576 2042 3632
rect 2098 3576 12622 3632
rect 12678 3576 12683 3632
rect 2037 3574 12683 3576
rect 2037 3571 2103 3574
rect 12617 3571 12683 3574
rect 13169 3634 13235 3637
rect 16246 3634 16252 3636
rect 13169 3632 16252 3634
rect 13169 3576 13174 3632
rect 13230 3576 16252 3632
rect 13169 3574 16252 3576
rect 13169 3571 13235 3574
rect 16246 3572 16252 3574
rect 16316 3572 16322 3636
rect 16665 3634 16731 3637
rect 17166 3634 17172 3636
rect 16665 3632 17172 3634
rect 16665 3576 16670 3632
rect 16726 3576 17172 3632
rect 16665 3574 17172 3576
rect 16665 3571 16731 3574
rect 17166 3572 17172 3574
rect 17236 3572 17242 3636
rect 18873 3634 18939 3637
rect 19200 3634 20000 3664
rect 18873 3632 20000 3634
rect 18873 3576 18878 3632
rect 18934 3576 20000 3632
rect 18873 3574 20000 3576
rect 18873 3571 18939 3574
rect 19200 3544 20000 3574
rect 0 3498 800 3528
rect 3509 3498 3575 3501
rect 6269 3498 6335 3501
rect 0 3496 3575 3498
rect 0 3440 3514 3496
rect 3570 3440 3575 3496
rect 0 3438 3575 3440
rect 0 3408 800 3438
rect 3509 3435 3575 3438
rect 4478 3496 6335 3498
rect 4478 3440 6274 3496
rect 6330 3440 6335 3496
rect 4478 3438 6335 3440
rect 1025 3362 1091 3365
rect 4478 3362 4538 3438
rect 6269 3435 6335 3438
rect 6913 3498 6979 3501
rect 8150 3498 8156 3500
rect 6913 3496 8156 3498
rect 6913 3440 6918 3496
rect 6974 3440 8156 3496
rect 6913 3438 8156 3440
rect 6913 3435 6979 3438
rect 8150 3436 8156 3438
rect 8220 3436 8226 3500
rect 8886 3436 8892 3500
rect 8956 3498 8962 3500
rect 13445 3498 13511 3501
rect 8956 3496 13511 3498
rect 8956 3440 13450 3496
rect 13506 3440 13511 3496
rect 8956 3438 13511 3440
rect 8956 3436 8962 3438
rect 13445 3435 13511 3438
rect 13670 3436 13676 3500
rect 13740 3498 13746 3500
rect 17217 3498 17283 3501
rect 13740 3496 17283 3498
rect 13740 3440 17222 3496
rect 17278 3440 17283 3496
rect 13740 3438 17283 3440
rect 13740 3436 13746 3438
rect 17217 3435 17283 3438
rect 1025 3360 4538 3362
rect 1025 3304 1030 3360
rect 1086 3304 4538 3360
rect 1025 3302 4538 3304
rect 6637 3362 6703 3365
rect 7925 3362 7991 3365
rect 6637 3360 7991 3362
rect 6637 3304 6642 3360
rect 6698 3304 7930 3360
rect 7986 3304 7991 3360
rect 6637 3302 7991 3304
rect 1025 3299 1091 3302
rect 6637 3299 6703 3302
rect 7925 3299 7991 3302
rect 10685 3362 10751 3365
rect 12065 3362 12131 3365
rect 10685 3360 12131 3362
rect 10685 3304 10690 3360
rect 10746 3304 12070 3360
rect 12126 3304 12131 3360
rect 10685 3302 12131 3304
rect 10685 3299 10751 3302
rect 12065 3299 12131 3302
rect 14774 3300 14780 3364
rect 14844 3362 14850 3364
rect 14844 3302 16682 3362
rect 14844 3300 14850 3302
rect 5392 3296 5712 3297
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 5392 3231 5712 3232
rect 9840 3296 10160 3297
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 9840 3231 10160 3232
rect 14288 3296 14608 3297
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 3231 14608 3232
rect 1342 3164 1348 3228
rect 1412 3226 1418 3228
rect 5809 3226 5875 3229
rect 7189 3226 7255 3229
rect 8201 3228 8267 3229
rect 8150 3226 8156 3228
rect 1412 3166 4722 3226
rect 1412 3164 1418 3166
rect 0 3090 800 3120
rect 3693 3090 3759 3093
rect 0 3088 3759 3090
rect 0 3032 3698 3088
rect 3754 3032 3759 3088
rect 0 3030 3759 3032
rect 4662 3090 4722 3166
rect 5809 3224 7255 3226
rect 5809 3168 5814 3224
rect 5870 3168 7194 3224
rect 7250 3168 7255 3224
rect 5809 3166 7255 3168
rect 8110 3166 8156 3226
rect 8220 3224 8267 3228
rect 8262 3168 8267 3224
rect 5809 3163 5875 3166
rect 7189 3163 7255 3166
rect 8150 3164 8156 3166
rect 8220 3164 8267 3168
rect 8201 3163 8267 3164
rect 10593 3226 10659 3229
rect 13537 3226 13603 3229
rect 10593 3224 13603 3226
rect 10593 3168 10598 3224
rect 10654 3168 13542 3224
rect 13598 3168 13603 3224
rect 10593 3166 13603 3168
rect 10593 3163 10659 3166
rect 13537 3163 13603 3166
rect 15377 3226 15443 3229
rect 15510 3226 15516 3228
rect 15377 3224 15516 3226
rect 15377 3168 15382 3224
rect 15438 3168 15516 3224
rect 15377 3166 15516 3168
rect 15377 3163 15443 3166
rect 15510 3164 15516 3166
rect 15580 3164 15586 3228
rect 15694 3164 15700 3228
rect 15764 3226 15770 3228
rect 16113 3226 16179 3229
rect 15764 3224 16179 3226
rect 15764 3168 16118 3224
rect 16174 3168 16179 3224
rect 15764 3166 16179 3168
rect 16622 3226 16682 3302
rect 19200 3226 20000 3256
rect 16622 3166 20000 3226
rect 15764 3164 15770 3166
rect 16113 3163 16179 3166
rect 19200 3136 20000 3166
rect 6729 3090 6795 3093
rect 4662 3088 6795 3090
rect 4662 3032 6734 3088
rect 6790 3032 6795 3088
rect 4662 3030 6795 3032
rect 0 3000 800 3030
rect 3693 3027 3759 3030
rect 6729 3027 6795 3030
rect 6913 3090 6979 3093
rect 12065 3090 12131 3093
rect 6913 3088 12131 3090
rect 6913 3032 6918 3088
rect 6974 3032 12070 3088
rect 12126 3032 12131 3088
rect 6913 3030 12131 3032
rect 6913 3027 6979 3030
rect 12065 3027 12131 3030
rect 14457 3090 14523 3093
rect 16205 3090 16271 3093
rect 14457 3088 16271 3090
rect 14457 3032 14462 3088
rect 14518 3032 16210 3088
rect 16266 3032 16271 3088
rect 14457 3030 16271 3032
rect 14457 3027 14523 3030
rect 16205 3027 16271 3030
rect 1393 2956 1459 2957
rect 1342 2954 1348 2956
rect 1302 2894 1348 2954
rect 1412 2952 1459 2956
rect 1454 2896 1459 2952
rect 1342 2892 1348 2894
rect 1412 2892 1459 2896
rect 1393 2891 1459 2892
rect 1761 2954 1827 2957
rect 10501 2954 10567 2957
rect 13997 2954 14063 2957
rect 1761 2952 10567 2954
rect 1761 2896 1766 2952
rect 1822 2896 10506 2952
rect 10562 2896 10567 2952
rect 1761 2894 10567 2896
rect 1761 2891 1827 2894
rect 10501 2891 10567 2894
rect 10734 2952 14063 2954
rect 10734 2896 14002 2952
rect 14058 2896 14063 2952
rect 10734 2894 14063 2896
rect 0 2818 800 2848
rect 2957 2818 3023 2821
rect 0 2816 3023 2818
rect 0 2760 2962 2816
rect 3018 2760 3023 2816
rect 0 2758 3023 2760
rect 0 2728 800 2758
rect 2957 2755 3023 2758
rect 3550 2756 3556 2820
rect 3620 2818 3626 2820
rect 3785 2818 3851 2821
rect 6913 2818 6979 2821
rect 3620 2816 6979 2818
rect 3620 2760 3790 2816
rect 3846 2760 6918 2816
rect 6974 2760 6979 2816
rect 3620 2758 6979 2760
rect 3620 2756 3626 2758
rect 3785 2755 3851 2758
rect 6913 2755 6979 2758
rect 7189 2818 7255 2821
rect 7414 2818 7420 2820
rect 7189 2816 7420 2818
rect 7189 2760 7194 2816
rect 7250 2760 7420 2816
rect 7189 2758 7420 2760
rect 7189 2755 7255 2758
rect 7414 2756 7420 2758
rect 7484 2756 7490 2820
rect 8150 2756 8156 2820
rect 8220 2818 8226 2820
rect 10734 2818 10794 2894
rect 13997 2891 14063 2894
rect 15469 2954 15535 2957
rect 15469 2952 17050 2954
rect 15469 2896 15474 2952
rect 15530 2896 17050 2952
rect 15469 2894 17050 2896
rect 15469 2891 15535 2894
rect 8220 2758 10794 2818
rect 14825 2818 14891 2821
rect 14958 2818 14964 2820
rect 14825 2816 14964 2818
rect 14825 2760 14830 2816
rect 14886 2760 14964 2816
rect 14825 2758 14964 2760
rect 8220 2756 8226 2758
rect 14825 2755 14891 2758
rect 14958 2756 14964 2758
rect 15028 2756 15034 2820
rect 16990 2818 17050 2894
rect 19200 2818 20000 2848
rect 16990 2758 20000 2818
rect 3168 2752 3488 2753
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2687 3488 2688
rect 7616 2752 7936 2753
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7616 2687 7936 2688
rect 12064 2752 12384 2753
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2687 12384 2688
rect 16512 2752 16832 2753
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 19200 2728 20000 2758
rect 16512 2687 16832 2688
rect 1158 2620 1164 2684
rect 1228 2682 1234 2684
rect 1761 2682 1827 2685
rect 1228 2680 1827 2682
rect 1228 2624 1766 2680
rect 1822 2624 1827 2680
rect 1228 2622 1827 2624
rect 1228 2620 1234 2622
rect 1761 2619 1827 2622
rect 3877 2682 3943 2685
rect 4102 2682 4108 2684
rect 3877 2680 4108 2682
rect 3877 2624 3882 2680
rect 3938 2624 4108 2680
rect 3877 2622 4108 2624
rect 3877 2619 3943 2622
rect 4102 2620 4108 2622
rect 4172 2620 4178 2684
rect 4337 2682 4403 2685
rect 6637 2682 6703 2685
rect 7097 2684 7163 2685
rect 7046 2682 7052 2684
rect 4337 2680 6703 2682
rect 4337 2624 4342 2680
rect 4398 2624 6642 2680
rect 6698 2624 6703 2680
rect 4337 2622 6703 2624
rect 7006 2622 7052 2682
rect 7116 2680 7163 2684
rect 7158 2624 7163 2680
rect 4337 2619 4403 2622
rect 6637 2619 6703 2622
rect 7046 2620 7052 2622
rect 7116 2620 7163 2624
rect 7097 2619 7163 2620
rect 8017 2682 8083 2685
rect 8017 2680 10794 2682
rect 8017 2624 8022 2680
rect 8078 2624 10794 2680
rect 8017 2622 10794 2624
rect 8017 2619 8083 2622
rect 974 2484 980 2548
rect 1044 2546 1050 2548
rect 6177 2546 6243 2549
rect 1044 2544 6243 2546
rect 1044 2488 6182 2544
rect 6238 2488 6243 2544
rect 1044 2486 6243 2488
rect 1044 2484 1050 2486
rect 6177 2483 6243 2486
rect 6637 2546 6703 2549
rect 10542 2546 10548 2548
rect 6637 2544 10548 2546
rect 6637 2488 6642 2544
rect 6698 2488 10548 2544
rect 6637 2486 10548 2488
rect 6637 2483 6703 2486
rect 10542 2484 10548 2486
rect 10612 2484 10618 2548
rect 10734 2546 10794 2622
rect 18045 2546 18111 2549
rect 10734 2544 18111 2546
rect 10734 2488 18050 2544
rect 18106 2488 18111 2544
rect 10734 2486 18111 2488
rect 18045 2483 18111 2486
rect 0 2410 800 2440
rect 18229 2410 18295 2413
rect 0 2408 18295 2410
rect 0 2352 18234 2408
rect 18290 2352 18295 2408
rect 0 2350 18295 2352
rect 0 2320 800 2350
rect 18229 2347 18295 2350
rect 18781 2410 18847 2413
rect 19200 2410 20000 2440
rect 18781 2408 20000 2410
rect 18781 2352 18786 2408
rect 18842 2352 20000 2408
rect 18781 2350 20000 2352
rect 18781 2347 18847 2350
rect 19200 2320 20000 2350
rect 4286 2212 4292 2276
rect 4356 2274 4362 2276
rect 4889 2274 4955 2277
rect 4356 2272 4955 2274
rect 4356 2216 4894 2272
rect 4950 2216 4955 2272
rect 4356 2214 4955 2216
rect 4356 2212 4362 2214
rect 4889 2211 4955 2214
rect 8477 2276 8543 2277
rect 8477 2272 8524 2276
rect 8588 2274 8594 2276
rect 8477 2216 8482 2272
rect 8477 2212 8524 2216
rect 8588 2214 8634 2274
rect 8588 2212 8594 2214
rect 8477 2211 8543 2212
rect 5392 2208 5712 2209
rect 0 2138 800 2168
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2143 5712 2144
rect 9840 2208 10160 2209
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2143 10160 2144
rect 14288 2208 14608 2209
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2143 14608 2144
rect 5257 2138 5323 2141
rect 0 2136 5323 2138
rect 0 2080 5262 2136
rect 5318 2080 5323 2136
rect 0 2078 5323 2080
rect 0 2048 800 2078
rect 5257 2075 5323 2078
rect 18321 2138 18387 2141
rect 19200 2138 20000 2168
rect 18321 2136 20000 2138
rect 18321 2080 18326 2136
rect 18382 2080 20000 2136
rect 18321 2078 20000 2080
rect 18321 2075 18387 2078
rect 19200 2048 20000 2078
rect 3417 2002 3483 2005
rect 11881 2002 11947 2005
rect 3417 2000 11947 2002
rect 3417 1944 3422 2000
rect 3478 1944 11886 2000
rect 11942 1944 11947 2000
rect 3417 1942 11947 1944
rect 3417 1939 3483 1942
rect 11881 1939 11947 1942
rect 0 1866 800 1896
rect 4061 1866 4127 1869
rect 0 1864 4127 1866
rect 0 1808 4066 1864
rect 4122 1808 4127 1864
rect 0 1806 4127 1808
rect 0 1776 800 1806
rect 4061 1803 4127 1806
rect 11830 1804 11836 1868
rect 11900 1866 11906 1868
rect 17953 1866 18019 1869
rect 11900 1864 18019 1866
rect 11900 1808 17958 1864
rect 18014 1808 18019 1864
rect 11900 1806 18019 1808
rect 11900 1804 11906 1806
rect 17953 1803 18019 1806
rect 5257 1730 5323 1733
rect 15929 1730 15995 1733
rect 5257 1728 15995 1730
rect 5257 1672 5262 1728
rect 5318 1672 15934 1728
rect 15990 1672 15995 1728
rect 5257 1670 15995 1672
rect 5257 1667 5323 1670
rect 15929 1667 15995 1670
rect 17493 1730 17559 1733
rect 19200 1730 20000 1760
rect 17493 1728 20000 1730
rect 17493 1672 17498 1728
rect 17554 1672 20000 1728
rect 17493 1670 20000 1672
rect 17493 1667 17559 1670
rect 19200 1640 20000 1670
rect 9489 1594 9555 1597
rect 17309 1594 17375 1597
rect 9489 1592 17375 1594
rect 9489 1536 9494 1592
rect 9550 1536 17314 1592
rect 17370 1536 17375 1592
rect 9489 1534 17375 1536
rect 9489 1531 9555 1534
rect 17309 1531 17375 1534
rect 0 1458 800 1488
rect 4061 1458 4127 1461
rect 0 1456 4127 1458
rect 0 1400 4066 1456
rect 4122 1400 4127 1456
rect 0 1398 4127 1400
rect 0 1368 800 1398
rect 4061 1395 4127 1398
rect 5809 1458 5875 1461
rect 12525 1458 12591 1461
rect 5809 1456 12591 1458
rect 5809 1400 5814 1456
rect 5870 1400 12530 1456
rect 12586 1400 12591 1456
rect 5809 1398 12591 1400
rect 5809 1395 5875 1398
rect 12525 1395 12591 1398
rect 15929 1322 15995 1325
rect 19200 1322 20000 1352
rect 15929 1320 20000 1322
rect 15929 1264 15934 1320
rect 15990 1264 20000 1320
rect 15929 1262 20000 1264
rect 15929 1259 15995 1262
rect 19200 1232 20000 1262
rect 0 1186 800 1216
rect 4061 1186 4127 1189
rect 0 1184 4127 1186
rect 0 1128 4066 1184
rect 4122 1128 4127 1184
rect 0 1126 4127 1128
rect 0 1096 800 1126
rect 4061 1123 4127 1126
rect 16941 914 17007 917
rect 19200 914 20000 944
rect 16941 912 20000 914
rect 16941 856 16946 912
rect 17002 856 20000 912
rect 16941 854 20000 856
rect 16941 851 17007 854
rect 19200 824 20000 854
rect 0 778 800 808
rect 3417 778 3483 781
rect 0 776 3483 778
rect 0 720 3422 776
rect 3478 720 3483 776
rect 0 718 3483 720
rect 0 688 800 718
rect 3417 715 3483 718
rect 0 506 800 536
rect 3693 506 3759 509
rect 0 504 3759 506
rect 0 448 3698 504
rect 3754 448 3759 504
rect 0 446 3759 448
rect 0 416 800 446
rect 3693 443 3759 446
rect 15837 506 15903 509
rect 19200 506 20000 536
rect 15837 504 20000 506
rect 15837 448 15842 504
rect 15898 448 20000 504
rect 15837 446 20000 448
rect 15837 443 15903 446
rect 19200 416 20000 446
rect 0 234 800 264
rect 1485 234 1551 237
rect 0 232 1551 234
rect 0 176 1490 232
rect 1546 176 1551 232
rect 0 174 1551 176
rect 0 144 800 174
rect 1485 171 1551 174
rect 15193 234 15259 237
rect 19200 234 20000 264
rect 15193 232 20000 234
rect 15193 176 15198 232
rect 15254 176 20000 232
rect 15193 174 20000 176
rect 15193 171 15259 174
rect 19200 144 20000 174
<< via3 >>
rect 980 15812 1044 15876
rect 12756 15812 12820 15876
rect 1164 15676 1228 15740
rect 9444 15676 9508 15740
rect 2636 15404 2700 15468
rect 12572 15404 12636 15468
rect 10916 14996 10980 15060
rect 16068 14860 16132 14924
rect 3176 14716 3240 14720
rect 3176 14660 3180 14716
rect 3180 14660 3236 14716
rect 3236 14660 3240 14716
rect 3176 14656 3240 14660
rect 3256 14716 3320 14720
rect 3256 14660 3260 14716
rect 3260 14660 3316 14716
rect 3316 14660 3320 14716
rect 3256 14656 3320 14660
rect 3336 14716 3400 14720
rect 3336 14660 3340 14716
rect 3340 14660 3396 14716
rect 3396 14660 3400 14716
rect 3336 14656 3400 14660
rect 3416 14716 3480 14720
rect 3416 14660 3420 14716
rect 3420 14660 3476 14716
rect 3476 14660 3480 14716
rect 3416 14656 3480 14660
rect 7624 14716 7688 14720
rect 7624 14660 7628 14716
rect 7628 14660 7684 14716
rect 7684 14660 7688 14716
rect 7624 14656 7688 14660
rect 7704 14716 7768 14720
rect 7704 14660 7708 14716
rect 7708 14660 7764 14716
rect 7764 14660 7768 14716
rect 7704 14656 7768 14660
rect 7784 14716 7848 14720
rect 7784 14660 7788 14716
rect 7788 14660 7844 14716
rect 7844 14660 7848 14716
rect 7784 14656 7848 14660
rect 7864 14716 7928 14720
rect 7864 14660 7868 14716
rect 7868 14660 7924 14716
rect 7924 14660 7928 14716
rect 7864 14656 7928 14660
rect 12072 14716 12136 14720
rect 12072 14660 12076 14716
rect 12076 14660 12132 14716
rect 12132 14660 12136 14716
rect 12072 14656 12136 14660
rect 12152 14716 12216 14720
rect 12152 14660 12156 14716
rect 12156 14660 12212 14716
rect 12212 14660 12216 14716
rect 12152 14656 12216 14660
rect 12232 14716 12296 14720
rect 12232 14660 12236 14716
rect 12236 14660 12292 14716
rect 12292 14660 12296 14716
rect 12232 14656 12296 14660
rect 12312 14716 12376 14720
rect 12312 14660 12316 14716
rect 12316 14660 12372 14716
rect 12372 14660 12376 14716
rect 12312 14656 12376 14660
rect 16520 14716 16584 14720
rect 16520 14660 16524 14716
rect 16524 14660 16580 14716
rect 16580 14660 16584 14716
rect 16520 14656 16584 14660
rect 16600 14716 16664 14720
rect 16600 14660 16604 14716
rect 16604 14660 16660 14716
rect 16660 14660 16664 14716
rect 16600 14656 16664 14660
rect 16680 14716 16744 14720
rect 16680 14660 16684 14716
rect 16684 14660 16740 14716
rect 16740 14660 16744 14716
rect 16680 14656 16744 14660
rect 16760 14716 16824 14720
rect 16760 14660 16764 14716
rect 16764 14660 16820 14716
rect 16820 14660 16824 14716
rect 16760 14656 16824 14660
rect 4476 14588 4540 14652
rect 10732 14588 10796 14652
rect 10364 14316 10428 14380
rect 16252 14180 16316 14244
rect 5400 14172 5464 14176
rect 5400 14116 5404 14172
rect 5404 14116 5460 14172
rect 5460 14116 5464 14172
rect 5400 14112 5464 14116
rect 5480 14172 5544 14176
rect 5480 14116 5484 14172
rect 5484 14116 5540 14172
rect 5540 14116 5544 14172
rect 5480 14112 5544 14116
rect 5560 14172 5624 14176
rect 5560 14116 5564 14172
rect 5564 14116 5620 14172
rect 5620 14116 5624 14172
rect 5560 14112 5624 14116
rect 5640 14172 5704 14176
rect 5640 14116 5644 14172
rect 5644 14116 5700 14172
rect 5700 14116 5704 14172
rect 5640 14112 5704 14116
rect 9848 14172 9912 14176
rect 9848 14116 9852 14172
rect 9852 14116 9908 14172
rect 9908 14116 9912 14172
rect 9848 14112 9912 14116
rect 9928 14172 9992 14176
rect 9928 14116 9932 14172
rect 9932 14116 9988 14172
rect 9988 14116 9992 14172
rect 9928 14112 9992 14116
rect 10008 14172 10072 14176
rect 10008 14116 10012 14172
rect 10012 14116 10068 14172
rect 10068 14116 10072 14172
rect 10008 14112 10072 14116
rect 10088 14172 10152 14176
rect 10088 14116 10092 14172
rect 10092 14116 10148 14172
rect 10148 14116 10152 14172
rect 10088 14112 10152 14116
rect 14296 14172 14360 14176
rect 14296 14116 14300 14172
rect 14300 14116 14356 14172
rect 14356 14116 14360 14172
rect 14296 14112 14360 14116
rect 14376 14172 14440 14176
rect 14376 14116 14380 14172
rect 14380 14116 14436 14172
rect 14436 14116 14440 14172
rect 14376 14112 14440 14116
rect 14456 14172 14520 14176
rect 14456 14116 14460 14172
rect 14460 14116 14516 14172
rect 14516 14116 14520 14172
rect 14456 14112 14520 14116
rect 14536 14172 14600 14176
rect 14536 14116 14540 14172
rect 14540 14116 14596 14172
rect 14596 14116 14600 14172
rect 14536 14112 14600 14116
rect 10548 14104 10612 14108
rect 10548 14048 10598 14104
rect 10598 14048 10612 14104
rect 10548 14044 10612 14048
rect 17356 14044 17420 14108
rect 14044 13772 14108 13836
rect 15516 13772 15580 13836
rect 3556 13636 3620 13700
rect 5028 13636 5092 13700
rect 3176 13628 3240 13632
rect 3176 13572 3180 13628
rect 3180 13572 3236 13628
rect 3236 13572 3240 13628
rect 3176 13568 3240 13572
rect 3256 13628 3320 13632
rect 3256 13572 3260 13628
rect 3260 13572 3316 13628
rect 3316 13572 3320 13628
rect 3256 13568 3320 13572
rect 3336 13628 3400 13632
rect 3336 13572 3340 13628
rect 3340 13572 3396 13628
rect 3396 13572 3400 13628
rect 3336 13568 3400 13572
rect 3416 13628 3480 13632
rect 3416 13572 3420 13628
rect 3420 13572 3476 13628
rect 3476 13572 3480 13628
rect 3416 13568 3480 13572
rect 7624 13628 7688 13632
rect 7624 13572 7628 13628
rect 7628 13572 7684 13628
rect 7684 13572 7688 13628
rect 7624 13568 7688 13572
rect 7704 13628 7768 13632
rect 7704 13572 7708 13628
rect 7708 13572 7764 13628
rect 7764 13572 7768 13628
rect 7704 13568 7768 13572
rect 7784 13628 7848 13632
rect 7784 13572 7788 13628
rect 7788 13572 7844 13628
rect 7844 13572 7848 13628
rect 7784 13568 7848 13572
rect 7864 13628 7928 13632
rect 7864 13572 7868 13628
rect 7868 13572 7924 13628
rect 7924 13572 7928 13628
rect 7864 13568 7928 13572
rect 12072 13628 12136 13632
rect 12072 13572 12076 13628
rect 12076 13572 12132 13628
rect 12132 13572 12136 13628
rect 12072 13568 12136 13572
rect 12152 13628 12216 13632
rect 12152 13572 12156 13628
rect 12156 13572 12212 13628
rect 12212 13572 12216 13628
rect 12152 13568 12216 13572
rect 12232 13628 12296 13632
rect 12232 13572 12236 13628
rect 12236 13572 12292 13628
rect 12292 13572 12296 13628
rect 12232 13568 12296 13572
rect 12312 13628 12376 13632
rect 12312 13572 12316 13628
rect 12316 13572 12372 13628
rect 12372 13572 12376 13628
rect 12312 13568 12376 13572
rect 16520 13628 16584 13632
rect 16520 13572 16524 13628
rect 16524 13572 16580 13628
rect 16580 13572 16584 13628
rect 16520 13568 16584 13572
rect 16600 13628 16664 13632
rect 16600 13572 16604 13628
rect 16604 13572 16660 13628
rect 16660 13572 16664 13628
rect 16600 13568 16664 13572
rect 16680 13628 16744 13632
rect 16680 13572 16684 13628
rect 16684 13572 16740 13628
rect 16740 13572 16744 13628
rect 16680 13568 16744 13572
rect 16760 13628 16824 13632
rect 16760 13572 16764 13628
rect 16764 13572 16820 13628
rect 16820 13572 16824 13628
rect 16760 13568 16824 13572
rect 14780 13500 14844 13564
rect 9444 13424 9508 13428
rect 9444 13368 9494 13424
rect 9494 13368 9508 13424
rect 9444 13364 9508 13368
rect 3556 13228 3620 13292
rect 3924 13228 3988 13292
rect 6684 13228 6748 13292
rect 11652 13228 11716 13292
rect 15700 13228 15764 13292
rect 2452 13092 2516 13156
rect 5400 13084 5464 13088
rect 5400 13028 5404 13084
rect 5404 13028 5460 13084
rect 5460 13028 5464 13084
rect 5400 13024 5464 13028
rect 5480 13084 5544 13088
rect 5480 13028 5484 13084
rect 5484 13028 5540 13084
rect 5540 13028 5544 13084
rect 5480 13024 5544 13028
rect 5560 13084 5624 13088
rect 5560 13028 5564 13084
rect 5564 13028 5620 13084
rect 5620 13028 5624 13084
rect 5560 13024 5624 13028
rect 5640 13084 5704 13088
rect 5640 13028 5644 13084
rect 5644 13028 5700 13084
rect 5700 13028 5704 13084
rect 5640 13024 5704 13028
rect 1348 12820 1412 12884
rect 3004 12880 3068 12884
rect 3004 12824 3054 12880
rect 3054 12824 3068 12880
rect 3004 12820 3068 12824
rect 4844 12880 4908 12884
rect 4844 12824 4894 12880
rect 4894 12824 4908 12880
rect 4844 12820 4908 12824
rect 5212 12820 5276 12884
rect 15332 13092 15396 13156
rect 9848 13084 9912 13088
rect 9848 13028 9852 13084
rect 9852 13028 9908 13084
rect 9908 13028 9912 13084
rect 9848 13024 9912 13028
rect 9928 13084 9992 13088
rect 9928 13028 9932 13084
rect 9932 13028 9988 13084
rect 9988 13028 9992 13084
rect 9928 13024 9992 13028
rect 10008 13084 10072 13088
rect 10008 13028 10012 13084
rect 10012 13028 10068 13084
rect 10068 13028 10072 13084
rect 10008 13024 10072 13028
rect 10088 13084 10152 13088
rect 10088 13028 10092 13084
rect 10092 13028 10148 13084
rect 10148 13028 10152 13084
rect 10088 13024 10152 13028
rect 14296 13084 14360 13088
rect 14296 13028 14300 13084
rect 14300 13028 14356 13084
rect 14356 13028 14360 13084
rect 14296 13024 14360 13028
rect 14376 13084 14440 13088
rect 14376 13028 14380 13084
rect 14380 13028 14436 13084
rect 14436 13028 14440 13084
rect 14376 13024 14440 13028
rect 14456 13084 14520 13088
rect 14456 13028 14460 13084
rect 14460 13028 14516 13084
rect 14516 13028 14520 13084
rect 14456 13024 14520 13028
rect 14536 13084 14600 13088
rect 14536 13028 14540 13084
rect 14540 13028 14596 13084
rect 14596 13028 14600 13084
rect 14536 13024 14600 13028
rect 13308 12956 13372 13020
rect 12940 12820 13004 12884
rect 13492 12820 13556 12884
rect 13676 12880 13740 12884
rect 13676 12824 13690 12880
rect 13690 12824 13740 12880
rect 13676 12820 13740 12824
rect 16988 12820 17052 12884
rect 8892 12684 8956 12748
rect 6316 12548 6380 12612
rect 6500 12548 6564 12612
rect 8156 12608 8220 12612
rect 8156 12552 8170 12608
rect 8170 12552 8220 12608
rect 8156 12548 8220 12552
rect 10548 12548 10612 12612
rect 11468 12548 11532 12612
rect 3176 12540 3240 12544
rect 3176 12484 3180 12540
rect 3180 12484 3236 12540
rect 3236 12484 3240 12540
rect 3176 12480 3240 12484
rect 3256 12540 3320 12544
rect 3256 12484 3260 12540
rect 3260 12484 3316 12540
rect 3316 12484 3320 12540
rect 3256 12480 3320 12484
rect 3336 12540 3400 12544
rect 3336 12484 3340 12540
rect 3340 12484 3396 12540
rect 3396 12484 3400 12540
rect 3336 12480 3400 12484
rect 3416 12540 3480 12544
rect 3416 12484 3420 12540
rect 3420 12484 3476 12540
rect 3476 12484 3480 12540
rect 3416 12480 3480 12484
rect 7624 12540 7688 12544
rect 7624 12484 7628 12540
rect 7628 12484 7684 12540
rect 7684 12484 7688 12540
rect 7624 12480 7688 12484
rect 7704 12540 7768 12544
rect 7704 12484 7708 12540
rect 7708 12484 7764 12540
rect 7764 12484 7768 12540
rect 7704 12480 7768 12484
rect 7784 12540 7848 12544
rect 7784 12484 7788 12540
rect 7788 12484 7844 12540
rect 7844 12484 7848 12540
rect 7784 12480 7848 12484
rect 7864 12540 7928 12544
rect 7864 12484 7868 12540
rect 7868 12484 7924 12540
rect 7924 12484 7928 12540
rect 7864 12480 7928 12484
rect 12072 12540 12136 12544
rect 12072 12484 12076 12540
rect 12076 12484 12132 12540
rect 12132 12484 12136 12540
rect 12072 12480 12136 12484
rect 12152 12540 12216 12544
rect 12152 12484 12156 12540
rect 12156 12484 12212 12540
rect 12212 12484 12216 12540
rect 12152 12480 12216 12484
rect 12232 12540 12296 12544
rect 12232 12484 12236 12540
rect 12236 12484 12292 12540
rect 12292 12484 12296 12540
rect 12232 12480 12296 12484
rect 12312 12540 12376 12544
rect 12312 12484 12316 12540
rect 12316 12484 12372 12540
rect 12372 12484 12376 12540
rect 12312 12480 12376 12484
rect 4108 12412 4172 12476
rect 7052 12472 7116 12476
rect 7052 12416 7066 12472
rect 7066 12416 7116 12472
rect 7052 12412 7116 12416
rect 7236 12276 7300 12340
rect 11100 12412 11164 12476
rect 15884 12548 15948 12612
rect 16520 12540 16584 12544
rect 16520 12484 16524 12540
rect 16524 12484 16580 12540
rect 16580 12484 16584 12540
rect 16520 12480 16584 12484
rect 16600 12540 16664 12544
rect 16600 12484 16604 12540
rect 16604 12484 16660 12540
rect 16660 12484 16664 12540
rect 16600 12480 16664 12484
rect 16680 12540 16744 12544
rect 16680 12484 16684 12540
rect 16684 12484 16740 12540
rect 16740 12484 16744 12540
rect 16680 12480 16744 12484
rect 16760 12540 16824 12544
rect 16760 12484 16764 12540
rect 16764 12484 16820 12540
rect 16820 12484 16824 12540
rect 16760 12480 16824 12484
rect 13492 12412 13556 12476
rect 14780 12412 14844 12476
rect 4108 12004 4172 12068
rect 8156 12004 8220 12068
rect 11284 12004 11348 12068
rect 13860 12064 13924 12068
rect 13860 12008 13874 12064
rect 13874 12008 13924 12064
rect 13860 12004 13924 12008
rect 5400 11996 5464 12000
rect 5400 11940 5404 11996
rect 5404 11940 5460 11996
rect 5460 11940 5464 11996
rect 5400 11936 5464 11940
rect 5480 11996 5544 12000
rect 5480 11940 5484 11996
rect 5484 11940 5540 11996
rect 5540 11940 5544 11996
rect 5480 11936 5544 11940
rect 5560 11996 5624 12000
rect 5560 11940 5564 11996
rect 5564 11940 5620 11996
rect 5620 11940 5624 11996
rect 5560 11936 5624 11940
rect 5640 11996 5704 12000
rect 5640 11940 5644 11996
rect 5644 11940 5700 11996
rect 5700 11940 5704 11996
rect 5640 11936 5704 11940
rect 9848 11996 9912 12000
rect 9848 11940 9852 11996
rect 9852 11940 9908 11996
rect 9908 11940 9912 11996
rect 9848 11936 9912 11940
rect 9928 11996 9992 12000
rect 9928 11940 9932 11996
rect 9932 11940 9988 11996
rect 9988 11940 9992 11996
rect 9928 11936 9992 11940
rect 10008 11996 10072 12000
rect 10008 11940 10012 11996
rect 10012 11940 10068 11996
rect 10068 11940 10072 11996
rect 10008 11936 10072 11940
rect 10088 11996 10152 12000
rect 10088 11940 10092 11996
rect 10092 11940 10148 11996
rect 10148 11940 10152 11996
rect 10088 11936 10152 11940
rect 2268 11868 2332 11932
rect 7420 11868 7484 11932
rect 14296 11996 14360 12000
rect 14296 11940 14300 11996
rect 14300 11940 14356 11996
rect 14356 11940 14360 11996
rect 14296 11936 14360 11940
rect 14376 11996 14440 12000
rect 14376 11940 14380 11996
rect 14380 11940 14436 11996
rect 14436 11940 14440 11996
rect 14376 11936 14440 11940
rect 14456 11996 14520 12000
rect 14456 11940 14460 11996
rect 14460 11940 14516 11996
rect 14516 11940 14520 11996
rect 14456 11936 14520 11940
rect 14536 11996 14600 12000
rect 14536 11940 14540 11996
rect 14540 11940 14596 11996
rect 14596 11940 14600 11996
rect 14536 11936 14600 11940
rect 13492 11868 13556 11932
rect 6868 11732 6932 11796
rect 9628 11732 9692 11796
rect 10732 11732 10796 11796
rect 11836 11732 11900 11796
rect 12572 11732 12636 11796
rect 15148 11732 15212 11796
rect 6132 11596 6196 11660
rect 10548 11460 10612 11524
rect 10916 11460 10980 11524
rect 12756 11460 12820 11524
rect 3176 11452 3240 11456
rect 3176 11396 3180 11452
rect 3180 11396 3236 11452
rect 3236 11396 3240 11452
rect 3176 11392 3240 11396
rect 3256 11452 3320 11456
rect 3256 11396 3260 11452
rect 3260 11396 3316 11452
rect 3316 11396 3320 11452
rect 3256 11392 3320 11396
rect 3336 11452 3400 11456
rect 3336 11396 3340 11452
rect 3340 11396 3396 11452
rect 3396 11396 3400 11452
rect 3336 11392 3400 11396
rect 3416 11452 3480 11456
rect 3416 11396 3420 11452
rect 3420 11396 3476 11452
rect 3476 11396 3480 11452
rect 3416 11392 3480 11396
rect 7624 11452 7688 11456
rect 7624 11396 7628 11452
rect 7628 11396 7684 11452
rect 7684 11396 7688 11452
rect 7624 11392 7688 11396
rect 7704 11452 7768 11456
rect 7704 11396 7708 11452
rect 7708 11396 7764 11452
rect 7764 11396 7768 11452
rect 7704 11392 7768 11396
rect 7784 11452 7848 11456
rect 7784 11396 7788 11452
rect 7788 11396 7844 11452
rect 7844 11396 7848 11452
rect 7784 11392 7848 11396
rect 7864 11452 7928 11456
rect 7864 11396 7868 11452
rect 7868 11396 7924 11452
rect 7924 11396 7928 11452
rect 7864 11392 7928 11396
rect 12072 11452 12136 11456
rect 12072 11396 12076 11452
rect 12076 11396 12132 11452
rect 12132 11396 12136 11452
rect 12072 11392 12136 11396
rect 12152 11452 12216 11456
rect 12152 11396 12156 11452
rect 12156 11396 12212 11452
rect 12212 11396 12216 11452
rect 12152 11392 12216 11396
rect 12232 11452 12296 11456
rect 12232 11396 12236 11452
rect 12236 11396 12292 11452
rect 12292 11396 12296 11452
rect 12232 11392 12296 11396
rect 12312 11452 12376 11456
rect 12312 11396 12316 11452
rect 12316 11396 12372 11452
rect 12372 11396 12376 11452
rect 12312 11392 12376 11396
rect 2084 11052 2148 11116
rect 5948 11188 6012 11252
rect 13124 11324 13188 11388
rect 14964 11460 15028 11524
rect 16520 11452 16584 11456
rect 16520 11396 16524 11452
rect 16524 11396 16580 11452
rect 16580 11396 16584 11452
rect 16520 11392 16584 11396
rect 16600 11452 16664 11456
rect 16600 11396 16604 11452
rect 16604 11396 16660 11452
rect 16660 11396 16664 11452
rect 16600 11392 16664 11396
rect 16680 11452 16744 11456
rect 16680 11396 16684 11452
rect 16684 11396 16740 11452
rect 16740 11396 16744 11452
rect 16680 11392 16744 11396
rect 16760 11452 16824 11456
rect 16760 11396 16764 11452
rect 16764 11396 16820 11452
rect 16820 11396 16824 11452
rect 16760 11392 16824 11396
rect 9444 11188 9508 11252
rect 8524 11052 8588 11116
rect 11652 11052 11716 11116
rect 5400 10908 5464 10912
rect 5400 10852 5404 10908
rect 5404 10852 5460 10908
rect 5460 10852 5464 10908
rect 5400 10848 5464 10852
rect 5480 10908 5544 10912
rect 5480 10852 5484 10908
rect 5484 10852 5540 10908
rect 5540 10852 5544 10908
rect 5480 10848 5544 10852
rect 5560 10908 5624 10912
rect 5560 10852 5564 10908
rect 5564 10852 5620 10908
rect 5620 10852 5624 10908
rect 5560 10848 5624 10852
rect 5640 10908 5704 10912
rect 5640 10852 5644 10908
rect 5644 10852 5700 10908
rect 5700 10852 5704 10908
rect 5640 10848 5704 10852
rect 9848 10908 9912 10912
rect 9848 10852 9852 10908
rect 9852 10852 9908 10908
rect 9908 10852 9912 10908
rect 9848 10848 9912 10852
rect 9928 10908 9992 10912
rect 9928 10852 9932 10908
rect 9932 10852 9988 10908
rect 9988 10852 9992 10908
rect 9928 10848 9992 10852
rect 10008 10908 10072 10912
rect 10008 10852 10012 10908
rect 10012 10852 10068 10908
rect 10068 10852 10072 10908
rect 10008 10848 10072 10852
rect 10088 10908 10152 10912
rect 10088 10852 10092 10908
rect 10092 10852 10148 10908
rect 10148 10852 10152 10908
rect 10088 10848 10152 10852
rect 14296 10908 14360 10912
rect 14296 10852 14300 10908
rect 14300 10852 14356 10908
rect 14356 10852 14360 10908
rect 14296 10848 14360 10852
rect 14376 10908 14440 10912
rect 14376 10852 14380 10908
rect 14380 10852 14436 10908
rect 14436 10852 14440 10908
rect 14376 10848 14440 10852
rect 14456 10908 14520 10912
rect 14456 10852 14460 10908
rect 14460 10852 14516 10908
rect 14516 10852 14520 10908
rect 14456 10848 14520 10852
rect 14536 10908 14600 10912
rect 14536 10852 14540 10908
rect 14540 10852 14596 10908
rect 14596 10852 14600 10908
rect 14536 10848 14600 10852
rect 2636 10780 2700 10844
rect 2820 10644 2884 10708
rect 3556 10644 3620 10708
rect 7236 10508 7300 10572
rect 11100 10508 11164 10572
rect 11652 10508 11716 10572
rect 13308 10508 13372 10572
rect 3176 10364 3240 10368
rect 3176 10308 3180 10364
rect 3180 10308 3236 10364
rect 3236 10308 3240 10364
rect 3176 10304 3240 10308
rect 3256 10364 3320 10368
rect 3256 10308 3260 10364
rect 3260 10308 3316 10364
rect 3316 10308 3320 10364
rect 3256 10304 3320 10308
rect 3336 10364 3400 10368
rect 3336 10308 3340 10364
rect 3340 10308 3396 10364
rect 3396 10308 3400 10364
rect 3336 10304 3400 10308
rect 3416 10364 3480 10368
rect 3416 10308 3420 10364
rect 3420 10308 3476 10364
rect 3476 10308 3480 10364
rect 3416 10304 3480 10308
rect 7624 10364 7688 10368
rect 7624 10308 7628 10364
rect 7628 10308 7684 10364
rect 7684 10308 7688 10364
rect 7624 10304 7688 10308
rect 7704 10364 7768 10368
rect 7704 10308 7708 10364
rect 7708 10308 7764 10364
rect 7764 10308 7768 10364
rect 7704 10304 7768 10308
rect 7784 10364 7848 10368
rect 7784 10308 7788 10364
rect 7788 10308 7844 10364
rect 7844 10308 7848 10364
rect 7784 10304 7848 10308
rect 7864 10364 7928 10368
rect 7864 10308 7868 10364
rect 7868 10308 7924 10364
rect 7924 10308 7928 10364
rect 7864 10304 7928 10308
rect 7420 10236 7484 10300
rect 612 10134 676 10198
rect 6684 9828 6748 9892
rect 7420 9828 7484 9892
rect 16068 10372 16132 10436
rect 12072 10364 12136 10368
rect 12072 10308 12076 10364
rect 12076 10308 12132 10364
rect 12132 10308 12136 10364
rect 12072 10304 12136 10308
rect 12152 10364 12216 10368
rect 12152 10308 12156 10364
rect 12156 10308 12212 10364
rect 12212 10308 12216 10364
rect 12152 10304 12216 10308
rect 12232 10364 12296 10368
rect 12232 10308 12236 10364
rect 12236 10308 12292 10364
rect 12292 10308 12296 10364
rect 12232 10304 12296 10308
rect 12312 10364 12376 10368
rect 12312 10308 12316 10364
rect 12316 10308 12372 10364
rect 12372 10308 12376 10364
rect 12312 10304 12376 10308
rect 16520 10364 16584 10368
rect 16520 10308 16524 10364
rect 16524 10308 16580 10364
rect 16580 10308 16584 10364
rect 16520 10304 16584 10308
rect 16600 10364 16664 10368
rect 16600 10308 16604 10364
rect 16604 10308 16660 10364
rect 16660 10308 16664 10364
rect 16600 10304 16664 10308
rect 16680 10364 16744 10368
rect 16680 10308 16684 10364
rect 16684 10308 16740 10364
rect 16740 10308 16744 10364
rect 16680 10304 16744 10308
rect 16760 10364 16824 10368
rect 16760 10308 16764 10364
rect 16764 10308 16820 10364
rect 16820 10308 16824 10364
rect 16760 10304 16824 10308
rect 11468 10296 11532 10300
rect 11468 10240 11518 10296
rect 11518 10240 11532 10296
rect 11468 10236 11532 10240
rect 11284 10100 11348 10164
rect 15332 10100 15396 10164
rect 5400 9820 5464 9824
rect 5400 9764 5404 9820
rect 5404 9764 5460 9820
rect 5460 9764 5464 9820
rect 5400 9760 5464 9764
rect 5480 9820 5544 9824
rect 5480 9764 5484 9820
rect 5484 9764 5540 9820
rect 5540 9764 5544 9820
rect 5480 9760 5544 9764
rect 5560 9820 5624 9824
rect 5560 9764 5564 9820
rect 5564 9764 5620 9820
rect 5620 9764 5624 9820
rect 5560 9760 5624 9764
rect 5640 9820 5704 9824
rect 5640 9764 5644 9820
rect 5644 9764 5700 9820
rect 5700 9764 5704 9820
rect 5640 9760 5704 9764
rect 4292 9692 4356 9756
rect 6500 9692 6564 9756
rect 9848 9820 9912 9824
rect 9848 9764 9852 9820
rect 9852 9764 9908 9820
rect 9908 9764 9912 9820
rect 9848 9760 9912 9764
rect 9928 9820 9992 9824
rect 9928 9764 9932 9820
rect 9932 9764 9988 9820
rect 9988 9764 9992 9820
rect 9928 9760 9992 9764
rect 10008 9820 10072 9824
rect 10008 9764 10012 9820
rect 10012 9764 10068 9820
rect 10068 9764 10072 9820
rect 10008 9760 10072 9764
rect 10088 9820 10152 9824
rect 10088 9764 10092 9820
rect 10092 9764 10148 9820
rect 10148 9764 10152 9820
rect 10088 9760 10152 9764
rect 8156 9692 8220 9756
rect 11652 9828 11716 9892
rect 14296 9820 14360 9824
rect 14296 9764 14300 9820
rect 14300 9764 14356 9820
rect 14356 9764 14360 9820
rect 14296 9760 14360 9764
rect 14376 9820 14440 9824
rect 14376 9764 14380 9820
rect 14380 9764 14436 9820
rect 14436 9764 14440 9820
rect 14376 9760 14440 9764
rect 14456 9820 14520 9824
rect 14456 9764 14460 9820
rect 14460 9764 14516 9820
rect 14516 9764 14520 9820
rect 14456 9760 14520 9764
rect 14536 9820 14600 9824
rect 14536 9764 14540 9820
rect 14540 9764 14596 9820
rect 14596 9764 14600 9820
rect 14536 9760 14600 9764
rect 11468 9692 11532 9756
rect 11836 9692 11900 9756
rect 16068 9692 16132 9756
rect 6132 9556 6196 9620
rect 14044 9420 14108 9484
rect 4108 9284 4172 9348
rect 3176 9276 3240 9280
rect 3176 9220 3180 9276
rect 3180 9220 3236 9276
rect 3236 9220 3240 9276
rect 3176 9216 3240 9220
rect 3256 9276 3320 9280
rect 3256 9220 3260 9276
rect 3260 9220 3316 9276
rect 3316 9220 3320 9276
rect 3256 9216 3320 9220
rect 3336 9276 3400 9280
rect 3336 9220 3340 9276
rect 3340 9220 3396 9276
rect 3396 9220 3400 9276
rect 3336 9216 3400 9220
rect 3416 9276 3480 9280
rect 3416 9220 3420 9276
rect 3420 9220 3476 9276
rect 3476 9220 3480 9276
rect 3416 9216 3480 9220
rect 7624 9276 7688 9280
rect 7624 9220 7628 9276
rect 7628 9220 7684 9276
rect 7684 9220 7688 9276
rect 7624 9216 7688 9220
rect 7704 9276 7768 9280
rect 7704 9220 7708 9276
rect 7708 9220 7764 9276
rect 7764 9220 7768 9276
rect 7704 9216 7768 9220
rect 7784 9276 7848 9280
rect 7784 9220 7788 9276
rect 7788 9220 7844 9276
rect 7844 9220 7848 9276
rect 7784 9216 7848 9220
rect 7864 9276 7928 9280
rect 7864 9220 7868 9276
rect 7868 9220 7924 9276
rect 7924 9220 7928 9276
rect 7864 9216 7928 9220
rect 12072 9276 12136 9280
rect 12072 9220 12076 9276
rect 12076 9220 12132 9276
rect 12132 9220 12136 9276
rect 12072 9216 12136 9220
rect 12152 9276 12216 9280
rect 12152 9220 12156 9276
rect 12156 9220 12212 9276
rect 12212 9220 12216 9276
rect 12152 9216 12216 9220
rect 12232 9276 12296 9280
rect 12232 9220 12236 9276
rect 12236 9220 12292 9276
rect 12292 9220 12296 9276
rect 12232 9216 12296 9220
rect 12312 9276 12376 9280
rect 12312 9220 12316 9276
rect 12316 9220 12372 9276
rect 12372 9220 12376 9276
rect 12312 9216 12376 9220
rect 16520 9276 16584 9280
rect 16520 9220 16524 9276
rect 16524 9220 16580 9276
rect 16580 9220 16584 9276
rect 16520 9216 16584 9220
rect 16600 9276 16664 9280
rect 16600 9220 16604 9276
rect 16604 9220 16660 9276
rect 16660 9220 16664 9276
rect 16600 9216 16664 9220
rect 16680 9276 16744 9280
rect 16680 9220 16684 9276
rect 16684 9220 16740 9276
rect 16740 9220 16744 9276
rect 16680 9216 16744 9220
rect 16760 9276 16824 9280
rect 16760 9220 16764 9276
rect 16764 9220 16820 9276
rect 16820 9220 16824 9276
rect 16760 9216 16824 9220
rect 7052 9148 7116 9212
rect 10732 9208 10796 9212
rect 10732 9152 10746 9208
rect 10746 9152 10796 9208
rect 10732 9148 10796 9152
rect 3740 9072 3804 9076
rect 3740 9016 3754 9072
rect 3754 9016 3804 9072
rect 3740 9012 3804 9016
rect 12940 9012 13004 9076
rect 13492 9012 13556 9076
rect 2820 8876 2884 8940
rect 6868 8876 6932 8940
rect 7420 8876 7484 8940
rect 13492 8876 13556 8940
rect 5400 8732 5464 8736
rect 5400 8676 5404 8732
rect 5404 8676 5460 8732
rect 5460 8676 5464 8732
rect 5400 8672 5464 8676
rect 5480 8732 5544 8736
rect 5480 8676 5484 8732
rect 5484 8676 5540 8732
rect 5540 8676 5544 8732
rect 5480 8672 5544 8676
rect 5560 8732 5624 8736
rect 5560 8676 5564 8732
rect 5564 8676 5620 8732
rect 5620 8676 5624 8732
rect 5560 8672 5624 8676
rect 5640 8732 5704 8736
rect 5640 8676 5644 8732
rect 5644 8676 5700 8732
rect 5700 8676 5704 8732
rect 5640 8672 5704 8676
rect 9848 8732 9912 8736
rect 9848 8676 9852 8732
rect 9852 8676 9908 8732
rect 9908 8676 9912 8732
rect 9848 8672 9912 8676
rect 9928 8732 9992 8736
rect 9928 8676 9932 8732
rect 9932 8676 9988 8732
rect 9988 8676 9992 8732
rect 9928 8672 9992 8676
rect 10008 8732 10072 8736
rect 10008 8676 10012 8732
rect 10012 8676 10068 8732
rect 10068 8676 10072 8732
rect 10008 8672 10072 8676
rect 10088 8732 10152 8736
rect 10088 8676 10092 8732
rect 10092 8676 10148 8732
rect 10148 8676 10152 8732
rect 10088 8672 10152 8676
rect 14296 8732 14360 8736
rect 14296 8676 14300 8732
rect 14300 8676 14356 8732
rect 14356 8676 14360 8732
rect 14296 8672 14360 8676
rect 14376 8732 14440 8736
rect 14376 8676 14380 8732
rect 14380 8676 14436 8732
rect 14436 8676 14440 8732
rect 14376 8672 14440 8676
rect 14456 8732 14520 8736
rect 14456 8676 14460 8732
rect 14460 8676 14516 8732
rect 14516 8676 14520 8732
rect 14456 8672 14520 8676
rect 14536 8732 14600 8736
rect 14536 8676 14540 8732
rect 14540 8676 14596 8732
rect 14596 8676 14600 8732
rect 14536 8672 14600 8676
rect 5212 8664 5276 8668
rect 5212 8608 5262 8664
rect 5262 8608 5276 8664
rect 5212 8604 5276 8608
rect 3740 8332 3804 8396
rect 3924 8392 3988 8396
rect 3924 8336 3974 8392
rect 3974 8336 3988 8392
rect 3924 8332 3988 8336
rect 8156 8332 8220 8396
rect 11836 8392 11900 8396
rect 11836 8336 11886 8392
rect 11886 8336 11900 8392
rect 11836 8332 11900 8336
rect 13676 8332 13740 8396
rect 15700 8332 15764 8396
rect 17172 8332 17236 8396
rect 2636 8256 2700 8260
rect 2636 8200 2650 8256
rect 2650 8200 2700 8256
rect 2636 8196 2700 8200
rect 2820 8256 2884 8260
rect 2820 8200 2834 8256
rect 2834 8200 2884 8256
rect 2820 8196 2884 8200
rect 3740 8196 3804 8260
rect 7420 8256 7484 8260
rect 7420 8200 7470 8256
rect 7470 8200 7484 8256
rect 7420 8196 7484 8200
rect 3176 8188 3240 8192
rect 3176 8132 3180 8188
rect 3180 8132 3236 8188
rect 3236 8132 3240 8188
rect 3176 8128 3240 8132
rect 3256 8188 3320 8192
rect 3256 8132 3260 8188
rect 3260 8132 3316 8188
rect 3316 8132 3320 8188
rect 3256 8128 3320 8132
rect 3336 8188 3400 8192
rect 3336 8132 3340 8188
rect 3340 8132 3396 8188
rect 3396 8132 3400 8188
rect 3336 8128 3400 8132
rect 3416 8188 3480 8192
rect 3416 8132 3420 8188
rect 3420 8132 3476 8188
rect 3476 8132 3480 8188
rect 3416 8128 3480 8132
rect 7624 8188 7688 8192
rect 7624 8132 7628 8188
rect 7628 8132 7684 8188
rect 7684 8132 7688 8188
rect 7624 8128 7688 8132
rect 7704 8188 7768 8192
rect 7704 8132 7708 8188
rect 7708 8132 7764 8188
rect 7764 8132 7768 8188
rect 7704 8128 7768 8132
rect 7784 8188 7848 8192
rect 7784 8132 7788 8188
rect 7788 8132 7844 8188
rect 7844 8132 7848 8188
rect 7784 8128 7848 8132
rect 7864 8188 7928 8192
rect 7864 8132 7868 8188
rect 7868 8132 7924 8188
rect 7924 8132 7928 8188
rect 7864 8128 7928 8132
rect 12072 8188 12136 8192
rect 12072 8132 12076 8188
rect 12076 8132 12132 8188
rect 12132 8132 12136 8188
rect 12072 8128 12136 8132
rect 12152 8188 12216 8192
rect 12152 8132 12156 8188
rect 12156 8132 12212 8188
rect 12212 8132 12216 8188
rect 12152 8128 12216 8132
rect 12232 8188 12296 8192
rect 12232 8132 12236 8188
rect 12236 8132 12292 8188
rect 12292 8132 12296 8188
rect 12232 8128 12296 8132
rect 12312 8188 12376 8192
rect 12312 8132 12316 8188
rect 12316 8132 12372 8188
rect 12372 8132 12376 8188
rect 12312 8128 12376 8132
rect 16520 8188 16584 8192
rect 16520 8132 16524 8188
rect 16524 8132 16580 8188
rect 16580 8132 16584 8188
rect 16520 8128 16584 8132
rect 16600 8188 16664 8192
rect 16600 8132 16604 8188
rect 16604 8132 16660 8188
rect 16660 8132 16664 8188
rect 16600 8128 16664 8132
rect 16680 8188 16744 8192
rect 16680 8132 16684 8188
rect 16684 8132 16740 8188
rect 16740 8132 16744 8188
rect 16680 8128 16744 8132
rect 16760 8188 16824 8192
rect 16760 8132 16764 8188
rect 16764 8132 16820 8188
rect 16820 8132 16824 8188
rect 16760 8128 16824 8132
rect 3556 8120 3620 8124
rect 3556 8064 3606 8120
rect 3606 8064 3620 8120
rect 3556 8060 3620 8064
rect 3924 8060 3988 8124
rect 5028 7788 5092 7852
rect 14044 7788 14108 7852
rect 4476 7652 4540 7716
rect 4108 7516 4172 7580
rect 5400 7644 5464 7648
rect 5400 7588 5404 7644
rect 5404 7588 5460 7644
rect 5460 7588 5464 7644
rect 5400 7584 5464 7588
rect 5480 7644 5544 7648
rect 5480 7588 5484 7644
rect 5484 7588 5540 7644
rect 5540 7588 5544 7644
rect 5480 7584 5544 7588
rect 5560 7644 5624 7648
rect 5560 7588 5564 7644
rect 5564 7588 5620 7644
rect 5620 7588 5624 7644
rect 5560 7584 5624 7588
rect 5640 7644 5704 7648
rect 5640 7588 5644 7644
rect 5644 7588 5700 7644
rect 5700 7588 5704 7644
rect 5640 7584 5704 7588
rect 9848 7644 9912 7648
rect 9848 7588 9852 7644
rect 9852 7588 9908 7644
rect 9908 7588 9912 7644
rect 9848 7584 9912 7588
rect 9928 7644 9992 7648
rect 9928 7588 9932 7644
rect 9932 7588 9988 7644
rect 9988 7588 9992 7644
rect 9928 7584 9992 7588
rect 10008 7644 10072 7648
rect 10008 7588 10012 7644
rect 10012 7588 10068 7644
rect 10068 7588 10072 7644
rect 10008 7584 10072 7588
rect 10088 7644 10152 7648
rect 10088 7588 10092 7644
rect 10092 7588 10148 7644
rect 10148 7588 10152 7644
rect 10088 7584 10152 7588
rect 14296 7644 14360 7648
rect 14296 7588 14300 7644
rect 14300 7588 14356 7644
rect 14356 7588 14360 7644
rect 14296 7584 14360 7588
rect 14376 7644 14440 7648
rect 14376 7588 14380 7644
rect 14380 7588 14436 7644
rect 14436 7588 14440 7644
rect 14376 7584 14440 7588
rect 14456 7644 14520 7648
rect 14456 7588 14460 7644
rect 14460 7588 14516 7644
rect 14516 7588 14520 7644
rect 14456 7584 14520 7588
rect 14536 7644 14600 7648
rect 14536 7588 14540 7644
rect 14540 7588 14596 7644
rect 14596 7588 14600 7644
rect 14536 7584 14600 7588
rect 4660 7576 4724 7580
rect 4660 7520 4674 7576
rect 4674 7520 4724 7576
rect 4660 7516 4724 7520
rect 15884 7576 15948 7580
rect 15884 7520 15934 7576
rect 15934 7520 15948 7576
rect 15884 7516 15948 7520
rect 3740 7304 3804 7308
rect 3740 7248 3754 7304
rect 3754 7248 3804 7304
rect 3740 7244 3804 7248
rect 3740 7168 3804 7172
rect 3740 7112 3790 7168
rect 3790 7112 3804 7168
rect 3740 7108 3804 7112
rect 4476 7108 4540 7172
rect 6132 7108 6196 7172
rect 9628 7244 9692 7308
rect 16988 7244 17052 7308
rect 15884 7108 15948 7172
rect 3176 7100 3240 7104
rect 3176 7044 3180 7100
rect 3180 7044 3236 7100
rect 3236 7044 3240 7100
rect 3176 7040 3240 7044
rect 3256 7100 3320 7104
rect 3256 7044 3260 7100
rect 3260 7044 3316 7100
rect 3316 7044 3320 7100
rect 3256 7040 3320 7044
rect 3336 7100 3400 7104
rect 3336 7044 3340 7100
rect 3340 7044 3396 7100
rect 3396 7044 3400 7100
rect 3336 7040 3400 7044
rect 3416 7100 3480 7104
rect 3416 7044 3420 7100
rect 3420 7044 3476 7100
rect 3476 7044 3480 7100
rect 3416 7040 3480 7044
rect 7624 7100 7688 7104
rect 7624 7044 7628 7100
rect 7628 7044 7684 7100
rect 7684 7044 7688 7100
rect 7624 7040 7688 7044
rect 7704 7100 7768 7104
rect 7704 7044 7708 7100
rect 7708 7044 7764 7100
rect 7764 7044 7768 7100
rect 7704 7040 7768 7044
rect 7784 7100 7848 7104
rect 7784 7044 7788 7100
rect 7788 7044 7844 7100
rect 7844 7044 7848 7100
rect 7784 7040 7848 7044
rect 7864 7100 7928 7104
rect 7864 7044 7868 7100
rect 7868 7044 7924 7100
rect 7924 7044 7928 7100
rect 7864 7040 7928 7044
rect 12072 7100 12136 7104
rect 12072 7044 12076 7100
rect 12076 7044 12132 7100
rect 12132 7044 12136 7100
rect 12072 7040 12136 7044
rect 12152 7100 12216 7104
rect 12152 7044 12156 7100
rect 12156 7044 12212 7100
rect 12212 7044 12216 7100
rect 12152 7040 12216 7044
rect 12232 7100 12296 7104
rect 12232 7044 12236 7100
rect 12236 7044 12292 7100
rect 12292 7044 12296 7100
rect 12232 7040 12296 7044
rect 12312 7100 12376 7104
rect 12312 7044 12316 7100
rect 12316 7044 12372 7100
rect 12372 7044 12376 7100
rect 12312 7040 12376 7044
rect 16520 7100 16584 7104
rect 16520 7044 16524 7100
rect 16524 7044 16580 7100
rect 16580 7044 16584 7100
rect 16520 7040 16584 7044
rect 16600 7100 16664 7104
rect 16600 7044 16604 7100
rect 16604 7044 16660 7100
rect 16660 7044 16664 7100
rect 16600 7040 16664 7044
rect 16680 7100 16744 7104
rect 16680 7044 16684 7100
rect 16684 7044 16740 7100
rect 16740 7044 16744 7100
rect 16680 7040 16744 7044
rect 16760 7100 16824 7104
rect 16760 7044 16764 7100
rect 16764 7044 16820 7100
rect 16820 7044 16824 7100
rect 16760 7040 16824 7044
rect 3004 6836 3068 6900
rect 4476 6836 4540 6900
rect 4844 6836 4908 6900
rect 11284 6972 11348 7036
rect 13124 6836 13188 6900
rect 14780 6972 14844 7036
rect 15700 6836 15764 6900
rect 17356 6836 17420 6900
rect 3556 6564 3620 6628
rect 3556 6292 3620 6356
rect 7052 6700 7116 6764
rect 5400 6556 5464 6560
rect 5400 6500 5404 6556
rect 5404 6500 5460 6556
rect 5460 6500 5464 6556
rect 5400 6496 5464 6500
rect 5480 6556 5544 6560
rect 5480 6500 5484 6556
rect 5484 6500 5540 6556
rect 5540 6500 5544 6556
rect 5480 6496 5544 6500
rect 5560 6556 5624 6560
rect 5560 6500 5564 6556
rect 5564 6500 5620 6556
rect 5620 6500 5624 6556
rect 5560 6496 5624 6500
rect 5640 6556 5704 6560
rect 5640 6500 5644 6556
rect 5644 6500 5700 6556
rect 5700 6500 5704 6556
rect 5640 6496 5704 6500
rect 7236 6428 7300 6492
rect 9848 6556 9912 6560
rect 9848 6500 9852 6556
rect 9852 6500 9908 6556
rect 9908 6500 9912 6556
rect 9848 6496 9912 6500
rect 9928 6556 9992 6560
rect 9928 6500 9932 6556
rect 9932 6500 9988 6556
rect 9988 6500 9992 6556
rect 9928 6496 9992 6500
rect 10008 6556 10072 6560
rect 10008 6500 10012 6556
rect 10012 6500 10068 6556
rect 10068 6500 10072 6556
rect 10008 6496 10072 6500
rect 10088 6556 10152 6560
rect 10088 6500 10092 6556
rect 10092 6500 10148 6556
rect 10148 6500 10152 6556
rect 10088 6496 10152 6500
rect 14296 6556 14360 6560
rect 14296 6500 14300 6556
rect 14300 6500 14356 6556
rect 14356 6500 14360 6556
rect 14296 6496 14360 6500
rect 14376 6556 14440 6560
rect 14376 6500 14380 6556
rect 14380 6500 14436 6556
rect 14436 6500 14440 6556
rect 14376 6496 14440 6500
rect 14456 6556 14520 6560
rect 14456 6500 14460 6556
rect 14460 6500 14516 6556
rect 14516 6500 14520 6556
rect 14456 6496 14520 6500
rect 14536 6556 14600 6560
rect 14536 6500 14540 6556
rect 14540 6500 14596 6556
rect 14596 6500 14600 6556
rect 14536 6496 14600 6500
rect 3924 6156 3988 6220
rect 6132 6156 6196 6220
rect 4660 6020 4724 6084
rect 3176 6012 3240 6016
rect 3176 5956 3180 6012
rect 3180 5956 3236 6012
rect 3236 5956 3240 6012
rect 3176 5952 3240 5956
rect 3256 6012 3320 6016
rect 3256 5956 3260 6012
rect 3260 5956 3316 6012
rect 3316 5956 3320 6012
rect 3256 5952 3320 5956
rect 3336 6012 3400 6016
rect 3336 5956 3340 6012
rect 3340 5956 3396 6012
rect 3396 5956 3400 6012
rect 3336 5952 3400 5956
rect 3416 6012 3480 6016
rect 3416 5956 3420 6012
rect 3420 5956 3476 6012
rect 3476 5956 3480 6012
rect 3416 5952 3480 5956
rect 7624 6012 7688 6016
rect 7624 5956 7628 6012
rect 7628 5956 7684 6012
rect 7684 5956 7688 6012
rect 7624 5952 7688 5956
rect 7704 6012 7768 6016
rect 7704 5956 7708 6012
rect 7708 5956 7764 6012
rect 7764 5956 7768 6012
rect 7704 5952 7768 5956
rect 7784 6012 7848 6016
rect 7784 5956 7788 6012
rect 7788 5956 7844 6012
rect 7844 5956 7848 6012
rect 7784 5952 7848 5956
rect 7864 6012 7928 6016
rect 7864 5956 7868 6012
rect 7868 5956 7924 6012
rect 7924 5956 7928 6012
rect 7864 5952 7928 5956
rect 12072 6012 12136 6016
rect 12072 5956 12076 6012
rect 12076 5956 12132 6012
rect 12132 5956 12136 6012
rect 12072 5952 12136 5956
rect 12152 6012 12216 6016
rect 12152 5956 12156 6012
rect 12156 5956 12212 6012
rect 12212 5956 12216 6012
rect 12152 5952 12216 5956
rect 12232 6012 12296 6016
rect 12232 5956 12236 6012
rect 12236 5956 12292 6012
rect 12292 5956 12296 6012
rect 12232 5952 12296 5956
rect 12312 6012 12376 6016
rect 12312 5956 12316 6012
rect 12316 5956 12372 6012
rect 12372 5956 12376 6012
rect 12312 5952 12376 5956
rect 2820 5884 2884 5948
rect 14964 5944 15028 5948
rect 14964 5888 15014 5944
rect 15014 5888 15028 5944
rect 14964 5884 15028 5888
rect 16520 6012 16584 6016
rect 16520 5956 16524 6012
rect 16524 5956 16580 6012
rect 16580 5956 16584 6012
rect 16520 5952 16584 5956
rect 16600 6012 16664 6016
rect 16600 5956 16604 6012
rect 16604 5956 16660 6012
rect 16660 5956 16664 6012
rect 16600 5952 16664 5956
rect 16680 6012 16744 6016
rect 16680 5956 16684 6012
rect 16684 5956 16740 6012
rect 16740 5956 16744 6012
rect 16680 5952 16744 5956
rect 16760 6012 16824 6016
rect 16760 5956 16764 6012
rect 16764 5956 16820 6012
rect 16820 5956 16824 6012
rect 16760 5952 16824 5956
rect 14964 5612 15028 5676
rect 5400 5468 5464 5472
rect 5400 5412 5404 5468
rect 5404 5412 5460 5468
rect 5460 5412 5464 5468
rect 5400 5408 5464 5412
rect 5480 5468 5544 5472
rect 5480 5412 5484 5468
rect 5484 5412 5540 5468
rect 5540 5412 5544 5468
rect 5480 5408 5544 5412
rect 5560 5468 5624 5472
rect 5560 5412 5564 5468
rect 5564 5412 5620 5468
rect 5620 5412 5624 5468
rect 5560 5408 5624 5412
rect 5640 5468 5704 5472
rect 5640 5412 5644 5468
rect 5644 5412 5700 5468
rect 5700 5412 5704 5468
rect 5640 5408 5704 5412
rect 9848 5468 9912 5472
rect 9848 5412 9852 5468
rect 9852 5412 9908 5468
rect 9908 5412 9912 5468
rect 9848 5408 9912 5412
rect 9928 5468 9992 5472
rect 9928 5412 9932 5468
rect 9932 5412 9988 5468
rect 9988 5412 9992 5468
rect 9928 5408 9992 5412
rect 10008 5468 10072 5472
rect 10008 5412 10012 5468
rect 10012 5412 10068 5468
rect 10068 5412 10072 5468
rect 10008 5408 10072 5412
rect 10088 5468 10152 5472
rect 10088 5412 10092 5468
rect 10092 5412 10148 5468
rect 10148 5412 10152 5468
rect 10088 5408 10152 5412
rect 5948 5340 6012 5404
rect 7236 5340 7300 5404
rect 14296 5468 14360 5472
rect 14296 5412 14300 5468
rect 14300 5412 14356 5468
rect 14356 5412 14360 5468
rect 14296 5408 14360 5412
rect 14376 5468 14440 5472
rect 14376 5412 14380 5468
rect 14380 5412 14436 5468
rect 14436 5412 14440 5468
rect 14376 5408 14440 5412
rect 14456 5468 14520 5472
rect 14456 5412 14460 5468
rect 14460 5412 14516 5468
rect 14516 5412 14520 5468
rect 14456 5408 14520 5412
rect 14536 5468 14600 5472
rect 14536 5412 14540 5468
rect 14540 5412 14596 5468
rect 14596 5412 14600 5468
rect 14536 5408 14600 5412
rect 10364 5068 10428 5132
rect 4108 4932 4172 4996
rect 3176 4924 3240 4928
rect 3176 4868 3180 4924
rect 3180 4868 3236 4924
rect 3236 4868 3240 4924
rect 3176 4864 3240 4868
rect 3256 4924 3320 4928
rect 3256 4868 3260 4924
rect 3260 4868 3316 4924
rect 3316 4868 3320 4924
rect 3256 4864 3320 4868
rect 3336 4924 3400 4928
rect 3336 4868 3340 4924
rect 3340 4868 3396 4924
rect 3396 4868 3400 4924
rect 3336 4864 3400 4868
rect 3416 4924 3480 4928
rect 3416 4868 3420 4924
rect 3420 4868 3476 4924
rect 3476 4868 3480 4924
rect 3416 4864 3480 4868
rect 7624 4924 7688 4928
rect 7624 4868 7628 4924
rect 7628 4868 7684 4924
rect 7684 4868 7688 4924
rect 7624 4864 7688 4868
rect 7704 4924 7768 4928
rect 7704 4868 7708 4924
rect 7708 4868 7764 4924
rect 7764 4868 7768 4924
rect 7704 4864 7768 4868
rect 7784 4924 7848 4928
rect 7784 4868 7788 4924
rect 7788 4868 7844 4924
rect 7844 4868 7848 4924
rect 7784 4864 7848 4868
rect 7864 4924 7928 4928
rect 7864 4868 7868 4924
rect 7868 4868 7924 4924
rect 7924 4868 7928 4924
rect 7864 4864 7928 4868
rect 12072 4924 12136 4928
rect 12072 4868 12076 4924
rect 12076 4868 12132 4924
rect 12132 4868 12136 4924
rect 12072 4864 12136 4868
rect 12152 4924 12216 4928
rect 12152 4868 12156 4924
rect 12156 4868 12212 4924
rect 12212 4868 12216 4924
rect 12152 4864 12216 4868
rect 12232 4924 12296 4928
rect 12232 4868 12236 4924
rect 12236 4868 12292 4924
rect 12292 4868 12296 4924
rect 12232 4864 12296 4868
rect 12312 4924 12376 4928
rect 12312 4868 12316 4924
rect 12316 4868 12372 4924
rect 12372 4868 12376 4924
rect 12312 4864 12376 4868
rect 16520 4924 16584 4928
rect 16520 4868 16524 4924
rect 16524 4868 16580 4924
rect 16580 4868 16584 4924
rect 16520 4864 16584 4868
rect 16600 4924 16664 4928
rect 16600 4868 16604 4924
rect 16604 4868 16660 4924
rect 16660 4868 16664 4924
rect 16600 4864 16664 4868
rect 16680 4924 16744 4928
rect 16680 4868 16684 4924
rect 16684 4868 16740 4924
rect 16740 4868 16744 4924
rect 16680 4864 16744 4868
rect 16760 4924 16824 4928
rect 16760 4868 16764 4924
rect 16764 4868 16820 4924
rect 16820 4868 16824 4924
rect 16760 4864 16824 4868
rect 2452 4856 2516 4860
rect 2452 4800 2466 4856
rect 2466 4800 2516 4856
rect 2452 4796 2516 4800
rect 6868 4796 6932 4860
rect 2268 4720 2332 4724
rect 2268 4664 2318 4720
rect 2318 4664 2332 4720
rect 2268 4660 2332 4664
rect 2636 4660 2700 4724
rect 10732 4388 10796 4452
rect 5400 4380 5464 4384
rect 5400 4324 5404 4380
rect 5404 4324 5460 4380
rect 5460 4324 5464 4380
rect 5400 4320 5464 4324
rect 5480 4380 5544 4384
rect 5480 4324 5484 4380
rect 5484 4324 5540 4380
rect 5540 4324 5544 4380
rect 5480 4320 5544 4324
rect 5560 4380 5624 4384
rect 5560 4324 5564 4380
rect 5564 4324 5620 4380
rect 5620 4324 5624 4380
rect 5560 4320 5624 4324
rect 5640 4380 5704 4384
rect 5640 4324 5644 4380
rect 5644 4324 5700 4380
rect 5700 4324 5704 4380
rect 5640 4320 5704 4324
rect 9848 4380 9912 4384
rect 9848 4324 9852 4380
rect 9852 4324 9908 4380
rect 9908 4324 9912 4380
rect 9848 4320 9912 4324
rect 9928 4380 9992 4384
rect 9928 4324 9932 4380
rect 9932 4324 9988 4380
rect 9988 4324 9992 4380
rect 9928 4320 9992 4324
rect 10008 4380 10072 4384
rect 10008 4324 10012 4380
rect 10012 4324 10068 4380
rect 10068 4324 10072 4380
rect 10008 4320 10072 4324
rect 10088 4380 10152 4384
rect 10088 4324 10092 4380
rect 10092 4324 10148 4380
rect 10148 4324 10152 4380
rect 10088 4320 10152 4324
rect 14296 4380 14360 4384
rect 14296 4324 14300 4380
rect 14300 4324 14356 4380
rect 14356 4324 14360 4380
rect 14296 4320 14360 4324
rect 14376 4380 14440 4384
rect 14376 4324 14380 4380
rect 14380 4324 14436 4380
rect 14436 4324 14440 4380
rect 14376 4320 14440 4324
rect 14456 4380 14520 4384
rect 14456 4324 14460 4380
rect 14460 4324 14516 4380
rect 14516 4324 14520 4380
rect 14456 4320 14520 4324
rect 14536 4380 14600 4384
rect 14536 4324 14540 4380
rect 14540 4324 14596 4380
rect 14596 4324 14600 4380
rect 14536 4320 14600 4324
rect 11652 4116 11716 4180
rect 3740 4040 3804 4044
rect 3740 3984 3790 4040
rect 3790 3984 3804 4040
rect 3740 3980 3804 3984
rect 15148 4040 15212 4044
rect 15148 3984 15162 4040
rect 15162 3984 15212 4040
rect 15148 3980 15212 3984
rect 2084 3844 2148 3908
rect 9628 3844 9692 3908
rect 13860 3844 13924 3908
rect 14780 3844 14844 3908
rect 3176 3836 3240 3840
rect 3176 3780 3180 3836
rect 3180 3780 3236 3836
rect 3236 3780 3240 3836
rect 3176 3776 3240 3780
rect 3256 3836 3320 3840
rect 3256 3780 3260 3836
rect 3260 3780 3316 3836
rect 3316 3780 3320 3836
rect 3256 3776 3320 3780
rect 3336 3836 3400 3840
rect 3336 3780 3340 3836
rect 3340 3780 3396 3836
rect 3396 3780 3400 3836
rect 3336 3776 3400 3780
rect 3416 3836 3480 3840
rect 3416 3780 3420 3836
rect 3420 3780 3476 3836
rect 3476 3780 3480 3836
rect 3416 3776 3480 3780
rect 7624 3836 7688 3840
rect 7624 3780 7628 3836
rect 7628 3780 7684 3836
rect 7684 3780 7688 3836
rect 7624 3776 7688 3780
rect 7704 3836 7768 3840
rect 7704 3780 7708 3836
rect 7708 3780 7764 3836
rect 7764 3780 7768 3836
rect 7704 3776 7768 3780
rect 7784 3836 7848 3840
rect 7784 3780 7788 3836
rect 7788 3780 7844 3836
rect 7844 3780 7848 3836
rect 7784 3776 7848 3780
rect 7864 3836 7928 3840
rect 7864 3780 7868 3836
rect 7868 3780 7924 3836
rect 7924 3780 7928 3836
rect 7864 3776 7928 3780
rect 12072 3836 12136 3840
rect 12072 3780 12076 3836
rect 12076 3780 12132 3836
rect 12132 3780 12136 3836
rect 12072 3776 12136 3780
rect 12152 3836 12216 3840
rect 12152 3780 12156 3836
rect 12156 3780 12212 3836
rect 12212 3780 12216 3836
rect 12152 3776 12216 3780
rect 12232 3836 12296 3840
rect 12232 3780 12236 3836
rect 12236 3780 12292 3836
rect 12292 3780 12296 3836
rect 12232 3776 12296 3780
rect 12312 3836 12376 3840
rect 12312 3780 12316 3836
rect 12316 3780 12372 3836
rect 12372 3780 12376 3836
rect 12312 3776 12376 3780
rect 16520 3836 16584 3840
rect 16520 3780 16524 3836
rect 16524 3780 16580 3836
rect 16580 3780 16584 3836
rect 16520 3776 16584 3780
rect 16600 3836 16664 3840
rect 16600 3780 16604 3836
rect 16604 3780 16660 3836
rect 16660 3780 16664 3836
rect 16600 3776 16664 3780
rect 16680 3836 16744 3840
rect 16680 3780 16684 3836
rect 16684 3780 16740 3836
rect 16740 3780 16744 3836
rect 16680 3776 16744 3780
rect 16760 3836 16824 3840
rect 16760 3780 16764 3836
rect 16764 3780 16820 3836
rect 16820 3780 16824 3836
rect 16760 3776 16824 3780
rect 7236 3708 7300 3772
rect 9444 3708 9508 3772
rect 14044 3708 14108 3772
rect 16252 3572 16316 3636
rect 17172 3572 17236 3636
rect 8156 3436 8220 3500
rect 8892 3436 8956 3500
rect 13676 3436 13740 3500
rect 14780 3300 14844 3364
rect 5400 3292 5464 3296
rect 5400 3236 5404 3292
rect 5404 3236 5460 3292
rect 5460 3236 5464 3292
rect 5400 3232 5464 3236
rect 5480 3292 5544 3296
rect 5480 3236 5484 3292
rect 5484 3236 5540 3292
rect 5540 3236 5544 3292
rect 5480 3232 5544 3236
rect 5560 3292 5624 3296
rect 5560 3236 5564 3292
rect 5564 3236 5620 3292
rect 5620 3236 5624 3292
rect 5560 3232 5624 3236
rect 5640 3292 5704 3296
rect 5640 3236 5644 3292
rect 5644 3236 5700 3292
rect 5700 3236 5704 3292
rect 5640 3232 5704 3236
rect 9848 3292 9912 3296
rect 9848 3236 9852 3292
rect 9852 3236 9908 3292
rect 9908 3236 9912 3292
rect 9848 3232 9912 3236
rect 9928 3292 9992 3296
rect 9928 3236 9932 3292
rect 9932 3236 9988 3292
rect 9988 3236 9992 3292
rect 9928 3232 9992 3236
rect 10008 3292 10072 3296
rect 10008 3236 10012 3292
rect 10012 3236 10068 3292
rect 10068 3236 10072 3292
rect 10008 3232 10072 3236
rect 10088 3292 10152 3296
rect 10088 3236 10092 3292
rect 10092 3236 10148 3292
rect 10148 3236 10152 3292
rect 10088 3232 10152 3236
rect 14296 3292 14360 3296
rect 14296 3236 14300 3292
rect 14300 3236 14356 3292
rect 14356 3236 14360 3292
rect 14296 3232 14360 3236
rect 14376 3292 14440 3296
rect 14376 3236 14380 3292
rect 14380 3236 14436 3292
rect 14436 3236 14440 3292
rect 14376 3232 14440 3236
rect 14456 3292 14520 3296
rect 14456 3236 14460 3292
rect 14460 3236 14516 3292
rect 14516 3236 14520 3292
rect 14456 3232 14520 3236
rect 14536 3292 14600 3296
rect 14536 3236 14540 3292
rect 14540 3236 14596 3292
rect 14596 3236 14600 3292
rect 14536 3232 14600 3236
rect 1348 3164 1412 3228
rect 8156 3224 8220 3228
rect 8156 3168 8206 3224
rect 8206 3168 8220 3224
rect 8156 3164 8220 3168
rect 15516 3164 15580 3228
rect 15700 3164 15764 3228
rect 1348 2952 1412 2956
rect 1348 2896 1398 2952
rect 1398 2896 1412 2952
rect 1348 2892 1412 2896
rect 3556 2756 3620 2820
rect 7420 2756 7484 2820
rect 8156 2756 8220 2820
rect 14964 2756 15028 2820
rect 3176 2748 3240 2752
rect 3176 2692 3180 2748
rect 3180 2692 3236 2748
rect 3236 2692 3240 2748
rect 3176 2688 3240 2692
rect 3256 2748 3320 2752
rect 3256 2692 3260 2748
rect 3260 2692 3316 2748
rect 3316 2692 3320 2748
rect 3256 2688 3320 2692
rect 3336 2748 3400 2752
rect 3336 2692 3340 2748
rect 3340 2692 3396 2748
rect 3396 2692 3400 2748
rect 3336 2688 3400 2692
rect 3416 2748 3480 2752
rect 3416 2692 3420 2748
rect 3420 2692 3476 2748
rect 3476 2692 3480 2748
rect 3416 2688 3480 2692
rect 7624 2748 7688 2752
rect 7624 2692 7628 2748
rect 7628 2692 7684 2748
rect 7684 2692 7688 2748
rect 7624 2688 7688 2692
rect 7704 2748 7768 2752
rect 7704 2692 7708 2748
rect 7708 2692 7764 2748
rect 7764 2692 7768 2748
rect 7704 2688 7768 2692
rect 7784 2748 7848 2752
rect 7784 2692 7788 2748
rect 7788 2692 7844 2748
rect 7844 2692 7848 2748
rect 7784 2688 7848 2692
rect 7864 2748 7928 2752
rect 7864 2692 7868 2748
rect 7868 2692 7924 2748
rect 7924 2692 7928 2748
rect 7864 2688 7928 2692
rect 12072 2748 12136 2752
rect 12072 2692 12076 2748
rect 12076 2692 12132 2748
rect 12132 2692 12136 2748
rect 12072 2688 12136 2692
rect 12152 2748 12216 2752
rect 12152 2692 12156 2748
rect 12156 2692 12212 2748
rect 12212 2692 12216 2748
rect 12152 2688 12216 2692
rect 12232 2748 12296 2752
rect 12232 2692 12236 2748
rect 12236 2692 12292 2748
rect 12292 2692 12296 2748
rect 12232 2688 12296 2692
rect 12312 2748 12376 2752
rect 12312 2692 12316 2748
rect 12316 2692 12372 2748
rect 12372 2692 12376 2748
rect 12312 2688 12376 2692
rect 16520 2748 16584 2752
rect 16520 2692 16524 2748
rect 16524 2692 16580 2748
rect 16580 2692 16584 2748
rect 16520 2688 16584 2692
rect 16600 2748 16664 2752
rect 16600 2692 16604 2748
rect 16604 2692 16660 2748
rect 16660 2692 16664 2748
rect 16600 2688 16664 2692
rect 16680 2748 16744 2752
rect 16680 2692 16684 2748
rect 16684 2692 16740 2748
rect 16740 2692 16744 2748
rect 16680 2688 16744 2692
rect 16760 2748 16824 2752
rect 16760 2692 16764 2748
rect 16764 2692 16820 2748
rect 16820 2692 16824 2748
rect 16760 2688 16824 2692
rect 1164 2620 1228 2684
rect 4108 2620 4172 2684
rect 7052 2680 7116 2684
rect 7052 2624 7102 2680
rect 7102 2624 7116 2680
rect 7052 2620 7116 2624
rect 980 2484 1044 2548
rect 10548 2484 10612 2548
rect 4292 2212 4356 2276
rect 8524 2272 8588 2276
rect 8524 2216 8538 2272
rect 8538 2216 8588 2272
rect 8524 2212 8588 2216
rect 5400 2204 5464 2208
rect 5400 2148 5404 2204
rect 5404 2148 5460 2204
rect 5460 2148 5464 2204
rect 5400 2144 5464 2148
rect 5480 2204 5544 2208
rect 5480 2148 5484 2204
rect 5484 2148 5540 2204
rect 5540 2148 5544 2204
rect 5480 2144 5544 2148
rect 5560 2204 5624 2208
rect 5560 2148 5564 2204
rect 5564 2148 5620 2204
rect 5620 2148 5624 2204
rect 5560 2144 5624 2148
rect 5640 2204 5704 2208
rect 5640 2148 5644 2204
rect 5644 2148 5700 2204
rect 5700 2148 5704 2204
rect 5640 2144 5704 2148
rect 9848 2204 9912 2208
rect 9848 2148 9852 2204
rect 9852 2148 9908 2204
rect 9908 2148 9912 2204
rect 9848 2144 9912 2148
rect 9928 2204 9992 2208
rect 9928 2148 9932 2204
rect 9932 2148 9988 2204
rect 9988 2148 9992 2204
rect 9928 2144 9992 2148
rect 10008 2204 10072 2208
rect 10008 2148 10012 2204
rect 10012 2148 10068 2204
rect 10068 2148 10072 2204
rect 10008 2144 10072 2148
rect 10088 2204 10152 2208
rect 10088 2148 10092 2204
rect 10092 2148 10148 2204
rect 10148 2148 10152 2204
rect 10088 2144 10152 2148
rect 14296 2204 14360 2208
rect 14296 2148 14300 2204
rect 14300 2148 14356 2204
rect 14356 2148 14360 2204
rect 14296 2144 14360 2148
rect 14376 2204 14440 2208
rect 14376 2148 14380 2204
rect 14380 2148 14436 2204
rect 14436 2148 14440 2204
rect 14376 2144 14440 2148
rect 14456 2204 14520 2208
rect 14456 2148 14460 2204
rect 14460 2148 14516 2204
rect 14516 2148 14520 2204
rect 14456 2144 14520 2148
rect 14536 2204 14600 2208
rect 14536 2148 14540 2204
rect 14540 2148 14596 2204
rect 14596 2148 14600 2204
rect 14536 2144 14600 2148
rect 11836 1804 11900 1868
<< metal4 >>
rect 979 15876 1045 15877
rect 979 15812 980 15876
rect 1044 15812 1045 15876
rect 979 15811 1045 15812
rect 12755 15876 12821 15877
rect 12755 15812 12756 15876
rect 12820 15812 12821 15876
rect 12755 15811 12821 15812
rect 611 10198 677 10199
rect 611 10134 612 10198
rect 676 10134 677 10198
rect 611 10133 677 10134
rect 614 5130 674 10133
rect 614 5070 858 5130
rect 798 2410 858 5070
rect 982 2549 1042 15811
rect 1163 15740 1229 15741
rect 1163 15676 1164 15740
rect 1228 15676 1229 15740
rect 1163 15675 1229 15676
rect 9443 15740 9509 15741
rect 9443 15676 9444 15740
rect 9508 15676 9509 15740
rect 9443 15675 9509 15676
rect 1166 2685 1226 15675
rect 2635 15468 2701 15469
rect 2635 15404 2636 15468
rect 2700 15404 2701 15468
rect 2635 15403 2701 15404
rect 2451 13156 2517 13157
rect 2451 13092 2452 13156
rect 2516 13092 2517 13156
rect 2451 13091 2517 13092
rect 1347 12884 1413 12885
rect 1347 12820 1348 12884
rect 1412 12820 1413 12884
rect 1347 12819 1413 12820
rect 1350 3229 1410 12819
rect 2267 11932 2333 11933
rect 2267 11868 2268 11932
rect 2332 11868 2333 11932
rect 2267 11867 2333 11868
rect 2083 11116 2149 11117
rect 2083 11052 2084 11116
rect 2148 11052 2149 11116
rect 2083 11051 2149 11052
rect 2086 3909 2146 11051
rect 2270 4725 2330 11867
rect 2454 4861 2514 13091
rect 2638 10845 2698 15403
rect 3168 14720 3488 14736
rect 3168 14656 3176 14720
rect 3240 14656 3256 14720
rect 3320 14656 3336 14720
rect 3400 14656 3416 14720
rect 3480 14656 3488 14720
rect 3168 13632 3488 14656
rect 4475 14652 4541 14653
rect 4475 14588 4476 14652
rect 4540 14588 4541 14652
rect 4475 14587 4541 14588
rect 3555 13700 3621 13701
rect 3555 13636 3556 13700
rect 3620 13636 3621 13700
rect 3555 13635 3621 13636
rect 3168 13568 3176 13632
rect 3240 13568 3256 13632
rect 3320 13568 3336 13632
rect 3400 13568 3416 13632
rect 3480 13568 3488 13632
rect 3003 12884 3069 12885
rect 3003 12820 3004 12884
rect 3068 12820 3069 12884
rect 3003 12819 3069 12820
rect 2635 10844 2701 10845
rect 2635 10780 2636 10844
rect 2700 10780 2701 10844
rect 2635 10779 2701 10780
rect 2819 10708 2885 10709
rect 2819 10644 2820 10708
rect 2884 10644 2885 10708
rect 2819 10643 2885 10644
rect 2822 8941 2882 10643
rect 2819 8940 2885 8941
rect 2819 8876 2820 8940
rect 2884 8876 2885 8940
rect 2819 8875 2885 8876
rect 2635 8260 2701 8261
rect 2635 8196 2636 8260
rect 2700 8196 2701 8260
rect 2635 8195 2701 8196
rect 2819 8260 2885 8261
rect 2819 8196 2820 8260
rect 2884 8196 2885 8260
rect 2819 8195 2885 8196
rect 2451 4860 2517 4861
rect 2451 4796 2452 4860
rect 2516 4796 2517 4860
rect 2451 4795 2517 4796
rect 2638 4725 2698 8195
rect 2822 5949 2882 8195
rect 3006 6901 3066 12819
rect 3168 12544 3488 13568
rect 3558 13293 3618 13635
rect 3555 13292 3621 13293
rect 3555 13228 3556 13292
rect 3620 13228 3621 13292
rect 3555 13227 3621 13228
rect 3923 13292 3989 13293
rect 3923 13228 3924 13292
rect 3988 13228 3989 13292
rect 3923 13227 3989 13228
rect 3168 12480 3176 12544
rect 3240 12480 3256 12544
rect 3320 12480 3336 12544
rect 3400 12480 3416 12544
rect 3480 12480 3488 12544
rect 3168 11456 3488 12480
rect 3168 11392 3176 11456
rect 3240 11392 3256 11456
rect 3320 11392 3336 11456
rect 3400 11392 3416 11456
rect 3480 11392 3488 11456
rect 3168 10368 3488 11392
rect 3558 10709 3618 13227
rect 3555 10708 3621 10709
rect 3555 10644 3556 10708
rect 3620 10644 3621 10708
rect 3555 10643 3621 10644
rect 3168 10304 3176 10368
rect 3240 10304 3256 10368
rect 3320 10304 3336 10368
rect 3400 10304 3416 10368
rect 3480 10304 3488 10368
rect 3168 9280 3488 10304
rect 3168 9216 3176 9280
rect 3240 9216 3256 9280
rect 3320 9216 3336 9280
rect 3400 9216 3416 9280
rect 3480 9216 3488 9280
rect 3168 8192 3488 9216
rect 3739 9076 3805 9077
rect 3739 9012 3740 9076
rect 3804 9012 3805 9076
rect 3739 9011 3805 9012
rect 3742 8397 3802 9011
rect 3926 8397 3986 13227
rect 4107 12476 4173 12477
rect 4107 12412 4108 12476
rect 4172 12412 4173 12476
rect 4107 12411 4173 12412
rect 4110 12069 4170 12411
rect 4107 12068 4173 12069
rect 4107 12004 4108 12068
rect 4172 12004 4173 12068
rect 4107 12003 4173 12004
rect 4110 9349 4170 12003
rect 4291 9756 4357 9757
rect 4291 9692 4292 9756
rect 4356 9692 4357 9756
rect 4291 9691 4357 9692
rect 4107 9348 4173 9349
rect 4107 9284 4108 9348
rect 4172 9284 4173 9348
rect 4107 9283 4173 9284
rect 3739 8396 3805 8397
rect 3739 8332 3740 8396
rect 3804 8332 3805 8396
rect 3739 8331 3805 8332
rect 3923 8396 3989 8397
rect 3923 8332 3924 8396
rect 3988 8332 3989 8396
rect 3923 8331 3989 8332
rect 3739 8260 3805 8261
rect 3739 8196 3740 8260
rect 3804 8196 3805 8260
rect 3739 8195 3805 8196
rect 3168 8128 3176 8192
rect 3240 8128 3256 8192
rect 3320 8128 3336 8192
rect 3400 8128 3416 8192
rect 3480 8128 3488 8192
rect 3168 7104 3488 8128
rect 3555 8124 3621 8125
rect 3555 8060 3556 8124
rect 3620 8060 3621 8124
rect 3555 8059 3621 8060
rect 3168 7040 3176 7104
rect 3240 7040 3256 7104
rect 3320 7040 3336 7104
rect 3400 7040 3416 7104
rect 3480 7040 3488 7104
rect 3003 6900 3069 6901
rect 3003 6836 3004 6900
rect 3068 6836 3069 6900
rect 3003 6835 3069 6836
rect 3168 6016 3488 7040
rect 3558 6629 3618 8059
rect 3742 7309 3802 8195
rect 3923 8124 3989 8125
rect 3923 8060 3924 8124
rect 3988 8060 3989 8124
rect 3923 8059 3989 8060
rect 3739 7308 3805 7309
rect 3739 7244 3740 7308
rect 3804 7244 3805 7308
rect 3739 7243 3805 7244
rect 3739 7172 3805 7173
rect 3739 7108 3740 7172
rect 3804 7108 3805 7172
rect 3739 7107 3805 7108
rect 3555 6628 3621 6629
rect 3555 6564 3556 6628
rect 3620 6564 3621 6628
rect 3555 6563 3621 6564
rect 3555 6356 3621 6357
rect 3555 6292 3556 6356
rect 3620 6292 3621 6356
rect 3555 6291 3621 6292
rect 3168 5952 3176 6016
rect 3240 5952 3256 6016
rect 3320 5952 3336 6016
rect 3400 5952 3416 6016
rect 3480 5952 3488 6016
rect 2819 5948 2885 5949
rect 2819 5884 2820 5948
rect 2884 5884 2885 5948
rect 2819 5883 2885 5884
rect 3168 4928 3488 5952
rect 3168 4864 3176 4928
rect 3240 4864 3256 4928
rect 3320 4864 3336 4928
rect 3400 4864 3416 4928
rect 3480 4864 3488 4928
rect 2267 4724 2333 4725
rect 2267 4660 2268 4724
rect 2332 4660 2333 4724
rect 2267 4659 2333 4660
rect 2635 4724 2701 4725
rect 2635 4660 2636 4724
rect 2700 4660 2701 4724
rect 2635 4659 2701 4660
rect 2083 3908 2149 3909
rect 2083 3844 2084 3908
rect 2148 3844 2149 3908
rect 2083 3843 2149 3844
rect 3168 3840 3488 4864
rect 3168 3776 3176 3840
rect 3240 3776 3256 3840
rect 3320 3776 3336 3840
rect 3400 3776 3416 3840
rect 3480 3776 3488 3840
rect 1347 3228 1413 3229
rect 1347 3164 1348 3228
rect 1412 3164 1413 3228
rect 1347 3163 1413 3164
rect 1347 2956 1413 2957
rect 1347 2892 1348 2956
rect 1412 2892 1413 2956
rect 1347 2891 1413 2892
rect 1163 2684 1229 2685
rect 1163 2620 1164 2684
rect 1228 2620 1229 2684
rect 1163 2619 1229 2620
rect 979 2548 1045 2549
rect 979 2484 980 2548
rect 1044 2484 1045 2548
rect 979 2483 1045 2484
rect 1350 2410 1410 2891
rect 798 2350 1410 2410
rect 3168 2752 3488 3776
rect 3558 2821 3618 6291
rect 3742 4045 3802 7107
rect 3926 6221 3986 8059
rect 4107 7580 4173 7581
rect 4107 7516 4108 7580
rect 4172 7516 4173 7580
rect 4107 7515 4173 7516
rect 3923 6220 3989 6221
rect 3923 6156 3924 6220
rect 3988 6156 3989 6220
rect 3923 6155 3989 6156
rect 4110 4997 4170 7515
rect 4107 4996 4173 4997
rect 4107 4932 4108 4996
rect 4172 4932 4173 4996
rect 4107 4931 4173 4932
rect 3739 4044 3805 4045
rect 3739 3980 3740 4044
rect 3804 3980 3805 4044
rect 3739 3979 3805 3980
rect 3555 2820 3621 2821
rect 3555 2756 3556 2820
rect 3620 2756 3621 2820
rect 3555 2755 3621 2756
rect 3168 2688 3176 2752
rect 3240 2688 3256 2752
rect 3320 2688 3336 2752
rect 3400 2688 3416 2752
rect 3480 2688 3488 2752
rect 3168 2128 3488 2688
rect 4110 2685 4170 4931
rect 4107 2684 4173 2685
rect 4107 2620 4108 2684
rect 4172 2620 4173 2684
rect 4107 2619 4173 2620
rect 4294 2277 4354 9691
rect 4478 7717 4538 14587
rect 5392 14176 5712 14736
rect 5392 14112 5400 14176
rect 5464 14112 5480 14176
rect 5544 14112 5560 14176
rect 5624 14112 5640 14176
rect 5704 14112 5712 14176
rect 5027 13700 5093 13701
rect 5027 13636 5028 13700
rect 5092 13636 5093 13700
rect 5027 13635 5093 13636
rect 4843 12884 4909 12885
rect 4843 12820 4844 12884
rect 4908 12820 4909 12884
rect 4843 12819 4909 12820
rect 4475 7716 4541 7717
rect 4475 7652 4476 7716
rect 4540 7652 4541 7716
rect 4475 7651 4541 7652
rect 4659 7580 4725 7581
rect 4659 7516 4660 7580
rect 4724 7516 4725 7580
rect 4659 7515 4725 7516
rect 4475 7172 4541 7173
rect 4475 7108 4476 7172
rect 4540 7108 4541 7172
rect 4475 7107 4541 7108
rect 4478 6901 4538 7107
rect 4475 6900 4541 6901
rect 4475 6836 4476 6900
rect 4540 6836 4541 6900
rect 4475 6835 4541 6836
rect 4662 6085 4722 7515
rect 4846 6901 4906 12819
rect 5030 7853 5090 13635
rect 5392 13088 5712 14112
rect 7616 14720 7936 14736
rect 7616 14656 7624 14720
rect 7688 14656 7704 14720
rect 7768 14656 7784 14720
rect 7848 14656 7864 14720
rect 7928 14656 7936 14720
rect 7616 13632 7936 14656
rect 7616 13568 7624 13632
rect 7688 13568 7704 13632
rect 7768 13568 7784 13632
rect 7848 13568 7864 13632
rect 7928 13568 7936 13632
rect 6683 13292 6749 13293
rect 6683 13228 6684 13292
rect 6748 13228 6749 13292
rect 6683 13227 6749 13228
rect 5392 13024 5400 13088
rect 5464 13024 5480 13088
rect 5544 13024 5560 13088
rect 5624 13024 5640 13088
rect 5704 13024 5712 13088
rect 5211 12884 5277 12885
rect 5211 12820 5212 12884
rect 5276 12820 5277 12884
rect 5211 12819 5277 12820
rect 5214 8669 5274 12819
rect 5392 12000 5712 13024
rect 6315 12612 6381 12613
rect 6315 12548 6316 12612
rect 6380 12548 6381 12612
rect 6315 12547 6381 12548
rect 6499 12612 6565 12613
rect 6499 12548 6500 12612
rect 6564 12548 6565 12612
rect 6499 12547 6565 12548
rect 5392 11936 5400 12000
rect 5464 11936 5480 12000
rect 5544 11936 5560 12000
rect 5624 11936 5640 12000
rect 5704 11936 5712 12000
rect 5392 10912 5712 11936
rect 6131 11660 6197 11661
rect 6131 11596 6132 11660
rect 6196 11596 6197 11660
rect 6131 11595 6197 11596
rect 5947 11252 6013 11253
rect 5947 11188 5948 11252
rect 6012 11188 6013 11252
rect 5947 11187 6013 11188
rect 5392 10848 5400 10912
rect 5464 10848 5480 10912
rect 5544 10848 5560 10912
rect 5624 10848 5640 10912
rect 5704 10848 5712 10912
rect 5392 9824 5712 10848
rect 5392 9760 5400 9824
rect 5464 9760 5480 9824
rect 5544 9760 5560 9824
rect 5624 9760 5640 9824
rect 5704 9760 5712 9824
rect 5392 8736 5712 9760
rect 5392 8672 5400 8736
rect 5464 8672 5480 8736
rect 5544 8672 5560 8736
rect 5624 8672 5640 8736
rect 5704 8672 5712 8736
rect 5211 8668 5277 8669
rect 5211 8604 5212 8668
rect 5276 8604 5277 8668
rect 5211 8603 5277 8604
rect 5027 7852 5093 7853
rect 5027 7788 5028 7852
rect 5092 7788 5093 7852
rect 5027 7787 5093 7788
rect 5392 7648 5712 8672
rect 5392 7584 5400 7648
rect 5464 7584 5480 7648
rect 5544 7584 5560 7648
rect 5624 7584 5640 7648
rect 5704 7584 5712 7648
rect 4843 6900 4909 6901
rect 4843 6836 4844 6900
rect 4908 6836 4909 6900
rect 4843 6835 4909 6836
rect 5392 6560 5712 7584
rect 5392 6496 5400 6560
rect 5464 6496 5480 6560
rect 5544 6496 5560 6560
rect 5624 6496 5640 6560
rect 5704 6496 5712 6560
rect 4659 6084 4725 6085
rect 4659 6020 4660 6084
rect 4724 6020 4725 6084
rect 4659 6019 4725 6020
rect 5392 5472 5712 6496
rect 5392 5408 5400 5472
rect 5464 5408 5480 5472
rect 5544 5408 5560 5472
rect 5624 5408 5640 5472
rect 5704 5408 5712 5472
rect 5392 4384 5712 5408
rect 5950 5405 6010 11187
rect 6134 9621 6194 11595
rect 6131 9620 6197 9621
rect 6131 9556 6132 9620
rect 6196 9556 6197 9620
rect 6131 9555 6197 9556
rect 6131 7172 6197 7173
rect 6131 7108 6132 7172
rect 6196 7170 6197 7172
rect 6318 7170 6378 12547
rect 6502 9757 6562 12547
rect 6686 9893 6746 13227
rect 7616 12544 7936 13568
rect 9446 13429 9506 15675
rect 12571 15468 12637 15469
rect 12571 15404 12572 15468
rect 12636 15404 12637 15468
rect 12571 15403 12637 15404
rect 10915 15060 10981 15061
rect 10915 14996 10916 15060
rect 10980 14996 10981 15060
rect 10915 14995 10981 14996
rect 9840 14176 10160 14736
rect 10731 14652 10797 14653
rect 10731 14588 10732 14652
rect 10796 14588 10797 14652
rect 10731 14587 10797 14588
rect 10363 14380 10429 14381
rect 10363 14316 10364 14380
rect 10428 14316 10429 14380
rect 10363 14315 10429 14316
rect 9840 14112 9848 14176
rect 9912 14112 9928 14176
rect 9992 14112 10008 14176
rect 10072 14112 10088 14176
rect 10152 14112 10160 14176
rect 9443 13428 9509 13429
rect 9443 13364 9444 13428
rect 9508 13364 9509 13428
rect 9443 13363 9509 13364
rect 9840 13088 10160 14112
rect 9840 13024 9848 13088
rect 9912 13024 9928 13088
rect 9992 13024 10008 13088
rect 10072 13024 10088 13088
rect 10152 13024 10160 13088
rect 8891 12748 8957 12749
rect 8891 12684 8892 12748
rect 8956 12684 8957 12748
rect 8891 12683 8957 12684
rect 8155 12612 8221 12613
rect 8155 12548 8156 12612
rect 8220 12548 8221 12612
rect 8155 12547 8221 12548
rect 7616 12480 7624 12544
rect 7688 12480 7704 12544
rect 7768 12480 7784 12544
rect 7848 12480 7864 12544
rect 7928 12480 7936 12544
rect 7051 12476 7117 12477
rect 7051 12412 7052 12476
rect 7116 12412 7117 12476
rect 7051 12411 7117 12412
rect 6867 11796 6933 11797
rect 6867 11732 6868 11796
rect 6932 11732 6933 11796
rect 6867 11731 6933 11732
rect 6683 9892 6749 9893
rect 6683 9828 6684 9892
rect 6748 9828 6749 9892
rect 6683 9827 6749 9828
rect 6499 9756 6565 9757
rect 6499 9692 6500 9756
rect 6564 9692 6565 9756
rect 6499 9691 6565 9692
rect 6870 8941 6930 11731
rect 7054 9213 7114 12411
rect 7235 12340 7301 12341
rect 7235 12276 7236 12340
rect 7300 12276 7301 12340
rect 7235 12275 7301 12276
rect 7238 10573 7298 12275
rect 7419 11932 7485 11933
rect 7419 11868 7420 11932
rect 7484 11868 7485 11932
rect 7419 11867 7485 11868
rect 7235 10572 7301 10573
rect 7235 10508 7236 10572
rect 7300 10508 7301 10572
rect 7235 10507 7301 10508
rect 7422 10301 7482 11867
rect 7616 11456 7936 12480
rect 8158 12069 8218 12547
rect 8155 12068 8221 12069
rect 8155 12004 8156 12068
rect 8220 12004 8221 12068
rect 8155 12003 8221 12004
rect 7616 11392 7624 11456
rect 7688 11392 7704 11456
rect 7768 11392 7784 11456
rect 7848 11392 7864 11456
rect 7928 11392 7936 11456
rect 7616 10368 7936 11392
rect 7616 10304 7624 10368
rect 7688 10304 7704 10368
rect 7768 10304 7784 10368
rect 7848 10304 7864 10368
rect 7928 10304 7936 10368
rect 7419 10300 7485 10301
rect 7419 10236 7420 10300
rect 7484 10236 7485 10300
rect 7419 10235 7485 10236
rect 7419 9892 7485 9893
rect 7419 9828 7420 9892
rect 7484 9828 7485 9892
rect 7419 9827 7485 9828
rect 7051 9212 7117 9213
rect 7051 9148 7052 9212
rect 7116 9210 7117 9212
rect 7116 9150 7298 9210
rect 7116 9148 7117 9150
rect 7051 9147 7117 9148
rect 6867 8940 6933 8941
rect 6867 8876 6868 8940
rect 6932 8876 6933 8940
rect 6867 8875 6933 8876
rect 6196 7110 6378 7170
rect 6196 7108 6197 7110
rect 6131 7107 6197 7108
rect 6134 6221 6194 7107
rect 6131 6220 6197 6221
rect 6131 6156 6132 6220
rect 6196 6156 6197 6220
rect 6131 6155 6197 6156
rect 5947 5404 6013 5405
rect 5947 5340 5948 5404
rect 6012 5340 6013 5404
rect 5947 5339 6013 5340
rect 6870 4861 6930 8875
rect 7051 6764 7117 6765
rect 7051 6700 7052 6764
rect 7116 6700 7117 6764
rect 7051 6699 7117 6700
rect 6867 4860 6933 4861
rect 6867 4796 6868 4860
rect 6932 4796 6933 4860
rect 6867 4795 6933 4796
rect 5392 4320 5400 4384
rect 5464 4320 5480 4384
rect 5544 4320 5560 4384
rect 5624 4320 5640 4384
rect 5704 4320 5712 4384
rect 5392 3296 5712 4320
rect 5392 3232 5400 3296
rect 5464 3232 5480 3296
rect 5544 3232 5560 3296
rect 5624 3232 5640 3296
rect 5704 3232 5712 3296
rect 4291 2276 4357 2277
rect 4291 2212 4292 2276
rect 4356 2212 4357 2276
rect 4291 2211 4357 2212
rect 5392 2208 5712 3232
rect 7054 2685 7114 6699
rect 7238 6493 7298 9150
rect 7422 8941 7482 9827
rect 7616 9280 7936 10304
rect 8158 9757 8218 12003
rect 8523 11116 8589 11117
rect 8523 11052 8524 11116
rect 8588 11052 8589 11116
rect 8523 11051 8589 11052
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 7616 9216 7624 9280
rect 7688 9216 7704 9280
rect 7768 9216 7784 9280
rect 7848 9216 7864 9280
rect 7928 9216 7936 9280
rect 7419 8940 7485 8941
rect 7419 8876 7420 8940
rect 7484 8876 7485 8940
rect 7419 8875 7485 8876
rect 7419 8260 7485 8261
rect 7419 8196 7420 8260
rect 7484 8196 7485 8260
rect 7419 8195 7485 8196
rect 7235 6492 7301 6493
rect 7235 6428 7236 6492
rect 7300 6428 7301 6492
rect 7235 6427 7301 6428
rect 7235 5404 7301 5405
rect 7235 5340 7236 5404
rect 7300 5340 7301 5404
rect 7235 5339 7301 5340
rect 7238 3773 7298 5339
rect 7235 3772 7301 3773
rect 7235 3708 7236 3772
rect 7300 3708 7301 3772
rect 7235 3707 7301 3708
rect 7422 2821 7482 8195
rect 7616 8192 7936 9216
rect 8155 8396 8221 8397
rect 8155 8332 8156 8396
rect 8220 8332 8221 8396
rect 8155 8331 8221 8332
rect 7616 8128 7624 8192
rect 7688 8128 7704 8192
rect 7768 8128 7784 8192
rect 7848 8128 7864 8192
rect 7928 8128 7936 8192
rect 7616 7104 7936 8128
rect 8158 7258 8218 8331
rect 7616 7040 7624 7104
rect 7688 7040 7704 7104
rect 7768 7040 7784 7104
rect 7848 7040 7864 7104
rect 7928 7040 7936 7104
rect 7616 6016 7936 7040
rect 7616 5952 7624 6016
rect 7688 5952 7704 6016
rect 7768 5952 7784 6016
rect 7848 5952 7864 6016
rect 7928 5952 7936 6016
rect 7616 4928 7936 5952
rect 7616 4864 7624 4928
rect 7688 4864 7704 4928
rect 7768 4864 7784 4928
rect 7848 4864 7864 4928
rect 7928 4864 7936 4928
rect 7616 3840 7936 4864
rect 7616 3776 7624 3840
rect 7688 3776 7704 3840
rect 7768 3776 7784 3840
rect 7848 3776 7864 3840
rect 7928 3776 7936 3840
rect 7419 2820 7485 2821
rect 7419 2756 7420 2820
rect 7484 2756 7485 2820
rect 7419 2755 7485 2756
rect 7616 2752 7936 3776
rect 8158 3501 8218 7022
rect 8155 3500 8221 3501
rect 8155 3436 8156 3500
rect 8220 3436 8221 3500
rect 8155 3435 8221 3436
rect 8155 3228 8221 3229
rect 8155 3164 8156 3228
rect 8220 3164 8221 3228
rect 8155 3163 8221 3164
rect 8158 2821 8218 3163
rect 8155 2820 8221 2821
rect 8155 2756 8156 2820
rect 8220 2756 8221 2820
rect 8155 2755 8221 2756
rect 7616 2688 7624 2752
rect 7688 2688 7704 2752
rect 7768 2688 7784 2752
rect 7848 2688 7864 2752
rect 7928 2688 7936 2752
rect 7051 2684 7117 2685
rect 7051 2620 7052 2684
rect 7116 2620 7117 2684
rect 7051 2619 7117 2620
rect 5392 2144 5400 2208
rect 5464 2144 5480 2208
rect 5544 2144 5560 2208
rect 5624 2144 5640 2208
rect 5704 2144 5712 2208
rect 5392 2128 5712 2144
rect 7616 2128 7936 2688
rect 8526 2277 8586 11051
rect 8894 3501 8954 12683
rect 9840 12000 10160 13024
rect 9840 11936 9848 12000
rect 9912 11936 9928 12000
rect 9992 11936 10008 12000
rect 10072 11936 10088 12000
rect 10152 11936 10160 12000
rect 9627 11796 9693 11797
rect 9627 11732 9628 11796
rect 9692 11732 9693 11796
rect 9627 11731 9693 11732
rect 9443 11252 9509 11253
rect 9443 11188 9444 11252
rect 9508 11188 9509 11252
rect 9443 11187 9509 11188
rect 9446 3773 9506 11187
rect 9630 7309 9690 11731
rect 9840 10912 10160 11936
rect 9840 10848 9848 10912
rect 9912 10848 9928 10912
rect 9992 10848 10008 10912
rect 10072 10848 10088 10912
rect 10152 10848 10160 10912
rect 9840 9824 10160 10848
rect 9840 9760 9848 9824
rect 9912 9760 9928 9824
rect 9992 9760 10008 9824
rect 10072 9760 10088 9824
rect 10152 9760 10160 9824
rect 9840 8736 10160 9760
rect 9840 8672 9848 8736
rect 9912 8672 9928 8736
rect 9992 8672 10008 8736
rect 10072 8672 10088 8736
rect 10152 8672 10160 8736
rect 9840 7648 10160 8672
rect 9840 7584 9848 7648
rect 9912 7584 9928 7648
rect 9992 7584 10008 7648
rect 10072 7584 10088 7648
rect 10152 7584 10160 7648
rect 9627 7308 9693 7309
rect 9627 7244 9628 7308
rect 9692 7244 9693 7308
rect 9627 7243 9693 7244
rect 9630 3909 9690 7243
rect 9840 6560 10160 7584
rect 9840 6496 9848 6560
rect 9912 6496 9928 6560
rect 9992 6496 10008 6560
rect 10072 6496 10088 6560
rect 10152 6496 10160 6560
rect 9840 5472 10160 6496
rect 9840 5408 9848 5472
rect 9912 5408 9928 5472
rect 9992 5408 10008 5472
rect 10072 5408 10088 5472
rect 10152 5408 10160 5472
rect 9840 4384 10160 5408
rect 10366 5133 10426 14315
rect 10547 14108 10613 14109
rect 10547 14044 10548 14108
rect 10612 14044 10613 14108
rect 10547 14043 10613 14044
rect 10550 12613 10610 14043
rect 10547 12612 10613 12613
rect 10547 12548 10548 12612
rect 10612 12548 10613 12612
rect 10547 12547 10613 12548
rect 10734 11797 10794 14587
rect 10731 11796 10797 11797
rect 10731 11732 10732 11796
rect 10796 11732 10797 11796
rect 10731 11731 10797 11732
rect 10918 11525 10978 14995
rect 12064 14720 12384 14736
rect 12064 14656 12072 14720
rect 12136 14656 12152 14720
rect 12216 14656 12232 14720
rect 12296 14656 12312 14720
rect 12376 14656 12384 14720
rect 12064 13632 12384 14656
rect 12064 13568 12072 13632
rect 12136 13568 12152 13632
rect 12216 13568 12232 13632
rect 12296 13568 12312 13632
rect 12376 13568 12384 13632
rect 11651 13292 11717 13293
rect 11651 13228 11652 13292
rect 11716 13228 11717 13292
rect 11651 13227 11717 13228
rect 11467 12612 11533 12613
rect 11467 12548 11468 12612
rect 11532 12548 11533 12612
rect 11467 12547 11533 12548
rect 11099 12476 11165 12477
rect 11099 12412 11100 12476
rect 11164 12412 11165 12476
rect 11099 12411 11165 12412
rect 10547 11524 10613 11525
rect 10547 11460 10548 11524
rect 10612 11460 10613 11524
rect 10547 11459 10613 11460
rect 10915 11524 10981 11525
rect 10915 11460 10916 11524
rect 10980 11460 10981 11524
rect 10915 11459 10981 11460
rect 10363 5132 10429 5133
rect 10363 5068 10364 5132
rect 10428 5068 10429 5132
rect 10363 5067 10429 5068
rect 9840 4320 9848 4384
rect 9912 4320 9928 4384
rect 9992 4320 10008 4384
rect 10072 4320 10088 4384
rect 10152 4320 10160 4384
rect 9627 3908 9693 3909
rect 9627 3844 9628 3908
rect 9692 3844 9693 3908
rect 9627 3843 9693 3844
rect 9443 3772 9509 3773
rect 9443 3708 9444 3772
rect 9508 3708 9509 3772
rect 9443 3707 9509 3708
rect 8891 3500 8957 3501
rect 8891 3436 8892 3500
rect 8956 3436 8957 3500
rect 8891 3435 8957 3436
rect 9840 3296 10160 4320
rect 9840 3232 9848 3296
rect 9912 3232 9928 3296
rect 9992 3232 10008 3296
rect 10072 3232 10088 3296
rect 10152 3232 10160 3296
rect 8523 2276 8589 2277
rect 8523 2212 8524 2276
rect 8588 2212 8589 2276
rect 8523 2211 8589 2212
rect 9840 2208 10160 3232
rect 10550 2549 10610 11459
rect 11102 10573 11162 12411
rect 11283 12068 11349 12069
rect 11283 12004 11284 12068
rect 11348 12004 11349 12068
rect 11283 12003 11349 12004
rect 11099 10572 11165 10573
rect 11099 10508 11100 10572
rect 11164 10508 11165 10572
rect 11099 10507 11165 10508
rect 11286 10165 11346 12003
rect 11470 10301 11530 12547
rect 11654 11117 11714 13227
rect 12064 12544 12384 13568
rect 12064 12480 12072 12544
rect 12136 12480 12152 12544
rect 12216 12480 12232 12544
rect 12296 12480 12312 12544
rect 12376 12480 12384 12544
rect 11835 11796 11901 11797
rect 11835 11732 11836 11796
rect 11900 11732 11901 11796
rect 11835 11731 11901 11732
rect 11651 11116 11717 11117
rect 11651 11052 11652 11116
rect 11716 11052 11717 11116
rect 11651 11051 11717 11052
rect 11651 10572 11717 10573
rect 11651 10508 11652 10572
rect 11716 10508 11717 10572
rect 11651 10507 11717 10508
rect 11467 10300 11533 10301
rect 11467 10236 11468 10300
rect 11532 10236 11533 10300
rect 11467 10235 11533 10236
rect 11283 10164 11349 10165
rect 11283 10100 11284 10164
rect 11348 10100 11349 10164
rect 11654 10162 11714 10507
rect 11283 10099 11349 10100
rect 11470 10102 11714 10162
rect 10731 9212 10797 9213
rect 10731 9148 10732 9212
rect 10796 9148 10797 9212
rect 10731 9147 10797 9148
rect 10734 4453 10794 9147
rect 11286 7037 11346 10099
rect 11470 9757 11530 10102
rect 11651 9892 11717 9893
rect 11651 9828 11652 9892
rect 11716 9828 11717 9892
rect 11651 9827 11717 9828
rect 11467 9756 11533 9757
rect 11467 9692 11468 9756
rect 11532 9692 11533 9756
rect 11467 9691 11533 9692
rect 11283 7036 11349 7037
rect 11283 6972 11284 7036
rect 11348 6972 11349 7036
rect 11283 6971 11349 6972
rect 10731 4452 10797 4453
rect 10731 4388 10732 4452
rect 10796 4388 10797 4452
rect 10731 4387 10797 4388
rect 11654 4181 11714 9827
rect 11838 9757 11898 11731
rect 12064 11456 12384 12480
rect 12574 11797 12634 15403
rect 12571 11796 12637 11797
rect 12571 11732 12572 11796
rect 12636 11732 12637 11796
rect 12571 11731 12637 11732
rect 12758 11525 12818 15811
rect 16067 14924 16133 14925
rect 16067 14860 16068 14924
rect 16132 14860 16133 14924
rect 16067 14859 16133 14860
rect 14288 14176 14608 14736
rect 14288 14112 14296 14176
rect 14360 14112 14376 14176
rect 14440 14112 14456 14176
rect 14520 14112 14536 14176
rect 14600 14112 14608 14176
rect 14043 13836 14109 13837
rect 14043 13772 14044 13836
rect 14108 13772 14109 13836
rect 14043 13771 14109 13772
rect 13307 13020 13373 13021
rect 13307 12956 13308 13020
rect 13372 12956 13373 13020
rect 13307 12955 13373 12956
rect 12939 12884 13005 12885
rect 12939 12820 12940 12884
rect 13004 12820 13005 12884
rect 12939 12819 13005 12820
rect 12755 11524 12821 11525
rect 12755 11460 12756 11524
rect 12820 11460 12821 11524
rect 12755 11459 12821 11460
rect 12064 11392 12072 11456
rect 12136 11392 12152 11456
rect 12216 11392 12232 11456
rect 12296 11392 12312 11456
rect 12376 11392 12384 11456
rect 12064 10368 12384 11392
rect 12064 10304 12072 10368
rect 12136 10304 12152 10368
rect 12216 10304 12232 10368
rect 12296 10304 12312 10368
rect 12376 10304 12384 10368
rect 11835 9756 11901 9757
rect 11835 9692 11836 9756
rect 11900 9692 11901 9756
rect 11835 9691 11901 9692
rect 12064 9280 12384 10304
rect 12064 9216 12072 9280
rect 12136 9216 12152 9280
rect 12216 9216 12232 9280
rect 12296 9216 12312 9280
rect 12376 9216 12384 9280
rect 11835 8396 11901 8397
rect 11835 8332 11836 8396
rect 11900 8332 11901 8396
rect 11835 8331 11901 8332
rect 11651 4180 11717 4181
rect 11651 4116 11652 4180
rect 11716 4116 11717 4180
rect 11651 4115 11717 4116
rect 10547 2548 10613 2549
rect 10547 2484 10548 2548
rect 10612 2484 10613 2548
rect 10547 2483 10613 2484
rect 9840 2144 9848 2208
rect 9912 2144 9928 2208
rect 9992 2144 10008 2208
rect 10072 2144 10088 2208
rect 10152 2144 10160 2208
rect 9840 2128 10160 2144
rect 11838 1869 11898 8331
rect 12064 8192 12384 9216
rect 12942 9077 13002 12819
rect 13123 11388 13189 11389
rect 13123 11324 13124 11388
rect 13188 11324 13189 11388
rect 13123 11323 13189 11324
rect 12939 9076 13005 9077
rect 12939 9012 12940 9076
rect 13004 9012 13005 9076
rect 12939 9011 13005 9012
rect 12064 8128 12072 8192
rect 12136 8128 12152 8192
rect 12216 8128 12232 8192
rect 12296 8128 12312 8192
rect 12376 8128 12384 8192
rect 12064 7104 12384 8128
rect 12064 7040 12072 7104
rect 12136 7040 12152 7104
rect 12216 7040 12232 7104
rect 12296 7040 12312 7104
rect 12376 7040 12384 7104
rect 12064 6016 12384 7040
rect 13126 6901 13186 11323
rect 13310 10573 13370 12955
rect 13491 12884 13557 12885
rect 13491 12820 13492 12884
rect 13556 12820 13557 12884
rect 13491 12819 13557 12820
rect 13675 12884 13741 12885
rect 13675 12820 13676 12884
rect 13740 12820 13741 12884
rect 13675 12819 13741 12820
rect 13494 12477 13554 12819
rect 13491 12476 13557 12477
rect 13491 12412 13492 12476
rect 13556 12412 13557 12476
rect 13491 12411 13557 12412
rect 13491 11932 13557 11933
rect 13491 11868 13492 11932
rect 13556 11868 13557 11932
rect 13491 11867 13557 11868
rect 13307 10572 13373 10573
rect 13307 10508 13308 10572
rect 13372 10508 13373 10572
rect 13307 10507 13373 10508
rect 13494 9077 13554 11867
rect 13491 9076 13557 9077
rect 13491 9012 13492 9076
rect 13556 9012 13557 9076
rect 13491 9011 13557 9012
rect 13491 8940 13557 8941
rect 13491 8876 13492 8940
rect 13556 8876 13557 8940
rect 13491 8875 13557 8876
rect 13494 7850 13554 8875
rect 13678 8397 13738 12819
rect 13859 12068 13925 12069
rect 13859 12004 13860 12068
rect 13924 12004 13925 12068
rect 13859 12003 13925 12004
rect 13675 8396 13741 8397
rect 13675 8332 13676 8396
rect 13740 8332 13741 8396
rect 13675 8331 13741 8332
rect 13494 7790 13738 7850
rect 13123 6900 13189 6901
rect 13123 6836 13124 6900
rect 13188 6836 13189 6900
rect 13123 6835 13189 6836
rect 12064 5952 12072 6016
rect 12136 5952 12152 6016
rect 12216 5952 12232 6016
rect 12296 5952 12312 6016
rect 12376 5952 12384 6016
rect 12064 4928 12384 5952
rect 12064 4864 12072 4928
rect 12136 4864 12152 4928
rect 12216 4864 12232 4928
rect 12296 4864 12312 4928
rect 12376 4864 12384 4928
rect 12064 3840 12384 4864
rect 12064 3776 12072 3840
rect 12136 3776 12152 3840
rect 12216 3776 12232 3840
rect 12296 3776 12312 3840
rect 12376 3776 12384 3840
rect 12064 2752 12384 3776
rect 13678 3501 13738 7790
rect 13862 3909 13922 12003
rect 14046 9485 14106 13771
rect 14288 13088 14608 14112
rect 15515 13836 15581 13837
rect 15515 13772 15516 13836
rect 15580 13772 15581 13836
rect 15515 13771 15581 13772
rect 14779 13564 14845 13565
rect 14779 13500 14780 13564
rect 14844 13500 14845 13564
rect 14779 13499 14845 13500
rect 14288 13024 14296 13088
rect 14360 13024 14376 13088
rect 14440 13024 14456 13088
rect 14520 13024 14536 13088
rect 14600 13024 14608 13088
rect 14288 12000 14608 13024
rect 14782 12477 14842 13499
rect 15331 13156 15397 13157
rect 15331 13092 15332 13156
rect 15396 13092 15397 13156
rect 15331 13091 15397 13092
rect 14779 12476 14845 12477
rect 14779 12412 14780 12476
rect 14844 12412 14845 12476
rect 14779 12411 14845 12412
rect 14288 11936 14296 12000
rect 14360 11936 14376 12000
rect 14440 11936 14456 12000
rect 14520 11936 14536 12000
rect 14600 11936 14608 12000
rect 14288 10912 14608 11936
rect 14288 10848 14296 10912
rect 14360 10848 14376 10912
rect 14440 10848 14456 10912
rect 14520 10848 14536 10912
rect 14600 10848 14608 10912
rect 14288 9824 14608 10848
rect 14288 9760 14296 9824
rect 14360 9760 14376 9824
rect 14440 9760 14456 9824
rect 14520 9760 14536 9824
rect 14600 9760 14608 9824
rect 14043 9484 14109 9485
rect 14043 9420 14044 9484
rect 14108 9420 14109 9484
rect 14043 9419 14109 9420
rect 14288 8736 14608 9760
rect 14288 8672 14296 8736
rect 14360 8672 14376 8736
rect 14440 8672 14456 8736
rect 14520 8672 14536 8736
rect 14600 8672 14608 8736
rect 14043 7852 14109 7853
rect 14043 7788 14044 7852
rect 14108 7788 14109 7852
rect 14043 7787 14109 7788
rect 13859 3908 13925 3909
rect 13859 3844 13860 3908
rect 13924 3844 13925 3908
rect 13859 3843 13925 3844
rect 14046 3773 14106 7787
rect 14288 7648 14608 8672
rect 14288 7584 14296 7648
rect 14360 7584 14376 7648
rect 14440 7584 14456 7648
rect 14520 7584 14536 7648
rect 14600 7584 14608 7648
rect 14288 6560 14608 7584
rect 14782 7037 14842 12411
rect 15147 11796 15213 11797
rect 15147 11732 15148 11796
rect 15212 11732 15213 11796
rect 15147 11731 15213 11732
rect 14963 11524 15029 11525
rect 14963 11460 14964 11524
rect 15028 11460 15029 11524
rect 14963 11459 15029 11460
rect 14779 7036 14845 7037
rect 14779 6972 14780 7036
rect 14844 6972 14845 7036
rect 14779 6971 14845 6972
rect 14288 6496 14296 6560
rect 14360 6496 14376 6560
rect 14440 6496 14456 6560
rect 14520 6496 14536 6560
rect 14600 6496 14608 6560
rect 14288 5472 14608 6496
rect 14966 5949 15026 11459
rect 14963 5948 15029 5949
rect 14963 5884 14964 5948
rect 15028 5884 15029 5948
rect 14963 5883 15029 5884
rect 14963 5676 15029 5677
rect 14963 5612 14964 5676
rect 15028 5612 15029 5676
rect 14963 5611 15029 5612
rect 14288 5408 14296 5472
rect 14360 5408 14376 5472
rect 14440 5408 14456 5472
rect 14520 5408 14536 5472
rect 14600 5408 14608 5472
rect 14288 4384 14608 5408
rect 14288 4320 14296 4384
rect 14360 4320 14376 4384
rect 14440 4320 14456 4384
rect 14520 4320 14536 4384
rect 14600 4320 14608 4384
rect 14043 3772 14109 3773
rect 14043 3708 14044 3772
rect 14108 3708 14109 3772
rect 14043 3707 14109 3708
rect 13675 3500 13741 3501
rect 13675 3436 13676 3500
rect 13740 3436 13741 3500
rect 13675 3435 13741 3436
rect 12064 2688 12072 2752
rect 12136 2688 12152 2752
rect 12216 2688 12232 2752
rect 12296 2688 12312 2752
rect 12376 2688 12384 2752
rect 12064 2128 12384 2688
rect 14288 3296 14608 4320
rect 14779 3908 14845 3909
rect 14779 3844 14780 3908
rect 14844 3844 14845 3908
rect 14779 3843 14845 3844
rect 14782 3365 14842 3843
rect 14779 3364 14845 3365
rect 14779 3300 14780 3364
rect 14844 3300 14845 3364
rect 14779 3299 14845 3300
rect 14288 3232 14296 3296
rect 14360 3232 14376 3296
rect 14440 3232 14456 3296
rect 14520 3232 14536 3296
rect 14600 3232 14608 3296
rect 14288 2208 14608 3232
rect 14966 2821 15026 5611
rect 15150 4045 15210 11731
rect 15334 10165 15394 13091
rect 15331 10164 15397 10165
rect 15331 10100 15332 10164
rect 15396 10100 15397 10164
rect 15331 10099 15397 10100
rect 15147 4044 15213 4045
rect 15147 3980 15148 4044
rect 15212 3980 15213 4044
rect 15147 3979 15213 3980
rect 15518 3229 15578 13771
rect 15699 13292 15765 13293
rect 15699 13228 15700 13292
rect 15764 13228 15765 13292
rect 15699 13227 15765 13228
rect 15702 8397 15762 13227
rect 15883 12612 15949 12613
rect 15883 12548 15884 12612
rect 15948 12548 15949 12612
rect 15883 12547 15949 12548
rect 15699 8396 15765 8397
rect 15699 8332 15700 8396
rect 15764 8332 15765 8396
rect 15699 8331 15765 8332
rect 15886 7581 15946 12547
rect 16070 10437 16130 14859
rect 16512 14720 16832 14736
rect 16512 14656 16520 14720
rect 16584 14656 16600 14720
rect 16664 14656 16680 14720
rect 16744 14656 16760 14720
rect 16824 14656 16832 14720
rect 16251 14244 16317 14245
rect 16251 14180 16252 14244
rect 16316 14180 16317 14244
rect 16251 14179 16317 14180
rect 16067 10436 16133 10437
rect 16067 10372 16068 10436
rect 16132 10372 16133 10436
rect 16067 10371 16133 10372
rect 16070 9757 16130 10371
rect 16067 9756 16133 9757
rect 16067 9692 16068 9756
rect 16132 9692 16133 9756
rect 16067 9691 16133 9692
rect 15883 7580 15949 7581
rect 15883 7516 15884 7580
rect 15948 7516 15949 7580
rect 15883 7515 15949 7516
rect 15699 6900 15765 6901
rect 15699 6836 15700 6900
rect 15764 6836 15765 6900
rect 15699 6835 15765 6836
rect 15702 3229 15762 6835
rect 16254 3637 16314 14179
rect 16512 13632 16832 14656
rect 17355 14108 17421 14109
rect 17355 14044 17356 14108
rect 17420 14044 17421 14108
rect 17355 14043 17421 14044
rect 16512 13568 16520 13632
rect 16584 13568 16600 13632
rect 16664 13568 16680 13632
rect 16744 13568 16760 13632
rect 16824 13568 16832 13632
rect 16512 12544 16832 13568
rect 16987 12884 17053 12885
rect 16987 12820 16988 12884
rect 17052 12820 17053 12884
rect 16987 12819 17053 12820
rect 16512 12480 16520 12544
rect 16584 12480 16600 12544
rect 16664 12480 16680 12544
rect 16744 12480 16760 12544
rect 16824 12480 16832 12544
rect 16512 11456 16832 12480
rect 16512 11392 16520 11456
rect 16584 11392 16600 11456
rect 16664 11392 16680 11456
rect 16744 11392 16760 11456
rect 16824 11392 16832 11456
rect 16512 10368 16832 11392
rect 16512 10304 16520 10368
rect 16584 10304 16600 10368
rect 16664 10304 16680 10368
rect 16744 10304 16760 10368
rect 16824 10304 16832 10368
rect 16512 9280 16832 10304
rect 16512 9216 16520 9280
rect 16584 9216 16600 9280
rect 16664 9216 16680 9280
rect 16744 9216 16760 9280
rect 16824 9216 16832 9280
rect 16512 8192 16832 9216
rect 16512 8128 16520 8192
rect 16584 8128 16600 8192
rect 16664 8128 16680 8192
rect 16744 8128 16760 8192
rect 16824 8128 16832 8192
rect 16512 7104 16832 8128
rect 16990 7309 17050 12819
rect 17171 8396 17237 8397
rect 17171 8332 17172 8396
rect 17236 8332 17237 8396
rect 17171 8331 17237 8332
rect 16987 7308 17053 7309
rect 16987 7244 16988 7308
rect 17052 7244 17053 7308
rect 16987 7243 17053 7244
rect 16512 7040 16520 7104
rect 16584 7040 16600 7104
rect 16664 7040 16680 7104
rect 16744 7040 16760 7104
rect 16824 7040 16832 7104
rect 16512 6016 16832 7040
rect 16512 5952 16520 6016
rect 16584 5952 16600 6016
rect 16664 5952 16680 6016
rect 16744 5952 16760 6016
rect 16824 5952 16832 6016
rect 16512 4928 16832 5952
rect 16512 4864 16520 4928
rect 16584 4864 16600 4928
rect 16664 4864 16680 4928
rect 16744 4864 16760 4928
rect 16824 4864 16832 4928
rect 16512 3840 16832 4864
rect 16512 3776 16520 3840
rect 16584 3776 16600 3840
rect 16664 3776 16680 3840
rect 16744 3776 16760 3840
rect 16824 3776 16832 3840
rect 16251 3636 16317 3637
rect 16251 3572 16252 3636
rect 16316 3572 16317 3636
rect 16251 3571 16317 3572
rect 15515 3228 15581 3229
rect 15515 3164 15516 3228
rect 15580 3164 15581 3228
rect 15515 3163 15581 3164
rect 15699 3228 15765 3229
rect 15699 3164 15700 3228
rect 15764 3164 15765 3228
rect 15699 3163 15765 3164
rect 14963 2820 15029 2821
rect 14963 2756 14964 2820
rect 15028 2756 15029 2820
rect 14963 2755 15029 2756
rect 14288 2144 14296 2208
rect 14360 2144 14376 2208
rect 14440 2144 14456 2208
rect 14520 2144 14536 2208
rect 14600 2144 14608 2208
rect 14288 2128 14608 2144
rect 16512 2752 16832 3776
rect 17174 3637 17234 8331
rect 17358 6901 17418 14043
rect 17355 6900 17421 6901
rect 17355 6836 17356 6900
rect 17420 6836 17421 6900
rect 17355 6835 17421 6836
rect 17171 3636 17237 3637
rect 17171 3572 17172 3636
rect 17236 3572 17237 3636
rect 17171 3571 17237 3572
rect 16512 2688 16520 2752
rect 16584 2688 16600 2752
rect 16664 2688 16680 2752
rect 16744 2688 16760 2752
rect 16824 2688 16832 2752
rect 16512 2128 16832 2688
rect 11835 1868 11901 1869
rect 11835 1804 11836 1868
rect 11900 1804 11901 1868
rect 11835 1803 11901 1804
<< via4 >>
rect 8070 7022 8306 7258
rect 15798 7172 16034 7258
rect 15798 7108 15884 7172
rect 15884 7108 15948 7172
rect 15948 7108 16034 7172
rect 15798 7022 16034 7108
<< metal5 >>
rect 8028 7258 16076 7300
rect 8028 7022 8070 7258
rect 8306 7022 15798 7258
rect 16034 7022 16076 7258
rect 8028 6980 16076 7022
use sky130_fd_sc_hd__diode_2  ANTENNA__36__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__37__A
timestamp 1649977179
transform 1 0 11776 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__40__A
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 17204 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__45__A
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform -1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__50__A
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__54__A
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__55__A
timestamp 1649977179
transform -1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__56__A
timestamp 1649977179
transform 1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform -1 0 13156 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform -1 0 14260 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform 1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform -1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 13984 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 14628 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_0_N_in_A
timestamp 1649977179
transform -1 0 12604 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 6992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 5704 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 8556 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 7820 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 6808 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 5336 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 5796 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 7360 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6440 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 5612 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 9476 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 7544 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 11408 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 12052 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 12604 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 12696 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 12512 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 12880 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 13248 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 11776 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 11960 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 17664 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 12236 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 12420 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 7084 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 6900 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 6256 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 7268 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 6072 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9752 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 9108 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9108 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 7912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 8188 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 3772 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A0
timestamp 1649977179
transform -1 0 8832 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 8280 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 5980 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 5520 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6992 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6992 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6992 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 6164 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5244 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6072 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 12604 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 9844 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5244 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12696 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 4600 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9476 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 6992 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 16560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10672 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 18584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11040 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_11.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 18584 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 16560 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 17664 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16560 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 14444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 18584 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10304 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11408 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9936 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 10764 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_ipin_15.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1649977179
transform 1 0 9476 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1649977179
transform -1 0 10120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater137_A
timestamp 1649977179
transform -1 0 5520 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_79
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_154
timestamp 1649977179
transform 1 0 15272 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_54
timestamp 1649977179
transform 1 0 6072 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_19
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_128
timestamp 1649977179
transform 1 0 12880 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_58
timestamp 1649977179
transform 1 0 6440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_130
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_157
timestamp 1649977179
transform 1 0 15548 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_30
timestamp 1649977179
transform 1 0 3864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_74
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_95
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_17
timestamp 1649977179
transform 1 0 2668 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_151
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_23
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_45
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_104
timestamp 1649977179
transform 1 0 10672 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_82
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_107
timestamp 1649977179
transform 1 0 10948 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_68
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_93 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_48
timestamp 1649977179
transform 1 0 5520 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_87 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_99 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_26
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_78
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_95
timestamp 1649977179
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_107
timestamp 1649977179
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_69
timestamp 1649977179
transform 1 0 7452 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1649977179
transform 1 0 9660 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_100
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_113
timestamp 1649977179
transform 1 0 11500 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_117
timestamp 1649977179
transform 1 0 11868 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 18860 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 16560 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _32_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform -1 0 13800 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 4784 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 13064 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform -1 0 7820 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 12420 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform -1 0 6440 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform -1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform -1 0 7452 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform -1 0 4232 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform -1 0 4416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform 1 0 4140 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 2024 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 5612 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 13984 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform 1 0 12328 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 5888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform -1 0 13248 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 8096 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform 1 0 13248 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 15640 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform 1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 18216 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 9476 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 14812 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform -1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_N_FTB01
timestamp 1649977179
transform -1 0 9844 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_S_FTB01
timestamp 1649977179
transform -1 0 14076 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_E_FTB01
timestamp 1649977179
transform -1 0 14812 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_W_FTB01
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_E_FTB01
timestamp 1649977179
transform 1 0 12420 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_W_FTB01
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_top_ipin_0.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11132 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_0_N_in
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_0_N_in
timestamp 1649977179
transform -1 0 14812 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_0_N_in
timestamp 1649977179
transform -1 0 17480 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 9660 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_top_ipin_0.prog_clk
timestamp 1649977179
transform 1 0 12972 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform -1 0 6900 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 6440 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform -1 0 6072 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform -1 0 3680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform -1 0 16376 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 5428 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform -1 0 17388 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 7452 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 8740 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 6532 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 3496 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 5152 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 8188 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform 1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform 1 0 3128 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform -1 0 2300 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1649977179
transform -1 0 2300 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform -1 0 2300 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 3220 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input15
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 3220 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 2300 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input23
timestamp 1649977179
transform 1 0 2300 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 18308 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform -1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 16744 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform -1 0 16192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform -1 0 18584 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform -1 0 17664 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 16560 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 15824 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 17664 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 13432 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 17388 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input39
timestamp 1649977179
transform 1 0 17664 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 15456 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1649977179
transform -1 0 15824 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 17664 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input44
timestamp 1649977179
transform -1 0 16560 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform -1 0 4324 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform -1 0 4600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform -1 0 4140 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2852 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3956 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 1472 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2852 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4048 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4600 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4600 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7820 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8372 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8004 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6256 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 6256 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5520 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 2852 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 3220 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 1472 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4232 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4600 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9476 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 7912 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8096 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10948 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 10396 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11316 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8188 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13064 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13340 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17020 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16284 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16468 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15916 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14444 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15640 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 16468 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13156 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 2484 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_0.mux_l2_in_3__145 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4600 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_1.mux_l2_in_3__146
timestamp 1649977179
transform -1 0 5336 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5336 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4600 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2668 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13156 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7544 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6716 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_2.mux_l2_in_3__153
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4416 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 4048 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_3.mux_l2_in_3__154
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3128 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 4784 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2024 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4416 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_4.mux_l2_in_3__155
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6992 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_5.mux_l2_in_3__140
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6808 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6164 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7176 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5244 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_6.mux_l2_in_3__141
timestamp 1649977179
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4784 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9476 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_7.mux_l2_in_3__142
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11592 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9476 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_8.mux_l2_in_3__143
timestamp 1649977179
transform -1 0 8464 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 8832 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 8188 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 7360 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_9.mux_l2_in_3__144
timestamp 1649977179
transform 1 0 16100 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9936 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_10.mux_l2_in_3__147
timestamp 1649977179
transform -1 0 12512 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12052 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6164 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15640 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15640 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 13156 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13984 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_11.mux_l2_in_3__148
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13156 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13432 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_12.mux_l2_in_3__149
timestamp 1649977179
transform 1 0 16284 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12788 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_13.mux_l2_in_3__150
timestamp 1649977179
transform -1 0 16928 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 16928 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16468 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16744 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 17572 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_14.mux_l2_in_3__151
timestamp 1649977179
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform -1 0 18308 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16744 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform 1 0 17480 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17572 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18032 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17388 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17112 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform 1 0 16560 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_ipin_15.mux_l2_in_3__152
timestamp 1649977179
transform -1 0 15364 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16376 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output51 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2668 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform 1 0 15916 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 3404 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 13432 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 11868 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform -1 0 12604 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 4140 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 3036 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 9476 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 4232 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 4508 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 6532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 5152 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 4324 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 8740 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 15732 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 6716 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 8188 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 13800 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform 1 0 18216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform 1 0 18216 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform 1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 18308 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 18216 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 18216 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 10396 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 13616 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 12972 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 12328 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 17112 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform -1 0 3036 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform -1 0 11592 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform -1 0 3404 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output117
timestamp 1649977179
transform -1 0 14536 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 16744 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 3036 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 14168 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 2668 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_W_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16560 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_N_FTB01
timestamp 1649977179
transform -1 0 15640 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_S_FTB01
timestamp 1649977179
transform -1 0 15088 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  prog_clk_2_E_FTB01
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_2_W_FTB01
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_E_FTB01
timestamp 1649977179
transform 1 0 14076 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_W_FTB01
timestamp 1649977179
transform 1 0 4416 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater124
timestamp 1649977179
transform -1 0 3864 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater125
timestamp 1649977179
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater126
timestamp 1649977179
transform -1 0 11408 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater127
timestamp 1649977179
transform -1 0 14904 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater128
timestamp 1649977179
transform 1 0 7912 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater129
timestamp 1649977179
transform -1 0 13800 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater130
timestamp 1649977179
transform -1 0 16652 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater131
timestamp 1649977179
transform 1 0 17388 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater132
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater133
timestamp 1649977179
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater134
timestamp 1649977179
transform 1 0 5520 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater135
timestamp 1649977179
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater136
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater137
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater138
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater139
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 406 592
<< labels >>
rlabel metal3 s 0 13608 800 13728 6 REGIN_FEEDTHROUGH
port 0 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 REGOUT_FEEDTHROUGH
port 1 nsew signal tristate
rlabel metal2 s 16670 0 16726 800 6 SC_IN_BOT
port 2 nsew signal input
rlabel metal2 s 1950 16400 2006 17200 6 SC_IN_TOP
port 3 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 SC_OUT_BOT
port 4 nsew signal tristate
rlabel metal2 s 5906 16400 5962 17200 6 SC_OUT_TOP
port 5 nsew signal tristate
rlabel metal4 s 5392 2128 5712 14736 6 VGND
port 6 nsew ground input
rlabel metal4 s 9840 2128 10160 14736 6 VGND
port 6 nsew ground input
rlabel metal4 s 14288 2128 14608 14736 6 VGND
port 6 nsew ground input
rlabel metal4 s 3168 2128 3488 14736 6 VPWR
port 7 nsew power input
rlabel metal4 s 7616 2128 7936 14736 6 VPWR
port 7 nsew power input
rlabel metal4 s 12064 2128 12384 14736 6 VPWR
port 7 nsew power input
rlabel metal4 s 16512 2128 16832 14736 6 VPWR
port 7 nsew power input
rlabel metal2 s 2134 0 2190 800 6 bottom_grid_pin_0_
port 8 nsew signal tristate
rlabel metal2 s 11242 0 11298 800 6 bottom_grid_pin_10_
port 9 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 bottom_grid_pin_11_
port 10 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 bottom_grid_pin_12_
port 11 nsew signal tristate
rlabel metal2 s 13910 0 13966 800 6 bottom_grid_pin_13_
port 12 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 bottom_grid_pin_14_
port 13 nsew signal tristate
rlabel metal2 s 15750 0 15806 800 6 bottom_grid_pin_15_
port 14 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 bottom_grid_pin_1_
port 15 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 bottom_grid_pin_2_
port 16 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 bottom_grid_pin_3_
port 17 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 bottom_grid_pin_4_
port 18 nsew signal tristate
rlabel metal2 s 6734 0 6790 800 6 bottom_grid_pin_5_
port 19 nsew signal tristate
rlabel metal2 s 7562 0 7618 800 6 bottom_grid_pin_6_
port 20 nsew signal tristate
rlabel metal2 s 8482 0 8538 800 6 bottom_grid_pin_7_
port 21 nsew signal tristate
rlabel metal2 s 9402 0 9458 800 6 bottom_grid_pin_8_
port 22 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 bottom_grid_pin_9_
port 23 nsew signal tristate
rlabel metal2 s 386 0 442 800 6 ccff_head
port 24 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 ccff_tail
port 25 nsew signal tristate
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[0]
port 26 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[10]
port 27 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[11]
port 28 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 chanx_left_in[12]
port 29 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[13]
port 30 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[14]
port 31 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[15]
port 32 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_in[16]
port 33 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 34 nsew signal input
rlabel metal3 s 0 12656 800 12776 6 chanx_left_in[18]
port 35 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 chanx_left_in[19]
port 36 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[1]
port 37 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[2]
port 38 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[3]
port 39 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[4]
port 40 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 chanx_left_in[5]
port 41 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 chanx_left_in[6]
port 42 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[7]
port 43 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 chanx_left_in[8]
port 44 nsew signal input
rlabel metal3 s 0 9664 800 9784 6 chanx_left_in[9]
port 45 nsew signal input
rlabel metal3 s 0 144 800 264 6 chanx_left_out[0]
port 46 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 chanx_left_out[10]
port 47 nsew signal tristate
rlabel metal3 s 0 3680 800 3800 6 chanx_left_out[11]
port 48 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 chanx_left_out[12]
port 49 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_out[13]
port 50 nsew signal tristate
rlabel metal3 s 0 4632 800 4752 6 chanx_left_out[14]
port 51 nsew signal tristate
rlabel metal3 s 0 5040 800 5160 6 chanx_left_out[15]
port 52 nsew signal tristate
rlabel metal3 s 0 5312 800 5432 6 chanx_left_out[16]
port 53 nsew signal tristate
rlabel metal3 s 0 5720 800 5840 6 chanx_left_out[17]
port 54 nsew signal tristate
rlabel metal3 s 0 5992 800 6112 6 chanx_left_out[18]
port 55 nsew signal tristate
rlabel metal3 s 0 6400 800 6520 6 chanx_left_out[19]
port 56 nsew signal tristate
rlabel metal3 s 0 416 800 536 6 chanx_left_out[1]
port 57 nsew signal tristate
rlabel metal3 s 0 688 800 808 6 chanx_left_out[2]
port 58 nsew signal tristate
rlabel metal3 s 0 1096 800 1216 6 chanx_left_out[3]
port 59 nsew signal tristate
rlabel metal3 s 0 1368 800 1488 6 chanx_left_out[4]
port 60 nsew signal tristate
rlabel metal3 s 0 1776 800 1896 6 chanx_left_out[5]
port 61 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 chanx_left_out[6]
port 62 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 chanx_left_out[7]
port 63 nsew signal tristate
rlabel metal3 s 0 2728 800 2848 6 chanx_left_out[8]
port 64 nsew signal tristate
rlabel metal3 s 0 3000 800 3120 6 chanx_left_out[9]
port 65 nsew signal tristate
rlabel metal3 s 19200 9664 20000 9784 6 chanx_right_in[0]
port 66 nsew signal input
rlabel metal3 s 19200 13472 20000 13592 6 chanx_right_in[10]
port 67 nsew signal input
rlabel metal3 s 19200 13744 20000 13864 6 chanx_right_in[11]
port 68 nsew signal input
rlabel metal3 s 19200 14152 20000 14272 6 chanx_right_in[12]
port 69 nsew signal input
rlabel metal3 s 19200 14560 20000 14680 6 chanx_right_in[13]
port 70 nsew signal input
rlabel metal3 s 19200 14968 20000 15088 6 chanx_right_in[14]
port 71 nsew signal input
rlabel metal3 s 19200 15376 20000 15496 6 chanx_right_in[15]
port 72 nsew signal input
rlabel metal3 s 19200 15648 20000 15768 6 chanx_right_in[16]
port 73 nsew signal input
rlabel metal3 s 19200 16056 20000 16176 6 chanx_right_in[17]
port 74 nsew signal input
rlabel metal3 s 19200 16464 20000 16584 6 chanx_right_in[18]
port 75 nsew signal input
rlabel metal3 s 19200 16872 20000 16992 6 chanx_right_in[19]
port 76 nsew signal input
rlabel metal3 s 19200 9936 20000 10056 6 chanx_right_in[1]
port 77 nsew signal input
rlabel metal3 s 19200 10344 20000 10464 6 chanx_right_in[2]
port 78 nsew signal input
rlabel metal3 s 19200 10752 20000 10872 6 chanx_right_in[3]
port 79 nsew signal input
rlabel metal3 s 19200 11160 20000 11280 6 chanx_right_in[4]
port 80 nsew signal input
rlabel metal3 s 19200 11568 20000 11688 6 chanx_right_in[5]
port 81 nsew signal input
rlabel metal3 s 19200 11840 20000 11960 6 chanx_right_in[6]
port 82 nsew signal input
rlabel metal3 s 19200 12248 20000 12368 6 chanx_right_in[7]
port 83 nsew signal input
rlabel metal3 s 19200 12656 20000 12776 6 chanx_right_in[8]
port 84 nsew signal input
rlabel metal3 s 19200 13064 20000 13184 6 chanx_right_in[9]
port 85 nsew signal input
rlabel metal3 s 19200 2048 20000 2168 6 chanx_right_out[0]
port 86 nsew signal tristate
rlabel metal3 s 19200 5856 20000 5976 6 chanx_right_out[10]
port 87 nsew signal tristate
rlabel metal3 s 19200 6128 20000 6248 6 chanx_right_out[11]
port 88 nsew signal tristate
rlabel metal3 s 19200 6536 20000 6656 6 chanx_right_out[12]
port 89 nsew signal tristate
rlabel metal3 s 19200 6944 20000 7064 6 chanx_right_out[13]
port 90 nsew signal tristate
rlabel metal3 s 19200 7352 20000 7472 6 chanx_right_out[14]
port 91 nsew signal tristate
rlabel metal3 s 19200 7760 20000 7880 6 chanx_right_out[15]
port 92 nsew signal tristate
rlabel metal3 s 19200 8032 20000 8152 6 chanx_right_out[16]
port 93 nsew signal tristate
rlabel metal3 s 19200 8440 20000 8560 6 chanx_right_out[17]
port 94 nsew signal tristate
rlabel metal3 s 19200 8848 20000 8968 6 chanx_right_out[18]
port 95 nsew signal tristate
rlabel metal3 s 19200 9256 20000 9376 6 chanx_right_out[19]
port 96 nsew signal tristate
rlabel metal3 s 19200 2320 20000 2440 6 chanx_right_out[1]
port 97 nsew signal tristate
rlabel metal3 s 19200 2728 20000 2848 6 chanx_right_out[2]
port 98 nsew signal tristate
rlabel metal3 s 19200 3136 20000 3256 6 chanx_right_out[3]
port 99 nsew signal tristate
rlabel metal3 s 19200 3544 20000 3664 6 chanx_right_out[4]
port 100 nsew signal tristate
rlabel metal3 s 19200 3952 20000 4072 6 chanx_right_out[5]
port 101 nsew signal tristate
rlabel metal3 s 19200 4224 20000 4344 6 chanx_right_out[6]
port 102 nsew signal tristate
rlabel metal3 s 19200 4632 20000 4752 6 chanx_right_out[7]
port 103 nsew signal tristate
rlabel metal3 s 19200 5040 20000 5160 6 chanx_right_out[8]
port 104 nsew signal tristate
rlabel metal3 s 19200 5448 20000 5568 6 chanx_right_out[9]
port 105 nsew signal tristate
rlabel metal2 s 9862 16400 9918 17200 6 clk_1_N_out
port 106 nsew signal tristate
rlabel metal2 s 18510 0 18566 800 6 clk_1_S_out
port 107 nsew signal tristate
rlabel metal3 s 0 16872 800 16992 6 clk_1_W_in
port 108 nsew signal input
rlabel metal3 s 19200 1640 20000 1760 6 clk_2_E_out
port 109 nsew signal tristate
rlabel metal3 s 0 16600 800 16720 6 clk_2_W_in
port 110 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 clk_2_W_out
port 111 nsew signal tristate
rlabel metal3 s 19200 1232 20000 1352 6 clk_3_E_out
port 112 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 clk_3_W_in
port 113 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 clk_3_W_out
port 114 nsew signal tristate
rlabel metal2 s 13910 16400 13966 17200 6 prog_clk_0_N_in
port 115 nsew signal input
rlabel metal2 s 17866 16400 17922 17200 6 prog_clk_0_W_out
port 116 nsew signal tristate
rlabel metal3 s 19200 824 20000 944 6 prog_clk_1_N_out
port 117 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 prog_clk_1_S_out
port 118 nsew signal tristate
rlabel metal3 s 0 15920 800 16040 6 prog_clk_1_W_in
port 119 nsew signal input
rlabel metal3 s 19200 416 20000 536 6 prog_clk_2_E_out
port 120 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 prog_clk_2_W_in
port 121 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 prog_clk_2_W_out
port 122 nsew signal tristate
rlabel metal3 s 19200 144 20000 264 6 prog_clk_3_E_out
port 123 nsew signal tristate
rlabel metal3 s 0 15240 800 15360 6 prog_clk_3_W_in
port 124 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 prog_clk_3_W_out
port 125 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 20000 17200
<< end >>
