magic
tech sky130A
magscale 1 2
timestamp 1650540980
<< viali >>
rect 5733 20553 5767 20587
rect 6653 20553 6687 20587
rect 8309 20553 8343 20587
rect 10333 20553 10367 20587
rect 11713 20553 11747 20587
rect 11989 20553 12023 20587
rect 12357 20553 12391 20587
rect 12725 20553 12759 20587
rect 13093 20553 13127 20587
rect 13461 20553 13495 20587
rect 13829 20553 13863 20587
rect 14289 20553 14323 20587
rect 14657 20553 14691 20587
rect 15025 20553 15059 20587
rect 15393 20553 15427 20587
rect 15761 20553 15795 20587
rect 16129 20553 16163 20587
rect 16497 20553 16531 20587
rect 19441 20553 19475 20587
rect 19717 20553 19751 20587
rect 20177 20553 20211 20587
rect 20545 20553 20579 20587
rect 21097 20553 21131 20587
rect 2513 20485 2547 20519
rect 4169 20485 4203 20519
rect 10057 20485 10091 20519
rect 19073 20485 19107 20519
rect 2237 20417 2271 20451
rect 3341 20417 3375 20451
rect 3617 20417 3651 20451
rect 3801 20417 3835 20451
rect 5825 20417 5859 20451
rect 6377 20417 6411 20451
rect 7021 20417 7055 20451
rect 7665 20417 7699 20451
rect 7941 20417 7975 20451
rect 8217 20417 8251 20451
rect 8677 20417 8711 20451
rect 10149 20417 10183 20451
rect 10517 20417 10551 20451
rect 11529 20417 11563 20451
rect 11805 20417 11839 20451
rect 12173 20417 12207 20451
rect 12541 20417 12575 20451
rect 12909 20417 12943 20451
rect 13277 20417 13311 20451
rect 13645 20417 13679 20451
rect 14105 20417 14139 20451
rect 14473 20417 14507 20451
rect 14841 20417 14875 20451
rect 15209 20417 15243 20451
rect 15577 20417 15611 20451
rect 15945 20417 15979 20451
rect 16313 20417 16347 20451
rect 16681 20417 16715 20451
rect 17049 20417 17083 20451
rect 19257 20417 19291 20451
rect 19876 20417 19910 20451
rect 19981 20417 20015 20451
rect 20361 20417 20395 20451
rect 20729 20417 20763 20451
rect 21281 20417 21315 20451
rect 1961 20349 1995 20383
rect 2697 20349 2731 20383
rect 4997 20349 5031 20383
rect 5273 20349 5307 20383
rect 5549 20349 5583 20383
rect 7113 20349 7147 20383
rect 7205 20349 7239 20383
rect 9597 20349 9631 20383
rect 9873 20349 9907 20383
rect 10793 20349 10827 20383
rect 6193 20281 6227 20315
rect 7757 20281 7791 20315
rect 16865 20281 16899 20315
rect 20913 20281 20947 20315
rect 3985 20213 4019 20247
rect 4261 20213 4295 20247
rect 6561 20213 6595 20247
rect 7481 20213 7515 20247
rect 8585 20213 8619 20247
rect 17233 20213 17267 20247
rect 17785 20213 17819 20247
rect 21465 20213 21499 20247
rect 1869 20009 1903 20043
rect 9045 20009 9079 20043
rect 10885 20009 10919 20043
rect 11161 20009 11195 20043
rect 12449 20009 12483 20043
rect 12817 20009 12851 20043
rect 13185 20009 13219 20043
rect 13461 20009 13495 20043
rect 13737 20009 13771 20043
rect 14657 20009 14691 20043
rect 15025 20009 15059 20043
rect 15393 20009 15427 20043
rect 16129 20009 16163 20043
rect 17601 20009 17635 20043
rect 18245 20009 18279 20043
rect 18889 20009 18923 20043
rect 20545 20009 20579 20043
rect 2697 19941 2731 19975
rect 8769 19941 8803 19975
rect 9505 19941 9539 19975
rect 12265 19941 12299 19975
rect 17233 19941 17267 19975
rect 17969 19941 18003 19975
rect 18521 19941 18555 19975
rect 3341 19873 3375 19907
rect 6837 19873 6871 19907
rect 7481 19873 7515 19907
rect 8309 19873 8343 19907
rect 11437 19873 11471 19907
rect 20913 19873 20947 19907
rect 1685 19805 1719 19839
rect 2053 19805 2087 19839
rect 2329 19805 2363 19839
rect 3617 19805 3651 19839
rect 5017 19805 5051 19839
rect 5273 19805 5307 19839
rect 6581 19805 6615 19839
rect 8217 19805 8251 19839
rect 8585 19805 8619 19839
rect 10701 19805 10735 19839
rect 10977 19805 11011 19839
rect 11529 19805 11563 19839
rect 12081 19805 12115 19839
rect 12633 19805 12667 19839
rect 13001 19805 13035 19839
rect 13277 19805 13311 19839
rect 13553 19805 13587 19839
rect 14381 19805 14415 19839
rect 14473 19805 14507 19839
rect 14841 19805 14875 19839
rect 15209 19805 15243 19839
rect 15761 19805 15795 19839
rect 16313 19805 16347 19839
rect 16497 19805 16531 19839
rect 16773 19805 16807 19839
rect 17049 19805 17083 19839
rect 17417 19805 17451 19839
rect 17785 19805 17819 19839
rect 18429 19805 18463 19839
rect 18705 19805 18739 19839
rect 19073 19805 19107 19839
rect 19717 19805 19751 19839
rect 19993 19805 20027 19839
rect 20349 19805 20383 19839
rect 20729 19805 20763 19839
rect 21281 19805 21315 19839
rect 2513 19737 2547 19771
rect 9137 19737 9171 19771
rect 9689 19737 9723 19771
rect 10057 19737 10091 19771
rect 10425 19737 10459 19771
rect 11621 19737 11655 19771
rect 13829 19737 13863 19771
rect 15485 19737 15519 19771
rect 19441 19737 19475 19771
rect 1501 19669 1535 19703
rect 2145 19669 2179 19703
rect 3893 19669 3927 19703
rect 5457 19669 5491 19703
rect 6929 19669 6963 19703
rect 7297 19669 7331 19703
rect 7389 19669 7423 19703
rect 7757 19669 7791 19703
rect 8125 19669 8159 19703
rect 9321 19669 9355 19703
rect 9965 19669 9999 19703
rect 10333 19669 10367 19703
rect 11989 19669 12023 19703
rect 14105 19669 14139 19703
rect 15945 19669 15979 19703
rect 16681 19669 16715 19703
rect 16957 19669 16991 19703
rect 19809 19669 19843 19703
rect 20177 19669 20211 19703
rect 21465 19669 21499 19703
rect 2237 19465 2271 19499
rect 2973 19465 3007 19499
rect 3433 19465 3467 19499
rect 5457 19465 5491 19499
rect 8309 19465 8343 19499
rect 9321 19465 9355 19499
rect 9597 19465 9631 19499
rect 9965 19465 9999 19499
rect 10425 19465 10459 19499
rect 11253 19465 11287 19499
rect 12909 19465 12943 19499
rect 13185 19465 13219 19499
rect 17049 19465 17083 19499
rect 17141 19465 17175 19499
rect 17601 19465 17635 19499
rect 17785 19465 17819 19499
rect 18245 19465 18279 19499
rect 18521 19465 18555 19499
rect 18797 19465 18831 19499
rect 19165 19465 19199 19499
rect 19625 19465 19659 19499
rect 5098 19397 5132 19431
rect 5825 19397 5859 19431
rect 8769 19397 8803 19431
rect 10057 19397 10091 19431
rect 10793 19397 10827 19431
rect 14197 19397 14231 19431
rect 21557 19397 21591 19431
rect 1685 19329 1719 19363
rect 2053 19329 2087 19363
rect 2421 19329 2455 19363
rect 2789 19329 2823 19363
rect 3341 19329 3375 19363
rect 5365 19329 5399 19363
rect 6653 19329 6687 19363
rect 7961 19329 7995 19363
rect 8677 19329 8711 19363
rect 9137 19329 9171 19363
rect 9413 19329 9447 19363
rect 10885 19329 10919 19363
rect 11785 19329 11819 19363
rect 13001 19329 13035 19363
rect 16865 19329 16899 19363
rect 17325 19329 17359 19363
rect 17417 19329 17451 19363
rect 17969 19329 18003 19363
rect 18061 19329 18095 19363
rect 18337 19329 18371 19363
rect 18613 19329 18647 19363
rect 19349 19329 19383 19363
rect 19441 19329 19475 19363
rect 3617 19261 3651 19295
rect 5917 19261 5951 19295
rect 6101 19261 6135 19295
rect 8217 19261 8251 19295
rect 8861 19261 8895 19295
rect 9873 19261 9907 19295
rect 10701 19261 10735 19295
rect 11529 19261 11563 19295
rect 14013 19261 14047 19295
rect 14565 19261 14599 19295
rect 14749 19261 14783 19295
rect 15301 19261 15335 19295
rect 19809 19261 19843 19295
rect 1869 19193 1903 19227
rect 2605 19193 2639 19227
rect 3893 19193 3927 19227
rect 13645 19193 13679 19227
rect 15393 19193 15427 19227
rect 1501 19125 1535 19159
rect 3985 19125 4019 19159
rect 6561 19125 6595 19159
rect 6837 19125 6871 19159
rect 13369 19125 13403 19159
rect 13461 19125 13495 19159
rect 13829 19125 13863 19159
rect 14381 19125 14415 19159
rect 15025 19125 15059 19159
rect 15577 19125 15611 19159
rect 15761 19125 15795 19159
rect 16405 19125 16439 19159
rect 16773 19125 16807 19159
rect 18981 19125 19015 19159
rect 1869 18921 1903 18955
rect 2237 18921 2271 18955
rect 2605 18921 2639 18955
rect 3985 18921 4019 18955
rect 5733 18921 5767 18955
rect 7481 18921 7515 18955
rect 8493 18921 8527 18955
rect 9229 18921 9263 18955
rect 9781 18921 9815 18955
rect 14381 18921 14415 18955
rect 14749 18921 14783 18955
rect 16589 18921 16623 18955
rect 17509 18921 17543 18955
rect 17877 18921 17911 18955
rect 18245 18921 18279 18955
rect 19073 18921 19107 18955
rect 19441 18921 19475 18955
rect 20545 18921 20579 18955
rect 8585 18853 8619 18887
rect 9137 18853 9171 18887
rect 9505 18853 9539 18887
rect 13645 18853 13679 18887
rect 17233 18853 17267 18887
rect 17969 18853 18003 18887
rect 19717 18853 19751 18887
rect 20085 18853 20119 18887
rect 3065 18785 3099 18819
rect 4721 18785 4755 18819
rect 4905 18785 4939 18819
rect 8125 18785 8159 18819
rect 11805 18785 11839 18819
rect 13277 18785 13311 18819
rect 1685 18717 1719 18751
rect 2053 18717 2087 18751
rect 2421 18717 2455 18751
rect 2789 18717 2823 18751
rect 3249 18717 3283 18751
rect 3801 18717 3835 18751
rect 5273 18717 5307 18751
rect 7113 18717 7147 18751
rect 8309 18717 8343 18751
rect 8769 18717 8803 18751
rect 8953 18717 8987 18751
rect 9413 18717 9447 18751
rect 9689 18717 9723 18751
rect 10894 18717 10928 18751
rect 11161 18717 11195 18751
rect 12072 18717 12106 18751
rect 14197 18717 14231 18751
rect 14565 18717 14599 18751
rect 16405 18717 16439 18751
rect 17693 18717 17727 18751
rect 18153 18717 18187 18751
rect 18429 18717 18463 18751
rect 18797 18717 18831 18751
rect 18889 18717 18923 18751
rect 19257 18717 19291 18751
rect 19901 18717 19935 18751
rect 20269 18717 20303 18751
rect 20361 18717 20395 18751
rect 20729 18717 20763 18751
rect 21281 18717 21315 18751
rect 3157 18649 3191 18683
rect 4629 18649 4663 18683
rect 5457 18649 5491 18683
rect 5641 18649 5675 18683
rect 6846 18649 6880 18683
rect 13461 18649 13495 18683
rect 13829 18649 13863 18683
rect 14841 18649 14875 18683
rect 21005 18649 21039 18683
rect 1501 18581 1535 18615
rect 3617 18581 3651 18615
rect 4169 18581 4203 18615
rect 4261 18581 4295 18615
rect 5089 18581 5123 18615
rect 7205 18581 7239 18615
rect 7849 18581 7883 18615
rect 7941 18581 7975 18615
rect 11253 18581 11287 18615
rect 11529 18581 11563 18615
rect 13185 18581 13219 18615
rect 17417 18581 17451 18615
rect 18613 18581 18647 18615
rect 21465 18581 21499 18615
rect 2789 18377 2823 18411
rect 3617 18377 3651 18411
rect 3985 18377 4019 18411
rect 5273 18377 5307 18411
rect 5825 18377 5859 18411
rect 6377 18377 6411 18411
rect 7205 18377 7239 18411
rect 7757 18377 7791 18411
rect 9781 18377 9815 18411
rect 10149 18377 10183 18411
rect 10609 18377 10643 18411
rect 10977 18377 11011 18411
rect 12725 18377 12759 18411
rect 12909 18377 12943 18411
rect 13277 18377 13311 18411
rect 13737 18377 13771 18411
rect 14657 18377 14691 18411
rect 14933 18377 14967 18411
rect 15209 18377 15243 18411
rect 15301 18377 15335 18411
rect 15945 18377 15979 18411
rect 18245 18377 18279 18411
rect 18521 18377 18555 18411
rect 19441 18377 19475 18411
rect 21097 18377 21131 18411
rect 2697 18309 2731 18343
rect 3525 18309 3559 18343
rect 4445 18309 4479 18343
rect 4905 18309 4939 18343
rect 5089 18309 5123 18343
rect 6837 18309 6871 18343
rect 11897 18309 11931 18343
rect 12541 18309 12575 18343
rect 14105 18309 14139 18343
rect 14381 18309 14415 18343
rect 14749 18309 14783 18343
rect 15485 18309 15519 18343
rect 18153 18309 18187 18343
rect 19809 18309 19843 18343
rect 1685 18241 1719 18275
rect 2053 18241 2087 18275
rect 4353 18241 4387 18275
rect 6745 18241 6779 18275
rect 7389 18241 7423 18275
rect 7849 18241 7883 18275
rect 8585 18241 8619 18275
rect 9405 18241 9439 18275
rect 9505 18241 9539 18275
rect 13093 18241 13127 18275
rect 13553 18241 13587 18275
rect 15761 18241 15795 18275
rect 17417 18241 17451 18275
rect 18705 18241 18739 18275
rect 19165 18241 19199 18275
rect 19257 18241 19291 18275
rect 19717 18241 19751 18275
rect 2973 18173 3007 18207
rect 3709 18173 3743 18207
rect 4629 18173 4663 18207
rect 5641 18173 5675 18207
rect 5733 18173 5767 18207
rect 6929 18173 6963 18207
rect 7665 18173 7699 18207
rect 8309 18173 8343 18207
rect 10241 18173 10275 18207
rect 10333 18173 10367 18207
rect 11069 18173 11103 18207
rect 11161 18173 11195 18207
rect 11989 18173 12023 18207
rect 12081 18173 12115 18207
rect 14289 18173 14323 18207
rect 6193 18105 6227 18139
rect 8217 18105 8251 18139
rect 17601 18105 17635 18139
rect 1501 18037 1535 18071
rect 1869 18037 1903 18071
rect 2145 18037 2179 18071
rect 2329 18037 2363 18071
rect 3157 18037 3191 18071
rect 9229 18037 9263 18071
rect 9689 18037 9723 18071
rect 11529 18037 11563 18071
rect 12449 18037 12483 18071
rect 13921 18037 13955 18071
rect 18797 18037 18831 18071
rect 18981 18037 19015 18071
rect 19533 18037 19567 18071
rect 1777 17833 1811 17867
rect 3801 17833 3835 17867
rect 4905 17833 4939 17867
rect 6929 17833 6963 17867
rect 7941 17833 7975 17867
rect 10609 17833 10643 17867
rect 11805 17833 11839 17867
rect 13461 17833 13495 17867
rect 16681 17833 16715 17867
rect 19257 17833 19291 17867
rect 19533 17833 19567 17867
rect 20269 17833 20303 17867
rect 2789 17765 2823 17799
rect 2881 17765 2915 17799
rect 4813 17765 4847 17799
rect 12449 17765 12483 17799
rect 13829 17765 13863 17799
rect 19993 17765 20027 17799
rect 2145 17697 2179 17731
rect 3525 17697 3559 17731
rect 4445 17697 4479 17731
rect 5365 17697 5399 17731
rect 6469 17697 6503 17731
rect 6653 17697 6687 17731
rect 7573 17697 7607 17731
rect 7757 17697 7791 17731
rect 8401 17697 8435 17731
rect 8493 17697 8527 17731
rect 11069 17697 11103 17731
rect 11161 17697 11195 17731
rect 11989 17697 12023 17731
rect 12909 17697 12943 17731
rect 15761 17697 15795 17731
rect 16865 17697 16899 17731
rect 1685 17629 1719 17663
rect 1961 17629 1995 17663
rect 2421 17629 2455 17663
rect 4261 17629 4295 17663
rect 4629 17629 4663 17663
rect 5089 17629 5123 17663
rect 5457 17629 5491 17663
rect 7297 17629 7331 17663
rect 8953 17629 8987 17663
rect 11621 17629 11655 17663
rect 12633 17629 12667 17663
rect 14105 17629 14139 17663
rect 14361 17629 14395 17663
rect 16497 17629 16531 17663
rect 19073 17629 19107 17663
rect 19441 17629 19475 17663
rect 19717 17629 19751 17663
rect 19809 17629 19843 17663
rect 20085 17629 20119 17663
rect 20361 17629 20395 17663
rect 20729 17629 20763 17663
rect 21281 17629 21315 17663
rect 3249 17561 3283 17595
rect 9198 17561 9232 17595
rect 13001 17561 13035 17595
rect 21005 17561 21039 17595
rect 1501 17493 1535 17527
rect 2329 17493 2363 17527
rect 3341 17493 3375 17527
rect 4169 17493 4203 17527
rect 5549 17493 5583 17527
rect 5917 17493 5951 17527
rect 6009 17493 6043 17527
rect 6377 17493 6411 17527
rect 7389 17493 7423 17527
rect 8309 17493 8343 17527
rect 10333 17493 10367 17527
rect 10517 17493 10551 17527
rect 10977 17493 11011 17527
rect 11437 17493 11471 17527
rect 12173 17493 12207 17527
rect 13093 17493 13127 17527
rect 13553 17493 13587 17527
rect 15485 17493 15519 17527
rect 15853 17493 15887 17527
rect 15945 17493 15979 17527
rect 16313 17493 16347 17527
rect 18889 17493 18923 17527
rect 20545 17493 20579 17527
rect 21465 17493 21499 17527
rect 4077 17289 4111 17323
rect 5641 17289 5675 17323
rect 7205 17289 7239 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 10517 17289 10551 17323
rect 10977 17289 11011 17323
rect 11805 17289 11839 17323
rect 12357 17289 12391 17323
rect 14197 17289 14231 17323
rect 14565 17289 14599 17323
rect 15761 17289 15795 17323
rect 16221 17289 16255 17323
rect 17141 17289 17175 17323
rect 19625 17289 19659 17323
rect 19901 17289 19935 17323
rect 20729 17289 20763 17323
rect 21189 17289 21223 17323
rect 2942 17221 2976 17255
rect 4436 17221 4470 17255
rect 7542 17221 7576 17255
rect 11897 17221 11931 17255
rect 14105 17221 14139 17255
rect 17049 17221 17083 17255
rect 1685 17153 1719 17187
rect 1961 17153 1995 17187
rect 2421 17153 2455 17187
rect 2697 17153 2731 17187
rect 4169 17153 4203 17187
rect 5825 17153 5859 17187
rect 6101 17153 6135 17187
rect 6837 17153 6871 17187
rect 8953 17153 8987 17187
rect 9229 17153 9263 17187
rect 9781 17153 9815 17187
rect 10609 17153 10643 17187
rect 13470 17153 13504 17187
rect 13737 17153 13771 17187
rect 14933 17153 14967 17187
rect 15393 17153 15427 17187
rect 16405 17153 16439 17187
rect 20085 17153 20119 17187
rect 20361 17153 20395 17187
rect 20637 17153 20671 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 21281 17153 21315 17187
rect 6653 17085 6687 17119
rect 6745 17085 6779 17119
rect 7297 17085 7331 17119
rect 9873 17085 9907 17119
rect 10057 17085 10091 17119
rect 10333 17085 10367 17119
rect 11713 17085 11747 17119
rect 14013 17085 14047 17119
rect 15117 17085 15151 17119
rect 15301 17085 15335 17119
rect 15853 17085 15887 17119
rect 17233 17085 17267 17119
rect 1869 17017 1903 17051
rect 5917 17017 5951 17051
rect 8677 17017 8711 17051
rect 8769 17017 8803 17051
rect 11253 17017 11287 17051
rect 14749 17017 14783 17051
rect 16681 17017 16715 17051
rect 1501 16949 1535 16983
rect 2145 16949 2179 16983
rect 2237 16949 2271 16983
rect 2605 16949 2639 16983
rect 5549 16949 5583 16983
rect 11069 16949 11103 16983
rect 12265 16949 12299 16983
rect 19441 16949 19475 16983
rect 19809 16949 19843 16983
rect 20177 16949 20211 16983
rect 20453 16949 20487 16983
rect 21465 16949 21499 16983
rect 3801 16745 3835 16779
rect 6469 16745 6503 16779
rect 10885 16745 10919 16779
rect 13553 16745 13587 16779
rect 17141 16745 17175 16779
rect 17325 16745 17359 16779
rect 21005 16745 21039 16779
rect 1869 16677 1903 16711
rect 6193 16677 6227 16711
rect 13093 16677 13127 16711
rect 15669 16677 15703 16711
rect 17785 16677 17819 16711
rect 17969 16677 18003 16711
rect 20729 16677 20763 16711
rect 3249 16609 3283 16643
rect 4445 16609 4479 16643
rect 5365 16609 5399 16643
rect 5457 16609 5491 16643
rect 7849 16609 7883 16643
rect 8585 16609 8619 16643
rect 9321 16609 9355 16643
rect 9505 16609 9539 16643
rect 11345 16609 11379 16643
rect 11529 16609 11563 16643
rect 11713 16609 11747 16643
rect 14289 16609 14323 16643
rect 17417 16609 17451 16643
rect 17693 16609 17727 16643
rect 19993 16609 20027 16643
rect 20177 16609 20211 16643
rect 1685 16541 1719 16575
rect 3525 16541 3559 16575
rect 3985 16541 4019 16575
rect 4261 16541 4295 16575
rect 4721 16541 4755 16575
rect 5549 16541 5583 16575
rect 6009 16541 6043 16575
rect 6285 16541 6319 16575
rect 8493 16541 8527 16575
rect 11253 16541 11287 16575
rect 15761 16541 15795 16575
rect 16017 16541 16051 16575
rect 20537 16541 20571 16575
rect 20821 16541 20855 16575
rect 21097 16541 21131 16575
rect 21281 16541 21315 16575
rect 2982 16473 3016 16507
rect 7582 16473 7616 16507
rect 9772 16473 9806 16507
rect 10977 16473 11011 16507
rect 11980 16473 12014 16507
rect 13369 16473 13403 16507
rect 14556 16473 14590 16507
rect 1501 16405 1535 16439
rect 3341 16405 3375 16439
rect 4077 16405 4111 16439
rect 4629 16405 4663 16439
rect 5089 16405 5123 16439
rect 5917 16405 5951 16439
rect 8033 16405 8067 16439
rect 8401 16405 8435 16439
rect 9045 16405 9079 16439
rect 13185 16405 13219 16439
rect 13921 16405 13955 16439
rect 14197 16405 14231 16439
rect 20361 16405 20395 16439
rect 21465 16405 21499 16439
rect 2145 16201 2179 16235
rect 2605 16201 2639 16235
rect 3985 16201 4019 16235
rect 4445 16201 4479 16235
rect 5273 16201 5307 16235
rect 5733 16201 5767 16235
rect 6193 16201 6227 16235
rect 7205 16201 7239 16235
rect 7665 16201 7699 16235
rect 8125 16201 8159 16235
rect 8769 16201 8803 16235
rect 10333 16201 10367 16235
rect 10609 16201 10643 16235
rect 12633 16201 12667 16235
rect 13001 16201 13035 16235
rect 13829 16201 13863 16235
rect 15025 16201 15059 16235
rect 15393 16201 15427 16235
rect 15853 16201 15887 16235
rect 16221 16201 16255 16235
rect 18153 16201 18187 16235
rect 19165 16201 19199 16235
rect 19901 16201 19935 16235
rect 20545 16201 20579 16235
rect 21005 16201 21039 16235
rect 5825 16133 5859 16167
rect 10425 16133 10459 16167
rect 14289 16133 14323 16167
rect 14933 16133 14967 16167
rect 16313 16133 16347 16167
rect 16948 16133 16982 16167
rect 18337 16133 18371 16167
rect 19717 16133 19751 16167
rect 21097 16133 21131 16167
rect 1685 16065 1719 16099
rect 2973 16065 3007 16099
rect 4813 16065 4847 16099
rect 6377 16065 6411 16099
rect 6837 16065 6871 16099
rect 7297 16065 7331 16099
rect 8953 16065 8987 16099
rect 9220 16065 9254 16099
rect 10977 16065 11011 16099
rect 11069 16065 11103 16099
rect 12541 16065 12575 16099
rect 13369 16065 13403 16099
rect 14197 16065 14231 16099
rect 16681 16065 16715 16099
rect 20729 16065 20763 16099
rect 20829 16065 20863 16099
rect 21281 16065 21315 16099
rect 1869 15997 1903 16031
rect 2053 15997 2087 16031
rect 3065 15997 3099 16031
rect 3249 15997 3283 16031
rect 4077 15997 4111 16031
rect 4169 15997 4203 16031
rect 4905 15997 4939 16031
rect 4997 15997 5031 16031
rect 5549 15997 5583 16031
rect 7021 15997 7055 16031
rect 8217 15997 8251 16031
rect 8309 15997 8343 16031
rect 11161 15997 11195 16031
rect 12725 15997 12759 16031
rect 13461 15997 13495 16031
rect 13553 15997 13587 16031
rect 14381 15997 14415 16031
rect 14841 15997 14875 16031
rect 15577 15997 15611 16031
rect 15761 15997 15795 16031
rect 19349 15997 19383 16031
rect 20085 15997 20119 16031
rect 3617 15929 3651 15963
rect 7757 15929 7791 15963
rect 20177 15929 20211 15963
rect 20361 15929 20395 15963
rect 1501 15861 1535 15895
rect 2513 15861 2547 15895
rect 3525 15861 3559 15895
rect 6561 15861 6595 15895
rect 8585 15861 8619 15895
rect 11529 15861 11563 15895
rect 11713 15861 11747 15895
rect 11897 15861 11931 15895
rect 12173 15861 12207 15895
rect 18061 15861 18095 15895
rect 18521 15861 18555 15895
rect 19533 15861 19567 15895
rect 21465 15861 21499 15895
rect 2237 15657 2271 15691
rect 3985 15657 4019 15691
rect 5457 15657 5491 15691
rect 8769 15657 8803 15691
rect 9413 15657 9447 15691
rect 10425 15657 10459 15691
rect 12265 15657 12299 15691
rect 13185 15657 13219 15691
rect 14473 15657 14507 15691
rect 15301 15657 15335 15691
rect 16681 15657 16715 15691
rect 17233 15657 17267 15691
rect 19073 15657 19107 15691
rect 19533 15657 19567 15691
rect 20177 15657 20211 15691
rect 20361 15657 20395 15691
rect 20821 15657 20855 15691
rect 8953 15589 8987 15623
rect 13093 15589 13127 15623
rect 17325 15589 17359 15623
rect 18705 15589 18739 15623
rect 3617 15521 3651 15555
rect 4537 15521 4571 15555
rect 7481 15521 7515 15555
rect 8217 15521 8251 15555
rect 10149 15521 10183 15555
rect 10977 15521 11011 15555
rect 11713 15521 11747 15555
rect 11805 15521 11839 15555
rect 12541 15521 12575 15555
rect 13737 15521 13771 15555
rect 14749 15521 14783 15555
rect 15485 15521 15519 15555
rect 18153 15521 18187 15555
rect 1685 15453 1719 15487
rect 2053 15453 2087 15487
rect 4169 15453 4203 15487
rect 4261 15453 4295 15487
rect 4813 15453 4847 15487
rect 6570 15453 6604 15487
rect 6837 15453 6871 15487
rect 7941 15453 7975 15487
rect 9137 15453 9171 15487
rect 9229 15453 9263 15487
rect 11897 15453 11931 15487
rect 14933 15453 14967 15487
rect 16221 15453 16255 15487
rect 16589 15453 16623 15487
rect 16865 15453 16899 15487
rect 17509 15453 17543 15487
rect 17601 15453 17635 15487
rect 18337 15453 18371 15487
rect 19993 15453 20027 15487
rect 20545 15453 20579 15487
rect 20637 15453 20671 15487
rect 20913 15453 20947 15487
rect 21281 15453 21315 15487
rect 3372 15385 3406 15419
rect 8401 15385 8435 15419
rect 11253 15385 11287 15419
rect 13553 15385 13587 15419
rect 14105 15385 14139 15419
rect 15761 15385 15795 15419
rect 16957 15385 16991 15419
rect 19625 15385 19659 15419
rect 1501 15317 1535 15351
rect 1869 15317 1903 15351
rect 3801 15317 3835 15351
rect 4445 15317 4479 15351
rect 6929 15317 6963 15351
rect 7297 15317 7331 15351
rect 7389 15317 7423 15351
rect 7757 15317 7791 15351
rect 8309 15317 8343 15351
rect 9597 15317 9631 15351
rect 9965 15317 9999 15351
rect 10057 15317 10091 15351
rect 10793 15317 10827 15351
rect 10885 15317 10919 15351
rect 12633 15317 12667 15351
rect 12725 15317 12759 15351
rect 13645 15317 13679 15351
rect 14841 15317 14875 15351
rect 15669 15317 15703 15351
rect 16129 15317 16163 15351
rect 16405 15317 16439 15351
rect 17785 15317 17819 15351
rect 18245 15317 18279 15351
rect 18797 15317 18831 15351
rect 19349 15317 19383 15351
rect 19901 15317 19935 15351
rect 21097 15317 21131 15351
rect 21465 15317 21499 15351
rect 1869 15113 1903 15147
rect 2421 15113 2455 15147
rect 2789 15113 2823 15147
rect 3985 15113 4019 15147
rect 4445 15113 4479 15147
rect 6193 15113 6227 15147
rect 6745 15113 6779 15147
rect 8401 15113 8435 15147
rect 8493 15113 8527 15147
rect 9965 15113 9999 15147
rect 10333 15113 10367 15147
rect 13001 15113 13035 15147
rect 14013 15113 14047 15147
rect 14933 15113 14967 15147
rect 15393 15113 15427 15147
rect 15853 15113 15887 15147
rect 20453 15113 20487 15147
rect 9606 15045 9640 15079
rect 11796 15045 11830 15079
rect 21097 15045 21131 15079
rect 1685 14977 1719 15011
rect 2053 14977 2087 15011
rect 2329 14977 2363 15011
rect 2605 14977 2639 15011
rect 3157 14977 3191 15011
rect 3617 14977 3651 15011
rect 4353 14977 4387 15011
rect 4813 14977 4847 15011
rect 5080 14977 5114 15011
rect 6929 14977 6963 15011
rect 7021 14977 7055 15011
rect 7277 14977 7311 15011
rect 10425 14977 10459 15011
rect 13369 14977 13403 15011
rect 15761 14977 15795 15011
rect 17805 14977 17839 15011
rect 18420 14977 18454 15011
rect 19993 14977 20027 15011
rect 20269 14977 20303 15011
rect 20545 14977 20579 15011
rect 20821 14977 20855 15011
rect 21281 14977 21315 15011
rect 3249 14909 3283 14943
rect 3433 14909 3467 14943
rect 4629 14909 4663 14943
rect 9873 14909 9907 14943
rect 10609 14909 10643 14943
rect 10793 14909 10827 14943
rect 11529 14909 11563 14943
rect 13461 14909 13495 14943
rect 13553 14909 13587 14943
rect 14749 14909 14783 14943
rect 14841 14909 14875 14943
rect 15945 14909 15979 14943
rect 16405 14909 16439 14943
rect 18061 14909 18095 14943
rect 18153 14909 18187 14943
rect 19809 14909 19843 14943
rect 2145 14841 2179 14875
rect 14197 14841 14231 14875
rect 15301 14841 15335 14875
rect 20177 14841 20211 14875
rect 20729 14841 20763 14875
rect 1501 14773 1535 14807
rect 6377 14773 6411 14807
rect 6653 14773 6687 14807
rect 11069 14773 11103 14807
rect 11345 14773 11379 14807
rect 12909 14773 12943 14807
rect 13829 14773 13863 14807
rect 14473 14773 14507 14807
rect 16681 14773 16715 14807
rect 19533 14773 19567 14807
rect 21005 14773 21039 14807
rect 21465 14773 21499 14807
rect 2789 14569 2823 14603
rect 3985 14569 4019 14603
rect 5181 14569 5215 14603
rect 6009 14569 6043 14603
rect 9965 14569 9999 14603
rect 11897 14569 11931 14603
rect 12265 14569 12299 14603
rect 13093 14569 13127 14603
rect 14105 14569 14139 14603
rect 18889 14569 18923 14603
rect 19993 14569 20027 14603
rect 20913 14569 20947 14603
rect 7113 14501 7147 14535
rect 13277 14501 13311 14535
rect 3433 14433 3467 14467
rect 4721 14433 4755 14467
rect 6561 14433 6595 14467
rect 7849 14433 7883 14467
rect 9413 14433 9447 14467
rect 10609 14433 10643 14467
rect 11345 14433 11379 14467
rect 12449 14433 12483 14467
rect 12633 14433 12667 14467
rect 17509 14433 17543 14467
rect 19349 14433 19383 14467
rect 20637 14433 20671 14467
rect 1685 14365 1719 14399
rect 1869 14365 1903 14399
rect 2329 14365 2363 14399
rect 2605 14365 2639 14399
rect 3801 14365 3835 14399
rect 5089 14365 5123 14399
rect 5733 14365 5767 14399
rect 6653 14365 6687 14399
rect 8309 14365 8343 14399
rect 8493 14365 8527 14399
rect 10517 14365 10551 14399
rect 10977 14365 11011 14399
rect 13461 14365 13495 14399
rect 13737 14365 13771 14399
rect 15485 14365 15519 14399
rect 16957 14365 16991 14399
rect 20453 14365 20487 14399
rect 21097 14365 21131 14399
rect 21281 14365 21315 14399
rect 5917 14297 5951 14331
rect 6745 14297 6779 14331
rect 8585 14297 8619 14331
rect 9597 14297 9631 14331
rect 15240 14297 15274 14331
rect 16712 14297 16746 14331
rect 17776 14297 17810 14331
rect 19625 14297 19659 14331
rect 1501 14229 1535 14263
rect 2053 14229 2087 14263
rect 2145 14229 2179 14263
rect 2421 14229 2455 14263
rect 3157 14229 3191 14263
rect 3249 14229 3283 14263
rect 4077 14229 4111 14263
rect 4445 14229 4479 14263
rect 4537 14229 4571 14263
rect 5549 14229 5583 14263
rect 6285 14229 6319 14263
rect 7205 14229 7239 14263
rect 7573 14229 7607 14263
rect 7665 14229 7699 14263
rect 8033 14229 8067 14263
rect 9137 14229 9171 14263
rect 9505 14229 9539 14263
rect 10057 14229 10091 14263
rect 10425 14229 10459 14263
rect 11437 14229 11471 14263
rect 11529 14229 11563 14263
rect 11989 14229 12023 14263
rect 12725 14229 12759 14263
rect 13553 14229 13587 14263
rect 13921 14229 13955 14263
rect 15577 14229 15611 14263
rect 17141 14229 17175 14263
rect 17417 14229 17451 14263
rect 18981 14229 19015 14263
rect 19533 14229 19567 14263
rect 20085 14229 20119 14263
rect 20545 14229 20579 14263
rect 21465 14229 21499 14263
rect 2329 14025 2363 14059
rect 5917 14025 5951 14059
rect 7205 14025 7239 14059
rect 7757 14025 7791 14059
rect 8769 14025 8803 14059
rect 9137 14025 9171 14059
rect 10333 14025 10367 14059
rect 10885 14025 10919 14059
rect 11253 14025 11287 14059
rect 11529 14025 11563 14059
rect 13553 14025 13587 14059
rect 15209 14025 15243 14059
rect 16037 14025 16071 14059
rect 17509 14025 17543 14059
rect 17969 14025 18003 14059
rect 18521 14025 18555 14059
rect 19349 14025 19383 14059
rect 19717 14025 19751 14059
rect 20821 14025 20855 14059
rect 21097 14025 21131 14059
rect 6101 13957 6135 13991
rect 6745 13957 6779 13991
rect 6837 13957 6871 13991
rect 8493 13957 8527 13991
rect 9229 13957 9263 13991
rect 9965 13957 9999 13991
rect 13369 13957 13403 13991
rect 16405 13957 16439 13991
rect 19809 13957 19843 13991
rect 1685 13889 1719 13923
rect 2053 13889 2087 13923
rect 2145 13889 2179 13923
rect 2605 13889 2639 13923
rect 2981 13893 3015 13927
rect 3332 13889 3366 13923
rect 4793 13889 4827 13923
rect 7665 13889 7699 13923
rect 9873 13889 9907 13923
rect 11897 13889 11931 13923
rect 12357 13889 12391 13923
rect 13737 13889 13771 13923
rect 14004 13889 14038 13923
rect 15577 13889 15611 13923
rect 16221 13889 16255 13923
rect 17233 13889 17267 13923
rect 18061 13889 18095 13923
rect 18889 13889 18923 13923
rect 20453 13889 20487 13923
rect 20637 13889 20671 13923
rect 20913 13889 20947 13923
rect 21281 13889 21315 13923
rect 3065 13821 3099 13855
rect 4537 13821 4571 13855
rect 6561 13821 6595 13855
rect 7849 13821 7883 13855
rect 9413 13821 9447 13855
rect 9689 13821 9723 13855
rect 10425 13821 10459 13855
rect 10701 13821 10735 13855
rect 11161 13821 11195 13855
rect 11989 13821 12023 13855
rect 12081 13821 12115 13855
rect 13001 13821 13035 13855
rect 13185 13821 13219 13855
rect 15669 13821 15703 13855
rect 15853 13821 15887 13855
rect 16681 13821 16715 13855
rect 17141 13821 17175 13855
rect 17877 13821 17911 13855
rect 18981 13821 19015 13855
rect 19165 13821 19199 13855
rect 19901 13821 19935 13855
rect 20177 13821 20211 13855
rect 1869 13753 1903 13787
rect 2421 13753 2455 13787
rect 8125 13753 8159 13787
rect 8309 13753 8343 13787
rect 15117 13753 15151 13787
rect 18429 13753 18463 13787
rect 1501 13685 1535 13719
rect 2789 13685 2823 13719
rect 4445 13685 4479 13719
rect 7297 13685 7331 13719
rect 12633 13685 12667 13719
rect 12817 13685 12851 13719
rect 16865 13685 16899 13719
rect 21465 13685 21499 13719
rect 2237 13481 2271 13515
rect 3893 13481 3927 13515
rect 4629 13481 4663 13515
rect 7021 13481 7055 13515
rect 9045 13481 9079 13515
rect 15117 13481 15151 13515
rect 16037 13481 16071 13515
rect 18061 13481 18095 13515
rect 19441 13481 19475 13515
rect 20729 13481 20763 13515
rect 21005 13481 21039 13515
rect 8493 13413 8527 13447
rect 13553 13413 13587 13447
rect 17049 13413 17083 13447
rect 17969 13413 18003 13447
rect 19349 13413 19383 13447
rect 19625 13413 19659 13447
rect 5181 13345 5215 13379
rect 5917 13345 5951 13379
rect 6009 13345 6043 13379
rect 6377 13345 6411 13379
rect 7113 13345 7147 13379
rect 9689 13345 9723 13379
rect 11621 13345 11655 13379
rect 14565 13345 14599 13379
rect 15853 13345 15887 13379
rect 16589 13345 16623 13379
rect 17417 13345 17451 13379
rect 18705 13345 18739 13379
rect 1685 13277 1719 13311
rect 2053 13277 2087 13311
rect 3617 13277 3651 13311
rect 5089 13277 5123 13311
rect 6653 13277 6687 13311
rect 7369 13277 7403 13311
rect 10149 13277 10183 13311
rect 11877 13277 11911 13311
rect 13737 13277 13771 13311
rect 14657 13277 14691 13311
rect 15669 13277 15703 13311
rect 16405 13277 16439 13311
rect 17509 13277 17543 13311
rect 20177 13277 20211 13311
rect 20545 13277 20579 13311
rect 20821 13277 20855 13311
rect 21097 13277 21131 13311
rect 21281 13277 21315 13311
rect 3350 13209 3384 13243
rect 3985 13209 4019 13243
rect 9137 13209 9171 13243
rect 9505 13209 9539 13243
rect 10416 13209 10450 13243
rect 13369 13209 13403 13243
rect 13829 13209 13863 13243
rect 14749 13209 14783 13243
rect 16497 13209 16531 13243
rect 18889 13209 18923 13243
rect 20453 13209 20487 13243
rect 1501 13141 1535 13175
rect 1869 13141 1903 13175
rect 4261 13141 4295 13175
rect 4997 13141 5031 13175
rect 5457 13141 5491 13175
rect 5825 13141 5859 13175
rect 6561 13141 6595 13175
rect 8677 13141 8711 13175
rect 9781 13141 9815 13175
rect 9965 13141 9999 13175
rect 11529 13141 11563 13175
rect 13001 13141 13035 13175
rect 13093 13141 13127 13175
rect 14197 13141 14231 13175
rect 15209 13141 15243 13175
rect 15577 13141 15611 13175
rect 16957 13141 16991 13175
rect 17601 13141 17635 13175
rect 18429 13141 18463 13175
rect 18521 13141 18555 13175
rect 19901 13141 19935 13175
rect 20085 13141 20119 13175
rect 21465 13141 21499 13175
rect 3433 12937 3467 12971
rect 4445 12937 4479 12971
rect 5917 12937 5951 12971
rect 6561 12937 6595 12971
rect 7665 12937 7699 12971
rect 8033 12937 8067 12971
rect 8125 12937 8159 12971
rect 10425 12937 10459 12971
rect 10885 12937 10919 12971
rect 11345 12937 11379 12971
rect 12265 12937 12299 12971
rect 12633 12937 12667 12971
rect 14105 12937 14139 12971
rect 15301 12937 15335 12971
rect 15761 12937 15795 12971
rect 16037 12937 16071 12971
rect 16681 12937 16715 12971
rect 19349 12937 19383 12971
rect 1869 12869 1903 12903
rect 9505 12869 9539 12903
rect 11529 12869 11563 12903
rect 12992 12869 13026 12903
rect 15393 12869 15427 12903
rect 17049 12869 17083 12903
rect 18144 12869 18178 12903
rect 19809 12869 19843 12903
rect 20637 12869 20671 12903
rect 1685 12801 1719 12835
rect 2217 12801 2251 12835
rect 3617 12801 3651 12835
rect 4077 12801 4111 12835
rect 4905 12801 4939 12835
rect 4997 12801 5031 12835
rect 5825 12801 5859 12835
rect 7205 12801 7239 12835
rect 8953 12801 8987 12835
rect 10977 12801 11011 12835
rect 12725 12801 12759 12835
rect 15945 12801 15979 12835
rect 17601 12801 17635 12835
rect 17877 12801 17911 12835
rect 19533 12801 19567 12835
rect 20821 12801 20855 12835
rect 21281 12801 21315 12835
rect 1961 12733 1995 12767
rect 3893 12733 3927 12767
rect 3985 12733 4019 12767
rect 5181 12733 5215 12767
rect 6101 12733 6135 12767
rect 7297 12733 7331 12767
rect 7389 12733 7423 12767
rect 8217 12733 8251 12767
rect 9045 12733 9079 12767
rect 9137 12733 9171 12767
rect 9781 12733 9815 12767
rect 10793 12733 10827 12767
rect 11989 12733 12023 12767
rect 12173 12733 12207 12767
rect 15209 12733 15243 12767
rect 16313 12733 16347 12767
rect 17141 12733 17175 12767
rect 17233 12733 17267 12767
rect 3341 12665 3375 12699
rect 4537 12665 4571 12699
rect 5457 12665 5491 12699
rect 14565 12665 14599 12699
rect 16405 12665 16439 12699
rect 19993 12665 20027 12699
rect 20453 12665 20487 12699
rect 21189 12665 21223 12699
rect 1501 12597 1535 12631
rect 6653 12597 6687 12631
rect 6837 12597 6871 12631
rect 8585 12597 8619 12631
rect 9597 12597 9631 12631
rect 10057 12597 10091 12631
rect 10241 12597 10275 12631
rect 11805 12597 11839 12631
rect 14197 12597 14231 12631
rect 14473 12597 14507 12631
rect 14749 12597 14783 12631
rect 17785 12597 17819 12631
rect 19257 12597 19291 12631
rect 19717 12597 19751 12631
rect 20269 12597 20303 12631
rect 21005 12597 21039 12631
rect 21465 12597 21499 12631
rect 1593 12393 1627 12427
rect 3249 12393 3283 12427
rect 3801 12393 3835 12427
rect 5365 12393 5399 12427
rect 7205 12393 7239 12427
rect 8033 12393 8067 12427
rect 11805 12393 11839 12427
rect 11897 12393 11931 12427
rect 13829 12393 13863 12427
rect 16773 12393 16807 12427
rect 19257 12393 19291 12427
rect 20269 12393 20303 12427
rect 21005 12393 21039 12427
rect 4721 12325 4755 12359
rect 8953 12325 8987 12359
rect 12817 12325 12851 12359
rect 13093 12325 13127 12359
rect 2973 12257 3007 12291
rect 4353 12257 4387 12291
rect 7757 12257 7791 12291
rect 8493 12257 8527 12291
rect 8585 12257 8619 12291
rect 10326 12257 10360 12291
rect 10425 12257 10459 12291
rect 12449 12257 12483 12291
rect 16589 12257 16623 12291
rect 17693 12257 17727 12291
rect 19809 12257 19843 12291
rect 3065 12189 3099 12223
rect 3525 12189 3559 12223
rect 4169 12189 4203 12223
rect 6754 12189 6788 12223
rect 7021 12189 7055 12223
rect 12265 12189 12299 12223
rect 13001 12189 13035 12223
rect 14565 12189 14599 12223
rect 14841 12189 14875 12223
rect 20085 12189 20119 12223
rect 20821 12189 20855 12223
rect 21281 12189 21315 12223
rect 2706 12121 2740 12155
rect 5089 12121 5123 12155
rect 10066 12121 10100 12155
rect 10692 12121 10726 12155
rect 13369 12121 13403 12155
rect 15086 12121 15120 12155
rect 16957 12121 16991 12155
rect 17960 12121 17994 12155
rect 19625 12121 19659 12155
rect 19717 12121 19751 12155
rect 21189 12121 21223 12155
rect 1501 12053 1535 12087
rect 3341 12053 3375 12087
rect 4261 12053 4295 12087
rect 4905 12053 4939 12087
rect 5457 12053 5491 12087
rect 5641 12053 5675 12087
rect 7573 12053 7607 12087
rect 7665 12053 7699 12087
rect 8401 12053 8435 12087
rect 12357 12053 12391 12087
rect 13461 12053 13495 12087
rect 14105 12053 14139 12087
rect 14381 12053 14415 12087
rect 16221 12053 16255 12087
rect 16405 12053 16439 12087
rect 17049 12053 17083 12087
rect 17233 12053 17267 12087
rect 17509 12053 17543 12087
rect 19073 12053 19107 12087
rect 20545 12053 20579 12087
rect 20729 12053 20763 12087
rect 21465 12053 21499 12087
rect 2789 11849 2823 11883
rect 3157 11849 3191 11883
rect 3617 11849 3651 11883
rect 4445 11849 4479 11883
rect 5457 11849 5491 11883
rect 8033 11849 8067 11883
rect 8861 11849 8895 11883
rect 10333 11849 10367 11883
rect 11345 11849 11379 11883
rect 11897 11849 11931 11883
rect 12265 11849 12299 11883
rect 12449 11849 12483 11883
rect 15301 11849 15335 11883
rect 18061 11849 18095 11883
rect 18981 11849 19015 11883
rect 19349 11849 19383 11883
rect 19809 11849 19843 11883
rect 20361 11849 20395 11883
rect 20637 11849 20671 11883
rect 5917 11781 5951 11815
rect 9321 11781 9355 11815
rect 9965 11781 9999 11815
rect 10885 11781 10919 11815
rect 12633 11781 12667 11815
rect 16405 11781 16439 11815
rect 2237 11713 2271 11747
rect 2421 11713 2455 11747
rect 3985 11713 4019 11747
rect 4629 11713 4663 11747
rect 5825 11713 5859 11747
rect 7490 11713 7524 11747
rect 7757 11713 7791 11747
rect 7941 11713 7975 11747
rect 8401 11713 8435 11747
rect 8493 11713 8527 11747
rect 9229 11713 9263 11747
rect 10517 11713 10551 11747
rect 10977 11713 11011 11747
rect 13277 11713 13311 11747
rect 13369 11713 13403 11747
rect 14953 11713 14987 11747
rect 15209 11713 15243 11747
rect 15669 11713 15703 11747
rect 15761 11713 15795 11747
rect 16681 11713 16715 11747
rect 16948 11713 16982 11747
rect 18521 11713 18555 11747
rect 19441 11713 19475 11747
rect 20177 11713 20211 11747
rect 20453 11713 20487 11747
rect 21281 11713 21315 11747
rect 1961 11645 1995 11679
rect 2605 11645 2639 11679
rect 3249 11645 3283 11679
rect 3341 11645 3375 11679
rect 4077 11645 4111 11679
rect 4169 11645 4203 11679
rect 5089 11645 5123 11679
rect 6101 11645 6135 11679
rect 8677 11645 8711 11679
rect 9413 11645 9447 11679
rect 9781 11645 9815 11679
rect 10793 11645 10827 11679
rect 11621 11645 11655 11679
rect 11805 11645 11839 11679
rect 13185 11645 13219 11679
rect 15853 11645 15887 11679
rect 18245 11645 18279 11679
rect 18429 11645 18463 11679
rect 19533 11645 19567 11679
rect 21557 11645 21591 11679
rect 13829 11577 13863 11611
rect 18889 11577 18923 11611
rect 4721 11509 4755 11543
rect 5181 11509 5215 11543
rect 6377 11509 6411 11543
rect 10149 11509 10183 11543
rect 12817 11509 12851 11543
rect 13737 11509 13771 11543
rect 16221 11509 16255 11543
rect 19993 11509 20027 11543
rect 2145 11305 2179 11339
rect 3617 11305 3651 11339
rect 4169 11305 4203 11339
rect 8585 11305 8619 11339
rect 9137 11305 9171 11339
rect 9873 11305 9907 11339
rect 11713 11305 11747 11339
rect 12541 11305 12575 11339
rect 15025 11305 15059 11339
rect 15485 11305 15519 11339
rect 18521 11305 18555 11339
rect 19533 11305 19567 11339
rect 20361 11305 20395 11339
rect 21005 11305 21039 11339
rect 21373 11305 21407 11339
rect 5825 11237 5859 11271
rect 9965 11237 9999 11271
rect 10885 11237 10919 11271
rect 12633 11237 12667 11271
rect 13001 11237 13035 11271
rect 14105 11237 14139 11271
rect 15577 11237 15611 11271
rect 17693 11237 17727 11271
rect 19349 11237 19383 11271
rect 20269 11237 20303 11271
rect 20821 11237 20855 11271
rect 1501 11169 1535 11203
rect 1685 11169 1719 11203
rect 2237 11169 2271 11203
rect 4813 11169 4847 11203
rect 5181 11169 5215 11203
rect 6377 11169 6411 11203
rect 10333 11169 10367 11203
rect 11161 11169 11195 11203
rect 11897 11169 11931 11203
rect 12081 11169 12115 11203
rect 13461 11169 13495 11203
rect 13553 11169 13587 11203
rect 13829 11169 13863 11203
rect 14657 11169 14691 11203
rect 16313 11169 16347 11203
rect 17969 11169 18003 11203
rect 3801 11101 3835 11135
rect 4629 11101 4663 11135
rect 6285 11101 6319 11135
rect 6745 11101 6779 11135
rect 8493 11101 8527 11135
rect 9413 11101 9447 11135
rect 9689 11101 9723 11135
rect 10517 11101 10551 11135
rect 12817 11101 12851 11135
rect 13369 11101 13403 11135
rect 14565 11101 14599 11135
rect 15209 11101 15243 11135
rect 16129 11101 16163 11135
rect 18613 11101 18647 11135
rect 19717 11101 19751 11135
rect 20085 11101 20119 11135
rect 20545 11101 20579 11135
rect 20637 11101 20671 11135
rect 21465 11101 21499 11135
rect 2504 11033 2538 11067
rect 4537 11033 4571 11067
rect 5365 11033 5399 11067
rect 6990 11033 7024 11067
rect 8309 11033 8343 11067
rect 9045 11033 9079 11067
rect 11345 11033 11379 11067
rect 12173 11033 12207 11067
rect 14473 11033 14507 11067
rect 16580 11033 16614 11067
rect 18153 11033 18187 11067
rect 19073 11033 19107 11067
rect 21097 11033 21131 11067
rect 1777 10965 1811 10999
rect 3985 10965 4019 10999
rect 5273 10965 5307 10999
rect 5733 10965 5767 10999
rect 6193 10965 6227 10999
rect 8125 10965 8159 10999
rect 10425 10965 10459 10999
rect 11253 10965 11287 10999
rect 15761 10965 15795 10999
rect 15945 10965 15979 10999
rect 18061 10965 18095 10999
rect 18797 10965 18831 10999
rect 19901 10965 19935 10999
rect 3801 10761 3835 10795
rect 4169 10761 4203 10795
rect 5457 10761 5491 10795
rect 6009 10761 6043 10795
rect 7389 10761 7423 10795
rect 7665 10761 7699 10795
rect 8217 10761 8251 10795
rect 8309 10761 8343 10795
rect 8953 10761 8987 10795
rect 11345 10761 11379 10795
rect 11713 10761 11747 10795
rect 12357 10761 12391 10795
rect 12541 10761 12575 10795
rect 14473 10761 14507 10795
rect 14841 10761 14875 10795
rect 15209 10761 15243 10795
rect 15669 10761 15703 10795
rect 16037 10761 16071 10795
rect 17049 10761 17083 10795
rect 17417 10761 17451 10795
rect 17785 10761 17819 10795
rect 18245 10761 18279 10795
rect 18337 10761 18371 10795
rect 18797 10761 18831 10795
rect 19165 10761 19199 10795
rect 19533 10761 19567 10795
rect 19993 10761 20027 10795
rect 20361 10761 20395 10795
rect 20453 10761 20487 10795
rect 1501 10693 1535 10727
rect 3249 10693 3283 10727
rect 3709 10693 3743 10727
rect 9781 10693 9815 10727
rect 13676 10693 13710 10727
rect 16957 10693 16991 10727
rect 18705 10693 18739 10727
rect 1777 10625 1811 10659
rect 2044 10625 2078 10659
rect 4629 10625 4663 10659
rect 6745 10625 6779 10659
rect 8677 10625 8711 10659
rect 9413 10625 9447 10659
rect 9965 10625 9999 10659
rect 10232 10625 10266 10659
rect 11897 10625 11931 10659
rect 14381 10625 14415 10659
rect 17877 10625 17911 10659
rect 21189 10625 21223 10659
rect 21281 10625 21315 10659
rect 3617 10557 3651 10591
rect 4721 10557 4755 10591
rect 4905 10557 4939 10591
rect 5549 10557 5583 10591
rect 5641 10557 5675 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 8401 10557 8435 10591
rect 9137 10557 9171 10591
rect 13921 10557 13955 10591
rect 14565 10557 14599 10591
rect 15301 10557 15335 10591
rect 15393 10557 15427 10591
rect 16129 10557 16163 10591
rect 16221 10557 16255 10591
rect 16865 10557 16899 10591
rect 17601 10557 17635 10591
rect 18889 10557 18923 10591
rect 19625 10557 19659 10591
rect 19717 10557 19751 10591
rect 20545 10557 20579 10591
rect 21465 10557 21499 10591
rect 4261 10489 4295 10523
rect 5089 10489 5123 10523
rect 6377 10489 6411 10523
rect 7297 10489 7331 10523
rect 1593 10421 1627 10455
rect 3157 10421 3191 10455
rect 7849 10421 7883 10455
rect 9229 10421 9263 10455
rect 9689 10421 9723 10455
rect 12081 10421 12115 10455
rect 12173 10421 12207 10455
rect 14013 10421 14047 10455
rect 20821 10421 20855 10455
rect 1869 10217 1903 10251
rect 3985 10217 4019 10251
rect 5181 10217 5215 10251
rect 10517 10217 10551 10251
rect 11897 10217 11931 10251
rect 12081 10217 12115 10251
rect 14105 10217 14139 10251
rect 14933 10217 14967 10251
rect 17325 10217 17359 10251
rect 18889 10217 18923 10251
rect 4077 10149 4111 10183
rect 6377 10149 6411 10183
rect 10609 10149 10643 10183
rect 11805 10149 11839 10183
rect 13921 10149 13955 10183
rect 18981 10149 19015 10183
rect 19257 10149 19291 10183
rect 21005 10149 21039 10183
rect 2513 10081 2547 10115
rect 3341 10081 3375 10115
rect 4629 10081 4663 10115
rect 6193 10081 6227 10115
rect 8401 10081 8435 10115
rect 9137 10081 9171 10115
rect 11161 10081 11195 10115
rect 12265 10081 12299 10115
rect 14657 10081 14691 10115
rect 15485 10081 15519 10115
rect 15945 10081 15979 10115
rect 16773 10081 16807 10115
rect 17509 10081 17543 10115
rect 20913 10081 20947 10115
rect 1501 10013 1535 10047
rect 3157 10013 3191 10047
rect 3801 10013 3835 10047
rect 4261 10013 4295 10047
rect 5457 10013 5491 10047
rect 6653 10013 6687 10047
rect 6929 10013 6963 10047
rect 8134 10013 8168 10047
rect 9045 10013 9079 10047
rect 12532 10013 12566 10047
rect 16129 10013 16163 10047
rect 16865 10013 16899 10047
rect 19441 10013 19475 10047
rect 21189 10013 21223 10047
rect 21465 10013 21499 10047
rect 1685 9945 1719 9979
rect 6009 9945 6043 9979
rect 8677 9945 8711 9979
rect 9382 9945 9416 9979
rect 10977 9945 11011 9979
rect 11437 9945 11471 9979
rect 17776 9945 17810 9979
rect 20646 9945 20680 9979
rect 2237 9877 2271 9911
rect 2329 9877 2363 9911
rect 2697 9877 2731 9911
rect 3065 9877 3099 9911
rect 3525 9877 3559 9911
rect 4721 9877 4755 9911
rect 4813 9877 4847 9911
rect 5273 9877 5307 9911
rect 5549 9877 5583 9911
rect 5917 9877 5951 9911
rect 6745 9877 6779 9911
rect 7021 9877 7055 9911
rect 8585 9877 8619 9911
rect 11069 9877 11103 9911
rect 13645 9877 13679 9911
rect 14473 9877 14507 9911
rect 14565 9877 14599 9911
rect 15301 9877 15335 9911
rect 15393 9877 15427 9911
rect 16037 9877 16071 9911
rect 16497 9877 16531 9911
rect 16957 9877 16991 9911
rect 19533 9877 19567 9911
rect 21373 9877 21407 9911
rect 2145 9673 2179 9707
rect 2605 9673 2639 9707
rect 4077 9673 4111 9707
rect 4537 9673 4571 9707
rect 4905 9673 4939 9707
rect 5825 9673 5859 9707
rect 6745 9673 6779 9707
rect 7389 9673 7423 9707
rect 10701 9673 10735 9707
rect 14565 9673 14599 9707
rect 15025 9673 15059 9707
rect 15393 9673 15427 9707
rect 15669 9673 15703 9707
rect 16773 9673 16807 9707
rect 17601 9673 17635 9707
rect 20637 9673 20671 9707
rect 20729 9673 20763 9707
rect 6561 9605 6595 9639
rect 8217 9605 8251 9639
rect 13369 9605 13403 9639
rect 16405 9605 16439 9639
rect 18061 9605 18095 9639
rect 1501 9537 1535 9571
rect 1777 9537 1811 9571
rect 2513 9537 2547 9571
rect 3801 9537 3835 9571
rect 4169 9537 4203 9571
rect 5733 9537 5767 9571
rect 8309 9537 8343 9571
rect 8861 9537 8895 9571
rect 9128 9537 9162 9571
rect 11345 9537 11379 9571
rect 12653 9537 12687 9571
rect 13277 9537 13311 9571
rect 14197 9537 14231 9571
rect 16221 9537 16255 9571
rect 17141 9537 17175 9571
rect 17969 9537 18003 9571
rect 18429 9537 18463 9571
rect 18613 9537 18647 9571
rect 19073 9537 19107 9571
rect 19524 9537 19558 9571
rect 21097 9537 21131 9571
rect 2697 9469 2731 9503
rect 4997 9469 5031 9503
rect 5089 9469 5123 9503
rect 5917 9469 5951 9503
rect 7481 9469 7515 9503
rect 7665 9469 7699 9503
rect 8401 9469 8435 9503
rect 10425 9469 10459 9503
rect 10609 9469 10643 9503
rect 12909 9469 12943 9503
rect 13185 9469 13219 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 16037 9469 16071 9503
rect 17233 9469 17267 9503
rect 17417 9469 17451 9503
rect 18245 9469 18279 9503
rect 19257 9469 19291 9503
rect 21189 9469 21223 9503
rect 21281 9469 21315 9503
rect 1961 9401 1995 9435
rect 5365 9401 5399 9435
rect 6377 9401 6411 9435
rect 15209 9401 15243 9435
rect 18889 9401 18923 9435
rect 1593 9333 1627 9367
rect 3571 9333 3605 9367
rect 4353 9333 4387 9367
rect 7021 9333 7055 9367
rect 7849 9333 7883 9367
rect 8677 9333 8711 9367
rect 10241 9333 10275 9367
rect 11069 9333 11103 9367
rect 11161 9333 11195 9367
rect 11529 9333 11563 9367
rect 13737 9333 13771 9367
rect 14657 9333 14691 9367
rect 14933 9333 14967 9367
rect 15761 9333 15795 9367
rect 18797 9333 18831 9367
rect 1961 9129 1995 9163
rect 2053 9129 2087 9163
rect 2881 9129 2915 9163
rect 3801 9129 3835 9163
rect 7573 9129 7607 9163
rect 9137 9129 9171 9163
rect 9413 9129 9447 9163
rect 10333 9129 10367 9163
rect 11989 9129 12023 9163
rect 12817 9129 12851 9163
rect 16589 9129 16623 9163
rect 17601 9129 17635 9163
rect 20729 9129 20763 9163
rect 4261 9061 4295 9095
rect 7297 9061 7331 9095
rect 12081 9061 12115 9095
rect 20637 9061 20671 9095
rect 2697 8993 2731 9027
rect 3341 8993 3375 9027
rect 3525 8993 3559 9027
rect 8125 8993 8159 9027
rect 8401 8993 8435 9027
rect 9781 8993 9815 9027
rect 10517 8993 10551 9027
rect 11345 8993 11379 9027
rect 13921 8993 13955 9027
rect 15945 8993 15979 9027
rect 17233 8993 17267 9027
rect 18521 8993 18555 9027
rect 19257 8993 19291 9027
rect 21281 8993 21315 9027
rect 1409 8925 1443 8959
rect 1777 8925 1811 8959
rect 3985 8925 4019 8959
rect 4077 8925 4111 8959
rect 4353 8925 4387 8959
rect 5825 8925 5859 8959
rect 7481 8925 7515 8959
rect 8769 8925 8803 8959
rect 10793 8925 10827 8959
rect 12449 8925 12483 8959
rect 13001 8925 13035 8959
rect 15229 8925 15263 8959
rect 15485 8925 15519 8959
rect 15761 8925 15795 8959
rect 17141 8925 17175 8959
rect 17877 8925 17911 8959
rect 17969 8925 18003 8959
rect 21189 8925 21223 8959
rect 4620 8857 4654 8891
rect 6092 8857 6126 8891
rect 13645 8857 13679 8891
rect 16221 8857 16255 8891
rect 18705 8857 18739 8891
rect 19524 8857 19558 8891
rect 1593 8789 1627 8823
rect 2421 8789 2455 8823
rect 2513 8789 2547 8823
rect 3249 8789 3283 8823
rect 5733 8789 5767 8823
rect 7205 8789 7239 8823
rect 7941 8789 7975 8823
rect 8033 8789 8067 8823
rect 8585 8789 8619 8823
rect 8953 8789 8987 8823
rect 9873 8789 9907 8823
rect 9965 8789 9999 8823
rect 10701 8789 10735 8823
rect 11161 8789 11195 8823
rect 11529 8789 11563 8823
rect 11621 8789 11655 8823
rect 12541 8789 12575 8823
rect 13093 8789 13127 8823
rect 13369 8789 13403 8823
rect 13553 8789 13587 8823
rect 14105 8789 14139 8823
rect 15577 8789 15611 8823
rect 16129 8789 16163 8823
rect 16681 8789 16715 8823
rect 17049 8789 17083 8823
rect 17693 8789 17727 8823
rect 18153 8789 18187 8823
rect 18613 8789 18647 8823
rect 19073 8789 19107 8823
rect 21097 8789 21131 8823
rect 2237 8585 2271 8619
rect 5181 8585 5215 8619
rect 6561 8585 6595 8619
rect 6929 8585 6963 8619
rect 7389 8585 7423 8619
rect 7849 8585 7883 8619
rect 8953 8585 8987 8619
rect 9413 8585 9447 8619
rect 9781 8585 9815 8619
rect 9965 8585 9999 8619
rect 10885 8585 10919 8619
rect 11345 8585 11379 8619
rect 11529 8585 11563 8619
rect 13369 8585 13403 8619
rect 13829 8585 13863 8619
rect 14197 8585 14231 8619
rect 14657 8585 14691 8619
rect 16681 8585 16715 8619
rect 17509 8585 17543 8619
rect 18613 8585 18647 8619
rect 19993 8585 20027 8619
rect 20959 8585 20993 8619
rect 1869 8517 1903 8551
rect 4068 8517 4102 8551
rect 10977 8517 11011 8551
rect 13461 8517 13495 8551
rect 15292 8517 15326 8551
rect 17141 8517 17175 8551
rect 18705 8517 18739 8551
rect 20545 8517 20579 8551
rect 2585 8449 2619 8483
rect 5273 8449 5307 8483
rect 5825 8449 5859 8483
rect 7757 8449 7791 8483
rect 8585 8449 8619 8483
rect 10425 8449 10459 8483
rect 12653 8449 12687 8483
rect 12909 8449 12943 8483
rect 14289 8449 14323 8483
rect 14841 8449 14875 8483
rect 17049 8449 17083 8483
rect 17877 8449 17911 8483
rect 17969 8449 18003 8483
rect 19625 8449 19659 8483
rect 1685 8381 1719 8415
rect 1777 8381 1811 8415
rect 2329 8381 2363 8415
rect 3801 8381 3835 8415
rect 5549 8381 5583 8415
rect 5733 8381 5767 8415
rect 7021 8381 7055 8415
rect 7113 8381 7147 8415
rect 7941 8381 7975 8415
rect 8401 8381 8435 8415
rect 8493 8381 8527 8415
rect 9137 8381 9171 8415
rect 9321 8381 9355 8415
rect 10057 8381 10091 8415
rect 10793 8381 10827 8415
rect 13553 8381 13587 8415
rect 14381 8381 14415 8415
rect 15025 8381 15059 8415
rect 17233 8381 17267 8415
rect 18061 8381 18095 8415
rect 18521 8381 18555 8415
rect 19349 8381 19383 8415
rect 19533 8381 19567 8415
rect 20269 8381 20303 8415
rect 20729 8381 20763 8415
rect 3709 8313 3743 8347
rect 10333 8313 10367 8347
rect 16405 8313 16439 8347
rect 19073 8313 19107 8347
rect 6193 8245 6227 8279
rect 6469 8245 6503 8279
rect 13001 8245 13035 8279
rect 20453 8245 20487 8279
rect 1777 8041 1811 8075
rect 3801 8041 3835 8075
rect 5457 8041 5491 8075
rect 8769 8041 8803 8075
rect 10333 8041 10367 8075
rect 10701 8041 10735 8075
rect 12449 8041 12483 8075
rect 14105 8041 14139 8075
rect 15577 8041 15611 8075
rect 19993 8041 20027 8075
rect 21373 8041 21407 8075
rect 4629 7973 4663 8007
rect 15485 7973 15519 8007
rect 17601 7973 17635 8007
rect 19073 7973 19107 8007
rect 3617 7905 3651 7939
rect 4353 7905 4387 7939
rect 5181 7905 5215 7939
rect 5917 7905 5951 7939
rect 6009 7905 6043 7939
rect 6837 7905 6871 7939
rect 7297 7905 7331 7939
rect 7481 7905 7515 7939
rect 8217 7905 8251 7939
rect 10977 7905 11011 7939
rect 13001 7905 13035 7939
rect 14657 7905 14691 7939
rect 16957 7905 16991 7939
rect 17233 7905 17267 7939
rect 17693 7905 17727 7939
rect 19441 7905 19475 7939
rect 19533 7905 19567 7939
rect 20177 7905 20211 7939
rect 1501 7837 1535 7871
rect 2890 7837 2924 7871
rect 3157 7837 3191 7871
rect 3249 7837 3283 7871
rect 4169 7837 4203 7871
rect 6745 7837 6779 7871
rect 8953 7837 8987 7871
rect 11244 7837 11278 7871
rect 12817 7837 12851 7871
rect 13277 7837 13311 7871
rect 14473 7837 14507 7871
rect 15117 7837 15151 7871
rect 15301 7837 15335 7871
rect 16690 7837 16724 7871
rect 17417 7837 17451 7871
rect 20453 7837 20487 7871
rect 21465 7837 21499 7871
rect 1685 7769 1719 7803
rect 4997 7769 5031 7803
rect 8401 7769 8435 7803
rect 9198 7769 9232 7803
rect 10517 7769 10551 7803
rect 13185 7769 13219 7803
rect 13737 7769 13771 7803
rect 17960 7769 17994 7803
rect 21097 7769 21131 7803
rect 3433 7701 3467 7735
rect 4261 7701 4295 7735
rect 5089 7701 5123 7735
rect 5825 7701 5859 7735
rect 6285 7701 6319 7735
rect 6653 7701 6687 7735
rect 7573 7701 7607 7735
rect 7941 7701 7975 7735
rect 8309 7701 8343 7735
rect 10885 7701 10919 7735
rect 12357 7701 12391 7735
rect 13645 7701 13679 7735
rect 14565 7701 14599 7735
rect 14933 7701 14967 7735
rect 19625 7701 19659 7735
rect 5365 7497 5399 7531
rect 5825 7497 5859 7531
rect 6377 7497 6411 7531
rect 6745 7497 6779 7531
rect 7665 7497 7699 7531
rect 9137 7497 9171 7531
rect 9597 7497 9631 7531
rect 10057 7497 10091 7531
rect 10885 7497 10919 7531
rect 11621 7497 11655 7531
rect 11989 7497 12023 7531
rect 12081 7497 12115 7531
rect 12725 7497 12759 7531
rect 12817 7497 12851 7531
rect 13277 7497 13311 7531
rect 13645 7497 13679 7531
rect 13737 7497 13771 7531
rect 14105 7497 14139 7531
rect 15577 7497 15611 7531
rect 16037 7497 16071 7531
rect 17233 7497 17267 7531
rect 18337 7497 18371 7531
rect 18797 7497 18831 7531
rect 19257 7497 19291 7531
rect 19717 7497 19751 7531
rect 20177 7497 20211 7531
rect 20821 7497 20855 7531
rect 21281 7497 21315 7531
rect 21373 7497 21407 7531
rect 1501 7429 1535 7463
rect 5917 7429 5951 7463
rect 6837 7429 6871 7463
rect 9505 7429 9539 7463
rect 2982 7361 3016 7395
rect 3249 7361 3283 7395
rect 3893 7361 3927 7395
rect 3985 7361 4019 7395
rect 4252 7361 4286 7395
rect 7297 7361 7331 7395
rect 7573 7361 7607 7395
rect 8778 7361 8812 7395
rect 9045 7361 9079 7395
rect 10977 7361 11011 7395
rect 14473 7361 14507 7395
rect 14565 7361 14599 7395
rect 15209 7361 15243 7395
rect 15761 7361 15795 7395
rect 16221 7361 16255 7395
rect 16497 7361 16531 7395
rect 16681 7361 16715 7395
rect 16957 7361 16991 7395
rect 17601 7361 17635 7395
rect 17693 7361 17727 7395
rect 18429 7361 18463 7395
rect 20085 7361 20119 7395
rect 20913 7361 20947 7395
rect 21557 7361 21591 7395
rect 3341 7293 3375 7327
rect 6009 7293 6043 7327
rect 6929 7293 6963 7327
rect 9689 7293 9723 7327
rect 10241 7293 10275 7327
rect 10793 7293 10827 7327
rect 12265 7293 12299 7327
rect 12541 7293 12575 7327
rect 13921 7293 13955 7327
rect 15025 7293 15059 7327
rect 15117 7293 15151 7327
rect 17785 7293 17819 7327
rect 18245 7293 18279 7327
rect 18981 7293 19015 7327
rect 19165 7293 19199 7327
rect 20269 7293 20303 7327
rect 20637 7293 20671 7327
rect 1685 7225 1719 7259
rect 5457 7225 5491 7259
rect 14289 7225 14323 7259
rect 16865 7225 16899 7259
rect 1869 7157 1903 7191
rect 3709 7157 3743 7191
rect 7389 7157 7423 7191
rect 11345 7157 11379 7191
rect 13185 7157 13219 7191
rect 14749 7157 14783 7191
rect 15945 7157 15979 7191
rect 16313 7157 16347 7191
rect 17141 7157 17175 7191
rect 19625 7157 19659 7191
rect 8953 6953 8987 6987
rect 13093 6953 13127 6987
rect 14381 6953 14415 6987
rect 20913 6953 20947 6987
rect 2881 6885 2915 6919
rect 7113 6885 7147 6919
rect 16773 6885 16807 6919
rect 18705 6885 18739 6919
rect 2145 6817 2179 6851
rect 2329 6817 2363 6851
rect 3525 6817 3559 6851
rect 3893 6817 3927 6851
rect 5733 6817 5767 6851
rect 7757 6817 7791 6851
rect 8217 6817 8251 6851
rect 8309 6817 8343 6851
rect 9505 6817 9539 6851
rect 10425 6817 10459 6851
rect 10977 6817 11011 6851
rect 11621 6817 11655 6851
rect 13553 6817 13587 6851
rect 13645 6817 13679 6851
rect 14473 6817 14507 6851
rect 16221 6817 16255 6851
rect 17325 6817 17359 6851
rect 17509 6817 17543 6851
rect 18245 6817 18279 6851
rect 21281 6817 21315 6851
rect 1501 6749 1535 6783
rect 1777 6749 1811 6783
rect 3249 6749 3283 6783
rect 3985 6749 4019 6783
rect 4261 6749 4295 6783
rect 4537 6749 4571 6783
rect 5181 6749 5215 6783
rect 5457 6749 5491 6783
rect 5989 6749 6023 6783
rect 7573 6749 7607 6783
rect 9321 6749 9355 6783
rect 10149 6749 10183 6783
rect 11161 6749 11195 6783
rect 13461 6749 13495 6783
rect 14197 6749 14231 6783
rect 18153 6749 18187 6783
rect 18521 6749 18555 6783
rect 19257 6749 19291 6783
rect 19533 6749 19567 6783
rect 21465 6749 21499 6783
rect 1685 6681 1719 6715
rect 3341 6681 3375 6715
rect 10609 6681 10643 6715
rect 11888 6681 11922 6715
rect 14740 6681 14774 6715
rect 16405 6681 16439 6715
rect 18981 6681 19015 6715
rect 19800 6681 19834 6715
rect 21005 6681 21039 6715
rect 1961 6613 1995 6647
rect 2421 6613 2455 6647
rect 2789 6613 2823 6647
rect 4169 6613 4203 6647
rect 5365 6613 5399 6647
rect 5641 6613 5675 6647
rect 7205 6613 7239 6647
rect 7665 6613 7699 6647
rect 8401 6613 8435 6647
rect 8769 6613 8803 6647
rect 9413 6613 9447 6647
rect 9781 6613 9815 6647
rect 10241 6613 10275 6647
rect 11069 6613 11103 6647
rect 11529 6613 11563 6647
rect 13001 6613 13035 6647
rect 15853 6613 15887 6647
rect 16313 6613 16347 6647
rect 16865 6613 16899 6647
rect 17233 6613 17267 6647
rect 17693 6613 17727 6647
rect 18061 6613 18095 6647
rect 18889 6613 18923 6647
rect 19441 6613 19475 6647
rect 1777 6409 1811 6443
rect 2329 6409 2363 6443
rect 2421 6409 2455 6443
rect 2789 6409 2823 6443
rect 3157 6409 3191 6443
rect 4261 6409 4295 6443
rect 5457 6409 5491 6443
rect 6377 6409 6411 6443
rect 6837 6409 6871 6443
rect 7205 6409 7239 6443
rect 8033 6409 8067 6443
rect 8953 6409 8987 6443
rect 9045 6409 9079 6443
rect 9781 6409 9815 6443
rect 10609 6409 10643 6443
rect 11529 6409 11563 6443
rect 13921 6409 13955 6443
rect 15117 6409 15151 6443
rect 17233 6409 17267 6443
rect 19073 6409 19107 6443
rect 20177 6409 20211 6443
rect 20637 6409 20671 6443
rect 1501 6341 1535 6375
rect 3249 6341 3283 6375
rect 5917 6341 5951 6375
rect 11989 6341 12023 6375
rect 12786 6341 12820 6375
rect 14197 6341 14231 6375
rect 14749 6341 14783 6375
rect 19533 6341 19567 6375
rect 3709 6273 3743 6307
rect 4169 6273 4203 6307
rect 4997 6273 5031 6307
rect 5825 6273 5859 6307
rect 6745 6273 6779 6307
rect 7389 6273 7423 6307
rect 7665 6273 7699 6307
rect 8125 6273 8159 6307
rect 10701 6273 10735 6307
rect 11161 6273 11195 6307
rect 11897 6273 11931 6307
rect 12449 6273 12483 6307
rect 12541 6273 12575 6307
rect 15669 6273 15703 6307
rect 16305 6273 16339 6307
rect 16681 6273 16715 6307
rect 17325 6273 17359 6307
rect 17601 6273 17635 6307
rect 18613 6273 18647 6307
rect 19441 6273 19475 6307
rect 20269 6273 20303 6307
rect 21005 6273 21039 6307
rect 1685 6205 1719 6239
rect 2605 6205 2639 6239
rect 3341 6205 3375 6239
rect 4353 6205 4387 6239
rect 5089 6205 5123 6239
rect 5273 6205 5307 6239
rect 6101 6205 6135 6239
rect 7021 6205 7055 6239
rect 7941 6205 7975 6239
rect 9229 6205 9263 6239
rect 9505 6205 9539 6239
rect 9689 6205 9723 6239
rect 10425 6205 10459 6239
rect 12081 6205 12115 6239
rect 14565 6205 14599 6239
rect 14657 6205 14691 6239
rect 15485 6205 15519 6239
rect 15577 6205 15611 6239
rect 18337 6205 18371 6239
rect 18521 6205 18555 6239
rect 19717 6205 19751 6239
rect 19993 6205 20027 6239
rect 20729 6205 20763 6239
rect 3801 6137 3835 6171
rect 14013 6137 14047 6171
rect 16037 6137 16071 6171
rect 18981 6137 19015 6171
rect 1961 6069 1995 6103
rect 4629 6069 4663 6103
rect 8493 6069 8527 6103
rect 8585 6069 8619 6103
rect 10149 6069 10183 6103
rect 11069 6069 11103 6103
rect 11345 6069 11379 6103
rect 16129 6069 16163 6103
rect 16497 6069 16531 6103
rect 16865 6069 16899 6103
rect 2145 5865 2179 5899
rect 4261 5865 4295 5899
rect 6101 5865 6135 5899
rect 6929 5865 6963 5899
rect 10609 5865 10643 5899
rect 10793 5865 10827 5899
rect 15025 5865 15059 5899
rect 17325 5865 17359 5899
rect 20637 5865 20671 5899
rect 20729 5865 20763 5899
rect 3985 5797 4019 5831
rect 14105 5797 14139 5831
rect 18429 5797 18463 5831
rect 18797 5797 18831 5831
rect 1593 5729 1627 5763
rect 1685 5729 1719 5763
rect 6745 5729 6779 5763
rect 7389 5729 7423 5763
rect 7573 5729 7607 5763
rect 7941 5729 7975 5763
rect 9229 5729 9263 5763
rect 11253 5729 11287 5763
rect 11437 5729 11471 5763
rect 11805 5729 11839 5763
rect 12633 5729 12667 5763
rect 14657 5729 14691 5763
rect 15117 5729 15151 5763
rect 16681 5729 16715 5763
rect 16865 5729 16899 5763
rect 18061 5729 18095 5763
rect 19257 5729 19291 5763
rect 21373 5729 21407 5763
rect 3361 5661 3395 5695
rect 3617 5661 3651 5695
rect 3801 5661 3835 5695
rect 5385 5661 5419 5695
rect 5641 5661 5675 5695
rect 5917 5661 5951 5695
rect 6561 5661 6595 5695
rect 8033 5661 8067 5695
rect 8125 5661 8159 5695
rect 8769 5661 8803 5695
rect 9137 5661 9171 5695
rect 11897 5661 11931 5695
rect 13461 5661 13495 5695
rect 13737 5661 13771 5695
rect 14565 5661 14599 5695
rect 15384 5661 15418 5695
rect 17785 5661 17819 5695
rect 18981 5661 19015 5695
rect 21097 5661 21131 5695
rect 7297 5593 7331 5627
rect 9496 5593 9530 5627
rect 11989 5593 12023 5627
rect 16957 5593 16991 5627
rect 18245 5593 18279 5627
rect 18613 5593 18647 5627
rect 19524 5593 19558 5627
rect 1777 5525 1811 5559
rect 2237 5525 2271 5559
rect 5733 5525 5767 5559
rect 6469 5525 6503 5559
rect 8493 5525 8527 5559
rect 8585 5525 8619 5559
rect 8953 5525 8987 5559
rect 11161 5525 11195 5559
rect 12357 5525 12391 5559
rect 12725 5525 12759 5559
rect 12817 5525 12851 5559
rect 13185 5525 13219 5559
rect 13277 5525 13311 5559
rect 13553 5525 13587 5559
rect 13921 5525 13955 5559
rect 14473 5525 14507 5559
rect 16497 5525 16531 5559
rect 17417 5525 17451 5559
rect 17877 5525 17911 5559
rect 21189 5525 21223 5559
rect 1593 5321 1627 5355
rect 3249 5321 3283 5355
rect 6193 5321 6227 5355
rect 8309 5321 8343 5355
rect 10425 5321 10459 5355
rect 10793 5321 10827 5355
rect 11253 5321 11287 5355
rect 11529 5321 11563 5355
rect 12173 5321 12207 5355
rect 14473 5321 14507 5355
rect 15301 5321 15335 5355
rect 15669 5321 15703 5355
rect 16037 5321 16071 5355
rect 16497 5321 16531 5355
rect 16957 5321 16991 5355
rect 17049 5321 17083 5355
rect 17509 5321 17543 5355
rect 17969 5321 18003 5355
rect 19809 5321 19843 5355
rect 20177 5321 20211 5355
rect 1501 5253 1535 5287
rect 7512 5253 7546 5287
rect 9312 5253 9346 5287
rect 10885 5253 10919 5287
rect 13746 5253 13780 5287
rect 16129 5253 16163 5287
rect 2136 5185 2170 5219
rect 3341 5185 3375 5219
rect 4077 5185 4111 5219
rect 4997 5185 5031 5219
rect 5549 5185 5583 5219
rect 6009 5185 6043 5219
rect 7757 5185 7791 5219
rect 8217 5185 8251 5219
rect 8861 5185 8895 5219
rect 9045 5185 9079 5219
rect 11713 5185 11747 5219
rect 14565 5185 14599 5219
rect 17877 5185 17911 5219
rect 18337 5185 18371 5219
rect 18604 5185 18638 5219
rect 20269 5185 20303 5219
rect 20729 5185 20763 5219
rect 1869 5117 1903 5151
rect 4169 5117 4203 5151
rect 4353 5117 4387 5151
rect 4537 5117 4571 5151
rect 5365 5117 5399 5151
rect 5457 5117 5491 5151
rect 8401 5117 8435 5151
rect 10609 5117 10643 5151
rect 11989 5117 12023 5151
rect 12081 5117 12115 5151
rect 14013 5117 14047 5151
rect 14657 5117 14691 5151
rect 15117 5117 15151 5151
rect 15209 5117 15243 5151
rect 15853 5117 15887 5151
rect 16773 5117 16807 5151
rect 18061 5117 18095 5151
rect 20453 5117 20487 5151
rect 21005 5117 21039 5151
rect 3709 5049 3743 5083
rect 17417 5049 17451 5083
rect 19717 5049 19751 5083
rect 3525 4981 3559 5015
rect 4813 4981 4847 5015
rect 5917 4981 5951 5015
rect 6377 4981 6411 5015
rect 7849 4981 7883 5015
rect 8677 4981 8711 5015
rect 12541 4981 12575 5015
rect 12633 4981 12667 5015
rect 14105 4981 14139 5015
rect 2881 4777 2915 4811
rect 4629 4777 4663 4811
rect 10057 4777 10091 4811
rect 13093 4777 13127 4811
rect 17049 4777 17083 4811
rect 19257 4777 19291 4811
rect 20453 4777 20487 4811
rect 21373 4777 21407 4811
rect 6009 4709 6043 4743
rect 7205 4709 7239 4743
rect 8953 4709 8987 4743
rect 11161 4709 11195 4743
rect 12173 4709 12207 4743
rect 15209 4709 15243 4743
rect 17141 4709 17175 4743
rect 3433 4641 3467 4675
rect 4353 4641 4387 4675
rect 5457 4641 5491 4675
rect 6101 4641 6135 4675
rect 7021 4641 7055 4675
rect 7665 4641 7699 4675
rect 7757 4641 7791 4675
rect 8585 4641 8619 4675
rect 9505 4641 9539 4675
rect 10241 4641 10275 4675
rect 10425 4641 10459 4675
rect 11437 4641 11471 4675
rect 11621 4641 11655 4675
rect 12449 4641 12483 4675
rect 12633 4641 12667 4675
rect 13645 4641 13679 4675
rect 13829 4641 13863 4675
rect 19901 4641 19935 4675
rect 20913 4641 20947 4675
rect 21097 4641 21131 4675
rect 2789 4573 2823 4607
rect 3249 4573 3283 4607
rect 4169 4573 4203 4607
rect 4813 4573 4847 4607
rect 5549 4573 5583 4607
rect 6377 4573 6411 4607
rect 10517 4573 10551 4607
rect 10977 4573 11011 4607
rect 13553 4573 13587 4607
rect 14381 4573 14415 4607
rect 14841 4573 14875 4607
rect 15025 4573 15059 4607
rect 15301 4573 15335 4607
rect 15669 4573 15703 4607
rect 15936 4573 15970 4607
rect 17693 4573 17727 4607
rect 20085 4573 20119 4607
rect 20269 4573 20303 4607
rect 21465 4573 21499 4607
rect 2544 4505 2578 4539
rect 4261 4505 4295 4539
rect 4905 4505 4939 4539
rect 5089 4505 5123 4539
rect 8401 4505 8435 4539
rect 9137 4505 9171 4539
rect 9689 4505 9723 4539
rect 17509 4505 17543 4539
rect 17960 4505 17994 4539
rect 19717 4505 19751 4539
rect 20821 4505 20855 4539
rect 1409 4437 1443 4471
rect 3341 4437 3375 4471
rect 3801 4437 3835 4471
rect 5641 4437 5675 4471
rect 7573 4437 7607 4471
rect 8033 4437 8067 4471
rect 8493 4437 8527 4471
rect 9597 4437 9631 4471
rect 10885 4437 10919 4471
rect 11713 4437 11747 4471
rect 12081 4437 12115 4471
rect 12725 4437 12759 4471
rect 13185 4437 13219 4471
rect 14289 4437 14323 4471
rect 14565 4437 14599 4471
rect 14657 4437 14691 4471
rect 15485 4437 15519 4471
rect 17417 4437 17451 4471
rect 19073 4437 19107 4471
rect 19625 4437 19659 4471
rect 3065 4233 3099 4267
rect 3525 4233 3559 4267
rect 4169 4233 4203 4267
rect 5733 4233 5767 4267
rect 9229 4233 9263 4267
rect 9597 4233 9631 4267
rect 11897 4233 11931 4267
rect 12817 4233 12851 4267
rect 13277 4233 13311 4267
rect 13737 4233 13771 4267
rect 14197 4233 14231 4267
rect 14565 4233 14599 4267
rect 15485 4233 15519 4267
rect 18889 4233 18923 4267
rect 19717 4233 19751 4267
rect 19809 4233 19843 4267
rect 20177 4233 20211 4267
rect 2697 4165 2731 4199
rect 4353 4165 4387 4199
rect 12909 4165 12943 4199
rect 13645 4165 13679 4199
rect 19349 4165 19383 4199
rect 1961 4097 1995 4131
rect 2237 4097 2271 4131
rect 2605 4097 2639 4131
rect 3433 4097 3467 4131
rect 4537 4097 4571 4131
rect 4997 4097 5031 4131
rect 5825 4097 5859 4131
rect 6469 4097 6503 4131
rect 6653 4097 6687 4131
rect 7104 4097 7138 4131
rect 8677 4097 8711 4131
rect 10425 4097 10459 4131
rect 10885 4097 10919 4131
rect 11161 4097 11195 4131
rect 15393 4097 15427 4131
rect 15945 4097 15979 4131
rect 16221 4097 16255 4131
rect 16948 4097 16982 4131
rect 18521 4097 18555 4131
rect 20729 4097 20763 4131
rect 2513 4029 2547 4063
rect 3249 4029 3283 4063
rect 5089 4029 5123 4063
rect 5273 4029 5307 4063
rect 5549 4029 5583 4063
rect 6837 4029 6871 4063
rect 8401 4029 8435 4063
rect 8585 4029 8619 4063
rect 9689 4029 9723 4063
rect 9781 4029 9815 4063
rect 10517 4029 10551 4063
rect 10701 4029 10735 4063
rect 11989 4029 12023 4063
rect 12081 4029 12115 4063
rect 12725 4029 12759 4063
rect 13461 4029 13495 4063
rect 14657 4029 14691 4063
rect 14749 4029 14783 4063
rect 15301 4029 15335 4063
rect 16681 4029 16715 4063
rect 18337 4029 18371 4063
rect 18429 4029 18463 4063
rect 19073 4029 19107 4063
rect 19257 4029 19291 4063
rect 20269 4029 20303 4063
rect 20361 4029 20395 4063
rect 21005 4029 21039 4063
rect 3893 3961 3927 3995
rect 6193 3961 6227 3995
rect 8217 3961 8251 3995
rect 10057 3961 10091 3995
rect 11069 3961 11103 3995
rect 16129 3961 16163 3995
rect 18061 3961 18095 3995
rect 4629 3893 4663 3927
rect 9045 3893 9079 3927
rect 11345 3893 11379 3927
rect 11529 3893 11563 3927
rect 12449 3893 12483 3927
rect 14105 3893 14139 3927
rect 15853 3893 15887 3927
rect 16405 3893 16439 3927
rect 5641 3689 5675 3723
rect 7849 3689 7883 3723
rect 8769 3689 8803 3723
rect 11713 3689 11747 3723
rect 13369 3689 13403 3723
rect 15669 3689 15703 3723
rect 18797 3689 18831 3723
rect 19257 3689 19291 3723
rect 11437 3621 11471 3655
rect 17969 3621 18003 3655
rect 21005 3621 21039 3655
rect 1961 3553 1995 3587
rect 4169 3553 4203 3587
rect 4261 3553 4295 3587
rect 5457 3553 5491 3587
rect 6101 3553 6135 3587
rect 6285 3553 6319 3587
rect 6469 3553 6503 3587
rect 8125 3553 8159 3587
rect 8309 3553 8343 3587
rect 9505 3553 9539 3587
rect 11161 3553 11195 3587
rect 11989 3553 12023 3587
rect 14565 3553 14599 3587
rect 14657 3553 14691 3587
rect 15117 3553 15151 3587
rect 16589 3553 16623 3587
rect 18153 3553 18187 3587
rect 18337 3553 18371 3587
rect 19717 3553 19751 3587
rect 19901 3553 19935 3587
rect 2237 3485 2271 3519
rect 2881 3485 2915 3519
rect 3157 3485 3191 3519
rect 3617 3485 3651 3519
rect 6009 3485 6043 3519
rect 11253 3485 11287 3519
rect 13461 3485 13495 3519
rect 13737 3485 13771 3519
rect 14473 3485 14507 3519
rect 15209 3485 15243 3519
rect 15761 3485 15795 3519
rect 16497 3485 16531 3519
rect 16856 3485 16890 3519
rect 19073 3485 19107 3519
rect 20085 3485 20119 3519
rect 20453 3485 20487 3519
rect 20821 3485 20855 3519
rect 21465 3485 21499 3519
rect 3433 3417 3467 3451
rect 4353 3417 4387 3451
rect 6736 3417 6770 3451
rect 10894 3417 10928 3451
rect 11805 3417 11839 3451
rect 12256 3417 12290 3451
rect 15301 3417 15335 3451
rect 16037 3417 16071 3451
rect 3893 3349 3927 3383
rect 4721 3349 4755 3383
rect 4813 3349 4847 3383
rect 5181 3349 5215 3383
rect 5273 3349 5307 3383
rect 8401 3349 8435 3383
rect 8953 3349 8987 3383
rect 9321 3349 9355 3383
rect 9413 3349 9447 3383
rect 9781 3349 9815 3383
rect 13645 3349 13679 3383
rect 13921 3349 13955 3383
rect 14105 3349 14139 3383
rect 15945 3349 15979 3383
rect 16313 3349 16347 3383
rect 18429 3349 18463 3383
rect 18889 3349 18923 3383
rect 19625 3349 19659 3383
rect 20269 3349 20303 3383
rect 20637 3349 20671 3383
rect 21373 3349 21407 3383
rect 6193 3145 6227 3179
rect 7205 3145 7239 3179
rect 7297 3145 7331 3179
rect 9689 3145 9723 3179
rect 9965 3145 9999 3179
rect 14933 3145 14967 3179
rect 16037 3145 16071 3179
rect 16405 3145 16439 3179
rect 18521 3145 18555 3179
rect 18981 3145 19015 3179
rect 19349 3145 19383 3179
rect 19717 3145 19751 3179
rect 2605 3077 2639 3111
rect 2789 3077 2823 3111
rect 4353 3077 4387 3111
rect 9781 3077 9815 3111
rect 11897 3077 11931 3111
rect 12449 3077 12483 3111
rect 12992 3077 13026 3111
rect 18061 3077 18095 3111
rect 20637 3077 20671 3111
rect 2237 3009 2271 3043
rect 4005 3009 4039 3043
rect 4261 3009 4295 3043
rect 4537 3009 4571 3043
rect 4804 3009 4838 3043
rect 6009 3009 6043 3043
rect 6653 3009 6687 3043
rect 8870 3009 8904 3043
rect 9137 3009 9171 3043
rect 9413 3009 9447 3043
rect 11089 3009 11123 3043
rect 12725 3009 12759 3043
rect 14381 3009 14415 3043
rect 14657 3009 14691 3043
rect 14749 3009 14783 3043
rect 15393 3009 15427 3043
rect 15761 3009 15795 3043
rect 15853 3009 15887 3043
rect 16221 3009 16255 3043
rect 16865 3009 16899 3043
rect 16957 3009 16991 3043
rect 17325 3009 17359 3043
rect 18889 3009 18923 3043
rect 20177 3009 20211 3043
rect 20729 3009 20763 3043
rect 1961 2941 1995 2975
rect 7113 2941 7147 2975
rect 11345 2941 11379 2975
rect 11989 2941 12023 2975
rect 12081 2941 12115 2975
rect 17785 2941 17819 2975
rect 17969 2941 18003 2975
rect 19165 2941 19199 2975
rect 19809 2941 19843 2975
rect 19901 2941 19935 2975
rect 21005 2941 21039 2975
rect 2881 2873 2915 2907
rect 7665 2873 7699 2907
rect 15209 2873 15243 2907
rect 15577 2873 15611 2907
rect 18429 2873 18463 2907
rect 2421 2805 2455 2839
rect 5917 2805 5951 2839
rect 6377 2805 6411 2839
rect 6745 2805 6779 2839
rect 7757 2805 7791 2839
rect 9321 2805 9355 2839
rect 11529 2805 11563 2839
rect 12541 2805 12575 2839
rect 14105 2805 14139 2839
rect 14197 2805 14231 2839
rect 14473 2805 14507 2839
rect 16681 2805 16715 2839
rect 17141 2805 17175 2839
rect 17509 2805 17543 2839
rect 20361 2805 20395 2839
rect 3387 2601 3421 2635
rect 9137 2601 9171 2635
rect 12357 2601 12391 2635
rect 13277 2601 13311 2635
rect 18797 2601 18831 2635
rect 19717 2601 19751 2635
rect 5181 2533 5215 2567
rect 10241 2533 10275 2567
rect 12265 2533 12299 2567
rect 13645 2533 13679 2567
rect 14565 2533 14599 2567
rect 15301 2533 15335 2567
rect 16773 2533 16807 2567
rect 17509 2533 17543 2567
rect 17785 2533 17819 2567
rect 2697 2465 2731 2499
rect 3617 2465 3651 2499
rect 5825 2465 5859 2499
rect 6929 2465 6963 2499
rect 9965 2465 9999 2499
rect 10793 2465 10827 2499
rect 11621 2465 11655 2499
rect 11805 2465 11839 2499
rect 12909 2465 12943 2499
rect 18199 2465 18233 2499
rect 18337 2465 18371 2499
rect 1777 2397 1811 2431
rect 2421 2397 2455 2431
rect 3801 2397 3835 2431
rect 4057 2397 4091 2431
rect 6101 2397 6135 2431
rect 7205 2397 7239 2431
rect 7941 2397 7975 2431
rect 8217 2397 8251 2431
rect 8677 2397 8711 2431
rect 9321 2397 9355 2431
rect 10609 2397 10643 2431
rect 10701 2397 10735 2431
rect 11253 2397 11287 2431
rect 11897 2397 11931 2431
rect 13461 2397 13495 2431
rect 13829 2397 13863 2431
rect 14105 2397 14139 2431
rect 14749 2397 14783 2431
rect 14841 2397 14875 2431
rect 15485 2397 15519 2431
rect 15853 2397 15887 2431
rect 15945 2397 15979 2431
rect 16497 2397 16531 2431
rect 16957 2397 16991 2431
rect 17325 2397 17359 2431
rect 17693 2397 17727 2431
rect 17969 2397 18003 2431
rect 18429 2397 18463 2431
rect 19073 2397 19107 2431
rect 19257 2397 19291 2431
rect 20361 2397 20395 2431
rect 20637 2397 20671 2431
rect 20729 2397 20763 2431
rect 21005 2397 21039 2431
rect 9873 2329 9907 2363
rect 11069 2329 11103 2363
rect 12817 2329 12851 2363
rect 1593 2261 1627 2295
rect 8309 2261 8343 2295
rect 8585 2261 8619 2295
rect 9413 2261 9447 2295
rect 9781 2261 9815 2295
rect 12725 2261 12759 2295
rect 14289 2261 14323 2295
rect 15025 2261 15059 2295
rect 15669 2261 15703 2295
rect 16129 2261 16163 2295
rect 16313 2261 16347 2295
rect 17141 2261 17175 2295
rect 18889 2261 18923 2295
rect 19441 2261 19475 2295
<< metal1 >>
rect 842 22040 848 22092
rect 900 22080 906 22092
rect 1026 22080 1032 22092
rect 900 22052 1032 22080
rect 900 22040 906 22052
rect 1026 22040 1032 22052
rect 1084 22040 1090 22092
rect 14 21632 20 21684
rect 72 21672 78 21684
rect 14274 21672 14280 21684
rect 72 21644 14280 21672
rect 72 21632 78 21644
rect 14274 21632 14280 21644
rect 14332 21632 14338 21684
rect 7558 21564 7564 21616
rect 7616 21604 7622 21616
rect 16206 21604 16212 21616
rect 7616 21576 16212 21604
rect 7616 21564 7622 21576
rect 16206 21564 16212 21576
rect 16264 21564 16270 21616
rect 1394 21496 1400 21548
rect 1452 21536 1458 21548
rect 2498 21536 2504 21548
rect 1452 21508 2504 21536
rect 1452 21496 1458 21508
rect 2498 21496 2504 21508
rect 2556 21496 2562 21548
rect 4706 21496 4712 21548
rect 4764 21536 4770 21548
rect 15654 21536 15660 21548
rect 4764 21508 15660 21536
rect 4764 21496 4770 21508
rect 15654 21496 15660 21508
rect 15712 21496 15718 21548
rect 2590 21428 2596 21480
rect 2648 21468 2654 21480
rect 16114 21468 16120 21480
rect 2648 21440 16120 21468
rect 2648 21428 2654 21440
rect 16114 21428 16120 21440
rect 16172 21428 16178 21480
rect 4798 21360 4804 21412
rect 4856 21400 4862 21412
rect 5074 21400 5080 21412
rect 4856 21372 5080 21400
rect 4856 21360 4862 21372
rect 5074 21360 5080 21372
rect 5132 21400 5138 21412
rect 12894 21400 12900 21412
rect 5132 21372 12900 21400
rect 5132 21360 5138 21372
rect 12894 21360 12900 21372
rect 12952 21360 12958 21412
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 17862 21332 17868 21344
rect 2832 21304 17868 21332
rect 2832 21292 2838 21304
rect 17862 21292 17868 21304
rect 17920 21292 17926 21344
rect 4062 21224 4068 21276
rect 4120 21264 4126 21276
rect 12158 21264 12164 21276
rect 4120 21236 12164 21264
rect 4120 21224 4126 21236
rect 12158 21224 12164 21236
rect 12216 21224 12222 21276
rect 3602 21156 3608 21208
rect 3660 21196 3666 21208
rect 13262 21196 13268 21208
rect 3660 21168 13268 21196
rect 3660 21156 3666 21168
rect 13262 21156 13268 21168
rect 13320 21156 13326 21208
rect 4430 21088 4436 21140
rect 4488 21128 4494 21140
rect 16022 21128 16028 21140
rect 4488 21100 16028 21128
rect 4488 21088 4494 21100
rect 16022 21088 16028 21100
rect 16080 21088 16086 21140
rect 2682 21020 2688 21072
rect 2740 21060 2746 21072
rect 7558 21060 7564 21072
rect 2740 21032 7564 21060
rect 2740 21020 2746 21032
rect 7558 21020 7564 21032
rect 7616 21020 7622 21072
rect 13078 21060 13084 21072
rect 12406 21032 13084 21060
rect 3326 20952 3332 21004
rect 3384 20992 3390 21004
rect 12406 20992 12434 21032
rect 13078 21020 13084 21032
rect 13136 21020 13142 21072
rect 3384 20964 12434 20992
rect 3384 20952 3390 20964
rect 3142 20884 3148 20936
rect 3200 20924 3206 20936
rect 11974 20924 11980 20936
rect 3200 20896 11980 20924
rect 3200 20884 3206 20896
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 12158 20884 12164 20936
rect 12216 20924 12222 20936
rect 14918 20924 14924 20936
rect 12216 20896 14924 20924
rect 12216 20884 12222 20896
rect 14918 20884 14924 20896
rect 14976 20884 14982 20936
rect 8202 20816 8208 20868
rect 8260 20856 8266 20868
rect 12986 20856 12992 20868
rect 8260 20828 12992 20856
rect 8260 20816 8266 20828
rect 12986 20816 12992 20828
rect 13044 20816 13050 20868
rect 934 20748 940 20800
rect 992 20788 998 20800
rect 3050 20788 3056 20800
rect 992 20760 3056 20788
rect 992 20748 998 20760
rect 3050 20748 3056 20760
rect 3108 20748 3114 20800
rect 4246 20748 4252 20800
rect 4304 20788 4310 20800
rect 10686 20788 10692 20800
rect 4304 20760 10692 20788
rect 4304 20748 4310 20760
rect 10686 20748 10692 20760
rect 10744 20748 10750 20800
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 5166 20584 5172 20596
rect 2516 20556 5172 20584
rect 2516 20525 2544 20556
rect 5166 20544 5172 20556
rect 5224 20544 5230 20596
rect 5721 20587 5779 20593
rect 5721 20553 5733 20587
rect 5767 20584 5779 20587
rect 6641 20587 6699 20593
rect 6641 20584 6653 20587
rect 5767 20556 6653 20584
rect 5767 20553 5779 20556
rect 5721 20547 5779 20553
rect 6641 20553 6653 20556
rect 6687 20553 6699 20587
rect 6641 20547 6699 20553
rect 6914 20544 6920 20596
rect 6972 20584 6978 20596
rect 7374 20584 7380 20596
rect 6972 20556 7380 20584
rect 6972 20544 6978 20556
rect 7374 20544 7380 20556
rect 7432 20584 7438 20596
rect 8202 20584 8208 20596
rect 7432 20556 8208 20584
rect 7432 20544 7438 20556
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 8297 20587 8355 20593
rect 8297 20553 8309 20587
rect 8343 20584 8355 20587
rect 8662 20584 8668 20596
rect 8343 20556 8668 20584
rect 8343 20553 8355 20556
rect 8297 20547 8355 20553
rect 8662 20544 8668 20556
rect 8720 20544 8726 20596
rect 9306 20544 9312 20596
rect 9364 20584 9370 20596
rect 10321 20587 10379 20593
rect 9364 20556 9996 20584
rect 9364 20544 9370 20556
rect 2501 20519 2559 20525
rect 2501 20485 2513 20519
rect 2547 20485 2559 20519
rect 2501 20479 2559 20485
rect 4157 20519 4215 20525
rect 4157 20485 4169 20519
rect 4203 20516 4215 20519
rect 5994 20516 6000 20528
rect 4203 20488 6000 20516
rect 4203 20485 4215 20488
rect 4157 20479 4215 20485
rect 5994 20476 6000 20488
rect 6052 20476 6058 20528
rect 9490 20516 9496 20528
rect 6196 20488 9496 20516
rect 1302 20408 1308 20460
rect 1360 20448 1366 20460
rect 2225 20451 2283 20457
rect 2225 20448 2237 20451
rect 1360 20420 2237 20448
rect 1360 20408 1366 20420
rect 2225 20417 2237 20420
rect 2271 20417 2283 20451
rect 3326 20448 3332 20460
rect 3287 20420 3332 20448
rect 2225 20411 2283 20417
rect 3326 20408 3332 20420
rect 3384 20408 3390 20460
rect 3602 20448 3608 20460
rect 3563 20420 3608 20448
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20448 3847 20451
rect 3835 20420 5396 20448
rect 3835 20417 3847 20420
rect 3789 20411 3847 20417
rect 1946 20380 1952 20392
rect 1907 20352 1952 20380
rect 1946 20340 1952 20352
rect 2004 20340 2010 20392
rect 2685 20383 2743 20389
rect 2685 20349 2697 20383
rect 2731 20380 2743 20383
rect 4614 20380 4620 20392
rect 2731 20352 4620 20380
rect 2731 20349 2743 20352
rect 2685 20343 2743 20349
rect 4614 20340 4620 20352
rect 4672 20340 4678 20392
rect 4982 20380 4988 20392
rect 4943 20352 4988 20380
rect 4982 20340 4988 20352
rect 5040 20340 5046 20392
rect 5261 20383 5319 20389
rect 5261 20349 5273 20383
rect 5307 20349 5319 20383
rect 5261 20343 5319 20349
rect 4338 20272 4344 20324
rect 4396 20312 4402 20324
rect 5276 20312 5304 20343
rect 4396 20284 5304 20312
rect 5368 20312 5396 20420
rect 5626 20408 5632 20460
rect 5684 20448 5690 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5684 20420 5825 20448
rect 5684 20408 5690 20420
rect 5813 20417 5825 20420
rect 5859 20417 5871 20451
rect 5813 20411 5871 20417
rect 5534 20380 5540 20392
rect 5495 20352 5540 20380
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 5810 20312 5816 20324
rect 5368 20284 5816 20312
rect 4396 20272 4402 20284
rect 3878 20204 3884 20256
rect 3936 20244 3942 20256
rect 3973 20247 4031 20253
rect 3973 20244 3985 20247
rect 3936 20216 3985 20244
rect 3936 20204 3942 20216
rect 3973 20213 3985 20216
rect 4019 20213 4031 20247
rect 3973 20207 4031 20213
rect 4249 20247 4307 20253
rect 4249 20213 4261 20247
rect 4295 20244 4307 20247
rect 4890 20244 4896 20256
rect 4295 20216 4896 20244
rect 4295 20213 4307 20216
rect 4249 20207 4307 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 5276 20244 5304 20284
rect 5810 20272 5816 20284
rect 5868 20272 5874 20324
rect 6196 20321 6224 20488
rect 9490 20476 9496 20488
rect 9548 20476 9554 20528
rect 6365 20451 6423 20457
rect 6365 20417 6377 20451
rect 6411 20448 6423 20451
rect 6822 20448 6828 20460
rect 6411 20420 6828 20448
rect 6411 20417 6423 20420
rect 6365 20411 6423 20417
rect 6822 20408 6828 20420
rect 6880 20408 6886 20460
rect 7009 20451 7067 20457
rect 7009 20417 7021 20451
rect 7055 20448 7067 20451
rect 7466 20448 7472 20460
rect 7055 20420 7472 20448
rect 7055 20417 7067 20420
rect 7009 20411 7067 20417
rect 7466 20408 7472 20420
rect 7524 20408 7530 20460
rect 7653 20451 7711 20457
rect 7653 20417 7665 20451
rect 7699 20417 7711 20451
rect 7653 20411 7711 20417
rect 6914 20340 6920 20392
rect 6972 20380 6978 20392
rect 7101 20383 7159 20389
rect 7101 20380 7113 20383
rect 6972 20352 7113 20380
rect 6972 20340 6978 20352
rect 7101 20349 7113 20352
rect 7147 20349 7159 20383
rect 7101 20343 7159 20349
rect 7193 20383 7251 20389
rect 7193 20349 7205 20383
rect 7239 20349 7251 20383
rect 7668 20380 7696 20411
rect 7834 20408 7840 20460
rect 7892 20448 7898 20460
rect 7929 20451 7987 20457
rect 7929 20448 7941 20451
rect 7892 20420 7941 20448
rect 7892 20408 7898 20420
rect 7929 20417 7941 20420
rect 7975 20417 7987 20451
rect 8202 20448 8208 20460
rect 8163 20420 8208 20448
rect 7929 20411 7987 20417
rect 8202 20408 8208 20420
rect 8260 20408 8266 20460
rect 8478 20408 8484 20460
rect 8536 20448 8542 20460
rect 8665 20451 8723 20457
rect 8665 20448 8677 20451
rect 8536 20420 8677 20448
rect 8536 20408 8542 20420
rect 8665 20417 8677 20420
rect 8711 20417 8723 20451
rect 8665 20411 8723 20417
rect 8938 20408 8944 20460
rect 8996 20448 9002 20460
rect 9674 20448 9680 20460
rect 8996 20420 9680 20448
rect 8996 20408 9002 20420
rect 9674 20408 9680 20420
rect 9732 20448 9738 20460
rect 9968 20448 9996 20556
rect 10321 20553 10333 20587
rect 10367 20584 10379 20587
rect 10870 20584 10876 20596
rect 10367 20556 10876 20584
rect 10367 20553 10379 20556
rect 10321 20547 10379 20553
rect 10870 20544 10876 20556
rect 10928 20544 10934 20596
rect 11701 20587 11759 20593
rect 11701 20553 11713 20587
rect 11747 20553 11759 20587
rect 11701 20547 11759 20553
rect 10045 20519 10103 20525
rect 10045 20485 10057 20519
rect 10091 20516 10103 20519
rect 10091 20488 10548 20516
rect 10091 20485 10103 20488
rect 10045 20479 10103 20485
rect 10520 20460 10548 20488
rect 10137 20451 10195 20457
rect 10137 20448 10149 20451
rect 9732 20420 9904 20448
rect 9968 20420 10149 20448
rect 9732 20408 9738 20420
rect 8018 20380 8024 20392
rect 7668 20352 8024 20380
rect 7193 20343 7251 20349
rect 6181 20315 6239 20321
rect 6181 20281 6193 20315
rect 6227 20281 6239 20315
rect 6181 20275 6239 20281
rect 6730 20272 6736 20324
rect 6788 20312 6794 20324
rect 7208 20312 7236 20343
rect 8018 20340 8024 20352
rect 8076 20340 8082 20392
rect 9122 20340 9128 20392
rect 9180 20380 9186 20392
rect 9876 20389 9904 20420
rect 10137 20417 10149 20420
rect 10183 20417 10195 20451
rect 10502 20448 10508 20460
rect 10463 20420 10508 20448
rect 10137 20411 10195 20417
rect 10502 20408 10508 20420
rect 10560 20408 10566 20460
rect 10686 20408 10692 20460
rect 10744 20448 10750 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 10744 20420 11529 20448
rect 10744 20408 10750 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 11716 20448 11744 20547
rect 11790 20544 11796 20596
rect 11848 20584 11854 20596
rect 11977 20587 12035 20593
rect 11977 20584 11989 20587
rect 11848 20556 11989 20584
rect 11848 20544 11854 20556
rect 11977 20553 11989 20556
rect 12023 20553 12035 20587
rect 11977 20547 12035 20553
rect 12066 20544 12072 20596
rect 12124 20584 12130 20596
rect 12345 20587 12403 20593
rect 12345 20584 12357 20587
rect 12124 20556 12357 20584
rect 12124 20544 12130 20556
rect 12345 20553 12357 20556
rect 12391 20553 12403 20587
rect 12345 20547 12403 20553
rect 12434 20544 12440 20596
rect 12492 20584 12498 20596
rect 12713 20587 12771 20593
rect 12713 20584 12725 20587
rect 12492 20556 12725 20584
rect 12492 20544 12498 20556
rect 12713 20553 12725 20556
rect 12759 20553 12771 20587
rect 12713 20547 12771 20553
rect 12802 20544 12808 20596
rect 12860 20584 12866 20596
rect 13081 20587 13139 20593
rect 13081 20584 13093 20587
rect 12860 20556 13093 20584
rect 12860 20544 12866 20556
rect 13081 20553 13093 20556
rect 13127 20553 13139 20587
rect 13081 20547 13139 20553
rect 13170 20544 13176 20596
rect 13228 20584 13234 20596
rect 13449 20587 13507 20593
rect 13449 20584 13461 20587
rect 13228 20556 13461 20584
rect 13228 20544 13234 20556
rect 13449 20553 13461 20556
rect 13495 20553 13507 20587
rect 13449 20547 13507 20553
rect 13538 20544 13544 20596
rect 13596 20584 13602 20596
rect 13817 20587 13875 20593
rect 13817 20584 13829 20587
rect 13596 20556 13829 20584
rect 13596 20544 13602 20556
rect 13817 20553 13829 20556
rect 13863 20553 13875 20587
rect 13817 20547 13875 20553
rect 13998 20544 14004 20596
rect 14056 20584 14062 20596
rect 14277 20587 14335 20593
rect 14277 20584 14289 20587
rect 14056 20556 14289 20584
rect 14056 20544 14062 20556
rect 14277 20553 14289 20556
rect 14323 20553 14335 20587
rect 14277 20547 14335 20553
rect 14366 20544 14372 20596
rect 14424 20584 14430 20596
rect 14645 20587 14703 20593
rect 14645 20584 14657 20587
rect 14424 20556 14657 20584
rect 14424 20544 14430 20556
rect 14645 20553 14657 20556
rect 14691 20553 14703 20587
rect 14645 20547 14703 20553
rect 14734 20544 14740 20596
rect 14792 20584 14798 20596
rect 15013 20587 15071 20593
rect 15013 20584 15025 20587
rect 14792 20556 15025 20584
rect 14792 20544 14798 20556
rect 15013 20553 15025 20556
rect 15059 20553 15071 20587
rect 15013 20547 15071 20553
rect 15194 20544 15200 20596
rect 15252 20584 15258 20596
rect 15381 20587 15439 20593
rect 15381 20584 15393 20587
rect 15252 20556 15393 20584
rect 15252 20544 15258 20556
rect 15381 20553 15393 20556
rect 15427 20553 15439 20587
rect 15381 20547 15439 20553
rect 15470 20544 15476 20596
rect 15528 20584 15534 20596
rect 15749 20587 15807 20593
rect 15749 20584 15761 20587
rect 15528 20556 15761 20584
rect 15528 20544 15534 20556
rect 15749 20553 15761 20556
rect 15795 20553 15807 20587
rect 15749 20547 15807 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16117 20587 16175 20593
rect 16117 20584 16129 20587
rect 15896 20556 16129 20584
rect 15896 20544 15902 20556
rect 16117 20553 16129 20556
rect 16163 20553 16175 20587
rect 16117 20547 16175 20553
rect 16485 20587 16543 20593
rect 16485 20553 16497 20587
rect 16531 20584 16543 20587
rect 17954 20584 17960 20596
rect 16531 20556 17960 20584
rect 16531 20553 16543 20556
rect 16485 20547 16543 20553
rect 17954 20544 17960 20556
rect 18012 20544 18018 20596
rect 18138 20544 18144 20596
rect 18196 20584 18202 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 18196 20556 19441 20584
rect 18196 20544 18202 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 19518 20544 19524 20596
rect 19576 20584 19582 20596
rect 19705 20587 19763 20593
rect 19705 20584 19717 20587
rect 19576 20556 19717 20584
rect 19576 20544 19582 20556
rect 19705 20553 19717 20556
rect 19751 20553 19763 20587
rect 19705 20547 19763 20553
rect 19794 20544 19800 20596
rect 19852 20544 19858 20596
rect 19978 20544 19984 20596
rect 20036 20544 20042 20596
rect 20165 20587 20223 20593
rect 20165 20553 20177 20587
rect 20211 20553 20223 20587
rect 20530 20584 20536 20596
rect 20491 20556 20536 20584
rect 20165 20547 20223 20553
rect 17494 20516 17500 20528
rect 17052 20488 17500 20516
rect 11793 20451 11851 20457
rect 11793 20448 11805 20451
rect 11716 20420 11805 20448
rect 11517 20411 11575 20417
rect 11793 20417 11805 20420
rect 11839 20417 11851 20451
rect 11793 20411 11851 20417
rect 11882 20408 11888 20460
rect 11940 20448 11946 20460
rect 12161 20451 12219 20457
rect 12161 20448 12173 20451
rect 11940 20420 12173 20448
rect 11940 20408 11946 20420
rect 12161 20417 12173 20420
rect 12207 20417 12219 20451
rect 12529 20451 12587 20457
rect 12529 20448 12541 20451
rect 12161 20411 12219 20417
rect 12406 20420 12541 20448
rect 9585 20383 9643 20389
rect 9585 20380 9597 20383
rect 9180 20352 9597 20380
rect 9180 20340 9186 20352
rect 9585 20349 9597 20352
rect 9631 20349 9643 20383
rect 9585 20343 9643 20349
rect 9861 20383 9919 20389
rect 9861 20349 9873 20383
rect 9907 20349 9919 20383
rect 10778 20380 10784 20392
rect 10739 20352 10784 20380
rect 9861 20343 9919 20349
rect 10778 20340 10784 20352
rect 10836 20340 10842 20392
rect 10870 20340 10876 20392
rect 10928 20380 10934 20392
rect 12406 20380 12434 20420
rect 12529 20417 12541 20420
rect 12575 20417 12587 20451
rect 12529 20411 12587 20417
rect 12802 20408 12808 20460
rect 12860 20448 12866 20460
rect 12897 20451 12955 20457
rect 12897 20448 12909 20451
rect 12860 20420 12909 20448
rect 12860 20408 12866 20420
rect 12897 20417 12909 20420
rect 12943 20417 12955 20451
rect 12897 20411 12955 20417
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 13228 20420 13277 20448
rect 13228 20408 13234 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20448 13691 20451
rect 13722 20448 13728 20460
rect 13679 20420 13728 20448
rect 13679 20417 13691 20420
rect 13633 20411 13691 20417
rect 13722 20408 13728 20420
rect 13780 20408 13786 20460
rect 14093 20451 14151 20457
rect 14093 20417 14105 20451
rect 14139 20417 14151 20451
rect 14458 20448 14464 20460
rect 14419 20420 14464 20448
rect 14093 20411 14151 20417
rect 10928 20352 12434 20380
rect 10928 20340 10934 20352
rect 13446 20340 13452 20392
rect 13504 20380 13510 20392
rect 14108 20380 14136 20411
rect 14458 20408 14464 20420
rect 14516 20408 14522 20460
rect 14642 20408 14648 20460
rect 14700 20448 14706 20460
rect 14829 20451 14887 20457
rect 14829 20448 14841 20451
rect 14700 20420 14841 20448
rect 14700 20408 14706 20420
rect 14829 20417 14841 20420
rect 14875 20417 14887 20451
rect 14829 20411 14887 20417
rect 15010 20408 15016 20460
rect 15068 20448 15074 20460
rect 15197 20451 15255 20457
rect 15197 20448 15209 20451
rect 15068 20420 15209 20448
rect 15068 20408 15074 20420
rect 15197 20417 15209 20420
rect 15243 20417 15255 20451
rect 15562 20448 15568 20460
rect 15523 20420 15568 20448
rect 15197 20411 15255 20417
rect 15562 20408 15568 20420
rect 15620 20408 15626 20460
rect 15930 20448 15936 20460
rect 15891 20420 15936 20448
rect 15930 20408 15936 20420
rect 15988 20408 15994 20460
rect 16301 20451 16359 20457
rect 16301 20417 16313 20451
rect 16347 20417 16359 20451
rect 16666 20448 16672 20460
rect 16627 20420 16672 20448
rect 16301 20411 16359 20417
rect 13504 20352 14136 20380
rect 16316 20380 16344 20411
rect 16666 20408 16672 20420
rect 16724 20408 16730 20460
rect 17052 20457 17080 20488
rect 17494 20476 17500 20488
rect 17552 20516 17558 20528
rect 18966 20516 18972 20528
rect 17552 20488 18972 20516
rect 17552 20476 17558 20488
rect 18966 20476 18972 20488
rect 19024 20476 19030 20528
rect 19061 20519 19119 20525
rect 19061 20485 19073 20519
rect 19107 20516 19119 20519
rect 19812 20516 19840 20544
rect 19107 20488 19840 20516
rect 19107 20485 19119 20488
rect 19061 20479 19119 20485
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17126 20408 17132 20460
rect 17184 20448 17190 20460
rect 19245 20451 19303 20457
rect 19245 20448 19257 20451
rect 17184 20420 19257 20448
rect 17184 20408 17190 20420
rect 19245 20417 19257 20420
rect 19291 20417 19303 20451
rect 19245 20411 19303 20417
rect 19518 20408 19524 20460
rect 19576 20408 19582 20460
rect 19996 20457 20024 20544
rect 20180 20516 20208 20547
rect 20530 20544 20536 20556
rect 20588 20544 20594 20596
rect 20898 20544 20904 20596
rect 20956 20584 20962 20596
rect 21085 20587 21143 20593
rect 21085 20584 21097 20587
rect 20956 20556 21097 20584
rect 20956 20544 20962 20556
rect 21085 20553 21097 20556
rect 21131 20553 21143 20587
rect 21085 20547 21143 20553
rect 21634 20516 21640 20528
rect 20180 20488 21640 20516
rect 21634 20476 21640 20488
rect 21692 20476 21698 20528
rect 19864 20451 19922 20457
rect 19864 20448 19876 20451
rect 19720 20420 19876 20448
rect 19426 20380 19432 20392
rect 16316 20352 19432 20380
rect 13504 20340 13510 20352
rect 19426 20340 19432 20352
rect 19484 20340 19490 20392
rect 6788 20284 7236 20312
rect 7745 20315 7803 20321
rect 6788 20272 6794 20284
rect 7745 20281 7757 20315
rect 7791 20312 7803 20315
rect 12618 20312 12624 20324
rect 7791 20284 8156 20312
rect 7791 20281 7803 20284
rect 7745 20275 7803 20281
rect 5350 20244 5356 20256
rect 5276 20216 5356 20244
rect 5350 20204 5356 20216
rect 5408 20204 5414 20256
rect 6454 20204 6460 20256
rect 6512 20244 6518 20256
rect 6549 20247 6607 20253
rect 6549 20244 6561 20247
rect 6512 20216 6561 20244
rect 6512 20204 6518 20216
rect 6549 20213 6561 20216
rect 6595 20213 6607 20247
rect 6549 20207 6607 20213
rect 6822 20204 6828 20256
rect 6880 20244 6886 20256
rect 7006 20244 7012 20256
rect 6880 20216 7012 20244
rect 6880 20204 6886 20216
rect 7006 20204 7012 20216
rect 7064 20244 7070 20256
rect 7374 20244 7380 20256
rect 7064 20216 7380 20244
rect 7064 20204 7070 20216
rect 7374 20204 7380 20216
rect 7432 20244 7438 20256
rect 7469 20247 7527 20253
rect 7469 20244 7481 20247
rect 7432 20216 7481 20244
rect 7432 20204 7438 20216
rect 7469 20213 7481 20216
rect 7515 20213 7527 20247
rect 8128 20244 8156 20284
rect 8404 20284 12624 20312
rect 8404 20244 8432 20284
rect 12618 20272 12624 20284
rect 12676 20272 12682 20324
rect 16574 20272 16580 20324
rect 16632 20312 16638 20324
rect 16853 20315 16911 20321
rect 16853 20312 16865 20315
rect 16632 20284 16865 20312
rect 16632 20272 16638 20284
rect 16853 20281 16865 20284
rect 16899 20281 16911 20315
rect 16853 20275 16911 20281
rect 18598 20272 18604 20324
rect 18656 20312 18662 20324
rect 19536 20312 19564 20408
rect 18656 20284 19564 20312
rect 18656 20272 18662 20284
rect 8570 20244 8576 20256
rect 8128 20216 8432 20244
rect 8531 20216 8576 20244
rect 7469 20207 7527 20213
rect 8570 20204 8576 20216
rect 8628 20204 8634 20256
rect 9398 20204 9404 20256
rect 9456 20244 9462 20256
rect 10502 20244 10508 20256
rect 9456 20216 10508 20244
rect 9456 20204 9462 20216
rect 10502 20204 10508 20216
rect 10560 20204 10566 20256
rect 10686 20204 10692 20256
rect 10744 20244 10750 20256
rect 12250 20244 12256 20256
rect 10744 20216 12256 20244
rect 10744 20204 10750 20216
rect 12250 20204 12256 20216
rect 12308 20204 12314 20256
rect 16022 20204 16028 20256
rect 16080 20244 16086 20256
rect 16390 20244 16396 20256
rect 16080 20216 16396 20244
rect 16080 20204 16086 20216
rect 16390 20204 16396 20216
rect 16448 20204 16454 20256
rect 17218 20244 17224 20256
rect 17179 20216 17224 20244
rect 17218 20204 17224 20216
rect 17276 20204 17282 20256
rect 17773 20247 17831 20253
rect 17773 20213 17785 20247
rect 17819 20244 17831 20247
rect 19610 20244 19616 20256
rect 17819 20216 19616 20244
rect 17819 20213 17831 20216
rect 17773 20207 17831 20213
rect 19610 20204 19616 20216
rect 19668 20204 19674 20256
rect 19720 20244 19748 20420
rect 19864 20417 19876 20420
rect 19910 20417 19922 20451
rect 19864 20411 19922 20417
rect 19969 20451 20027 20457
rect 19969 20417 19981 20451
rect 20015 20417 20027 20451
rect 20346 20448 20352 20460
rect 20307 20420 20352 20448
rect 19969 20411 20027 20417
rect 20346 20408 20352 20420
rect 20404 20408 20410 20460
rect 20717 20451 20775 20457
rect 20717 20417 20729 20451
rect 20763 20417 20775 20451
rect 20717 20411 20775 20417
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20448 21327 20451
rect 21358 20448 21364 20460
rect 21315 20420 21364 20448
rect 21315 20417 21327 20420
rect 21269 20411 21327 20417
rect 20162 20272 20168 20324
rect 20220 20312 20226 20324
rect 20732 20312 20760 20411
rect 21358 20408 21364 20420
rect 21416 20408 21422 20460
rect 20220 20284 20760 20312
rect 20901 20315 20959 20321
rect 20220 20272 20226 20284
rect 20901 20281 20913 20315
rect 20947 20312 20959 20315
rect 20990 20312 20996 20324
rect 20947 20284 20996 20312
rect 20947 20281 20959 20284
rect 20901 20275 20959 20281
rect 20990 20272 20996 20284
rect 21048 20272 21054 20324
rect 21082 20244 21088 20256
rect 19720 20216 21088 20244
rect 21082 20204 21088 20216
rect 21140 20204 21146 20256
rect 21450 20244 21456 20256
rect 21411 20216 21456 20244
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 1578 20000 1584 20052
rect 1636 20040 1642 20052
rect 1857 20043 1915 20049
rect 1857 20040 1869 20043
rect 1636 20012 1869 20040
rect 1636 20000 1642 20012
rect 1857 20009 1869 20012
rect 1903 20009 1915 20043
rect 1857 20003 1915 20009
rect 3344 20012 7052 20040
rect 2682 19972 2688 19984
rect 2643 19944 2688 19972
rect 2682 19932 2688 19944
rect 2740 19932 2746 19984
rect 3344 19913 3372 20012
rect 3602 19932 3608 19984
rect 3660 19932 3666 19984
rect 3786 19932 3792 19984
rect 3844 19972 3850 19984
rect 3970 19972 3976 19984
rect 3844 19944 3976 19972
rect 3844 19932 3850 19944
rect 3970 19932 3976 19944
rect 4028 19932 4034 19984
rect 3329 19907 3387 19913
rect 1688 19876 2774 19904
rect 1486 19796 1492 19848
rect 1544 19796 1550 19848
rect 1688 19845 1716 19876
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19805 1731 19839
rect 2038 19836 2044 19848
rect 1999 19808 2044 19836
rect 1673 19799 1731 19805
rect 2038 19796 2044 19808
rect 2096 19796 2102 19848
rect 2317 19839 2375 19845
rect 2317 19805 2329 19839
rect 2363 19805 2375 19839
rect 2317 19799 2375 19805
rect 1504 19768 1532 19796
rect 2332 19768 2360 19799
rect 1504 19740 2360 19768
rect 2501 19771 2559 19777
rect 2501 19737 2513 19771
rect 2547 19737 2559 19771
rect 2746 19768 2774 19876
rect 3329 19873 3341 19907
rect 3375 19873 3387 19907
rect 3620 19904 3648 19932
rect 4062 19904 4068 19916
rect 3620 19876 4068 19904
rect 3329 19867 3387 19873
rect 4062 19864 4068 19876
rect 4120 19864 4126 19916
rect 5534 19904 5540 19916
rect 5184 19876 5540 19904
rect 3234 19796 3240 19848
rect 3292 19836 3298 19848
rect 3605 19839 3663 19845
rect 3605 19836 3617 19839
rect 3292 19808 3617 19836
rect 3292 19796 3298 19808
rect 3605 19805 3617 19808
rect 3651 19836 3663 19839
rect 3694 19836 3700 19848
rect 3651 19808 3700 19836
rect 3651 19805 3663 19808
rect 3605 19799 3663 19805
rect 3694 19796 3700 19808
rect 3752 19796 3758 19848
rect 5005 19839 5063 19845
rect 5005 19805 5017 19839
rect 5051 19836 5063 19839
rect 5184 19836 5212 19876
rect 5534 19864 5540 19876
rect 5592 19904 5598 19916
rect 6822 19904 6828 19916
rect 5592 19876 5672 19904
rect 6783 19876 6828 19904
rect 5592 19864 5598 19876
rect 5051 19808 5212 19836
rect 5261 19839 5319 19845
rect 5051 19805 5063 19808
rect 5005 19799 5063 19805
rect 5261 19805 5273 19839
rect 5307 19836 5319 19839
rect 5442 19836 5448 19848
rect 5307 19808 5448 19836
rect 5307 19805 5319 19808
rect 5261 19799 5319 19805
rect 5442 19796 5448 19808
rect 5500 19796 5506 19848
rect 5534 19768 5540 19780
rect 2746 19740 5540 19768
rect 2501 19731 2559 19737
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2133 19703 2191 19709
rect 2133 19700 2145 19703
rect 1728 19672 2145 19700
rect 1728 19660 1734 19672
rect 2133 19669 2145 19672
rect 2179 19669 2191 19703
rect 2516 19700 2544 19731
rect 5534 19728 5540 19740
rect 5592 19728 5598 19780
rect 3326 19700 3332 19712
rect 2516 19672 3332 19700
rect 2133 19663 2191 19669
rect 3326 19660 3332 19672
rect 3384 19700 3390 19712
rect 3786 19700 3792 19712
rect 3384 19672 3792 19700
rect 3384 19660 3390 19672
rect 3786 19660 3792 19672
rect 3844 19660 3850 19712
rect 3881 19703 3939 19709
rect 3881 19669 3893 19703
rect 3927 19700 3939 19703
rect 4890 19700 4896 19712
rect 3927 19672 4896 19700
rect 3927 19669 3939 19672
rect 3881 19663 3939 19669
rect 4890 19660 4896 19672
rect 4948 19660 4954 19712
rect 5445 19703 5503 19709
rect 5445 19669 5457 19703
rect 5491 19700 5503 19703
rect 5644 19700 5672 19876
rect 6822 19864 6828 19876
rect 6880 19864 6886 19916
rect 6569 19839 6627 19845
rect 6569 19805 6581 19839
rect 6615 19836 6627 19839
rect 6730 19836 6736 19848
rect 6615 19808 6736 19836
rect 6615 19805 6627 19808
rect 6569 19799 6627 19805
rect 6730 19796 6736 19808
rect 6788 19796 6794 19848
rect 7024 19836 7052 20012
rect 7558 20000 7564 20052
rect 7616 20040 7622 20052
rect 9033 20043 9091 20049
rect 7616 20012 8892 20040
rect 7616 20000 7622 20012
rect 7098 19932 7104 19984
rect 7156 19972 7162 19984
rect 8757 19975 8815 19981
rect 7156 19944 8524 19972
rect 7156 19932 7162 19944
rect 7469 19907 7527 19913
rect 7469 19873 7481 19907
rect 7515 19873 7527 19907
rect 8294 19904 8300 19916
rect 8255 19876 8300 19904
rect 7469 19867 7527 19873
rect 7098 19836 7104 19848
rect 7024 19808 7104 19836
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 6822 19728 6828 19780
rect 6880 19768 6886 19780
rect 7484 19768 7512 19867
rect 8294 19864 8300 19876
rect 8352 19864 8358 19916
rect 7742 19796 7748 19848
rect 7800 19836 7806 19848
rect 8205 19839 8263 19845
rect 8205 19836 8217 19839
rect 7800 19808 8217 19836
rect 7800 19796 7806 19808
rect 8205 19805 8217 19808
rect 8251 19805 8263 19839
rect 8205 19799 8263 19805
rect 6880 19740 7512 19768
rect 6880 19728 6886 19740
rect 7926 19728 7932 19780
rect 7984 19768 7990 19780
rect 8496 19768 8524 19944
rect 8757 19941 8769 19975
rect 8803 19941 8815 19975
rect 8864 19972 8892 20012
rect 9033 20009 9045 20043
rect 9079 20040 9091 20043
rect 10686 20040 10692 20052
rect 9079 20012 10692 20040
rect 9079 20009 9091 20012
rect 9033 20003 9091 20009
rect 10686 20000 10692 20012
rect 10744 20000 10750 20052
rect 10870 20040 10876 20052
rect 10831 20012 10876 20040
rect 10870 20000 10876 20012
rect 10928 20000 10934 20052
rect 11149 20043 11207 20049
rect 11149 20009 11161 20043
rect 11195 20040 11207 20043
rect 11882 20040 11888 20052
rect 11195 20012 11888 20040
rect 11195 20009 11207 20012
rect 11149 20003 11207 20009
rect 11882 20000 11888 20012
rect 11940 20000 11946 20052
rect 12434 20000 12440 20052
rect 12492 20040 12498 20052
rect 12802 20040 12808 20052
rect 12492 20012 12537 20040
rect 12763 20012 12808 20040
rect 12492 20000 12498 20012
rect 12802 20000 12808 20012
rect 12860 20000 12866 20052
rect 13170 20040 13176 20052
rect 13131 20012 13176 20040
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 13446 20040 13452 20052
rect 13407 20012 13452 20040
rect 13446 20000 13452 20012
rect 13504 20000 13510 20052
rect 13722 20040 13728 20052
rect 13683 20012 13728 20040
rect 13722 20000 13728 20012
rect 13780 20000 13786 20052
rect 14642 20040 14648 20052
rect 14603 20012 14648 20040
rect 14642 20000 14648 20012
rect 14700 20000 14706 20052
rect 15010 20040 15016 20052
rect 14971 20012 15016 20040
rect 15010 20000 15016 20012
rect 15068 20000 15074 20052
rect 15381 20043 15439 20049
rect 15381 20009 15393 20043
rect 15427 20040 15439 20043
rect 15930 20040 15936 20052
rect 15427 20012 15936 20040
rect 15427 20009 15439 20012
rect 15381 20003 15439 20009
rect 15930 20000 15936 20012
rect 15988 20000 15994 20052
rect 16114 20040 16120 20052
rect 16075 20012 16120 20040
rect 16114 20000 16120 20012
rect 16172 20000 16178 20052
rect 17034 20000 17040 20052
rect 17092 20040 17098 20052
rect 17589 20043 17647 20049
rect 17589 20040 17601 20043
rect 17092 20012 17601 20040
rect 17092 20000 17098 20012
rect 17589 20009 17601 20012
rect 17635 20009 17647 20043
rect 17589 20003 17647 20009
rect 17770 20000 17776 20052
rect 17828 20040 17834 20052
rect 18233 20043 18291 20049
rect 18233 20040 18245 20043
rect 17828 20012 18245 20040
rect 17828 20000 17834 20012
rect 18233 20009 18245 20012
rect 18279 20009 18291 20043
rect 18690 20040 18696 20052
rect 18233 20003 18291 20009
rect 18432 20012 18696 20040
rect 9493 19975 9551 19981
rect 9493 19972 9505 19975
rect 8864 19944 9505 19972
rect 8757 19935 8815 19941
rect 9493 19941 9505 19944
rect 9539 19941 9551 19975
rect 9493 19935 9551 19941
rect 8772 19904 8800 19935
rect 11238 19932 11244 19984
rect 11296 19972 11302 19984
rect 12253 19975 12311 19981
rect 12253 19972 12265 19975
rect 11296 19944 12265 19972
rect 11296 19932 11302 19944
rect 12253 19941 12265 19944
rect 12299 19941 12311 19975
rect 12253 19935 12311 19941
rect 12342 19932 12348 19984
rect 12400 19972 12406 19984
rect 15838 19972 15844 19984
rect 12400 19944 15844 19972
rect 12400 19932 12406 19944
rect 15838 19932 15844 19944
rect 15896 19932 15902 19984
rect 16942 19932 16948 19984
rect 17000 19972 17006 19984
rect 17221 19975 17279 19981
rect 17221 19972 17233 19975
rect 17000 19944 17233 19972
rect 17000 19932 17006 19944
rect 17221 19941 17233 19944
rect 17267 19941 17279 19975
rect 17221 19935 17279 19941
rect 17402 19932 17408 19984
rect 17460 19972 17466 19984
rect 17957 19975 18015 19981
rect 17957 19972 17969 19975
rect 17460 19944 17969 19972
rect 17460 19932 17466 19944
rect 17957 19941 17969 19944
rect 18003 19941 18015 19975
rect 17957 19935 18015 19941
rect 11425 19907 11483 19913
rect 8772 19876 10824 19904
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 8754 19836 8760 19848
rect 8619 19808 8760 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 8754 19796 8760 19808
rect 8812 19796 8818 19848
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 10689 19839 10747 19845
rect 10689 19836 10701 19839
rect 9640 19808 10701 19836
rect 9640 19796 9646 19808
rect 10689 19805 10701 19808
rect 10735 19805 10747 19839
rect 10689 19799 10747 19805
rect 9122 19768 9128 19780
rect 7984 19740 8432 19768
rect 8496 19740 9128 19768
rect 7984 19728 7990 19740
rect 6914 19700 6920 19712
rect 5491 19672 5672 19700
rect 6875 19672 6920 19700
rect 5491 19669 5503 19672
rect 5445 19663 5503 19669
rect 6914 19660 6920 19672
rect 6972 19660 6978 19712
rect 7282 19700 7288 19712
rect 7243 19672 7288 19700
rect 7282 19660 7288 19672
rect 7340 19660 7346 19712
rect 7377 19703 7435 19709
rect 7377 19669 7389 19703
rect 7423 19700 7435 19703
rect 7745 19703 7803 19709
rect 7745 19700 7757 19703
rect 7423 19672 7757 19700
rect 7423 19669 7435 19672
rect 7377 19663 7435 19669
rect 7745 19669 7757 19672
rect 7791 19669 7803 19703
rect 8110 19700 8116 19712
rect 8071 19672 8116 19700
rect 7745 19663 7803 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 8404 19700 8432 19740
rect 9122 19728 9128 19740
rect 9180 19728 9186 19780
rect 9398 19728 9404 19780
rect 9456 19768 9462 19780
rect 9677 19771 9735 19777
rect 9677 19768 9689 19771
rect 9456 19740 9689 19768
rect 9456 19728 9462 19740
rect 9677 19737 9689 19740
rect 9723 19737 9735 19771
rect 9677 19731 9735 19737
rect 9766 19728 9772 19780
rect 9824 19768 9830 19780
rect 10045 19771 10103 19777
rect 10045 19768 10057 19771
rect 9824 19740 10057 19768
rect 9824 19728 9830 19740
rect 10045 19737 10057 19740
rect 10091 19737 10103 19771
rect 10045 19731 10103 19737
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10413 19771 10471 19777
rect 10413 19768 10425 19771
rect 10192 19740 10425 19768
rect 10192 19728 10198 19740
rect 10413 19737 10425 19740
rect 10459 19737 10471 19771
rect 10796 19768 10824 19876
rect 11425 19873 11437 19907
rect 11471 19904 11483 19907
rect 11698 19904 11704 19916
rect 11471 19876 11704 19904
rect 11471 19873 11483 19876
rect 11425 19867 11483 19873
rect 11698 19864 11704 19876
rect 11756 19864 11762 19916
rect 13354 19904 13360 19916
rect 13004 19876 13360 19904
rect 10962 19836 10968 19848
rect 10923 19808 10968 19836
rect 10962 19796 10968 19808
rect 11020 19796 11026 19848
rect 11054 19796 11060 19848
rect 11112 19836 11118 19848
rect 11517 19839 11575 19845
rect 11517 19836 11529 19839
rect 11112 19808 11529 19836
rect 11112 19796 11118 19808
rect 11517 19805 11529 19808
rect 11563 19805 11575 19839
rect 12069 19839 12127 19845
rect 12069 19836 12081 19839
rect 11517 19799 11575 19805
rect 11716 19808 12081 19836
rect 10796 19740 11192 19768
rect 10413 19731 10471 19737
rect 9214 19700 9220 19712
rect 8404 19672 9220 19700
rect 9214 19660 9220 19672
rect 9272 19700 9278 19712
rect 9309 19703 9367 19709
rect 9309 19700 9321 19703
rect 9272 19672 9321 19700
rect 9272 19660 9278 19672
rect 9309 19669 9321 19672
rect 9355 19669 9367 19703
rect 9950 19700 9956 19712
rect 9911 19672 9956 19700
rect 9309 19663 9367 19669
rect 9950 19660 9956 19672
rect 10008 19660 10014 19712
rect 10318 19700 10324 19712
rect 10279 19672 10324 19700
rect 10318 19660 10324 19672
rect 10376 19660 10382 19712
rect 11164 19700 11192 19740
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 11609 19771 11667 19777
rect 11609 19768 11621 19771
rect 11296 19740 11621 19768
rect 11296 19728 11302 19740
rect 11609 19737 11621 19740
rect 11655 19737 11667 19771
rect 11609 19731 11667 19737
rect 11716 19700 11744 19808
rect 12069 19805 12081 19808
rect 12115 19805 12127 19839
rect 12069 19799 12127 19805
rect 12434 19796 12440 19848
rect 12492 19836 12498 19848
rect 13004 19845 13032 19876
rect 13354 19864 13360 19876
rect 13412 19864 13418 19916
rect 18432 19904 18460 20012
rect 18690 20000 18696 20012
rect 18748 20000 18754 20052
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 20346 20040 20352 20052
rect 18984 20012 20352 20040
rect 18509 19975 18567 19981
rect 18509 19941 18521 19975
rect 18555 19941 18567 19975
rect 18509 19935 18567 19941
rect 16316 19876 18460 19904
rect 12621 19839 12679 19845
rect 12621 19836 12633 19839
rect 12492 19808 12633 19836
rect 12492 19796 12498 19808
rect 12621 19805 12633 19808
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 12989 19839 13047 19845
rect 12989 19805 13001 19839
rect 13035 19805 13047 19839
rect 12989 19799 13047 19805
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 13228 19808 13277 19836
rect 13228 19796 13234 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 13541 19839 13599 19845
rect 13541 19805 13553 19839
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 14369 19839 14427 19845
rect 14369 19805 14381 19839
rect 14415 19836 14427 19839
rect 14461 19839 14519 19845
rect 14461 19836 14473 19839
rect 14415 19808 14473 19836
rect 14415 19805 14427 19808
rect 14369 19799 14427 19805
rect 14461 19805 14473 19808
rect 14507 19805 14519 19839
rect 14826 19836 14832 19848
rect 14787 19808 14832 19836
rect 14461 19799 14519 19805
rect 11882 19728 11888 19780
rect 11940 19768 11946 19780
rect 11940 19740 12296 19768
rect 11940 19728 11946 19740
rect 11164 19672 11744 19700
rect 11977 19703 12035 19709
rect 11977 19669 11989 19703
rect 12023 19700 12035 19703
rect 12158 19700 12164 19712
rect 12023 19672 12164 19700
rect 12023 19669 12035 19672
rect 11977 19663 12035 19669
rect 12158 19660 12164 19672
rect 12216 19660 12222 19712
rect 12268 19700 12296 19740
rect 12342 19728 12348 19780
rect 12400 19768 12406 19780
rect 13556 19768 13584 19799
rect 13817 19771 13875 19777
rect 13817 19768 13829 19771
rect 12400 19740 13829 19768
rect 12400 19728 12406 19740
rect 13817 19737 13829 19740
rect 13863 19737 13875 19771
rect 14476 19768 14504 19799
rect 14826 19796 14832 19808
rect 14884 19796 14890 19848
rect 15194 19836 15200 19848
rect 15155 19808 15200 19836
rect 15194 19796 15200 19808
rect 15252 19796 15258 19848
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19836 15807 19839
rect 15930 19836 15936 19848
rect 15795 19808 15936 19836
rect 15795 19805 15807 19808
rect 15749 19799 15807 19805
rect 15930 19796 15936 19808
rect 15988 19796 15994 19848
rect 16316 19845 16344 19876
rect 16301 19839 16359 19845
rect 16301 19805 16313 19839
rect 16347 19805 16359 19839
rect 16301 19799 16359 19805
rect 16390 19796 16396 19848
rect 16448 19836 16454 19848
rect 16485 19839 16543 19845
rect 16485 19836 16497 19839
rect 16448 19808 16497 19836
rect 16448 19796 16454 19808
rect 16485 19805 16497 19808
rect 16531 19805 16543 19839
rect 16666 19836 16672 19848
rect 16485 19799 16543 19805
rect 16592 19808 16672 19836
rect 14550 19768 14556 19780
rect 14476 19740 14556 19768
rect 13817 19731 13875 19737
rect 14550 19728 14556 19740
rect 14608 19728 14614 19780
rect 14844 19768 14872 19796
rect 15473 19771 15531 19777
rect 15473 19768 15485 19771
rect 14844 19740 15485 19768
rect 15473 19737 15485 19740
rect 15519 19737 15531 19771
rect 16592 19768 16620 19808
rect 16666 19796 16672 19808
rect 16724 19796 16730 19848
rect 16761 19839 16819 19845
rect 16761 19805 16773 19839
rect 16807 19836 16819 19839
rect 16942 19836 16948 19848
rect 16807 19808 16948 19836
rect 16807 19805 16819 19808
rect 16761 19799 16819 19805
rect 16942 19796 16948 19808
rect 17000 19796 17006 19848
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17402 19836 17408 19848
rect 17363 19808 17408 19836
rect 17037 19799 17095 19805
rect 17052 19768 17080 19799
rect 17402 19796 17408 19808
rect 17460 19796 17466 19848
rect 17586 19796 17592 19848
rect 17644 19836 17650 19848
rect 17773 19839 17831 19845
rect 17773 19836 17785 19839
rect 17644 19808 17785 19836
rect 17644 19796 17650 19808
rect 17773 19805 17785 19808
rect 17819 19805 17831 19839
rect 17773 19799 17831 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19836 18475 19839
rect 18524 19836 18552 19935
rect 18782 19932 18788 19984
rect 18840 19972 18846 19984
rect 18984 19972 19012 20012
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20530 20040 20536 20052
rect 20491 20012 20536 20040
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 18840 19944 19012 19972
rect 18840 19932 18846 19944
rect 19058 19932 19064 19984
rect 19116 19972 19122 19984
rect 19116 19944 20576 19972
rect 19116 19932 19122 19944
rect 20548 19916 20576 19944
rect 19610 19864 19616 19916
rect 19668 19864 19674 19916
rect 20530 19864 20536 19916
rect 20588 19864 20594 19916
rect 20806 19864 20812 19916
rect 20864 19904 20870 19916
rect 20901 19907 20959 19913
rect 20901 19904 20913 19907
rect 20864 19876 20913 19904
rect 20864 19864 20870 19876
rect 20901 19873 20913 19876
rect 20947 19873 20959 19907
rect 20901 19867 20959 19873
rect 18463 19808 18552 19836
rect 18693 19839 18751 19845
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18874 19836 18880 19848
rect 18739 19808 18880 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18874 19796 18880 19808
rect 18932 19796 18938 19848
rect 19061 19839 19119 19845
rect 19061 19805 19073 19839
rect 19107 19805 19119 19839
rect 19628 19836 19656 19864
rect 20346 19845 20352 19848
rect 19705 19839 19763 19845
rect 19705 19836 19717 19839
rect 19628 19808 19717 19836
rect 19061 19799 19119 19805
rect 19705 19805 19717 19808
rect 19751 19805 19763 19839
rect 19705 19799 19763 19805
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19805 20039 19839
rect 19981 19799 20039 19805
rect 20337 19839 20352 19845
rect 20337 19805 20349 19839
rect 20337 19799 20352 19805
rect 15473 19731 15531 19737
rect 15948 19740 16620 19768
rect 16684 19740 17080 19768
rect 15948 19709 15976 19740
rect 16684 19709 16712 19740
rect 18598 19728 18604 19780
rect 18656 19768 18662 19780
rect 19076 19768 19104 19799
rect 19426 19768 19432 19780
rect 18656 19740 19104 19768
rect 19387 19740 19432 19768
rect 18656 19728 18662 19740
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 19996 19768 20024 19799
rect 20346 19796 20352 19799
rect 20404 19796 20410 19848
rect 20714 19836 20720 19848
rect 20675 19808 20720 19836
rect 20714 19796 20720 19808
rect 20772 19796 20778 19848
rect 21266 19836 21272 19848
rect 21227 19808 21272 19836
rect 21266 19796 21272 19808
rect 21324 19796 21330 19848
rect 22002 19768 22008 19780
rect 19536 19740 20024 19768
rect 20180 19740 22008 19768
rect 14093 19703 14151 19709
rect 14093 19700 14105 19703
rect 12268 19672 14105 19700
rect 14093 19669 14105 19672
rect 14139 19669 14151 19703
rect 14093 19663 14151 19669
rect 15933 19703 15991 19709
rect 15933 19669 15945 19703
rect 15979 19669 15991 19703
rect 15933 19663 15991 19669
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19669 16727 19703
rect 16669 19663 16727 19669
rect 16945 19703 17003 19709
rect 16945 19669 16957 19703
rect 16991 19700 17003 19703
rect 17126 19700 17132 19712
rect 16991 19672 17132 19700
rect 16991 19669 17003 19672
rect 16945 19663 17003 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 18506 19660 18512 19712
rect 18564 19700 18570 19712
rect 19536 19700 19564 19740
rect 18564 19672 19564 19700
rect 18564 19660 18570 19672
rect 19610 19660 19616 19712
rect 19668 19700 19674 19712
rect 20180 19709 20208 19740
rect 22002 19728 22008 19740
rect 22060 19728 22066 19780
rect 19797 19703 19855 19709
rect 19797 19700 19809 19703
rect 19668 19672 19809 19700
rect 19668 19660 19674 19672
rect 19797 19669 19809 19672
rect 19843 19669 19855 19703
rect 19797 19663 19855 19669
rect 20165 19703 20223 19709
rect 20165 19669 20177 19703
rect 20211 19669 20223 19703
rect 20165 19663 20223 19669
rect 21453 19703 21511 19709
rect 21453 19669 21465 19703
rect 21499 19700 21511 19703
rect 21542 19700 21548 19712
rect 21499 19672 21548 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 21542 19660 21548 19672
rect 21600 19660 21606 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 2225 19499 2283 19505
rect 2225 19465 2237 19499
rect 2271 19465 2283 19499
rect 2225 19459 2283 19465
rect 2240 19428 2268 19459
rect 2590 19456 2596 19508
rect 2648 19496 2654 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 2648 19468 2973 19496
rect 2648 19456 2654 19468
rect 2961 19465 2973 19468
rect 3007 19465 3019 19499
rect 2961 19459 3019 19465
rect 3421 19499 3479 19505
rect 3421 19465 3433 19499
rect 3467 19496 3479 19499
rect 5445 19499 5503 19505
rect 3467 19468 5396 19496
rect 3467 19465 3479 19468
rect 3421 19459 3479 19465
rect 2866 19428 2872 19440
rect 2240 19400 2872 19428
rect 2866 19388 2872 19400
rect 2924 19388 2930 19440
rect 3970 19428 3976 19440
rect 3620 19400 3976 19428
rect 1673 19363 1731 19369
rect 1673 19329 1685 19363
rect 1719 19360 1731 19363
rect 1946 19360 1952 19372
rect 1719 19332 1952 19360
rect 1719 19329 1731 19332
rect 1673 19323 1731 19329
rect 1946 19320 1952 19332
rect 2004 19320 2010 19372
rect 2038 19320 2044 19372
rect 2096 19360 2102 19372
rect 2096 19332 2141 19360
rect 2096 19320 2102 19332
rect 2314 19320 2320 19372
rect 2372 19360 2378 19372
rect 2409 19363 2467 19369
rect 2409 19360 2421 19363
rect 2372 19332 2421 19360
rect 2372 19320 2378 19332
rect 2409 19329 2421 19332
rect 2455 19329 2467 19363
rect 2409 19323 2467 19329
rect 2498 19320 2504 19372
rect 2556 19360 2562 19372
rect 2556 19332 2636 19360
rect 2556 19320 2562 19332
rect 1854 19224 1860 19236
rect 1815 19196 1860 19224
rect 1854 19184 1860 19196
rect 1912 19184 1918 19236
rect 2608 19233 2636 19332
rect 2774 19320 2780 19372
rect 2832 19360 2838 19372
rect 2832 19332 2877 19360
rect 2832 19320 2838 19332
rect 3234 19320 3240 19372
rect 3292 19360 3298 19372
rect 3329 19363 3387 19369
rect 3329 19360 3341 19363
rect 3292 19332 3341 19360
rect 3292 19320 3298 19332
rect 3329 19329 3341 19332
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 2866 19252 2872 19304
rect 2924 19292 2930 19304
rect 3510 19292 3516 19304
rect 2924 19264 3516 19292
rect 2924 19252 2930 19264
rect 3510 19252 3516 19264
rect 3568 19252 3574 19304
rect 3620 19301 3648 19400
rect 3970 19388 3976 19400
rect 4028 19388 4034 19440
rect 4890 19388 4896 19440
rect 4948 19428 4954 19440
rect 5086 19431 5144 19437
rect 5086 19428 5098 19431
rect 4948 19400 5098 19428
rect 4948 19388 4954 19400
rect 5086 19397 5098 19400
rect 5132 19397 5144 19431
rect 5368 19428 5396 19468
rect 5445 19465 5457 19499
rect 5491 19496 5503 19499
rect 5626 19496 5632 19508
rect 5491 19468 5632 19496
rect 5491 19465 5503 19468
rect 5445 19459 5503 19465
rect 5626 19456 5632 19468
rect 5684 19456 5690 19508
rect 5736 19468 7236 19496
rect 5736 19428 5764 19468
rect 5368 19400 5764 19428
rect 5813 19431 5871 19437
rect 5086 19391 5144 19397
rect 5813 19397 5825 19431
rect 5859 19428 5871 19431
rect 5902 19428 5908 19440
rect 5859 19400 5908 19428
rect 5859 19397 5871 19400
rect 5813 19391 5871 19397
rect 5902 19388 5908 19400
rect 5960 19388 5966 19440
rect 7006 19428 7012 19440
rect 6380 19400 7012 19428
rect 3694 19320 3700 19372
rect 3752 19360 3758 19372
rect 5353 19363 5411 19369
rect 3752 19332 5304 19360
rect 3752 19320 3758 19332
rect 3605 19295 3663 19301
rect 3605 19261 3617 19295
rect 3651 19261 3663 19295
rect 4062 19292 4068 19304
rect 3605 19255 3663 19261
rect 3804 19264 4068 19292
rect 2593 19227 2651 19233
rect 2593 19193 2605 19227
rect 2639 19193 2651 19227
rect 2593 19187 2651 19193
rect 2958 19184 2964 19236
rect 3016 19224 3022 19236
rect 3804 19224 3832 19264
rect 4062 19252 4068 19264
rect 4120 19252 4126 19304
rect 5276 19292 5304 19332
rect 5353 19329 5365 19363
rect 5399 19360 5411 19363
rect 5442 19360 5448 19372
rect 5399 19332 5448 19360
rect 5399 19329 5411 19332
rect 5353 19323 5411 19329
rect 5442 19320 5448 19332
rect 5500 19360 5506 19372
rect 6380 19360 6408 19400
rect 7006 19388 7012 19400
rect 7064 19388 7070 19440
rect 7208 19428 7236 19468
rect 7282 19456 7288 19508
rect 7340 19496 7346 19508
rect 8297 19499 8355 19505
rect 8297 19496 8309 19499
rect 7340 19468 8309 19496
rect 7340 19456 7346 19468
rect 8297 19465 8309 19468
rect 8343 19465 8355 19499
rect 9306 19496 9312 19508
rect 9267 19468 9312 19496
rect 8297 19459 8355 19465
rect 9306 19456 9312 19468
rect 9364 19456 9370 19508
rect 9582 19496 9588 19508
rect 9543 19468 9588 19496
rect 9582 19456 9588 19468
rect 9640 19456 9646 19508
rect 9858 19456 9864 19508
rect 9916 19496 9922 19508
rect 9953 19499 10011 19505
rect 9953 19496 9965 19499
rect 9916 19468 9965 19496
rect 9916 19456 9922 19468
rect 9953 19465 9965 19468
rect 9999 19465 10011 19499
rect 9953 19459 10011 19465
rect 10413 19499 10471 19505
rect 10413 19465 10425 19499
rect 10459 19496 10471 19499
rect 11054 19496 11060 19508
rect 10459 19468 11060 19496
rect 10459 19465 10471 19468
rect 10413 19459 10471 19465
rect 11054 19456 11060 19468
rect 11112 19456 11118 19508
rect 11238 19496 11244 19508
rect 11199 19468 11244 19496
rect 11238 19456 11244 19468
rect 11296 19456 11302 19508
rect 11698 19456 11704 19508
rect 11756 19496 11762 19508
rect 12434 19496 12440 19508
rect 11756 19468 12440 19496
rect 11756 19456 11762 19468
rect 12434 19456 12440 19468
rect 12492 19496 12498 19508
rect 12897 19499 12955 19505
rect 12897 19496 12909 19499
rect 12492 19468 12909 19496
rect 12492 19456 12498 19468
rect 12897 19465 12909 19468
rect 12943 19465 12955 19499
rect 13170 19496 13176 19508
rect 13131 19468 13176 19496
rect 12897 19459 12955 19465
rect 13170 19456 13176 19468
rect 13228 19456 13234 19508
rect 17037 19499 17095 19505
rect 17037 19465 17049 19499
rect 17083 19465 17095 19499
rect 17037 19459 17095 19465
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17310 19496 17316 19508
rect 17175 19468 17316 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 8757 19431 8815 19437
rect 8757 19428 8769 19431
rect 7208 19400 8769 19428
rect 5500 19332 6408 19360
rect 5500 19320 5506 19332
rect 6454 19320 6460 19372
rect 6512 19360 6518 19372
rect 6638 19360 6644 19372
rect 6512 19332 6644 19360
rect 6512 19320 6518 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 7208 19360 7236 19400
rect 8757 19397 8769 19400
rect 8803 19428 8815 19431
rect 10045 19431 10103 19437
rect 8803 19400 9996 19428
rect 8803 19397 8815 19400
rect 8757 19391 8815 19397
rect 7024 19332 7236 19360
rect 7949 19363 8007 19369
rect 7024 19304 7052 19332
rect 7949 19329 7961 19363
rect 7995 19360 8007 19363
rect 8294 19360 8300 19372
rect 7995 19332 8300 19360
rect 7995 19329 8007 19332
rect 7949 19323 8007 19329
rect 8294 19320 8300 19332
rect 8352 19320 8358 19372
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8665 19363 8723 19369
rect 8665 19360 8677 19363
rect 8628 19332 8677 19360
rect 8628 19320 8634 19332
rect 8665 19329 8677 19332
rect 8711 19329 8723 19363
rect 9122 19360 9128 19372
rect 9083 19332 9128 19360
rect 8665 19323 8723 19329
rect 9122 19320 9128 19332
rect 9180 19320 9186 19372
rect 9401 19363 9459 19369
rect 9401 19329 9413 19363
rect 9447 19329 9459 19363
rect 9968 19360 9996 19400
rect 10045 19397 10057 19431
rect 10091 19428 10103 19431
rect 10134 19428 10140 19440
rect 10091 19400 10140 19428
rect 10091 19397 10103 19400
rect 10045 19391 10103 19397
rect 10134 19388 10140 19400
rect 10192 19388 10198 19440
rect 10778 19428 10784 19440
rect 10739 19400 10784 19428
rect 10778 19388 10784 19400
rect 10836 19388 10842 19440
rect 11146 19388 11152 19440
rect 11204 19428 11210 19440
rect 11882 19428 11888 19440
rect 11204 19400 11888 19428
rect 11204 19388 11210 19400
rect 11882 19388 11888 19400
rect 11940 19388 11946 19440
rect 12250 19388 12256 19440
rect 12308 19428 12314 19440
rect 14185 19431 14243 19437
rect 14185 19428 14197 19431
rect 12308 19400 14197 19428
rect 12308 19388 12314 19400
rect 14185 19397 14197 19400
rect 14231 19397 14243 19431
rect 17052 19428 17080 19459
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 17586 19496 17592 19508
rect 17547 19468 17592 19496
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 17773 19499 17831 19505
rect 17773 19465 17785 19499
rect 17819 19496 17831 19499
rect 17862 19496 17868 19508
rect 17819 19468 17868 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 17862 19456 17868 19468
rect 17920 19456 17926 19508
rect 18233 19499 18291 19505
rect 18233 19465 18245 19499
rect 18279 19465 18291 19499
rect 18506 19496 18512 19508
rect 18467 19468 18512 19496
rect 18233 19459 18291 19465
rect 18138 19428 18144 19440
rect 17052 19400 18144 19428
rect 14185 19391 14243 19397
rect 10226 19360 10232 19372
rect 9968 19332 10232 19360
rect 9401 19323 9459 19329
rect 5902 19292 5908 19304
rect 5276 19264 5396 19292
rect 5863 19264 5908 19292
rect 3016 19196 3832 19224
rect 3881 19227 3939 19233
rect 3016 19184 3022 19196
rect 3881 19193 3893 19227
rect 3927 19224 3939 19227
rect 4154 19224 4160 19236
rect 3927 19196 4160 19224
rect 3927 19193 3939 19196
rect 3881 19187 3939 19193
rect 4154 19184 4160 19196
rect 4212 19184 4218 19236
rect 5368 19224 5396 19264
rect 5902 19252 5908 19264
rect 5960 19252 5966 19304
rect 6086 19252 6092 19304
rect 6144 19292 6150 19304
rect 6730 19292 6736 19304
rect 6144 19264 6736 19292
rect 6144 19252 6150 19264
rect 6730 19252 6736 19264
rect 6788 19252 6794 19304
rect 7006 19252 7012 19304
rect 7064 19252 7070 19304
rect 8205 19295 8263 19301
rect 8205 19261 8217 19295
rect 8251 19261 8263 19295
rect 8205 19255 8263 19261
rect 8849 19295 8907 19301
rect 8849 19261 8861 19295
rect 8895 19261 8907 19295
rect 9416 19292 9444 19323
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 10870 19360 10876 19372
rect 10831 19332 10876 19360
rect 10870 19320 10876 19332
rect 10928 19320 10934 19372
rect 11773 19363 11831 19369
rect 11773 19360 11785 19363
rect 10980 19332 11785 19360
rect 9490 19292 9496 19304
rect 9416 19264 9496 19292
rect 8849 19255 8907 19261
rect 6362 19224 6368 19236
rect 5368 19196 6368 19224
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 8220 19168 8248 19255
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 8864 19224 8892 19255
rect 9490 19252 9496 19264
rect 9548 19252 9554 19304
rect 9861 19295 9919 19301
rect 9861 19261 9873 19295
rect 9907 19261 9919 19295
rect 9861 19255 9919 19261
rect 10689 19295 10747 19301
rect 10689 19261 10701 19295
rect 10735 19292 10747 19295
rect 10980 19292 11008 19332
rect 11773 19329 11785 19332
rect 11819 19329 11831 19363
rect 11773 19323 11831 19329
rect 12158 19320 12164 19372
rect 12216 19360 12222 19372
rect 12989 19363 13047 19369
rect 12989 19360 13001 19363
rect 12216 19332 13001 19360
rect 12216 19320 12222 19332
rect 12989 19329 13001 19332
rect 13035 19329 13047 19363
rect 12989 19323 13047 19329
rect 13630 19320 13636 19372
rect 13688 19360 13694 19372
rect 17328 19369 17356 19400
rect 18138 19388 18144 19400
rect 18196 19388 18202 19440
rect 18248 19428 18276 19459
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 18782 19496 18788 19508
rect 18743 19468 18788 19496
rect 18782 19456 18788 19468
rect 18840 19456 18846 19508
rect 19150 19496 19156 19508
rect 19111 19468 19156 19496
rect 19150 19456 19156 19468
rect 19208 19456 19214 19508
rect 19242 19456 19248 19508
rect 19300 19496 19306 19508
rect 19613 19499 19671 19505
rect 19613 19496 19625 19499
rect 19300 19468 19625 19496
rect 19300 19456 19306 19468
rect 19613 19465 19625 19468
rect 19659 19465 19671 19499
rect 19613 19459 19671 19465
rect 18248 19400 19288 19428
rect 16853 19363 16911 19369
rect 13688 19332 14136 19360
rect 13688 19320 13694 19332
rect 11514 19292 11520 19304
rect 10735 19264 11008 19292
rect 11475 19264 11520 19292
rect 10735 19261 10747 19264
rect 10689 19255 10747 19261
rect 8352 19196 8892 19224
rect 9876 19224 9904 19255
rect 10318 19224 10324 19236
rect 9876 19196 10324 19224
rect 8352 19184 8358 19196
rect 10318 19184 10324 19196
rect 10376 19224 10382 19236
rect 10704 19224 10732 19255
rect 11514 19252 11520 19264
rect 11572 19252 11578 19304
rect 12526 19252 12532 19304
rect 12584 19292 12590 19304
rect 14001 19295 14059 19301
rect 14001 19292 14013 19295
rect 12584 19264 14013 19292
rect 12584 19252 12590 19264
rect 14001 19261 14013 19264
rect 14047 19261 14059 19295
rect 14108 19292 14136 19332
rect 16853 19329 16865 19363
rect 16899 19329 16911 19363
rect 16853 19323 16911 19329
rect 17313 19363 17371 19369
rect 17313 19329 17325 19363
rect 17359 19329 17371 19363
rect 17313 19323 17371 19329
rect 17405 19363 17463 19369
rect 17405 19329 17417 19363
rect 17451 19329 17463 19363
rect 17954 19360 17960 19372
rect 17915 19332 17960 19360
rect 17405 19323 17463 19329
rect 14553 19295 14611 19301
rect 14553 19292 14565 19295
rect 14108 19264 14565 19292
rect 14001 19255 14059 19261
rect 14553 19261 14565 19264
rect 14599 19261 14611 19295
rect 14734 19292 14740 19304
rect 14695 19264 14740 19292
rect 14553 19255 14611 19261
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 15286 19292 15292 19304
rect 15199 19264 15292 19292
rect 15286 19252 15292 19264
rect 15344 19292 15350 19304
rect 16298 19292 16304 19304
rect 15344 19264 16304 19292
rect 15344 19252 15350 19264
rect 16298 19252 16304 19264
rect 16356 19252 16362 19304
rect 10376 19196 10732 19224
rect 10376 19184 10382 19196
rect 13538 19184 13544 19236
rect 13596 19224 13602 19236
rect 13633 19227 13691 19233
rect 13633 19224 13645 19227
rect 13596 19196 13645 19224
rect 13596 19184 13602 19196
rect 13633 19193 13645 19196
rect 13679 19193 13691 19227
rect 13633 19187 13691 19193
rect 13722 19184 13728 19236
rect 13780 19224 13786 19236
rect 15381 19227 15439 19233
rect 15381 19224 15393 19227
rect 13780 19196 15393 19224
rect 13780 19184 13786 19196
rect 15381 19193 15393 19196
rect 15427 19193 15439 19227
rect 15930 19224 15936 19236
rect 15381 19187 15439 19193
rect 15580 19196 15936 19224
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 3970 19156 3976 19168
rect 3931 19128 3976 19156
rect 3970 19116 3976 19128
rect 4028 19116 4034 19168
rect 6546 19116 6552 19168
rect 6604 19156 6610 19168
rect 6822 19156 6828 19168
rect 6604 19128 6649 19156
rect 6783 19128 6828 19156
rect 6604 19116 6610 19128
rect 6822 19116 6828 19128
rect 6880 19116 6886 19168
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 7926 19156 7932 19168
rect 6972 19128 7932 19156
rect 6972 19116 6978 19128
rect 7926 19116 7932 19128
rect 7984 19116 7990 19168
rect 8018 19116 8024 19168
rect 8076 19156 8082 19168
rect 8202 19156 8208 19168
rect 8076 19128 8208 19156
rect 8076 19116 8082 19128
rect 8202 19116 8208 19128
rect 8260 19116 8266 19168
rect 8478 19116 8484 19168
rect 8536 19156 8542 19168
rect 12250 19156 12256 19168
rect 8536 19128 12256 19156
rect 8536 19116 8542 19128
rect 12250 19116 12256 19128
rect 12308 19116 12314 19168
rect 12434 19116 12440 19168
rect 12492 19156 12498 19168
rect 12618 19156 12624 19168
rect 12492 19128 12624 19156
rect 12492 19116 12498 19128
rect 12618 19116 12624 19128
rect 12676 19116 12682 19168
rect 13354 19156 13360 19168
rect 13315 19128 13360 19156
rect 13354 19116 13360 19128
rect 13412 19116 13418 19168
rect 13446 19116 13452 19168
rect 13504 19156 13510 19168
rect 13814 19156 13820 19168
rect 13504 19128 13549 19156
rect 13775 19128 13820 19156
rect 13504 19116 13510 19128
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 14366 19156 14372 19168
rect 14327 19128 14372 19156
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 15010 19156 15016 19168
rect 14971 19128 15016 19156
rect 15010 19116 15016 19128
rect 15068 19116 15074 19168
rect 15286 19116 15292 19168
rect 15344 19156 15350 19168
rect 15580 19165 15608 19196
rect 15930 19184 15936 19196
rect 15988 19184 15994 19236
rect 16868 19224 16896 19323
rect 17420 19292 17448 19323
rect 17954 19320 17960 19332
rect 18012 19320 18018 19372
rect 18049 19363 18107 19369
rect 18049 19329 18061 19363
rect 18095 19360 18107 19363
rect 18230 19360 18236 19372
rect 18095 19332 18236 19360
rect 18095 19329 18107 19332
rect 18049 19323 18107 19329
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18325 19363 18383 19369
rect 18325 19329 18337 19363
rect 18371 19329 18383 19363
rect 18325 19323 18383 19329
rect 17586 19292 17592 19304
rect 17420 19264 17592 19292
rect 17586 19252 17592 19264
rect 17644 19252 17650 19304
rect 17972 19292 18000 19320
rect 18340 19292 18368 19323
rect 18414 19320 18420 19372
rect 18472 19360 18478 19372
rect 18601 19363 18659 19369
rect 18601 19360 18613 19363
rect 18472 19332 18613 19360
rect 18472 19320 18478 19332
rect 18601 19329 18613 19332
rect 18647 19360 18659 19363
rect 18966 19360 18972 19372
rect 18647 19332 18972 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18966 19320 18972 19332
rect 19024 19320 19030 19372
rect 17972 19264 18368 19292
rect 19260 19292 19288 19400
rect 19352 19400 19656 19428
rect 19352 19369 19380 19400
rect 19628 19372 19656 19400
rect 20898 19388 20904 19440
rect 20956 19428 20962 19440
rect 21545 19431 21603 19437
rect 21545 19428 21557 19431
rect 20956 19400 21557 19428
rect 20956 19388 20962 19400
rect 21545 19397 21557 19400
rect 21591 19397 21603 19431
rect 21545 19391 21603 19397
rect 19337 19363 19395 19369
rect 19337 19329 19349 19363
rect 19383 19329 19395 19363
rect 19337 19323 19395 19329
rect 19429 19363 19487 19369
rect 19429 19329 19441 19363
rect 19475 19360 19487 19363
rect 19518 19360 19524 19372
rect 19475 19332 19524 19360
rect 19475 19329 19487 19332
rect 19429 19323 19487 19329
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 19610 19320 19616 19372
rect 19668 19320 19674 19372
rect 19794 19292 19800 19304
rect 19260 19264 19656 19292
rect 19755 19264 19800 19292
rect 17310 19224 17316 19236
rect 16868 19196 17316 19224
rect 17310 19184 17316 19196
rect 17368 19224 17374 19236
rect 19334 19224 19340 19236
rect 17368 19196 19340 19224
rect 17368 19184 17374 19196
rect 19334 19184 19340 19196
rect 19392 19184 19398 19236
rect 19628 19224 19656 19264
rect 19794 19252 19800 19264
rect 19852 19252 19858 19304
rect 20346 19224 20352 19236
rect 19628 19196 20352 19224
rect 20346 19184 20352 19196
rect 20404 19184 20410 19236
rect 15565 19159 15623 19165
rect 15565 19156 15577 19159
rect 15344 19128 15577 19156
rect 15344 19116 15350 19128
rect 15565 19125 15577 19128
rect 15611 19125 15623 19159
rect 15746 19156 15752 19168
rect 15707 19128 15752 19156
rect 15565 19119 15623 19125
rect 15746 19116 15752 19128
rect 15804 19116 15810 19168
rect 16390 19156 16396 19168
rect 16351 19128 16396 19156
rect 16390 19116 16396 19128
rect 16448 19116 16454 19168
rect 16761 19159 16819 19165
rect 16761 19125 16773 19159
rect 16807 19156 16819 19159
rect 17034 19156 17040 19168
rect 16807 19128 17040 19156
rect 16807 19125 16819 19128
rect 16761 19119 16819 19125
rect 17034 19116 17040 19128
rect 17092 19116 17098 19168
rect 18782 19116 18788 19168
rect 18840 19156 18846 19168
rect 18969 19159 19027 19165
rect 18969 19156 18981 19159
rect 18840 19128 18981 19156
rect 18840 19116 18846 19128
rect 18969 19125 18981 19128
rect 19015 19156 19027 19159
rect 21174 19156 21180 19168
rect 19015 19128 21180 19156
rect 19015 19125 19027 19128
rect 18969 19119 19027 19125
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1762 18912 1768 18964
rect 1820 18952 1826 18964
rect 1857 18955 1915 18961
rect 1857 18952 1869 18955
rect 1820 18924 1869 18952
rect 1820 18912 1826 18924
rect 1857 18921 1869 18924
rect 1903 18921 1915 18955
rect 2222 18952 2228 18964
rect 2183 18924 2228 18952
rect 1857 18915 1915 18921
rect 2222 18912 2228 18924
rect 2280 18912 2286 18964
rect 2406 18912 2412 18964
rect 2464 18952 2470 18964
rect 2593 18955 2651 18961
rect 2593 18952 2605 18955
rect 2464 18924 2605 18952
rect 2464 18912 2470 18924
rect 2593 18921 2605 18924
rect 2639 18921 2651 18955
rect 3418 18952 3424 18964
rect 2593 18915 2651 18921
rect 2792 18924 3424 18952
rect 842 18844 848 18896
rect 900 18884 906 18896
rect 1118 18884 1124 18896
rect 900 18856 1124 18884
rect 900 18844 906 18856
rect 1118 18844 1124 18856
rect 1176 18844 1182 18896
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 2041 18751 2099 18757
rect 2041 18717 2053 18751
rect 2087 18748 2099 18751
rect 2314 18748 2320 18760
rect 2087 18720 2320 18748
rect 2087 18717 2099 18720
rect 2041 18711 2099 18717
rect 2314 18708 2320 18720
rect 2372 18708 2378 18760
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 2682 18748 2688 18760
rect 2455 18720 2688 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 2682 18708 2688 18720
rect 2740 18708 2746 18760
rect 2792 18757 2820 18924
rect 3418 18912 3424 18924
rect 3476 18912 3482 18964
rect 3973 18955 4031 18961
rect 3973 18921 3985 18955
rect 4019 18952 4031 18955
rect 4246 18952 4252 18964
rect 4019 18924 4252 18952
rect 4019 18921 4031 18924
rect 3973 18915 4031 18921
rect 4246 18912 4252 18924
rect 4304 18912 4310 18964
rect 5721 18955 5779 18961
rect 5721 18921 5733 18955
rect 5767 18952 5779 18955
rect 6086 18952 6092 18964
rect 5767 18924 6092 18952
rect 5767 18921 5779 18924
rect 5721 18915 5779 18921
rect 6086 18912 6092 18924
rect 6144 18912 6150 18964
rect 6730 18952 6736 18964
rect 6196 18924 6736 18952
rect 3694 18844 3700 18896
rect 3752 18884 3758 18896
rect 5350 18884 5356 18896
rect 3752 18856 5356 18884
rect 3752 18844 3758 18856
rect 5350 18844 5356 18856
rect 5408 18844 5414 18896
rect 6196 18884 6224 18924
rect 6730 18912 6736 18924
rect 6788 18952 6794 18964
rect 7282 18952 7288 18964
rect 6788 18924 7288 18952
rect 6788 18912 6794 18924
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 7466 18952 7472 18964
rect 7427 18924 7472 18952
rect 7466 18912 7472 18924
rect 7524 18912 7530 18964
rect 8110 18952 8116 18964
rect 7576 18924 8116 18952
rect 6104 18856 6224 18884
rect 3053 18819 3111 18825
rect 3053 18785 3065 18819
rect 3099 18816 3111 18819
rect 3099 18788 4016 18816
rect 3099 18785 3111 18788
rect 3053 18779 3111 18785
rect 3988 18760 4016 18788
rect 4522 18776 4528 18828
rect 4580 18816 4586 18828
rect 4709 18819 4767 18825
rect 4709 18816 4721 18819
rect 4580 18788 4721 18816
rect 4580 18776 4586 18788
rect 4709 18785 4721 18788
rect 4755 18785 4767 18819
rect 4890 18816 4896 18828
rect 4851 18788 4896 18816
rect 4709 18779 4767 18785
rect 4890 18776 4896 18788
rect 4948 18776 4954 18828
rect 6104 18816 6132 18856
rect 7576 18816 7604 18924
rect 8110 18912 8116 18924
rect 8168 18912 8174 18964
rect 8478 18952 8484 18964
rect 8439 18924 8484 18952
rect 8478 18912 8484 18924
rect 8536 18912 8542 18964
rect 8662 18912 8668 18964
rect 8720 18952 8726 18964
rect 9217 18955 9275 18961
rect 9217 18952 9229 18955
rect 8720 18924 9229 18952
rect 8720 18912 8726 18924
rect 9217 18921 9229 18924
rect 9263 18921 9275 18955
rect 9217 18915 9275 18921
rect 9769 18955 9827 18961
rect 9769 18921 9781 18955
rect 9815 18952 9827 18955
rect 9858 18952 9864 18964
rect 9815 18924 9864 18952
rect 9815 18921 9827 18924
rect 9769 18915 9827 18921
rect 9858 18912 9864 18924
rect 9916 18912 9922 18964
rect 10226 18912 10232 18964
rect 10284 18912 10290 18964
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 13814 18952 13820 18964
rect 10560 18924 13820 18952
rect 10560 18912 10566 18924
rect 13814 18912 13820 18924
rect 13872 18912 13878 18964
rect 14369 18955 14427 18961
rect 14369 18921 14381 18955
rect 14415 18952 14427 18955
rect 14458 18952 14464 18964
rect 14415 18924 14464 18952
rect 14415 18921 14427 18924
rect 14369 18915 14427 18921
rect 14458 18912 14464 18924
rect 14516 18912 14522 18964
rect 14737 18955 14795 18961
rect 14737 18921 14749 18955
rect 14783 18952 14795 18955
rect 15562 18952 15568 18964
rect 14783 18924 15568 18952
rect 14783 18921 14795 18924
rect 14737 18915 14795 18921
rect 15562 18912 15568 18924
rect 15620 18912 15626 18964
rect 16577 18955 16635 18961
rect 16577 18921 16589 18955
rect 16623 18952 16635 18955
rect 17402 18952 17408 18964
rect 16623 18924 17408 18952
rect 16623 18921 16635 18924
rect 16577 18915 16635 18921
rect 17402 18912 17408 18924
rect 17460 18912 17466 18964
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17865 18955 17923 18961
rect 17552 18924 17597 18952
rect 17552 18912 17558 18924
rect 17865 18921 17877 18955
rect 17911 18952 17923 18955
rect 18046 18952 18052 18964
rect 17911 18924 18052 18952
rect 17911 18921 17923 18924
rect 17865 18915 17923 18921
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 18230 18952 18236 18964
rect 18191 18924 18236 18952
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 19058 18952 19064 18964
rect 19019 18924 19064 18952
rect 19058 18912 19064 18924
rect 19116 18912 19122 18964
rect 19429 18955 19487 18961
rect 19429 18921 19441 18955
rect 19475 18952 19487 18955
rect 19978 18952 19984 18964
rect 19475 18924 19984 18952
rect 19475 18921 19487 18924
rect 19429 18915 19487 18921
rect 19978 18912 19984 18924
rect 20036 18912 20042 18964
rect 20438 18912 20444 18964
rect 20496 18952 20502 18964
rect 20533 18955 20591 18961
rect 20533 18952 20545 18955
rect 20496 18924 20545 18952
rect 20496 18912 20502 18924
rect 20533 18921 20545 18924
rect 20579 18921 20591 18955
rect 20533 18915 20591 18921
rect 5368 18788 6132 18816
rect 7024 18788 7604 18816
rect 8036 18856 8248 18884
rect 2777 18751 2835 18757
rect 2777 18717 2789 18751
rect 2823 18717 2835 18751
rect 2777 18711 2835 18717
rect 3237 18751 3295 18757
rect 3237 18717 3249 18751
rect 3283 18748 3295 18751
rect 3694 18748 3700 18760
rect 3283 18720 3700 18748
rect 3283 18717 3295 18720
rect 3237 18711 3295 18717
rect 3694 18708 3700 18720
rect 3752 18708 3758 18760
rect 3789 18751 3847 18757
rect 3789 18717 3801 18751
rect 3835 18748 3847 18751
rect 3878 18748 3884 18760
rect 3835 18720 3884 18748
rect 3835 18717 3847 18720
rect 3789 18711 3847 18717
rect 3878 18708 3884 18720
rect 3936 18708 3942 18760
rect 3970 18708 3976 18760
rect 4028 18748 4034 18760
rect 5261 18751 5319 18757
rect 5261 18748 5273 18751
rect 4028 18720 5273 18748
rect 4028 18708 4034 18720
rect 5261 18717 5273 18720
rect 5307 18717 5319 18751
rect 5261 18711 5319 18717
rect 3145 18683 3203 18689
rect 3145 18649 3157 18683
rect 3191 18680 3203 18683
rect 4617 18683 4675 18689
rect 3191 18652 4292 18680
rect 3191 18649 3203 18652
rect 3145 18643 3203 18649
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 3602 18612 3608 18624
rect 3563 18584 3608 18612
rect 3602 18572 3608 18584
rect 3660 18572 3666 18624
rect 4154 18612 4160 18624
rect 4115 18584 4160 18612
rect 4154 18572 4160 18584
rect 4212 18572 4218 18624
rect 4264 18621 4292 18652
rect 4617 18649 4629 18683
rect 4663 18680 4675 18683
rect 5368 18680 5396 18788
rect 6454 18708 6460 18760
rect 6512 18748 6518 18760
rect 7024 18748 7052 18788
rect 8036 18760 8064 18856
rect 8113 18819 8171 18825
rect 8113 18785 8125 18819
rect 8159 18785 8171 18819
rect 8113 18779 8171 18785
rect 6512 18720 7052 18748
rect 7101 18751 7159 18757
rect 6512 18708 6518 18720
rect 7101 18717 7113 18751
rect 7147 18748 7159 18751
rect 7374 18748 7380 18760
rect 7147 18720 7380 18748
rect 7147 18717 7159 18720
rect 7101 18711 7159 18717
rect 7374 18708 7380 18720
rect 7432 18708 7438 18760
rect 8018 18708 8024 18760
rect 8076 18708 8082 18760
rect 4663 18652 5396 18680
rect 4663 18649 4675 18652
rect 4617 18643 4675 18649
rect 5442 18640 5448 18692
rect 5500 18680 5506 18692
rect 5629 18683 5687 18689
rect 5500 18652 5545 18680
rect 5500 18640 5506 18652
rect 5629 18649 5641 18683
rect 5675 18680 5687 18683
rect 5718 18680 5724 18692
rect 5675 18652 5724 18680
rect 5675 18649 5687 18652
rect 5629 18643 5687 18649
rect 5718 18640 5724 18652
rect 5776 18640 5782 18692
rect 6178 18640 6184 18692
rect 6236 18680 6242 18692
rect 6730 18680 6736 18692
rect 6236 18652 6736 18680
rect 6236 18640 6242 18652
rect 6730 18640 6736 18652
rect 6788 18640 6794 18692
rect 6822 18640 6828 18692
rect 6880 18689 6886 18692
rect 6880 18680 6892 18689
rect 8128 18680 8156 18779
rect 8220 18748 8248 18856
rect 8386 18844 8392 18896
rect 8444 18884 8450 18896
rect 8573 18887 8631 18893
rect 8573 18884 8585 18887
rect 8444 18856 8585 18884
rect 8444 18844 8450 18856
rect 8573 18853 8585 18856
rect 8619 18853 8631 18887
rect 8573 18847 8631 18853
rect 8680 18856 8984 18884
rect 8680 18816 8708 18856
rect 8404 18788 8708 18816
rect 8404 18760 8432 18788
rect 8297 18751 8355 18757
rect 8297 18748 8309 18751
rect 8220 18720 8309 18748
rect 8297 18717 8309 18720
rect 8343 18717 8355 18751
rect 8297 18711 8355 18717
rect 8386 18708 8392 18760
rect 8444 18708 8450 18760
rect 8956 18757 8984 18856
rect 9122 18844 9128 18896
rect 9180 18884 9186 18896
rect 9493 18887 9551 18893
rect 9180 18856 9225 18884
rect 9180 18844 9186 18856
rect 9493 18853 9505 18887
rect 9539 18884 9551 18887
rect 10244 18884 10272 18912
rect 9539 18856 10272 18884
rect 9539 18853 9551 18856
rect 9493 18847 9551 18853
rect 12986 18844 12992 18896
rect 13044 18884 13050 18896
rect 13633 18887 13691 18893
rect 13633 18884 13645 18887
rect 13044 18856 13645 18884
rect 13044 18844 13050 18856
rect 13633 18853 13645 18856
rect 13679 18853 13691 18887
rect 13633 18847 13691 18853
rect 13722 18844 13728 18896
rect 13780 18884 13786 18896
rect 15286 18884 15292 18896
rect 13780 18856 15292 18884
rect 13780 18844 13786 18856
rect 15286 18844 15292 18856
rect 15344 18844 15350 18896
rect 17221 18887 17279 18893
rect 17221 18853 17233 18887
rect 17267 18884 17279 18887
rect 17310 18884 17316 18896
rect 17267 18856 17316 18884
rect 17267 18853 17279 18856
rect 17221 18847 17279 18853
rect 17310 18844 17316 18856
rect 17368 18844 17374 18896
rect 17954 18884 17960 18896
rect 17867 18856 17960 18884
rect 17954 18844 17960 18856
rect 18012 18884 18018 18896
rect 18874 18884 18880 18896
rect 18012 18856 18880 18884
rect 18012 18844 18018 18856
rect 18874 18844 18880 18856
rect 18932 18844 18938 18896
rect 19702 18884 19708 18896
rect 19663 18856 19708 18884
rect 19702 18844 19708 18856
rect 19760 18844 19766 18896
rect 19886 18844 19892 18896
rect 19944 18844 19950 18896
rect 20073 18887 20131 18893
rect 20073 18853 20085 18887
rect 20119 18884 20131 18887
rect 22738 18884 22744 18896
rect 20119 18856 22744 18884
rect 20119 18853 20131 18856
rect 20073 18847 20131 18853
rect 22738 18844 22744 18856
rect 22796 18844 22802 18896
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11624 18788 11805 18816
rect 11624 18760 11652 18788
rect 11793 18785 11805 18788
rect 11839 18785 11851 18819
rect 11793 18779 11851 18785
rect 12802 18776 12808 18828
rect 12860 18816 12866 18828
rect 13170 18816 13176 18828
rect 12860 18788 13176 18816
rect 12860 18776 12866 18788
rect 13170 18776 13176 18788
rect 13228 18816 13234 18828
rect 13265 18819 13323 18825
rect 13265 18816 13277 18819
rect 13228 18788 13277 18816
rect 13228 18776 13234 18788
rect 13265 18785 13277 18788
rect 13311 18785 13323 18819
rect 19904 18816 19932 18844
rect 13265 18779 13323 18785
rect 18156 18788 19932 18816
rect 8757 18751 8815 18757
rect 8757 18717 8769 18751
rect 8803 18717 8815 18751
rect 8757 18711 8815 18717
rect 8941 18751 8999 18757
rect 8941 18717 8953 18751
rect 8987 18717 8999 18751
rect 8941 18711 8999 18717
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18744 9459 18751
rect 9490 18744 9496 18760
rect 9447 18717 9496 18744
rect 9401 18716 9496 18717
rect 9401 18711 9459 18716
rect 6880 18652 8156 18680
rect 8772 18680 8800 18711
rect 9490 18708 9496 18716
rect 9548 18708 9554 18760
rect 9677 18751 9735 18757
rect 9677 18717 9689 18751
rect 9723 18748 9735 18751
rect 9766 18748 9772 18760
rect 9723 18720 9772 18748
rect 9723 18717 9735 18720
rect 9677 18711 9735 18717
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 10318 18708 10324 18760
rect 10376 18748 10382 18760
rect 10882 18751 10940 18757
rect 10882 18748 10894 18751
rect 10376 18720 10894 18748
rect 10376 18708 10382 18720
rect 10882 18717 10894 18720
rect 10928 18717 10940 18751
rect 10882 18711 10940 18717
rect 11149 18751 11207 18757
rect 11149 18717 11161 18751
rect 11195 18748 11207 18751
rect 11606 18748 11612 18760
rect 11195 18720 11612 18748
rect 11195 18717 11207 18720
rect 11149 18711 11207 18717
rect 11606 18708 11612 18720
rect 11664 18708 11670 18760
rect 12060 18751 12118 18757
rect 12060 18717 12072 18751
rect 12106 18748 12118 18751
rect 12526 18748 12532 18760
rect 12106 18720 12532 18748
rect 12106 18717 12118 18720
rect 12060 18711 12118 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 14185 18751 14243 18757
rect 14185 18748 14197 18751
rect 12820 18720 14197 18748
rect 10962 18680 10968 18692
rect 8772 18652 10968 18680
rect 6880 18643 6892 18652
rect 6880 18640 6886 18643
rect 10962 18640 10968 18652
rect 11020 18640 11026 18692
rect 12820 18680 12848 18720
rect 14185 18717 14197 18720
rect 14231 18717 14243 18751
rect 14550 18748 14556 18760
rect 14511 18720 14556 18748
rect 14185 18711 14243 18717
rect 13449 18683 13507 18689
rect 13449 18680 13461 18683
rect 11072 18652 11376 18680
rect 4249 18615 4307 18621
rect 4249 18581 4261 18615
rect 4295 18581 4307 18615
rect 4249 18575 4307 18581
rect 4798 18572 4804 18624
rect 4856 18612 4862 18624
rect 5077 18615 5135 18621
rect 5077 18612 5089 18615
rect 4856 18584 5089 18612
rect 4856 18572 4862 18584
rect 5077 18581 5089 18584
rect 5123 18581 5135 18615
rect 5077 18575 5135 18581
rect 5810 18572 5816 18624
rect 5868 18612 5874 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 5868 18584 7205 18612
rect 5868 18572 5874 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7834 18612 7840 18624
rect 7795 18584 7840 18612
rect 7193 18575 7251 18581
rect 7834 18572 7840 18584
rect 7892 18572 7898 18624
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8018 18612 8024 18624
rect 7975 18584 8024 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8018 18572 8024 18584
rect 8076 18572 8082 18624
rect 8110 18572 8116 18624
rect 8168 18612 8174 18624
rect 10134 18612 10140 18624
rect 8168 18584 10140 18612
rect 8168 18572 8174 18584
rect 10134 18572 10140 18584
rect 10192 18572 10198 18624
rect 10686 18572 10692 18624
rect 10744 18612 10750 18624
rect 11072 18612 11100 18652
rect 11238 18612 11244 18624
rect 10744 18584 11100 18612
rect 11199 18584 11244 18612
rect 10744 18572 10750 18584
rect 11238 18572 11244 18584
rect 11296 18572 11302 18624
rect 11348 18612 11376 18652
rect 12360 18652 12848 18680
rect 12912 18652 13461 18680
rect 11517 18615 11575 18621
rect 11517 18612 11529 18615
rect 11348 18584 11529 18612
rect 11517 18581 11529 18584
rect 11563 18612 11575 18615
rect 12360 18612 12388 18652
rect 11563 18584 12388 18612
rect 11563 18581 11575 18584
rect 11517 18575 11575 18581
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 12912 18612 12940 18652
rect 13449 18649 13461 18652
rect 13495 18649 13507 18683
rect 13814 18680 13820 18692
rect 13775 18652 13820 18680
rect 13449 18643 13507 18649
rect 13814 18640 13820 18652
rect 13872 18640 13878 18692
rect 14200 18680 14228 18711
rect 14550 18708 14556 18720
rect 14608 18708 14614 18760
rect 15930 18708 15936 18760
rect 15988 18748 15994 18760
rect 16393 18751 16451 18757
rect 16393 18748 16405 18751
rect 15988 18720 16405 18748
rect 15988 18708 15994 18720
rect 16393 18717 16405 18720
rect 16439 18717 16451 18751
rect 16393 18711 16451 18717
rect 17218 18708 17224 18760
rect 17276 18748 17282 18760
rect 18156 18757 18184 18788
rect 20438 18776 20444 18828
rect 20496 18816 20502 18828
rect 20496 18788 21312 18816
rect 20496 18776 20502 18788
rect 17681 18751 17739 18757
rect 17681 18748 17693 18751
rect 17276 18720 17693 18748
rect 17276 18708 17282 18720
rect 17681 18717 17693 18720
rect 17727 18717 17739 18751
rect 17681 18711 17739 18717
rect 18141 18751 18199 18757
rect 18141 18717 18153 18751
rect 18187 18748 18199 18751
rect 18230 18748 18236 18760
rect 18187 18720 18236 18748
rect 18187 18717 18199 18720
rect 18141 18711 18199 18717
rect 14829 18683 14887 18689
rect 14829 18680 14841 18683
rect 14200 18652 14841 18680
rect 14829 18649 14841 18652
rect 14875 18649 14887 18683
rect 17696 18680 17724 18711
rect 18230 18708 18236 18720
rect 18288 18708 18294 18760
rect 18417 18751 18475 18757
rect 18417 18717 18429 18751
rect 18463 18717 18475 18751
rect 18782 18748 18788 18760
rect 18743 18720 18788 18748
rect 18417 18711 18475 18717
rect 18432 18680 18460 18711
rect 18782 18708 18788 18720
rect 18840 18708 18846 18760
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 18932 18720 18977 18748
rect 18932 18708 18938 18720
rect 19058 18708 19064 18760
rect 19116 18748 19122 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19116 18720 19257 18748
rect 19116 18708 19122 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19886 18748 19892 18760
rect 19847 18720 19892 18748
rect 19245 18711 19303 18717
rect 19886 18708 19892 18720
rect 19944 18708 19950 18760
rect 20257 18751 20315 18757
rect 20257 18717 20269 18751
rect 20303 18717 20315 18751
rect 20257 18711 20315 18717
rect 17696 18652 18460 18680
rect 20272 18680 20300 18711
rect 20346 18708 20352 18760
rect 20404 18748 20410 18760
rect 20714 18748 20720 18760
rect 20404 18720 20449 18748
rect 20675 18720 20720 18748
rect 20404 18708 20410 18720
rect 20714 18708 20720 18720
rect 20772 18708 20778 18760
rect 21284 18757 21312 18788
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18717 21327 18751
rect 21269 18711 21327 18717
rect 20806 18680 20812 18692
rect 20272 18652 20812 18680
rect 14829 18643 14887 18649
rect 20806 18640 20812 18652
rect 20864 18640 20870 18692
rect 20990 18680 20996 18692
rect 20951 18652 20996 18680
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 13170 18612 13176 18624
rect 12492 18584 12940 18612
rect 13131 18584 13176 18612
rect 12492 18572 12498 18584
rect 13170 18572 13176 18584
rect 13228 18572 13234 18624
rect 17402 18612 17408 18624
rect 17363 18584 17408 18612
rect 17402 18572 17408 18584
rect 17460 18572 17466 18624
rect 18322 18572 18328 18624
rect 18380 18612 18386 18624
rect 18601 18615 18659 18621
rect 18601 18612 18613 18615
rect 18380 18584 18613 18612
rect 18380 18572 18386 18584
rect 18601 18581 18613 18584
rect 18647 18612 18659 18615
rect 18690 18612 18696 18624
rect 18647 18584 18696 18612
rect 18647 18581 18659 18584
rect 18601 18575 18659 18581
rect 18690 18572 18696 18584
rect 18748 18572 18754 18624
rect 21450 18612 21456 18624
rect 21411 18584 21456 18612
rect 21450 18572 21456 18584
rect 21508 18572 21514 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 2590 18368 2596 18420
rect 2648 18408 2654 18420
rect 2777 18411 2835 18417
rect 2777 18408 2789 18411
rect 2648 18380 2789 18408
rect 2648 18368 2654 18380
rect 2777 18377 2789 18380
rect 2823 18377 2835 18411
rect 3602 18408 3608 18420
rect 3563 18380 3608 18408
rect 2777 18371 2835 18377
rect 3602 18368 3608 18380
rect 3660 18368 3666 18420
rect 3973 18411 4031 18417
rect 3973 18377 3985 18411
rect 4019 18377 4031 18411
rect 3973 18371 4031 18377
rect 2685 18343 2743 18349
rect 2685 18309 2697 18343
rect 2731 18340 2743 18343
rect 2866 18340 2872 18352
rect 2731 18312 2872 18340
rect 2731 18309 2743 18312
rect 2685 18303 2743 18309
rect 2866 18300 2872 18312
rect 2924 18300 2930 18352
rect 3513 18343 3571 18349
rect 3513 18309 3525 18343
rect 3559 18340 3571 18343
rect 3988 18340 4016 18371
rect 4062 18368 4068 18420
rect 4120 18408 4126 18420
rect 5261 18411 5319 18417
rect 5261 18408 5273 18411
rect 4120 18380 5273 18408
rect 4120 18368 4126 18380
rect 5261 18377 5273 18380
rect 5307 18377 5319 18411
rect 5810 18408 5816 18420
rect 5771 18380 5816 18408
rect 5261 18371 5319 18377
rect 4430 18340 4436 18352
rect 3559 18312 4016 18340
rect 4391 18312 4436 18340
rect 3559 18309 3571 18312
rect 3513 18303 3571 18309
rect 4430 18300 4436 18312
rect 4488 18300 4494 18352
rect 4706 18300 4712 18352
rect 4764 18340 4770 18352
rect 4893 18343 4951 18349
rect 4893 18340 4905 18343
rect 4764 18312 4905 18340
rect 4764 18300 4770 18312
rect 4893 18309 4905 18312
rect 4939 18309 4951 18343
rect 5074 18340 5080 18352
rect 5035 18312 5080 18340
rect 4893 18303 4951 18309
rect 5074 18300 5080 18312
rect 5132 18300 5138 18352
rect 5276 18340 5304 18371
rect 5810 18368 5816 18380
rect 5868 18368 5874 18420
rect 5902 18368 5908 18420
rect 5960 18408 5966 18420
rect 6365 18411 6423 18417
rect 6365 18408 6377 18411
rect 5960 18380 6377 18408
rect 5960 18368 5966 18380
rect 6365 18377 6377 18380
rect 6411 18377 6423 18411
rect 7190 18408 7196 18420
rect 6365 18371 6423 18377
rect 6757 18380 7052 18408
rect 7151 18380 7196 18408
rect 6757 18340 6785 18380
rect 5276 18312 6785 18340
rect 6825 18343 6883 18349
rect 6825 18309 6837 18343
rect 6871 18340 6883 18343
rect 6914 18340 6920 18352
rect 6871 18312 6920 18340
rect 6871 18309 6883 18312
rect 6825 18303 6883 18309
rect 6914 18300 6920 18312
rect 6972 18300 6978 18352
rect 7024 18340 7052 18380
rect 7190 18368 7196 18380
rect 7248 18368 7254 18420
rect 7282 18368 7288 18420
rect 7340 18408 7346 18420
rect 7650 18408 7656 18420
rect 7340 18380 7656 18408
rect 7340 18368 7346 18380
rect 7650 18368 7656 18380
rect 7708 18408 7714 18420
rect 7745 18411 7803 18417
rect 7745 18408 7757 18411
rect 7708 18380 7757 18408
rect 7708 18368 7714 18380
rect 7745 18377 7757 18380
rect 7791 18377 7803 18411
rect 7745 18371 7803 18377
rect 7926 18368 7932 18420
rect 7984 18368 7990 18420
rect 9769 18411 9827 18417
rect 8036 18380 9720 18408
rect 7944 18340 7972 18368
rect 7024 18312 7972 18340
rect 1670 18272 1676 18284
rect 1631 18244 1676 18272
rect 1670 18232 1676 18244
rect 1728 18232 1734 18284
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18272 2099 18275
rect 4062 18272 4068 18284
rect 2087 18244 4068 18272
rect 2087 18241 2099 18244
rect 2041 18235 2099 18241
rect 4062 18232 4068 18244
rect 4120 18232 4126 18284
rect 4341 18275 4399 18281
rect 4341 18241 4353 18275
rect 4387 18272 4399 18275
rect 5442 18272 5448 18284
rect 4387 18244 5448 18272
rect 4387 18241 4399 18244
rect 4341 18235 4399 18241
rect 2498 18164 2504 18216
rect 2556 18204 2562 18216
rect 2961 18207 3019 18213
rect 2961 18204 2973 18207
rect 2556 18176 2973 18204
rect 2556 18164 2562 18176
rect 2961 18173 2973 18176
rect 3007 18204 3019 18207
rect 3697 18207 3755 18213
rect 3697 18204 3709 18207
rect 3007 18176 3709 18204
rect 3007 18173 3019 18176
rect 2961 18167 3019 18173
rect 3697 18173 3709 18176
rect 3743 18173 3755 18207
rect 3697 18167 3755 18173
rect 566 18096 572 18148
rect 624 18136 630 18148
rect 4540 18136 4568 18244
rect 5442 18232 5448 18244
rect 5500 18232 5506 18284
rect 5644 18244 6684 18272
rect 4617 18207 4675 18213
rect 4617 18173 4629 18207
rect 4663 18204 4675 18207
rect 4798 18204 4804 18216
rect 4663 18176 4804 18204
rect 4663 18173 4675 18176
rect 4617 18167 4675 18173
rect 4798 18164 4804 18176
rect 4856 18164 4862 18216
rect 4890 18164 4896 18216
rect 4948 18204 4954 18216
rect 5166 18204 5172 18216
rect 4948 18176 5172 18204
rect 4948 18164 4954 18176
rect 5166 18164 5172 18176
rect 5224 18164 5230 18216
rect 5258 18164 5264 18216
rect 5316 18204 5322 18216
rect 5644 18213 5672 18244
rect 5629 18207 5687 18213
rect 5316 18176 5580 18204
rect 5316 18164 5322 18176
rect 4706 18136 4712 18148
rect 624 18108 4292 18136
rect 4540 18108 4712 18136
rect 624 18096 630 18108
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 1854 18068 1860 18080
rect 1815 18040 1860 18068
rect 1854 18028 1860 18040
rect 1912 18028 1918 18080
rect 2130 18068 2136 18080
rect 2091 18040 2136 18068
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 2314 18068 2320 18080
rect 2275 18040 2320 18068
rect 2314 18028 2320 18040
rect 2372 18028 2378 18080
rect 2774 18028 2780 18080
rect 2832 18068 2838 18080
rect 3145 18071 3203 18077
rect 3145 18068 3157 18071
rect 2832 18040 3157 18068
rect 2832 18028 2838 18040
rect 3145 18037 3157 18040
rect 3191 18037 3203 18071
rect 4264 18068 4292 18108
rect 4706 18096 4712 18108
rect 4764 18096 4770 18148
rect 5552 18136 5580 18176
rect 5629 18173 5641 18207
rect 5675 18173 5687 18207
rect 5629 18167 5687 18173
rect 5718 18164 5724 18216
rect 5776 18204 5782 18216
rect 6656 18204 6684 18244
rect 6730 18232 6736 18284
rect 6788 18272 6794 18284
rect 6788 18244 6833 18272
rect 6788 18232 6794 18244
rect 7006 18232 7012 18284
rect 7064 18272 7070 18284
rect 7377 18275 7435 18281
rect 7377 18272 7389 18275
rect 7064 18244 7389 18272
rect 7064 18232 7070 18244
rect 7377 18241 7389 18244
rect 7423 18241 7435 18275
rect 7377 18235 7435 18241
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 7837 18275 7895 18281
rect 7837 18272 7849 18275
rect 7524 18244 7849 18272
rect 7524 18232 7530 18244
rect 7837 18241 7849 18244
rect 7883 18241 7895 18275
rect 7837 18235 7895 18241
rect 6822 18204 6828 18216
rect 5776 18176 5821 18204
rect 5920 18176 6316 18204
rect 6656 18176 6828 18204
rect 5776 18164 5782 18176
rect 5920 18136 5948 18176
rect 5552 18108 5948 18136
rect 5994 18096 6000 18148
rect 6052 18136 6058 18148
rect 6181 18139 6239 18145
rect 6181 18136 6193 18139
rect 6052 18108 6193 18136
rect 6052 18096 6058 18108
rect 6181 18105 6193 18108
rect 6227 18105 6239 18139
rect 6288 18136 6316 18176
rect 6822 18164 6828 18176
rect 6880 18204 6886 18216
rect 6917 18207 6975 18213
rect 6917 18204 6929 18207
rect 6880 18176 6929 18204
rect 6880 18164 6886 18176
rect 6917 18173 6929 18176
rect 6963 18173 6975 18207
rect 7650 18204 7656 18216
rect 7611 18176 7656 18204
rect 6917 18167 6975 18173
rect 7650 18164 7656 18176
rect 7708 18164 7714 18216
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 8036 18204 8064 18380
rect 8294 18300 8300 18352
rect 8352 18340 8358 18352
rect 8352 18312 8616 18340
rect 8352 18300 8358 18312
rect 8110 18232 8116 18284
rect 8168 18272 8174 18284
rect 8588 18281 8616 18312
rect 8754 18300 8760 18352
rect 8812 18340 8818 18352
rect 9030 18340 9036 18352
rect 8812 18312 9036 18340
rect 8812 18300 8818 18312
rect 9030 18300 9036 18312
rect 9088 18300 9094 18352
rect 9692 18340 9720 18380
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 9950 18408 9956 18420
rect 9815 18380 9956 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 9950 18368 9956 18380
rect 10008 18368 10014 18420
rect 10137 18411 10195 18417
rect 10137 18377 10149 18411
rect 10183 18408 10195 18411
rect 10502 18408 10508 18420
rect 10183 18380 10508 18408
rect 10183 18377 10195 18380
rect 10137 18371 10195 18377
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 10597 18411 10655 18417
rect 10597 18377 10609 18411
rect 10643 18408 10655 18411
rect 10870 18408 10876 18420
rect 10643 18380 10876 18408
rect 10643 18377 10655 18380
rect 10597 18371 10655 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 12434 18408 12440 18420
rect 11020 18380 11065 18408
rect 11164 18380 12440 18408
rect 11020 18368 11026 18380
rect 11164 18340 11192 18380
rect 12434 18368 12440 18380
rect 12492 18368 12498 18420
rect 12710 18408 12716 18420
rect 12671 18380 12716 18408
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 12894 18408 12900 18420
rect 12855 18380 12900 18408
rect 12894 18368 12900 18380
rect 12952 18368 12958 18420
rect 13262 18408 13268 18420
rect 13223 18380 13268 18408
rect 13262 18368 13268 18380
rect 13320 18368 13326 18420
rect 13538 18368 13544 18420
rect 13596 18368 13602 18420
rect 13725 18411 13783 18417
rect 13725 18377 13737 18411
rect 13771 18408 13783 18411
rect 14550 18408 14556 18420
rect 13771 18380 14556 18408
rect 13771 18377 13783 18380
rect 13725 18371 13783 18377
rect 14550 18368 14556 18380
rect 14608 18368 14614 18420
rect 14642 18368 14648 18420
rect 14700 18408 14706 18420
rect 14918 18408 14924 18420
rect 14700 18380 14745 18408
rect 14879 18380 14924 18408
rect 14700 18368 14706 18380
rect 14918 18368 14924 18380
rect 14976 18368 14982 18420
rect 15194 18408 15200 18420
rect 15155 18380 15200 18408
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15930 18408 15936 18420
rect 15344 18380 15389 18408
rect 15891 18380 15936 18408
rect 15344 18368 15350 18380
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16390 18368 16396 18420
rect 16448 18408 16454 18420
rect 17586 18408 17592 18420
rect 16448 18380 17592 18408
rect 16448 18368 16454 18380
rect 17586 18368 17592 18380
rect 17644 18368 17650 18420
rect 18230 18408 18236 18420
rect 18191 18380 18236 18408
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 18506 18408 18512 18420
rect 18467 18380 18512 18408
rect 18506 18368 18512 18380
rect 18564 18368 18570 18420
rect 19429 18411 19487 18417
rect 19429 18377 19441 18411
rect 19475 18408 19487 18411
rect 19518 18408 19524 18420
rect 19475 18380 19524 18408
rect 19475 18377 19487 18380
rect 19429 18371 19487 18377
rect 19518 18368 19524 18380
rect 19576 18368 19582 18420
rect 20714 18368 20720 18420
rect 20772 18408 20778 18420
rect 21085 18411 21143 18417
rect 21085 18408 21097 18411
rect 20772 18380 21097 18408
rect 20772 18368 20778 18380
rect 21085 18377 21097 18380
rect 21131 18377 21143 18411
rect 21085 18371 21143 18377
rect 9692 18312 11192 18340
rect 11422 18300 11428 18352
rect 11480 18340 11486 18352
rect 11885 18343 11943 18349
rect 11885 18340 11897 18343
rect 11480 18312 11897 18340
rect 11480 18300 11486 18312
rect 11885 18309 11897 18312
rect 11931 18309 11943 18343
rect 12526 18340 12532 18352
rect 12487 18312 12532 18340
rect 11885 18303 11943 18309
rect 12526 18300 12532 18312
rect 12584 18300 12590 18352
rect 13556 18340 13584 18368
rect 13188 18312 13584 18340
rect 14093 18343 14151 18349
rect 8573 18275 8631 18281
rect 8168 18244 8524 18272
rect 8168 18232 8174 18244
rect 7800 18176 8064 18204
rect 7800 18164 7806 18176
rect 8294 18164 8300 18216
rect 8352 18204 8358 18216
rect 8496 18204 8524 18244
rect 8573 18241 8585 18275
rect 8619 18272 8631 18275
rect 8662 18272 8668 18284
rect 8619 18244 8668 18272
rect 8619 18241 8631 18244
rect 8573 18235 8631 18241
rect 8662 18232 8668 18244
rect 8720 18232 8726 18284
rect 9393 18275 9451 18281
rect 9393 18241 9405 18275
rect 9439 18241 9451 18275
rect 9393 18235 9451 18241
rect 9493 18275 9551 18281
rect 9493 18241 9505 18275
rect 9539 18272 9551 18275
rect 9582 18272 9588 18284
rect 9539 18244 9588 18272
rect 9539 18241 9551 18244
rect 9493 18235 9551 18241
rect 8754 18204 8760 18216
rect 8352 18176 8397 18204
rect 8496 18176 8760 18204
rect 8352 18164 8358 18176
rect 8754 18164 8760 18176
rect 8812 18164 8818 18216
rect 9048 18176 9260 18204
rect 8110 18136 8116 18148
rect 6288 18108 8116 18136
rect 6181 18099 6239 18105
rect 8110 18096 8116 18108
rect 8168 18096 8174 18148
rect 8205 18139 8263 18145
rect 8205 18105 8217 18139
rect 8251 18136 8263 18139
rect 9048 18136 9076 18176
rect 8251 18108 9076 18136
rect 9232 18136 9260 18176
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 9416 18204 9444 18235
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 13081 18275 13139 18281
rect 13081 18272 13093 18275
rect 10695 18244 13093 18272
rect 9364 18176 9444 18204
rect 10229 18207 10287 18213
rect 9364 18164 9370 18176
rect 10229 18173 10241 18207
rect 10275 18173 10287 18207
rect 10229 18167 10287 18173
rect 10244 18136 10272 18167
rect 10318 18164 10324 18216
rect 10376 18204 10382 18216
rect 10376 18176 10421 18204
rect 10376 18164 10382 18176
rect 10502 18164 10508 18216
rect 10560 18204 10566 18216
rect 10695 18204 10723 18244
rect 13081 18241 13093 18244
rect 13127 18241 13139 18275
rect 13081 18235 13139 18241
rect 11054 18204 11060 18216
rect 10560 18176 10723 18204
rect 11015 18176 11060 18204
rect 10560 18164 10566 18176
rect 11054 18164 11060 18176
rect 11112 18164 11118 18216
rect 11149 18207 11207 18213
rect 11149 18173 11161 18207
rect 11195 18173 11207 18207
rect 11974 18204 11980 18216
rect 11935 18176 11980 18204
rect 11149 18167 11207 18173
rect 9232 18108 10272 18136
rect 10336 18136 10364 18164
rect 11164 18136 11192 18167
rect 11974 18164 11980 18176
rect 12032 18164 12038 18216
rect 12069 18207 12127 18213
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 10336 18108 11192 18136
rect 8251 18105 8263 18108
rect 8205 18099 8263 18105
rect 11238 18096 11244 18148
rect 11296 18136 11302 18148
rect 12084 18136 12112 18167
rect 11296 18108 12112 18136
rect 11296 18096 11302 18108
rect 12342 18096 12348 18148
rect 12400 18136 12406 18148
rect 13188 18136 13216 18312
rect 14093 18309 14105 18343
rect 14139 18340 14151 18343
rect 14274 18340 14280 18352
rect 14139 18312 14280 18340
rect 14139 18309 14151 18312
rect 14093 18303 14151 18309
rect 14274 18300 14280 18312
rect 14332 18300 14338 18352
rect 14366 18300 14372 18352
rect 14424 18340 14430 18352
rect 14734 18340 14740 18352
rect 14424 18312 14469 18340
rect 14695 18312 14740 18340
rect 14424 18300 14430 18312
rect 14734 18300 14740 18312
rect 14792 18300 14798 18352
rect 15378 18300 15384 18352
rect 15436 18340 15442 18352
rect 15473 18343 15531 18349
rect 15473 18340 15485 18343
rect 15436 18312 15485 18340
rect 15436 18300 15442 18312
rect 15473 18309 15485 18312
rect 15519 18309 15531 18343
rect 15473 18303 15531 18309
rect 18141 18343 18199 18349
rect 18141 18309 18153 18343
rect 18187 18340 18199 18343
rect 19794 18340 19800 18352
rect 18187 18312 19472 18340
rect 19755 18312 19800 18340
rect 18187 18309 18199 18312
rect 18141 18303 18199 18309
rect 13538 18272 13544 18284
rect 13499 18244 13544 18272
rect 13538 18232 13544 18244
rect 13596 18232 13602 18284
rect 15749 18275 15807 18281
rect 15749 18241 15761 18275
rect 15795 18272 15807 18275
rect 16942 18272 16948 18284
rect 15795 18244 16948 18272
rect 15795 18241 15807 18244
rect 15749 18235 15807 18241
rect 16942 18232 16948 18244
rect 17000 18232 17006 18284
rect 17402 18272 17408 18284
rect 17363 18244 17408 18272
rect 17402 18232 17408 18244
rect 17460 18232 17466 18284
rect 18690 18272 18696 18284
rect 18651 18244 18696 18272
rect 18690 18232 18696 18244
rect 18748 18232 18754 18284
rect 19058 18232 19064 18284
rect 19116 18272 19122 18284
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 19116 18244 19165 18272
rect 19116 18232 19122 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19153 18235 19211 18241
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18241 19303 18275
rect 19444 18272 19472 18312
rect 19794 18300 19800 18312
rect 19852 18300 19858 18352
rect 19705 18275 19763 18281
rect 19705 18272 19717 18275
rect 19444 18244 19717 18272
rect 19245 18235 19303 18241
rect 19705 18241 19717 18244
rect 19751 18272 19763 18275
rect 20254 18272 20260 18284
rect 19751 18244 20260 18272
rect 19751 18241 19763 18244
rect 19705 18235 19763 18241
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14550 18204 14556 18216
rect 14323 18176 14556 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 14550 18164 14556 18176
rect 14608 18164 14614 18216
rect 18782 18164 18788 18216
rect 18840 18204 18846 18216
rect 19260 18204 19288 18235
rect 20254 18232 20260 18244
rect 20312 18232 20318 18284
rect 18840 18176 19288 18204
rect 18840 18164 18846 18176
rect 12400 18108 13216 18136
rect 12400 18096 12406 18108
rect 13446 18096 13452 18148
rect 13504 18136 13510 18148
rect 16390 18136 16396 18148
rect 13504 18108 16396 18136
rect 13504 18096 13510 18108
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 17589 18139 17647 18145
rect 17589 18105 17601 18139
rect 17635 18136 17647 18139
rect 21358 18136 21364 18148
rect 17635 18108 21364 18136
rect 17635 18105 17647 18108
rect 17589 18099 17647 18105
rect 21358 18096 21364 18108
rect 21416 18096 21422 18148
rect 4890 18068 4896 18080
rect 4264 18040 4896 18068
rect 3145 18031 3203 18037
rect 4890 18028 4896 18040
rect 4948 18028 4954 18080
rect 5442 18028 5448 18080
rect 5500 18068 5506 18080
rect 9217 18071 9275 18077
rect 9217 18068 9229 18071
rect 5500 18040 9229 18068
rect 5500 18028 5506 18040
rect 9217 18037 9229 18040
rect 9263 18037 9275 18071
rect 9217 18031 9275 18037
rect 9677 18071 9735 18077
rect 9677 18037 9689 18071
rect 9723 18068 9735 18071
rect 9858 18068 9864 18080
rect 9723 18040 9864 18068
rect 9723 18037 9735 18040
rect 9677 18031 9735 18037
rect 9858 18028 9864 18040
rect 9916 18068 9922 18080
rect 10962 18068 10968 18080
rect 9916 18040 10968 18068
rect 9916 18028 9922 18040
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11517 18071 11575 18077
rect 11517 18068 11529 18071
rect 11112 18040 11529 18068
rect 11112 18028 11118 18040
rect 11517 18037 11529 18040
rect 11563 18037 11575 18071
rect 11517 18031 11575 18037
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 12437 18071 12495 18077
rect 12437 18068 12449 18071
rect 12032 18040 12449 18068
rect 12032 18028 12038 18040
rect 12437 18037 12449 18040
rect 12483 18037 12495 18071
rect 12437 18031 12495 18037
rect 13909 18071 13967 18077
rect 13909 18037 13921 18071
rect 13955 18068 13967 18071
rect 14274 18068 14280 18080
rect 13955 18040 14280 18068
rect 13955 18037 13967 18040
rect 13909 18031 13967 18037
rect 14274 18028 14280 18040
rect 14332 18068 14338 18080
rect 15010 18068 15016 18080
rect 14332 18040 15016 18068
rect 14332 18028 14338 18040
rect 15010 18028 15016 18040
rect 15068 18028 15074 18080
rect 18782 18068 18788 18080
rect 18743 18040 18788 18068
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 18966 18068 18972 18080
rect 18927 18040 18972 18068
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 19518 18068 19524 18080
rect 19479 18040 19524 18068
rect 19518 18028 19524 18040
rect 19576 18028 19582 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 1765 17867 1823 17873
rect 1765 17864 1777 17867
rect 1728 17836 1777 17864
rect 1728 17824 1734 17836
rect 1765 17833 1777 17836
rect 1811 17833 1823 17867
rect 1765 17827 1823 17833
rect 2038 17824 2044 17876
rect 2096 17864 2102 17876
rect 3326 17864 3332 17876
rect 2096 17836 3332 17864
rect 2096 17824 2102 17836
rect 3326 17824 3332 17836
rect 3384 17824 3390 17876
rect 3789 17867 3847 17873
rect 3789 17833 3801 17867
rect 3835 17864 3847 17867
rect 3878 17864 3884 17876
rect 3835 17836 3884 17864
rect 3835 17833 3847 17836
rect 3789 17827 3847 17833
rect 3878 17824 3884 17836
rect 3936 17824 3942 17876
rect 4062 17824 4068 17876
rect 4120 17864 4126 17876
rect 4893 17867 4951 17873
rect 4893 17864 4905 17867
rect 4120 17836 4200 17864
rect 4120 17824 4126 17836
rect 2777 17799 2835 17805
rect 2777 17765 2789 17799
rect 2823 17765 2835 17799
rect 2777 17759 2835 17765
rect 1762 17688 1768 17740
rect 1820 17728 1826 17740
rect 2133 17731 2191 17737
rect 2133 17728 2145 17731
rect 1820 17700 2145 17728
rect 1820 17688 1826 17700
rect 2133 17697 2145 17700
rect 2179 17697 2191 17731
rect 2682 17728 2688 17740
rect 2133 17691 2191 17697
rect 2240 17700 2688 17728
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17629 1731 17663
rect 1673 17623 1731 17629
rect 1949 17663 2007 17669
rect 1949 17629 1961 17663
rect 1995 17660 2007 17663
rect 2240 17660 2268 17700
rect 2682 17688 2688 17700
rect 2740 17688 2746 17740
rect 2792 17728 2820 17759
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 4172 17796 4200 17836
rect 4724 17836 4905 17864
rect 4724 17796 4752 17836
rect 4893 17833 4905 17836
rect 4939 17833 4951 17867
rect 4893 17827 4951 17833
rect 5350 17824 5356 17876
rect 5408 17824 5414 17876
rect 6270 17864 6276 17876
rect 5644 17836 6276 17864
rect 2924 17768 2969 17796
rect 4172 17768 4752 17796
rect 4801 17799 4859 17805
rect 2924 17756 2930 17768
rect 4801 17765 4813 17799
rect 4847 17796 4859 17799
rect 5368 17796 5396 17824
rect 5644 17796 5672 17836
rect 6270 17824 6276 17836
rect 6328 17824 6334 17876
rect 6914 17864 6920 17876
rect 6875 17836 6920 17864
rect 6914 17824 6920 17836
rect 6972 17824 6978 17876
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 7929 17867 7987 17873
rect 7929 17864 7941 17867
rect 7892 17836 7941 17864
rect 7892 17824 7898 17836
rect 7929 17833 7941 17836
rect 7975 17833 7987 17867
rect 7929 17827 7987 17833
rect 8294 17824 8300 17876
rect 8352 17864 8358 17876
rect 8478 17864 8484 17876
rect 8352 17836 8484 17864
rect 8352 17824 8358 17836
rect 8478 17824 8484 17836
rect 8536 17824 8542 17876
rect 9858 17864 9864 17876
rect 8680 17836 9864 17864
rect 8570 17796 8576 17808
rect 4847 17768 5304 17796
rect 5368 17768 5672 17796
rect 7576 17768 8576 17796
rect 4847 17765 4859 17768
rect 4801 17759 4859 17765
rect 3513 17731 3571 17737
rect 2792 17700 3464 17728
rect 1995 17632 2268 17660
rect 1995 17629 2007 17632
rect 1949 17623 2007 17629
rect 1688 17592 1716 17623
rect 2314 17620 2320 17672
rect 2372 17660 2378 17672
rect 2409 17663 2467 17669
rect 2409 17660 2421 17663
rect 2372 17632 2421 17660
rect 2372 17620 2378 17632
rect 2409 17629 2421 17632
rect 2455 17629 2467 17663
rect 2409 17623 2467 17629
rect 3326 17620 3332 17672
rect 3384 17620 3390 17672
rect 3436 17660 3464 17700
rect 3513 17697 3525 17731
rect 3559 17728 3571 17731
rect 3970 17728 3976 17740
rect 3559 17700 3976 17728
rect 3559 17697 3571 17700
rect 3513 17691 3571 17697
rect 3970 17688 3976 17700
rect 4028 17688 4034 17740
rect 4430 17728 4436 17740
rect 4391 17700 4436 17728
rect 4430 17688 4436 17700
rect 4488 17688 4494 17740
rect 4249 17663 4307 17669
rect 4249 17660 4261 17663
rect 3436 17632 4261 17660
rect 4249 17629 4261 17632
rect 4295 17629 4307 17663
rect 4614 17660 4620 17672
rect 4575 17632 4620 17660
rect 4249 17623 4307 17629
rect 4614 17620 4620 17632
rect 4672 17620 4678 17672
rect 5074 17660 5080 17672
rect 5035 17632 5080 17660
rect 5074 17620 5080 17632
rect 5132 17620 5138 17672
rect 2038 17592 2044 17604
rect 1688 17564 2044 17592
rect 2038 17552 2044 17564
rect 2096 17552 2102 17604
rect 2774 17592 2780 17604
rect 2332 17564 2780 17592
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2332 17533 2360 17564
rect 2774 17552 2780 17564
rect 2832 17552 2838 17604
rect 3237 17595 3295 17601
rect 3237 17561 3249 17595
rect 3283 17561 3295 17595
rect 3344 17592 3372 17620
rect 5276 17592 5304 17768
rect 5350 17688 5356 17740
rect 5408 17728 5414 17740
rect 6457 17731 6515 17737
rect 6457 17728 6469 17731
rect 5408 17700 5453 17728
rect 5736 17700 6469 17728
rect 5408 17688 5414 17700
rect 5442 17660 5448 17672
rect 5403 17632 5448 17660
rect 5442 17620 5448 17632
rect 5500 17620 5506 17672
rect 5626 17620 5632 17672
rect 5684 17660 5690 17672
rect 5736 17660 5764 17700
rect 6457 17697 6469 17700
rect 6503 17697 6515 17731
rect 6457 17691 6515 17697
rect 6641 17731 6699 17737
rect 6641 17697 6653 17731
rect 6687 17728 6699 17731
rect 6822 17728 6828 17740
rect 6687 17700 6828 17728
rect 6687 17697 6699 17700
rect 6641 17691 6699 17697
rect 6822 17688 6828 17700
rect 6880 17688 6886 17740
rect 7576 17737 7604 17768
rect 8570 17756 8576 17768
rect 8628 17756 8634 17808
rect 7561 17731 7619 17737
rect 7561 17697 7573 17731
rect 7607 17697 7619 17731
rect 7742 17728 7748 17740
rect 7703 17700 7748 17728
rect 7561 17691 7619 17697
rect 7742 17688 7748 17700
rect 7800 17728 7806 17740
rect 7926 17728 7932 17740
rect 7800 17700 7932 17728
rect 7800 17688 7806 17700
rect 7926 17688 7932 17700
rect 7984 17728 7990 17740
rect 8389 17731 8447 17737
rect 8389 17728 8401 17731
rect 7984 17700 8401 17728
rect 7984 17688 7990 17700
rect 8389 17697 8401 17700
rect 8435 17697 8447 17731
rect 8389 17691 8447 17697
rect 8478 17688 8484 17740
rect 8536 17728 8542 17740
rect 8536 17700 8581 17728
rect 8536 17688 8542 17700
rect 7006 17660 7012 17672
rect 5684 17632 5764 17660
rect 6104 17632 7012 17660
rect 5684 17620 5690 17632
rect 6104 17592 6132 17632
rect 7006 17620 7012 17632
rect 7064 17620 7070 17672
rect 7282 17660 7288 17672
rect 7243 17632 7288 17660
rect 7282 17620 7288 17632
rect 7340 17620 7346 17672
rect 8680 17660 8708 17836
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 10042 17824 10048 17876
rect 10100 17864 10106 17876
rect 10597 17867 10655 17873
rect 10597 17864 10609 17867
rect 10100 17836 10609 17864
rect 10100 17824 10106 17836
rect 10597 17833 10609 17836
rect 10643 17833 10655 17867
rect 10597 17827 10655 17833
rect 10686 17824 10692 17876
rect 10744 17864 10750 17876
rect 11793 17867 11851 17873
rect 11793 17864 11805 17867
rect 10744 17836 11805 17864
rect 10744 17824 10750 17836
rect 11793 17833 11805 17836
rect 11839 17833 11851 17867
rect 11793 17827 11851 17833
rect 11882 17824 11888 17876
rect 11940 17864 11946 17876
rect 13354 17864 13360 17876
rect 11940 17836 13360 17864
rect 11940 17824 11946 17836
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 13449 17867 13507 17873
rect 13449 17833 13461 17867
rect 13495 17864 13507 17867
rect 13538 17864 13544 17876
rect 13495 17836 13544 17864
rect 13495 17833 13507 17836
rect 13449 17827 13507 17833
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 16669 17867 16727 17873
rect 13648 17836 16620 17864
rect 10134 17756 10140 17808
rect 10192 17796 10198 17808
rect 10192 17768 11284 17796
rect 10192 17756 10198 17768
rect 9950 17688 9956 17740
rect 10008 17728 10014 17740
rect 10870 17728 10876 17740
rect 10008 17700 10876 17728
rect 10008 17688 10014 17700
rect 10870 17688 10876 17700
rect 10928 17688 10934 17740
rect 11054 17728 11060 17740
rect 11015 17700 11060 17728
rect 11054 17688 11060 17700
rect 11112 17688 11118 17740
rect 11149 17731 11207 17737
rect 11149 17697 11161 17731
rect 11195 17697 11207 17731
rect 11256 17728 11284 17768
rect 11698 17756 11704 17808
rect 11756 17796 11762 17808
rect 12437 17799 12495 17805
rect 12437 17796 12449 17799
rect 11756 17768 12449 17796
rect 11756 17756 11762 17768
rect 12437 17765 12449 17768
rect 12483 17765 12495 17799
rect 12437 17759 12495 17765
rect 12986 17756 12992 17808
rect 13044 17796 13050 17808
rect 13648 17796 13676 17836
rect 13814 17796 13820 17808
rect 13044 17768 13676 17796
rect 13775 17768 13820 17796
rect 13044 17756 13050 17768
rect 13814 17756 13820 17768
rect 13872 17756 13878 17808
rect 16592 17796 16620 17836
rect 16669 17833 16681 17867
rect 16715 17864 16727 17867
rect 17402 17864 17408 17876
rect 16715 17836 17408 17864
rect 16715 17833 16727 17836
rect 16669 17827 16727 17833
rect 17402 17824 17408 17836
rect 17460 17824 17466 17876
rect 19058 17824 19064 17876
rect 19116 17864 19122 17876
rect 19245 17867 19303 17873
rect 19245 17864 19257 17867
rect 19116 17836 19257 17864
rect 19116 17824 19122 17836
rect 19245 17833 19257 17836
rect 19291 17833 19303 17867
rect 19245 17827 19303 17833
rect 19521 17867 19579 17873
rect 19521 17833 19533 17867
rect 19567 17864 19579 17867
rect 19610 17864 19616 17876
rect 19567 17836 19616 17864
rect 19567 17833 19579 17836
rect 19521 17827 19579 17833
rect 19610 17824 19616 17836
rect 19668 17824 19674 17876
rect 20070 17864 20076 17876
rect 19720 17836 20076 17864
rect 18046 17796 18052 17808
rect 16592 17768 18052 17796
rect 18046 17756 18052 17768
rect 18104 17756 18110 17808
rect 11977 17731 12035 17737
rect 11977 17728 11989 17731
rect 11256 17700 11989 17728
rect 11149 17691 11207 17697
rect 11977 17697 11989 17700
rect 12023 17697 12035 17731
rect 12897 17731 12955 17737
rect 12897 17728 12909 17731
rect 11977 17691 12035 17697
rect 12452 17700 12909 17728
rect 7585 17632 8708 17660
rect 8941 17663 8999 17669
rect 3344 17564 5120 17592
rect 5276 17564 6132 17592
rect 3237 17555 3295 17561
rect 2317 17527 2375 17533
rect 2317 17493 2329 17527
rect 2363 17493 2375 17527
rect 2317 17487 2375 17493
rect 2590 17484 2596 17536
rect 2648 17524 2654 17536
rect 3252 17524 3280 17555
rect 5092 17536 5120 17564
rect 6270 17552 6276 17604
rect 6328 17592 6334 17604
rect 7585 17592 7613 17632
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9490 17660 9496 17672
rect 8987 17632 9496 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9490 17620 9496 17632
rect 9548 17620 9554 17672
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 11164 17660 11192 17691
rect 10376 17632 11192 17660
rect 10376 17620 10382 17632
rect 11238 17620 11244 17672
rect 11296 17620 11302 17672
rect 11422 17620 11428 17672
rect 11480 17660 11486 17672
rect 11609 17663 11667 17669
rect 11609 17660 11621 17663
rect 11480 17632 11621 17660
rect 11480 17620 11486 17632
rect 11609 17629 11621 17632
rect 11655 17629 11667 17663
rect 11609 17623 11667 17629
rect 6328 17564 7613 17592
rect 6328 17552 6334 17564
rect 2648 17496 3280 17524
rect 3329 17527 3387 17533
rect 2648 17484 2654 17496
rect 3329 17493 3341 17527
rect 3375 17524 3387 17527
rect 3970 17524 3976 17536
rect 3375 17496 3976 17524
rect 3375 17493 3387 17496
rect 3329 17487 3387 17493
rect 3970 17484 3976 17496
rect 4028 17484 4034 17536
rect 4154 17524 4160 17536
rect 4115 17496 4160 17524
rect 4154 17484 4160 17496
rect 4212 17484 4218 17536
rect 5074 17484 5080 17536
rect 5132 17484 5138 17536
rect 5537 17527 5595 17533
rect 5537 17493 5549 17527
rect 5583 17524 5595 17527
rect 5718 17524 5724 17536
rect 5583 17496 5724 17524
rect 5583 17493 5595 17496
rect 5537 17487 5595 17493
rect 5718 17484 5724 17496
rect 5776 17484 5782 17536
rect 5902 17524 5908 17536
rect 5863 17496 5908 17524
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6380 17533 6408 17564
rect 7650 17552 7656 17604
rect 7708 17592 7714 17604
rect 9186 17595 9244 17601
rect 9186 17592 9198 17595
rect 7708 17564 9198 17592
rect 7708 17552 7714 17564
rect 9186 17561 9198 17564
rect 9232 17592 9244 17595
rect 10870 17592 10876 17604
rect 9232 17564 10876 17592
rect 9232 17561 9244 17564
rect 9186 17555 9244 17561
rect 10870 17552 10876 17564
rect 10928 17592 10934 17604
rect 11256 17592 11284 17620
rect 10928 17564 11284 17592
rect 11440 17564 12296 17592
rect 10928 17552 10934 17564
rect 6365 17527 6423 17533
rect 6052 17496 6097 17524
rect 6052 17484 6058 17496
rect 6365 17493 6377 17527
rect 6411 17493 6423 17527
rect 6365 17487 6423 17493
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 7377 17527 7435 17533
rect 7377 17524 7389 17527
rect 7340 17496 7389 17524
rect 7340 17484 7346 17496
rect 7377 17493 7389 17496
rect 7423 17493 7435 17527
rect 7377 17487 7435 17493
rect 7742 17484 7748 17536
rect 7800 17524 7806 17536
rect 8297 17527 8355 17533
rect 8297 17524 8309 17527
rect 7800 17496 8309 17524
rect 7800 17484 7806 17496
rect 8297 17493 8309 17496
rect 8343 17493 8355 17527
rect 10318 17524 10324 17536
rect 10279 17496 10324 17524
rect 8297 17487 8355 17493
rect 10318 17484 10324 17496
rect 10376 17484 10382 17536
rect 10502 17524 10508 17536
rect 10463 17496 10508 17524
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 10686 17484 10692 17536
rect 10744 17524 10750 17536
rect 11440 17533 11468 17564
rect 10965 17527 11023 17533
rect 10965 17524 10977 17527
rect 10744 17496 10977 17524
rect 10744 17484 10750 17496
rect 10965 17493 10977 17496
rect 11011 17524 11023 17527
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 11011 17496 11437 17524
rect 11011 17493 11023 17496
rect 10965 17487 11023 17493
rect 11425 17493 11437 17496
rect 11471 17493 11483 17527
rect 12158 17524 12164 17536
rect 12119 17496 12164 17524
rect 11425 17487 11483 17493
rect 12158 17484 12164 17496
rect 12216 17484 12222 17536
rect 12268 17524 12296 17564
rect 12342 17552 12348 17604
rect 12400 17592 12406 17604
rect 12452 17592 12480 17700
rect 12897 17697 12909 17700
rect 12943 17728 12955 17731
rect 15749 17731 15807 17737
rect 12943 17700 14228 17728
rect 12943 17697 12955 17700
rect 12897 17691 12955 17697
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17660 12679 17663
rect 13722 17660 13728 17672
rect 12667 17632 13728 17660
rect 12667 17629 12679 17632
rect 12621 17623 12679 17629
rect 13722 17620 13728 17632
rect 13780 17660 13786 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13780 17632 14105 17660
rect 13780 17620 13786 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14200 17660 14228 17700
rect 15749 17697 15761 17731
rect 15795 17728 15807 17731
rect 16022 17728 16028 17740
rect 15795 17700 16028 17728
rect 15795 17697 15807 17700
rect 15749 17691 15807 17697
rect 16022 17688 16028 17700
rect 16080 17688 16086 17740
rect 16850 17728 16856 17740
rect 16811 17700 16856 17728
rect 16850 17688 16856 17700
rect 16908 17688 16914 17740
rect 19610 17728 19616 17740
rect 19444 17700 19616 17728
rect 14349 17663 14407 17669
rect 14349 17660 14361 17663
rect 14200 17632 14361 17660
rect 14093 17623 14151 17629
rect 14349 17629 14361 17632
rect 14395 17629 14407 17663
rect 14349 17623 14407 17629
rect 16485 17663 16543 17669
rect 16485 17629 16497 17663
rect 16531 17660 16543 17663
rect 17034 17660 17040 17672
rect 16531 17632 17040 17660
rect 16531 17629 16543 17632
rect 16485 17623 16543 17629
rect 17034 17620 17040 17632
rect 17092 17620 17098 17672
rect 18690 17620 18696 17672
rect 18748 17660 18754 17672
rect 19058 17660 19064 17672
rect 18748 17632 19064 17660
rect 18748 17620 18754 17632
rect 19058 17620 19064 17632
rect 19116 17620 19122 17672
rect 19444 17669 19472 17700
rect 19610 17688 19616 17700
rect 19668 17728 19674 17740
rect 19720 17728 19748 17836
rect 20070 17824 20076 17836
rect 20128 17824 20134 17876
rect 20257 17867 20315 17873
rect 20257 17833 20269 17867
rect 20303 17864 20315 17867
rect 20438 17864 20444 17876
rect 20303 17836 20444 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 20438 17824 20444 17836
rect 20496 17824 20502 17876
rect 19981 17799 20039 17805
rect 19981 17765 19993 17799
rect 20027 17796 20039 17799
rect 21266 17796 21272 17808
rect 20027 17768 21272 17796
rect 20027 17765 20039 17768
rect 19981 17759 20039 17765
rect 21266 17756 21272 17768
rect 21324 17756 21330 17808
rect 19668 17700 19748 17728
rect 19668 17688 19674 17700
rect 19429 17663 19487 17669
rect 19429 17629 19441 17663
rect 19475 17629 19487 17663
rect 19702 17660 19708 17672
rect 19663 17632 19708 17660
rect 19429 17623 19487 17629
rect 19702 17620 19708 17632
rect 19760 17620 19766 17672
rect 19794 17620 19800 17672
rect 19852 17660 19858 17672
rect 20070 17660 20076 17672
rect 19852 17632 19897 17660
rect 20031 17632 20076 17660
rect 19852 17620 19858 17632
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20346 17660 20352 17672
rect 20307 17632 20352 17660
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20714 17660 20720 17672
rect 20675 17632 20720 17660
rect 20714 17620 20720 17632
rect 20772 17620 20778 17672
rect 21082 17620 21088 17672
rect 21140 17660 21146 17672
rect 21269 17663 21327 17669
rect 21269 17660 21281 17663
rect 21140 17632 21281 17660
rect 21140 17620 21146 17632
rect 21269 17629 21281 17632
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 12400 17564 12480 17592
rect 12989 17595 13047 17601
rect 12400 17552 12406 17564
rect 12989 17561 13001 17595
rect 13035 17592 13047 17595
rect 13814 17592 13820 17604
rect 13035 17564 13820 17592
rect 13035 17561 13047 17564
rect 12989 17555 13047 17561
rect 13814 17552 13820 17564
rect 13872 17552 13878 17604
rect 16206 17552 16212 17604
rect 16264 17592 16270 17604
rect 16264 17564 20852 17592
rect 16264 17552 16270 17564
rect 12526 17524 12532 17536
rect 12268 17496 12532 17524
rect 12526 17484 12532 17496
rect 12584 17484 12590 17536
rect 13078 17484 13084 17536
rect 13136 17524 13142 17536
rect 13136 17496 13181 17524
rect 13136 17484 13142 17496
rect 13262 17484 13268 17536
rect 13320 17524 13326 17536
rect 13541 17527 13599 17533
rect 13541 17524 13553 17527
rect 13320 17496 13553 17524
rect 13320 17484 13326 17496
rect 13541 17493 13553 17496
rect 13587 17493 13599 17527
rect 13541 17487 13599 17493
rect 15102 17484 15108 17536
rect 15160 17524 15166 17536
rect 15473 17527 15531 17533
rect 15473 17524 15485 17527
rect 15160 17496 15485 17524
rect 15160 17484 15166 17496
rect 15473 17493 15485 17496
rect 15519 17493 15531 17527
rect 15473 17487 15531 17493
rect 15562 17484 15568 17536
rect 15620 17524 15626 17536
rect 15841 17527 15899 17533
rect 15841 17524 15853 17527
rect 15620 17496 15853 17524
rect 15620 17484 15626 17496
rect 15841 17493 15853 17496
rect 15887 17493 15899 17527
rect 15841 17487 15899 17493
rect 15930 17484 15936 17536
rect 15988 17524 15994 17536
rect 16298 17524 16304 17536
rect 15988 17496 16033 17524
rect 16259 17496 16304 17524
rect 15988 17484 15994 17496
rect 16298 17484 16304 17496
rect 16356 17484 16362 17536
rect 18138 17484 18144 17536
rect 18196 17524 18202 17536
rect 18877 17527 18935 17533
rect 18877 17524 18889 17527
rect 18196 17496 18889 17524
rect 18196 17484 18202 17496
rect 18877 17493 18889 17496
rect 18923 17493 18935 17527
rect 20530 17524 20536 17536
rect 20491 17496 20536 17524
rect 18877 17487 18935 17493
rect 20530 17484 20536 17496
rect 20588 17484 20594 17536
rect 20824 17524 20852 17564
rect 20898 17552 20904 17604
rect 20956 17592 20962 17604
rect 20993 17595 21051 17601
rect 20993 17592 21005 17595
rect 20956 17564 21005 17592
rect 20956 17552 20962 17564
rect 20993 17561 21005 17564
rect 21039 17561 21051 17595
rect 22646 17592 22652 17604
rect 20993 17555 21051 17561
rect 21284 17564 22652 17592
rect 21284 17524 21312 17564
rect 22646 17552 22652 17564
rect 22704 17552 22710 17604
rect 21450 17524 21456 17536
rect 20824 17496 21312 17524
rect 21411 17496 21456 17524
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 1762 17280 1768 17332
rect 1820 17320 1826 17332
rect 4065 17323 4123 17329
rect 1820 17292 2774 17320
rect 1820 17280 1826 17292
rect 2746 17252 2774 17292
rect 4065 17289 4077 17323
rect 4111 17289 4123 17323
rect 5629 17323 5687 17329
rect 5629 17320 5641 17323
rect 4065 17283 4123 17289
rect 5460 17292 5641 17320
rect 2930 17255 2988 17261
rect 2930 17252 2942 17255
rect 2746 17224 2942 17252
rect 2930 17221 2942 17224
rect 2976 17221 2988 17255
rect 4080 17252 4108 17283
rect 4430 17261 4436 17264
rect 4424 17252 4436 17261
rect 4080 17224 4436 17252
rect 2930 17215 2988 17221
rect 4424 17215 4436 17224
rect 4430 17212 4436 17215
rect 4488 17212 4494 17264
rect 5074 17212 5080 17264
rect 5132 17252 5138 17264
rect 5460 17252 5488 17292
rect 5629 17289 5641 17292
rect 5675 17289 5687 17323
rect 5629 17283 5687 17289
rect 5718 17280 5724 17332
rect 5776 17320 5782 17332
rect 5776 17292 6224 17320
rect 5776 17280 5782 17292
rect 6196 17264 6224 17292
rect 6546 17280 6552 17332
rect 6604 17320 6610 17332
rect 7098 17320 7104 17332
rect 6604 17292 7104 17320
rect 6604 17280 6610 17292
rect 7098 17280 7104 17292
rect 7156 17280 7162 17332
rect 7193 17323 7251 17329
rect 7193 17289 7205 17323
rect 7239 17320 7251 17323
rect 8386 17320 8392 17332
rect 7239 17292 8392 17320
rect 7239 17289 7251 17292
rect 7193 17283 7251 17289
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 8662 17280 8668 17332
rect 8720 17320 8726 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8720 17292 9045 17320
rect 8720 17280 8726 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9033 17283 9091 17289
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10502 17320 10508 17332
rect 10008 17292 10508 17320
rect 10008 17280 10014 17292
rect 10502 17280 10508 17292
rect 10560 17280 10566 17332
rect 10778 17280 10784 17332
rect 10836 17320 10842 17332
rect 10965 17323 11023 17329
rect 10965 17320 10977 17323
rect 10836 17292 10977 17320
rect 10836 17280 10842 17292
rect 10965 17289 10977 17292
rect 11011 17289 11023 17323
rect 10965 17283 11023 17289
rect 11793 17323 11851 17329
rect 11793 17289 11805 17323
rect 11839 17289 11851 17323
rect 12342 17320 12348 17332
rect 12303 17292 12348 17320
rect 11793 17283 11851 17289
rect 5132 17224 5488 17252
rect 5736 17224 5948 17252
rect 5132 17212 5138 17224
rect 5736 17196 5764 17224
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 1854 17144 1860 17196
rect 1912 17184 1918 17196
rect 1949 17187 2007 17193
rect 1949 17184 1961 17187
rect 1912 17156 1961 17184
rect 1912 17144 1918 17156
rect 1949 17153 1961 17156
rect 1995 17153 2007 17187
rect 2406 17184 2412 17196
rect 2367 17156 2412 17184
rect 1949 17147 2007 17153
rect 2406 17144 2412 17156
rect 2464 17144 2470 17196
rect 2685 17187 2743 17193
rect 2685 17153 2697 17187
rect 2731 17184 2743 17187
rect 3234 17184 3240 17196
rect 2731 17156 3240 17184
rect 2731 17153 2743 17156
rect 2685 17147 2743 17153
rect 3234 17144 3240 17156
rect 3292 17184 3298 17196
rect 4157 17187 4215 17193
rect 4157 17184 4169 17187
rect 3292 17156 4169 17184
rect 3292 17144 3298 17156
rect 4157 17153 4169 17156
rect 4203 17153 4215 17187
rect 5718 17184 5724 17196
rect 4157 17147 4215 17153
rect 4264 17156 5724 17184
rect 4264 17116 4292 17156
rect 5718 17144 5724 17156
rect 5776 17144 5782 17196
rect 5813 17188 5871 17193
rect 5920 17188 5948 17224
rect 6178 17212 6184 17264
rect 6236 17212 6242 17264
rect 7530 17255 7588 17261
rect 7530 17252 7542 17255
rect 6656 17224 7542 17252
rect 5813 17187 5948 17188
rect 5813 17153 5825 17187
rect 5859 17160 5948 17187
rect 6089 17187 6147 17193
rect 5859 17153 5871 17160
rect 5813 17147 5871 17153
rect 6089 17153 6101 17187
rect 6135 17184 6147 17187
rect 6362 17184 6368 17196
rect 6135 17156 6368 17184
rect 6135 17153 6147 17156
rect 6089 17147 6147 17153
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 4172 17088 4292 17116
rect 1857 17051 1915 17057
rect 1857 17017 1869 17051
rect 1903 17048 1915 17051
rect 1946 17048 1952 17060
rect 1903 17020 1952 17048
rect 1903 17017 1915 17020
rect 1857 17011 1915 17017
rect 1946 17008 1952 17020
rect 2004 17008 2010 17060
rect 1486 16980 1492 16992
rect 1447 16952 1492 16980
rect 1486 16940 1492 16952
rect 1544 16940 1550 16992
rect 2130 16980 2136 16992
rect 2091 16952 2136 16980
rect 2130 16940 2136 16952
rect 2188 16940 2194 16992
rect 2222 16940 2228 16992
rect 2280 16980 2286 16992
rect 2593 16983 2651 16989
rect 2280 16952 2325 16980
rect 2280 16940 2286 16952
rect 2593 16949 2605 16983
rect 2639 16980 2651 16983
rect 4172 16980 4200 17088
rect 5534 17076 5540 17128
rect 5592 17116 5598 17128
rect 5592 17088 5948 17116
rect 5592 17076 5598 17088
rect 5920 17057 5948 17088
rect 6454 17076 6460 17128
rect 6512 17116 6518 17128
rect 6656 17125 6684 17224
rect 7530 17221 7542 17224
rect 7576 17221 7588 17255
rect 7530 17215 7588 17221
rect 8202 17212 8208 17264
rect 8260 17212 8266 17264
rect 8294 17212 8300 17264
rect 8352 17252 8358 17264
rect 9122 17252 9128 17264
rect 8352 17224 9128 17252
rect 8352 17212 8358 17224
rect 9122 17212 9128 17224
rect 9180 17212 9186 17264
rect 11808 17252 11836 17283
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 14185 17323 14243 17329
rect 14185 17320 14197 17323
rect 12492 17292 14197 17320
rect 12492 17280 12498 17292
rect 14185 17289 14197 17292
rect 14231 17289 14243 17323
rect 14185 17283 14243 17289
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17320 14611 17323
rect 15562 17320 15568 17332
rect 14599 17292 15568 17320
rect 14599 17289 14611 17292
rect 14553 17283 14611 17289
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 15749 17323 15807 17329
rect 15749 17289 15761 17323
rect 15795 17320 15807 17323
rect 16206 17320 16212 17332
rect 15795 17292 16068 17320
rect 16167 17292 16212 17320
rect 15795 17289 15807 17292
rect 15749 17283 15807 17289
rect 11072 17224 11836 17252
rect 11885 17255 11943 17261
rect 6825 17187 6883 17193
rect 6825 17153 6837 17187
rect 6871 17184 6883 17187
rect 7374 17184 7380 17196
rect 6871 17156 7380 17184
rect 6871 17153 6883 17156
rect 6825 17147 6883 17153
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 8220 17184 8248 17212
rect 7892 17156 8340 17184
rect 7892 17144 7898 17156
rect 6641 17119 6699 17125
rect 6641 17116 6653 17119
rect 6512 17088 6653 17116
rect 6512 17076 6518 17088
rect 6641 17085 6653 17088
rect 6687 17085 6699 17119
rect 6641 17079 6699 17085
rect 6730 17076 6736 17128
rect 6788 17116 6794 17128
rect 7285 17119 7343 17125
rect 6788 17088 6833 17116
rect 6788 17076 6794 17088
rect 7285 17085 7297 17119
rect 7331 17085 7343 17119
rect 8312 17116 8340 17156
rect 8662 17144 8668 17196
rect 8720 17184 8726 17196
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8720 17156 8953 17184
rect 8720 17144 8726 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 9214 17184 9220 17196
rect 9175 17156 9220 17184
rect 8941 17147 8999 17153
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9766 17184 9772 17196
rect 9727 17156 9772 17184
rect 9766 17144 9772 17156
rect 9824 17144 9830 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 10686 17184 10692 17196
rect 10643 17156 10692 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 10686 17144 10692 17156
rect 10744 17144 10750 17196
rect 10962 17144 10968 17196
rect 11020 17184 11026 17196
rect 11072 17184 11100 17224
rect 11885 17221 11897 17255
rect 11931 17221 11943 17255
rect 11885 17215 11943 17221
rect 11900 17184 11928 17215
rect 12066 17212 12072 17264
rect 12124 17252 12130 17264
rect 12986 17252 12992 17264
rect 12124 17224 12992 17252
rect 12124 17212 12130 17224
rect 12986 17212 12992 17224
rect 13044 17212 13050 17264
rect 13354 17212 13360 17264
rect 13412 17252 13418 17264
rect 14093 17255 14151 17261
rect 14093 17252 14105 17255
rect 13412 17224 14105 17252
rect 13412 17212 13418 17224
rect 14093 17221 14105 17224
rect 14139 17221 14151 17255
rect 14093 17215 14151 17221
rect 14642 17212 14648 17264
rect 14700 17252 14706 17264
rect 16040 17252 16068 17292
rect 16206 17280 16212 17292
rect 16264 17280 16270 17332
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 17129 17323 17187 17329
rect 17129 17320 17141 17323
rect 16356 17292 17141 17320
rect 16356 17280 16362 17292
rect 17129 17289 17141 17292
rect 17175 17289 17187 17323
rect 19610 17320 19616 17332
rect 19571 17292 19616 17320
rect 17129 17283 17187 17289
rect 19610 17280 19616 17292
rect 19668 17280 19674 17332
rect 19886 17320 19892 17332
rect 19847 17292 19892 17320
rect 19886 17280 19892 17292
rect 19944 17280 19950 17332
rect 20717 17323 20775 17329
rect 20717 17289 20729 17323
rect 20763 17320 20775 17323
rect 20806 17320 20812 17332
rect 20763 17292 20812 17320
rect 20763 17289 20775 17292
rect 20717 17283 20775 17289
rect 20806 17280 20812 17292
rect 20864 17280 20870 17332
rect 21177 17323 21235 17329
rect 21177 17289 21189 17323
rect 21223 17320 21235 17323
rect 22370 17320 22376 17332
rect 21223 17292 22376 17320
rect 21223 17289 21235 17292
rect 21177 17283 21235 17289
rect 22370 17280 22376 17292
rect 22428 17280 22434 17332
rect 17037 17255 17095 17261
rect 17037 17252 17049 17255
rect 14700 17224 15700 17252
rect 16040 17224 17049 17252
rect 14700 17212 14706 17224
rect 12710 17184 12716 17196
rect 11020 17156 11100 17184
rect 11164 17156 11928 17184
rect 12406 17156 12716 17184
rect 11020 17144 11026 17156
rect 8312 17088 8800 17116
rect 7285 17079 7343 17085
rect 5905 17051 5963 17057
rect 5905 17017 5917 17051
rect 5951 17017 5963 17051
rect 5905 17011 5963 17017
rect 2639 16952 4200 16980
rect 2639 16949 2651 16952
rect 2593 16943 2651 16949
rect 4430 16940 4436 16992
rect 4488 16980 4494 16992
rect 5537 16983 5595 16989
rect 5537 16980 5549 16983
rect 4488 16952 5549 16980
rect 4488 16940 4494 16952
rect 5537 16949 5549 16952
rect 5583 16980 5595 16983
rect 7098 16980 7104 16992
rect 5583 16952 7104 16980
rect 5583 16949 5595 16952
rect 5537 16943 5595 16949
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 7300 16980 7328 17079
rect 8478 17008 8484 17060
rect 8536 17048 8542 17060
rect 8772 17057 8800 17088
rect 9122 17076 9128 17128
rect 9180 17116 9186 17128
rect 9861 17119 9919 17125
rect 9861 17116 9873 17119
rect 9180 17088 9873 17116
rect 9180 17076 9186 17088
rect 9861 17085 9873 17088
rect 9907 17085 9919 17119
rect 10042 17116 10048 17128
rect 10003 17088 10048 17116
rect 9861 17079 9919 17085
rect 10042 17076 10048 17088
rect 10100 17076 10106 17128
rect 10318 17116 10324 17128
rect 10279 17088 10324 17116
rect 10318 17076 10324 17088
rect 10376 17076 10382 17128
rect 8665 17051 8723 17057
rect 8665 17048 8677 17051
rect 8536 17020 8677 17048
rect 8536 17008 8542 17020
rect 8665 17017 8677 17020
rect 8711 17017 8723 17051
rect 8665 17011 8723 17017
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17017 8815 17051
rect 8757 17011 8815 17017
rect 8846 17008 8852 17060
rect 8904 17048 8910 17060
rect 11164 17048 11192 17156
rect 11701 17119 11759 17125
rect 11701 17085 11713 17119
rect 11747 17085 11759 17119
rect 11701 17079 11759 17085
rect 8904 17020 11192 17048
rect 8904 17008 8910 17020
rect 11238 17008 11244 17060
rect 11296 17048 11302 17060
rect 11716 17048 11744 17079
rect 12406 17048 12434 17156
rect 12710 17144 12716 17156
rect 12768 17184 12774 17196
rect 13170 17184 13176 17196
rect 12768 17156 13176 17184
rect 12768 17144 12774 17156
rect 13170 17144 13176 17156
rect 13228 17144 13234 17196
rect 13446 17144 13452 17196
rect 13504 17193 13510 17196
rect 13504 17184 13516 17193
rect 13722 17184 13728 17196
rect 13504 17156 13549 17184
rect 13683 17156 13728 17184
rect 13504 17147 13516 17156
rect 13504 17144 13510 17147
rect 13722 17144 13728 17156
rect 13780 17144 13786 17196
rect 14921 17187 14979 17193
rect 14921 17153 14933 17187
rect 14967 17184 14979 17187
rect 15194 17184 15200 17196
rect 14967 17156 15200 17184
rect 14967 17153 14979 17156
rect 14921 17147 14979 17153
rect 15194 17144 15200 17156
rect 15252 17144 15258 17196
rect 15378 17184 15384 17196
rect 15339 17156 15384 17184
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15672 17184 15700 17224
rect 17037 17221 17049 17224
rect 17083 17221 17095 17255
rect 17037 17215 17095 17221
rect 18874 17212 18880 17264
rect 18932 17252 18938 17264
rect 18932 17224 20392 17252
rect 18932 17212 18938 17224
rect 15764 17184 15976 17188
rect 16390 17184 16396 17196
rect 15672 17160 15976 17184
rect 15672 17156 15792 17160
rect 13740 17116 13768 17144
rect 14001 17119 14059 17125
rect 13740 17088 13952 17116
rect 11296 17020 11341 17048
rect 11716 17020 12434 17048
rect 13924 17048 13952 17088
rect 14001 17085 14013 17119
rect 14047 17116 14059 17119
rect 15010 17116 15016 17128
rect 14047 17088 15016 17116
rect 14047 17085 14059 17088
rect 14001 17079 14059 17085
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15105 17119 15163 17125
rect 15105 17085 15117 17119
rect 15151 17085 15163 17119
rect 15286 17116 15292 17128
rect 15247 17088 15292 17116
rect 15105 17079 15163 17085
rect 14274 17048 14280 17060
rect 13924 17020 14280 17048
rect 11296 17008 11302 17020
rect 14274 17008 14280 17020
rect 14332 17048 14338 17060
rect 14737 17051 14795 17057
rect 14737 17048 14749 17051
rect 14332 17020 14749 17048
rect 14332 17008 14338 17020
rect 14737 17017 14749 17020
rect 14783 17017 14795 17051
rect 15120 17048 15148 17079
rect 15286 17076 15292 17088
rect 15344 17076 15350 17128
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17085 15899 17119
rect 15948 17116 15976 17160
rect 16351 17156 16396 17184
rect 16390 17144 16396 17156
rect 16448 17144 16454 17196
rect 19426 17184 19432 17196
rect 17144 17156 19432 17184
rect 17144 17116 17172 17156
rect 19426 17144 19432 17156
rect 19484 17144 19490 17196
rect 19518 17144 19524 17196
rect 19576 17184 19582 17196
rect 20364 17193 20392 17224
rect 20456 17224 20944 17252
rect 20073 17187 20131 17193
rect 20073 17184 20085 17187
rect 19576 17156 20085 17184
rect 19576 17144 19582 17156
rect 20073 17153 20085 17156
rect 20119 17153 20131 17187
rect 20073 17147 20131 17153
rect 20349 17187 20407 17193
rect 20349 17153 20361 17187
rect 20395 17153 20407 17187
rect 20349 17147 20407 17153
rect 15948 17088 17172 17116
rect 15841 17079 15899 17085
rect 15654 17048 15660 17060
rect 15120 17020 15660 17048
rect 14737 17011 14795 17017
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 8570 16980 8576 16992
rect 7300 16952 8576 16980
rect 8570 16940 8576 16952
rect 8628 16940 8634 16992
rect 10134 16940 10140 16992
rect 10192 16980 10198 16992
rect 10686 16980 10692 16992
rect 10192 16952 10692 16980
rect 10192 16940 10198 16952
rect 10686 16940 10692 16952
rect 10744 16980 10750 16992
rect 11057 16983 11115 16989
rect 11057 16980 11069 16983
rect 10744 16952 11069 16980
rect 10744 16940 10750 16952
rect 11057 16949 11069 16952
rect 11103 16980 11115 16983
rect 12066 16980 12072 16992
rect 11103 16952 12072 16980
rect 11103 16949 11115 16952
rect 11057 16943 11115 16949
rect 12066 16940 12072 16952
rect 12124 16940 12130 16992
rect 12250 16980 12256 16992
rect 12211 16952 12256 16980
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 12342 16940 12348 16992
rect 12400 16980 12406 16992
rect 14642 16980 14648 16992
rect 12400 16952 14648 16980
rect 12400 16940 12406 16952
rect 14642 16940 14648 16952
rect 14700 16940 14706 16992
rect 14918 16940 14924 16992
rect 14976 16980 14982 16992
rect 15856 16980 15884 17079
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 17276 17088 17321 17116
rect 17276 17076 17282 17088
rect 19058 17076 19064 17128
rect 19116 17116 19122 17128
rect 20456 17116 20484 17224
rect 20916 17193 20944 17224
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20901 17187 20959 17193
rect 20901 17153 20913 17187
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 19116 17088 20484 17116
rect 19116 17076 19122 17088
rect 16669 17051 16727 17057
rect 16669 17017 16681 17051
rect 16715 17048 16727 17051
rect 16942 17048 16948 17060
rect 16715 17020 16948 17048
rect 16715 17017 16727 17020
rect 16669 17011 16727 17017
rect 16942 17008 16948 17020
rect 17000 17008 17006 17060
rect 18506 17008 18512 17060
rect 18564 17048 18570 17060
rect 20640 17048 20668 17147
rect 20990 17144 20996 17196
rect 21048 17184 21054 17196
rect 21266 17184 21272 17196
rect 21048 17156 21093 17184
rect 21227 17156 21272 17184
rect 21048 17144 21054 17156
rect 21266 17144 21272 17156
rect 21324 17144 21330 17196
rect 18564 17020 20668 17048
rect 18564 17008 18570 17020
rect 14976 16952 15884 16980
rect 14976 16940 14982 16952
rect 16390 16940 16396 16992
rect 16448 16980 16454 16992
rect 17126 16980 17132 16992
rect 16448 16952 17132 16980
rect 16448 16940 16454 16952
rect 17126 16940 17132 16952
rect 17184 16940 17190 16992
rect 19429 16983 19487 16989
rect 19429 16949 19441 16983
rect 19475 16980 19487 16983
rect 19610 16980 19616 16992
rect 19475 16952 19616 16980
rect 19475 16949 19487 16952
rect 19429 16943 19487 16949
rect 19610 16940 19616 16952
rect 19668 16940 19674 16992
rect 19794 16940 19800 16992
rect 19852 16980 19858 16992
rect 20070 16980 20076 16992
rect 19852 16952 20076 16980
rect 19852 16940 19858 16952
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20441 16983 20499 16989
rect 20220 16952 20265 16980
rect 20220 16940 20226 16952
rect 20441 16949 20453 16983
rect 20487 16980 20499 16983
rect 20622 16980 20628 16992
rect 20487 16952 20628 16980
rect 20487 16949 20499 16952
rect 20441 16943 20499 16949
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 21450 16980 21456 16992
rect 21411 16952 21456 16980
rect 21450 16940 21456 16952
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1670 16736 1676 16788
rect 1728 16776 1734 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 1728 16748 3801 16776
rect 1728 16736 1734 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 3789 16739 3847 16745
rect 5350 16736 5356 16788
rect 5408 16776 5414 16788
rect 6454 16776 6460 16788
rect 5408 16748 6316 16776
rect 6415 16748 6460 16776
rect 5408 16736 5414 16748
rect 1762 16668 1768 16720
rect 1820 16708 1826 16720
rect 1857 16711 1915 16717
rect 1857 16708 1869 16711
rect 1820 16680 1869 16708
rect 1820 16668 1826 16680
rect 1857 16677 1869 16680
rect 1903 16677 1915 16711
rect 5626 16708 5632 16720
rect 1857 16671 1915 16677
rect 3896 16680 4752 16708
rect 3234 16640 3240 16652
rect 3195 16612 3240 16640
rect 3234 16600 3240 16612
rect 3292 16600 3298 16652
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2222 16572 2228 16584
rect 1719 16544 2228 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 3513 16575 3571 16581
rect 2746 16544 3096 16572
rect 2038 16464 2044 16516
rect 2096 16504 2102 16516
rect 2746 16504 2774 16544
rect 2958 16504 2964 16516
rect 3016 16513 3022 16516
rect 2096 16476 2774 16504
rect 2928 16476 2964 16504
rect 2096 16464 2102 16476
rect 2958 16464 2964 16476
rect 3016 16467 3028 16513
rect 3068 16504 3096 16544
rect 3513 16541 3525 16575
rect 3559 16572 3571 16575
rect 3896 16572 3924 16680
rect 4430 16640 4436 16652
rect 4391 16612 4436 16640
rect 4430 16600 4436 16612
rect 4488 16600 4494 16652
rect 4724 16640 4752 16680
rect 5368 16680 5632 16708
rect 5368 16649 5396 16680
rect 5626 16668 5632 16680
rect 5684 16668 5690 16720
rect 5994 16668 6000 16720
rect 6052 16668 6058 16720
rect 6178 16708 6184 16720
rect 6139 16680 6184 16708
rect 6178 16668 6184 16680
rect 6236 16668 6242 16720
rect 6288 16708 6316 16748
rect 6454 16736 6460 16748
rect 6512 16736 6518 16788
rect 9398 16736 9404 16788
rect 9456 16776 9462 16788
rect 10870 16776 10876 16788
rect 9456 16748 10456 16776
rect 10831 16748 10876 16776
rect 9456 16736 9462 16748
rect 6822 16708 6828 16720
rect 6288 16680 6828 16708
rect 6822 16668 6828 16680
rect 6880 16668 6886 16720
rect 7926 16668 7932 16720
rect 7984 16708 7990 16720
rect 8846 16708 8852 16720
rect 7984 16680 8852 16708
rect 7984 16668 7990 16680
rect 8846 16668 8852 16680
rect 8904 16668 8910 16720
rect 10428 16708 10456 16748
rect 10870 16736 10876 16748
rect 10928 16736 10934 16788
rect 12342 16776 12348 16788
rect 10980 16748 12348 16776
rect 10980 16708 11008 16748
rect 12342 16736 12348 16748
rect 12400 16736 12406 16788
rect 12434 16736 12440 16788
rect 12492 16776 12498 16788
rect 13538 16776 13544 16788
rect 12492 16748 13400 16776
rect 13499 16748 13544 16776
rect 12492 16736 12498 16748
rect 10428 16680 11008 16708
rect 13081 16711 13139 16717
rect 13081 16677 13093 16711
rect 13127 16677 13139 16711
rect 13372 16708 13400 16748
rect 13538 16736 13544 16748
rect 13596 16736 13602 16788
rect 17129 16779 17187 16785
rect 14292 16748 17080 16776
rect 14292 16708 14320 16748
rect 15654 16708 15660 16720
rect 13372 16680 14320 16708
rect 15567 16680 15660 16708
rect 13081 16671 13139 16677
rect 5353 16643 5411 16649
rect 4724 16612 4844 16640
rect 3559 16544 3924 16572
rect 3559 16541 3571 16544
rect 3513 16535 3571 16541
rect 3970 16532 3976 16584
rect 4028 16572 4034 16584
rect 4249 16575 4307 16581
rect 4028 16544 4073 16572
rect 4028 16532 4034 16544
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 4706 16572 4712 16584
rect 4295 16544 4384 16572
rect 4667 16544 4712 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 3068 16476 4108 16504
rect 3016 16464 3022 16467
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 1670 16396 1676 16448
rect 1728 16436 1734 16448
rect 4080 16445 4108 16476
rect 3329 16439 3387 16445
rect 3329 16436 3341 16439
rect 1728 16408 3341 16436
rect 1728 16396 1734 16408
rect 3329 16405 3341 16408
rect 3375 16405 3387 16439
rect 3329 16399 3387 16405
rect 4065 16439 4123 16445
rect 4065 16405 4077 16439
rect 4111 16405 4123 16439
rect 4065 16399 4123 16405
rect 4246 16396 4252 16448
rect 4304 16436 4310 16448
rect 4356 16436 4384 16544
rect 4706 16532 4712 16544
rect 4764 16532 4770 16584
rect 4816 16504 4844 16612
rect 5353 16609 5365 16643
rect 5399 16609 5411 16643
rect 5353 16603 5411 16609
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 6012 16640 6040 16668
rect 7834 16640 7840 16652
rect 5491 16612 6040 16640
rect 7795 16612 7840 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 7834 16600 7840 16612
rect 7892 16600 7898 16652
rect 8570 16640 8576 16652
rect 8531 16612 8576 16640
rect 8570 16600 8576 16612
rect 8628 16600 8634 16652
rect 9309 16643 9367 16649
rect 9309 16640 9321 16643
rect 8680 16612 9321 16640
rect 5537 16575 5595 16581
rect 5537 16541 5549 16575
rect 5583 16572 5595 16575
rect 5902 16572 5908 16584
rect 5583 16544 5908 16572
rect 5583 16541 5595 16544
rect 5537 16535 5595 16541
rect 5902 16532 5908 16544
rect 5960 16532 5966 16584
rect 5994 16532 6000 16584
rect 6052 16572 6058 16584
rect 6270 16572 6276 16584
rect 6052 16544 6097 16572
rect 6231 16544 6276 16572
rect 6052 16532 6058 16544
rect 6270 16532 6276 16544
rect 6328 16532 6334 16584
rect 6362 16532 6368 16584
rect 6420 16572 6426 16584
rect 7006 16572 7012 16584
rect 6420 16544 7012 16572
rect 6420 16532 6426 16544
rect 7006 16532 7012 16544
rect 7064 16532 7070 16584
rect 7282 16532 7288 16584
rect 7340 16572 7346 16584
rect 8478 16572 8484 16584
rect 7340 16544 8248 16572
rect 8439 16544 8484 16572
rect 7340 16532 7346 16544
rect 8220 16516 8248 16544
rect 8478 16532 8484 16544
rect 8536 16572 8542 16584
rect 8680 16572 8708 16612
rect 9309 16609 9321 16612
rect 9355 16609 9367 16643
rect 9490 16640 9496 16652
rect 9451 16612 9496 16640
rect 9309 16603 9367 16609
rect 9490 16600 9496 16612
rect 9548 16600 9554 16652
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11333 16643 11391 16649
rect 11333 16640 11345 16643
rect 11204 16612 11345 16640
rect 11204 16600 11210 16612
rect 11333 16609 11345 16612
rect 11379 16609 11391 16643
rect 11514 16640 11520 16652
rect 11475 16612 11520 16640
rect 11333 16603 11391 16609
rect 11514 16600 11520 16612
rect 11572 16600 11578 16652
rect 11698 16640 11704 16652
rect 11659 16612 11704 16640
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 13096 16640 13124 16671
rect 15654 16668 15660 16680
rect 15712 16668 15718 16720
rect 17052 16708 17080 16748
rect 17129 16745 17141 16779
rect 17175 16776 17187 16779
rect 17218 16776 17224 16788
rect 17175 16748 17224 16776
rect 17175 16745 17187 16748
rect 17129 16739 17187 16745
rect 17218 16736 17224 16748
rect 17276 16736 17282 16788
rect 17310 16736 17316 16788
rect 17368 16776 17374 16788
rect 17368 16748 17413 16776
rect 17368 16736 17374 16748
rect 18690 16736 18696 16788
rect 18748 16776 18754 16788
rect 20162 16776 20168 16788
rect 18748 16748 20168 16776
rect 18748 16736 18754 16748
rect 20162 16736 20168 16748
rect 20220 16736 20226 16788
rect 20993 16779 21051 16785
rect 20456 16748 20677 16776
rect 17494 16708 17500 16720
rect 17052 16680 17500 16708
rect 17494 16668 17500 16680
rect 17552 16668 17558 16720
rect 17770 16708 17776 16720
rect 17731 16680 17776 16708
rect 17770 16668 17776 16680
rect 17828 16668 17834 16720
rect 17954 16708 17960 16720
rect 17915 16680 17960 16708
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 18598 16668 18604 16720
rect 18656 16708 18662 16720
rect 20254 16708 20260 16720
rect 18656 16680 20260 16708
rect 18656 16668 18662 16680
rect 20254 16668 20260 16680
rect 20312 16668 20318 16720
rect 13538 16640 13544 16652
rect 13096 16612 13544 16640
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 14274 16640 14280 16652
rect 14235 16612 14280 16640
rect 14274 16600 14280 16612
rect 14332 16600 14338 16652
rect 15672 16640 15700 16668
rect 15672 16612 15884 16640
rect 8536 16544 8708 16572
rect 8536 16532 8542 16544
rect 10502 16532 10508 16584
rect 10560 16572 10566 16584
rect 11238 16572 11244 16584
rect 10560 16544 11244 16572
rect 10560 16532 10566 16544
rect 11238 16532 11244 16544
rect 11296 16532 11302 16584
rect 12986 16532 12992 16584
rect 13044 16572 13050 16584
rect 13630 16572 13636 16584
rect 13044 16544 13636 16572
rect 13044 16532 13050 16544
rect 13630 16532 13636 16544
rect 13688 16532 13694 16584
rect 15749 16575 15807 16581
rect 15749 16541 15761 16575
rect 15795 16541 15807 16575
rect 15856 16572 15884 16612
rect 17310 16600 17316 16652
rect 17368 16640 17374 16652
rect 17405 16643 17463 16649
rect 17405 16640 17417 16643
rect 17368 16612 17417 16640
rect 17368 16600 17374 16612
rect 17405 16609 17417 16612
rect 17451 16609 17463 16643
rect 17405 16603 17463 16609
rect 17681 16643 17739 16649
rect 17681 16609 17693 16643
rect 17727 16640 17739 16643
rect 17862 16640 17868 16652
rect 17727 16612 17868 16640
rect 17727 16609 17739 16612
rect 17681 16603 17739 16609
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 19978 16640 19984 16652
rect 19939 16612 19984 16640
rect 19978 16600 19984 16612
rect 20036 16600 20042 16652
rect 20165 16643 20223 16649
rect 20165 16609 20177 16643
rect 20211 16640 20223 16643
rect 20456 16640 20484 16748
rect 20211 16612 20484 16640
rect 20649 16640 20677 16748
rect 20993 16745 21005 16779
rect 21039 16776 21051 16779
rect 21266 16776 21272 16788
rect 21039 16748 21272 16776
rect 21039 16745 21051 16748
rect 20993 16739 21051 16745
rect 21266 16736 21272 16748
rect 21324 16736 21330 16788
rect 20717 16711 20775 16717
rect 20717 16677 20729 16711
rect 20763 16708 20775 16711
rect 21082 16708 21088 16720
rect 20763 16680 21088 16708
rect 20763 16677 20775 16680
rect 20717 16671 20775 16677
rect 21082 16668 21088 16680
rect 21140 16668 21146 16720
rect 21726 16640 21732 16652
rect 20649 16612 21732 16640
rect 20211 16609 20223 16612
rect 20165 16603 20223 16609
rect 21726 16600 21732 16612
rect 21784 16600 21790 16652
rect 16022 16581 16028 16584
rect 16005 16575 16028 16581
rect 16005 16572 16017 16575
rect 15856 16544 16017 16572
rect 15749 16535 15807 16541
rect 16005 16541 16017 16544
rect 16005 16535 16028 16541
rect 5442 16504 5448 16516
rect 4816 16476 5448 16504
rect 5442 16464 5448 16476
rect 5500 16464 5506 16516
rect 7570 16507 7628 16513
rect 7570 16504 7582 16507
rect 5552 16476 7582 16504
rect 5552 16448 5580 16476
rect 7570 16473 7582 16476
rect 7616 16504 7628 16507
rect 8110 16504 8116 16516
rect 7616 16476 8116 16504
rect 7616 16473 7628 16476
rect 7570 16467 7628 16473
rect 8110 16464 8116 16476
rect 8168 16464 8174 16516
rect 8202 16464 8208 16516
rect 8260 16504 8266 16516
rect 9760 16507 9818 16513
rect 8260 16476 9168 16504
rect 8260 16464 8266 16476
rect 4304 16408 4384 16436
rect 4304 16396 4310 16408
rect 4522 16396 4528 16448
rect 4580 16436 4586 16448
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 4580 16408 4629 16436
rect 4580 16396 4586 16408
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 5074 16436 5080 16448
rect 5035 16408 5080 16436
rect 4617 16399 4675 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5534 16396 5540 16448
rect 5592 16396 5598 16448
rect 5902 16436 5908 16448
rect 5863 16408 5908 16436
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 8018 16436 8024 16448
rect 7979 16408 8024 16436
rect 8018 16396 8024 16408
rect 8076 16396 8082 16448
rect 8386 16436 8392 16448
rect 8347 16408 8392 16436
rect 8386 16396 8392 16408
rect 8444 16436 8450 16448
rect 9033 16439 9091 16445
rect 9033 16436 9045 16439
rect 8444 16408 9045 16436
rect 8444 16396 8450 16408
rect 9033 16405 9045 16408
rect 9079 16405 9091 16439
rect 9140 16436 9168 16476
rect 9760 16473 9772 16507
rect 9806 16504 9818 16507
rect 10042 16504 10048 16516
rect 9806 16476 10048 16504
rect 9806 16473 9818 16476
rect 9760 16467 9818 16473
rect 10042 16464 10048 16476
rect 10100 16504 10106 16516
rect 10318 16504 10324 16516
rect 10100 16476 10324 16504
rect 10100 16464 10106 16476
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 10965 16507 11023 16513
rect 10965 16504 10977 16507
rect 10836 16476 10977 16504
rect 10836 16464 10842 16476
rect 10965 16473 10977 16476
rect 11011 16473 11023 16507
rect 10965 16467 11023 16473
rect 11968 16507 12026 16513
rect 11968 16473 11980 16507
rect 12014 16504 12026 16507
rect 12434 16504 12440 16516
rect 12014 16476 12440 16504
rect 12014 16473 12026 16476
rect 11968 16467 12026 16473
rect 12434 16464 12440 16476
rect 12492 16464 12498 16516
rect 12618 16464 12624 16516
rect 12676 16504 12682 16516
rect 13357 16507 13415 16513
rect 13357 16504 13369 16507
rect 12676 16476 13369 16504
rect 12676 16464 12682 16476
rect 13357 16473 13369 16476
rect 13403 16473 13415 16507
rect 13357 16467 13415 16473
rect 14544 16507 14602 16513
rect 14544 16473 14556 16507
rect 14590 16504 14602 16507
rect 15102 16504 15108 16516
rect 14590 16476 15108 16504
rect 14590 16473 14602 16476
rect 14544 16467 14602 16473
rect 15102 16464 15108 16476
rect 15160 16464 15166 16516
rect 15194 16464 15200 16516
rect 15252 16504 15258 16516
rect 15764 16504 15792 16535
rect 16022 16532 16028 16535
rect 16080 16532 16086 16584
rect 19886 16572 19892 16584
rect 17144 16544 19892 16572
rect 16942 16504 16948 16516
rect 15252 16476 16948 16504
rect 15252 16464 15258 16476
rect 16942 16464 16948 16476
rect 17000 16464 17006 16516
rect 10686 16436 10692 16448
rect 9140 16408 10692 16436
rect 9033 16399 9091 16405
rect 10686 16396 10692 16408
rect 10744 16436 10750 16448
rect 11882 16436 11888 16448
rect 10744 16408 11888 16436
rect 10744 16396 10750 16408
rect 11882 16396 11888 16408
rect 11940 16396 11946 16448
rect 12802 16396 12808 16448
rect 12860 16436 12866 16448
rect 13173 16439 13231 16445
rect 13173 16436 13185 16439
rect 12860 16408 13185 16436
rect 12860 16396 12866 16408
rect 13173 16405 13185 16408
rect 13219 16436 13231 16439
rect 13722 16436 13728 16448
rect 13219 16408 13728 16436
rect 13219 16405 13231 16408
rect 13173 16399 13231 16405
rect 13722 16396 13728 16408
rect 13780 16396 13786 16448
rect 13906 16436 13912 16448
rect 13867 16408 13912 16436
rect 13906 16396 13912 16408
rect 13964 16396 13970 16448
rect 14185 16439 14243 16445
rect 14185 16405 14197 16439
rect 14231 16436 14243 16439
rect 14366 16436 14372 16448
rect 14231 16408 14372 16436
rect 14231 16405 14243 16408
rect 14185 16399 14243 16405
rect 14366 16396 14372 16408
rect 14424 16396 14430 16448
rect 14734 16396 14740 16448
rect 14792 16436 14798 16448
rect 17144 16436 17172 16544
rect 19886 16532 19892 16544
rect 19944 16532 19950 16584
rect 20525 16575 20583 16581
rect 20525 16572 20537 16575
rect 20364 16544 20537 16572
rect 18046 16464 18052 16516
rect 18104 16504 18110 16516
rect 20162 16504 20168 16516
rect 18104 16476 20168 16504
rect 18104 16464 18110 16476
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 14792 16408 17172 16436
rect 14792 16396 14798 16408
rect 17494 16396 17500 16448
rect 17552 16436 17558 16448
rect 18414 16436 18420 16448
rect 17552 16408 18420 16436
rect 17552 16396 17558 16408
rect 18414 16396 18420 16408
rect 18472 16396 18478 16448
rect 18874 16396 18880 16448
rect 18932 16436 18938 16448
rect 20364 16445 20392 16544
rect 20525 16541 20537 16544
rect 20571 16541 20583 16575
rect 20806 16572 20812 16584
rect 20767 16544 20812 16572
rect 20525 16535 20583 16541
rect 20806 16532 20812 16544
rect 20864 16572 20870 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20864 16544 21097 16572
rect 20864 16532 20870 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21266 16572 21272 16584
rect 21227 16544 21272 16572
rect 21085 16535 21143 16541
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 20349 16439 20407 16445
rect 20349 16436 20361 16439
rect 18932 16408 20361 16436
rect 18932 16396 18938 16408
rect 20349 16405 20361 16408
rect 20395 16405 20407 16439
rect 21450 16436 21456 16448
rect 21411 16408 21456 16436
rect 20349 16399 20407 16405
rect 21450 16396 21456 16408
rect 21508 16396 21514 16448
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 2133 16235 2191 16241
rect 2133 16201 2145 16235
rect 2179 16232 2191 16235
rect 2593 16235 2651 16241
rect 2593 16232 2605 16235
rect 2179 16204 2605 16232
rect 2179 16201 2191 16204
rect 2133 16195 2191 16201
rect 2593 16201 2605 16204
rect 2639 16201 2651 16235
rect 2593 16195 2651 16201
rect 2958 16192 2964 16244
rect 3016 16192 3022 16244
rect 3973 16235 4031 16241
rect 3973 16201 3985 16235
rect 4019 16232 4031 16235
rect 4433 16235 4491 16241
rect 4433 16232 4445 16235
rect 4019 16204 4445 16232
rect 4019 16201 4031 16204
rect 3973 16195 4031 16201
rect 4433 16201 4445 16204
rect 4479 16201 4491 16235
rect 4433 16195 4491 16201
rect 4890 16192 4896 16244
rect 4948 16232 4954 16244
rect 5258 16232 5264 16244
rect 4948 16204 5264 16232
rect 4948 16192 4954 16204
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 5721 16235 5779 16241
rect 5721 16201 5733 16235
rect 5767 16232 5779 16235
rect 5902 16232 5908 16244
rect 5767 16204 5908 16232
rect 5767 16201 5779 16204
rect 5721 16195 5779 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6181 16235 6239 16241
rect 6181 16201 6193 16235
rect 6227 16232 6239 16235
rect 6730 16232 6736 16244
rect 6227 16204 6736 16232
rect 6227 16201 6239 16204
rect 6181 16195 6239 16201
rect 6730 16192 6736 16204
rect 6788 16192 6794 16244
rect 7190 16232 7196 16244
rect 7151 16204 7196 16232
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7653 16235 7711 16241
rect 7653 16201 7665 16235
rect 7699 16232 7711 16235
rect 8113 16235 8171 16241
rect 8113 16232 8125 16235
rect 7699 16204 8125 16232
rect 7699 16201 7711 16204
rect 7653 16195 7711 16201
rect 8113 16201 8125 16204
rect 8159 16201 8171 16235
rect 8113 16195 8171 16201
rect 8202 16192 8208 16244
rect 8260 16232 8266 16244
rect 8757 16235 8815 16241
rect 8757 16232 8769 16235
rect 8260 16204 8769 16232
rect 8260 16192 8266 16204
rect 8757 16201 8769 16204
rect 8803 16201 8815 16235
rect 10318 16232 10324 16244
rect 8757 16195 8815 16201
rect 8884 16204 10180 16232
rect 10279 16204 10324 16232
rect 2222 16124 2228 16176
rect 2280 16164 2286 16176
rect 2406 16164 2412 16176
rect 2280 16136 2412 16164
rect 2280 16124 2286 16136
rect 2406 16124 2412 16136
rect 2464 16164 2470 16176
rect 2976 16164 3004 16192
rect 5813 16167 5871 16173
rect 2464 16136 3280 16164
rect 2464 16124 2470 16136
rect 1670 16096 1676 16108
rect 1631 16068 1676 16096
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 2958 16096 2964 16108
rect 2919 16068 2964 16096
rect 2958 16056 2964 16068
rect 3016 16056 3022 16108
rect 3252 16096 3280 16136
rect 5813 16133 5825 16167
rect 5859 16164 5871 16167
rect 5859 16136 5948 16164
rect 5859 16133 5871 16136
rect 5813 16127 5871 16133
rect 5920 16108 5948 16136
rect 6086 16124 6092 16176
rect 6144 16164 6150 16176
rect 8884 16164 8912 16204
rect 9490 16164 9496 16176
rect 6144 16136 8912 16164
rect 8956 16136 9496 16164
rect 6144 16124 6150 16136
rect 3252 16068 4200 16096
rect 1762 15988 1768 16040
rect 1820 16028 1826 16040
rect 1857 16031 1915 16037
rect 1857 16028 1869 16031
rect 1820 16000 1869 16028
rect 1820 15988 1826 16000
rect 1857 15997 1869 16000
rect 1903 15997 1915 16031
rect 1857 15991 1915 15997
rect 2041 16031 2099 16037
rect 2041 15997 2053 16031
rect 2087 15997 2099 16031
rect 3050 16028 3056 16040
rect 3011 16000 3056 16028
rect 2041 15991 2099 15997
rect 2056 15960 2084 15991
rect 3050 15988 3056 16000
rect 3108 15988 3114 16040
rect 3252 16037 3280 16068
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 15997 3295 16031
rect 4062 16028 4068 16040
rect 4023 16000 4068 16028
rect 3237 15991 3295 15997
rect 4062 15988 4068 16000
rect 4120 15988 4126 16040
rect 4172 16037 4200 16068
rect 4338 16056 4344 16108
rect 4396 16096 4402 16108
rect 4801 16099 4859 16105
rect 4801 16096 4813 16099
rect 4396 16068 4813 16096
rect 4396 16056 4402 16068
rect 4801 16065 4813 16068
rect 4847 16096 4859 16099
rect 4847 16068 5212 16096
rect 4847 16065 4859 16068
rect 4801 16059 4859 16065
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 15997 4215 16031
rect 4890 16028 4896 16040
rect 4851 16000 4896 16028
rect 4157 15991 4215 15997
rect 4890 15988 4896 16000
rect 4948 15988 4954 16040
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 15997 5043 16031
rect 5184 16028 5212 16068
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 5316 16068 5764 16096
rect 5316 16056 5322 16068
rect 5350 16028 5356 16040
rect 5184 16000 5356 16028
rect 4985 15991 5043 15997
rect 3605 15963 3663 15969
rect 3605 15960 3617 15963
rect 2056 15932 3617 15960
rect 3605 15929 3617 15932
rect 3651 15929 3663 15963
rect 3605 15923 3663 15929
rect 3970 15920 3976 15972
rect 4028 15960 4034 15972
rect 4028 15932 4752 15960
rect 4028 15920 4034 15932
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 2498 15892 2504 15904
rect 2459 15864 2504 15892
rect 2498 15852 2504 15864
rect 2556 15852 2562 15904
rect 3513 15895 3571 15901
rect 3513 15861 3525 15895
rect 3559 15892 3571 15895
rect 4338 15892 4344 15904
rect 3559 15864 4344 15892
rect 3559 15861 3571 15864
rect 3513 15855 3571 15861
rect 4338 15852 4344 15864
rect 4396 15852 4402 15904
rect 4724 15892 4752 15932
rect 4798 15920 4804 15972
rect 4856 15960 4862 15972
rect 5000 15960 5028 15991
rect 5350 15988 5356 16000
rect 5408 15988 5414 16040
rect 5534 16028 5540 16040
rect 5495 16000 5540 16028
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 5736 16028 5764 16068
rect 5902 16056 5908 16108
rect 5960 16056 5966 16108
rect 6365 16099 6423 16105
rect 6365 16096 6377 16099
rect 6012 16068 6377 16096
rect 6012 16028 6040 16068
rect 6365 16065 6377 16068
rect 6411 16065 6423 16099
rect 6365 16059 6423 16065
rect 6825 16099 6883 16105
rect 6825 16065 6837 16099
rect 6871 16096 6883 16099
rect 7285 16099 7343 16105
rect 7285 16096 7297 16099
rect 6871 16068 7297 16096
rect 6871 16065 6883 16068
rect 6825 16059 6883 16065
rect 7285 16065 7297 16068
rect 7331 16065 7343 16099
rect 7285 16059 7343 16065
rect 8110 16056 8116 16108
rect 8168 16096 8174 16108
rect 8956 16105 8984 16136
rect 9490 16124 9496 16136
rect 9548 16124 9554 16176
rect 10152 16164 10180 16204
rect 10318 16192 10324 16204
rect 10376 16192 10382 16244
rect 10594 16232 10600 16244
rect 10555 16204 10600 16232
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 11238 16192 11244 16244
rect 11296 16232 11302 16244
rect 12618 16232 12624 16244
rect 11296 16204 12624 16232
rect 11296 16192 11302 16204
rect 12618 16192 12624 16204
rect 12676 16192 12682 16244
rect 12989 16235 13047 16241
rect 12989 16201 13001 16235
rect 13035 16232 13047 16235
rect 13078 16232 13084 16244
rect 13035 16204 13084 16232
rect 13035 16201 13047 16204
rect 12989 16195 13047 16201
rect 13078 16192 13084 16204
rect 13136 16192 13142 16244
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 13906 16192 13912 16244
rect 13964 16232 13970 16244
rect 15013 16235 15071 16241
rect 15013 16232 15025 16235
rect 13964 16204 15025 16232
rect 13964 16192 13970 16204
rect 15013 16201 15025 16204
rect 15059 16201 15071 16235
rect 15013 16195 15071 16201
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15381 16235 15439 16241
rect 15381 16232 15393 16235
rect 15344 16204 15393 16232
rect 15344 16192 15350 16204
rect 15381 16201 15393 16204
rect 15427 16201 15439 16235
rect 15381 16195 15439 16201
rect 15654 16192 15660 16244
rect 15712 16232 15718 16244
rect 15841 16235 15899 16241
rect 15841 16232 15853 16235
rect 15712 16204 15853 16232
rect 15712 16192 15718 16204
rect 15841 16201 15853 16204
rect 15887 16201 15899 16235
rect 15841 16195 15899 16201
rect 10413 16167 10471 16173
rect 10413 16164 10425 16167
rect 10152 16136 10425 16164
rect 10413 16133 10425 16136
rect 10459 16164 10471 16167
rect 12158 16164 12164 16176
rect 10459 16136 12164 16164
rect 10459 16133 10471 16136
rect 10413 16127 10471 16133
rect 12158 16124 12164 16136
rect 12216 16124 12222 16176
rect 12342 16124 12348 16176
rect 12400 16164 12406 16176
rect 14277 16167 14335 16173
rect 14277 16164 14289 16167
rect 12400 16136 14289 16164
rect 12400 16124 12406 16136
rect 14277 16133 14289 16136
rect 14323 16133 14335 16167
rect 14277 16127 14335 16133
rect 14366 16124 14372 16176
rect 14424 16164 14430 16176
rect 14826 16164 14832 16176
rect 14424 16136 14832 16164
rect 14424 16124 14430 16136
rect 14826 16124 14832 16136
rect 14884 16164 14890 16176
rect 14921 16167 14979 16173
rect 14921 16164 14933 16167
rect 14884 16136 14933 16164
rect 14884 16124 14890 16136
rect 14921 16133 14933 16136
rect 14967 16133 14979 16167
rect 15856 16164 15884 16195
rect 15930 16192 15936 16244
rect 15988 16232 15994 16244
rect 16209 16235 16267 16241
rect 16209 16232 16221 16235
rect 15988 16204 16221 16232
rect 15988 16192 15994 16204
rect 16209 16201 16221 16204
rect 16255 16201 16267 16235
rect 16209 16195 16267 16201
rect 17218 16192 17224 16244
rect 17276 16192 17282 16244
rect 18046 16192 18052 16244
rect 18104 16232 18110 16244
rect 18141 16235 18199 16241
rect 18141 16232 18153 16235
rect 18104 16204 18153 16232
rect 18104 16192 18110 16204
rect 18141 16201 18153 16204
rect 18187 16232 18199 16235
rect 18230 16232 18236 16244
rect 18187 16204 18236 16232
rect 18187 16201 18199 16204
rect 18141 16195 18199 16201
rect 18230 16192 18236 16204
rect 18288 16192 18294 16244
rect 19150 16232 19156 16244
rect 19111 16204 19156 16232
rect 19150 16192 19156 16204
rect 19208 16192 19214 16244
rect 19886 16232 19892 16244
rect 19847 16204 19892 16232
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 20346 16192 20352 16244
rect 20404 16232 20410 16244
rect 20533 16235 20591 16241
rect 20533 16232 20545 16235
rect 20404 16204 20545 16232
rect 20404 16192 20410 16204
rect 20533 16201 20545 16204
rect 20579 16201 20591 16235
rect 20533 16195 20591 16201
rect 20993 16235 21051 16241
rect 20993 16201 21005 16235
rect 21039 16232 21051 16235
rect 21039 16204 21312 16232
rect 21039 16201 21051 16204
rect 20993 16195 21051 16201
rect 16301 16167 16359 16173
rect 16301 16164 16313 16167
rect 15856 16136 16313 16164
rect 14921 16127 14979 16133
rect 16301 16133 16313 16136
rect 16347 16133 16359 16167
rect 16301 16127 16359 16133
rect 16936 16167 16994 16173
rect 16936 16133 16948 16167
rect 16982 16164 16994 16167
rect 17236 16164 17264 16192
rect 18322 16164 18328 16176
rect 16982 16136 17264 16164
rect 18283 16136 18328 16164
rect 16982 16133 16994 16136
rect 16936 16127 16994 16133
rect 18322 16124 18328 16136
rect 18380 16124 18386 16176
rect 19705 16167 19763 16173
rect 19705 16133 19717 16167
rect 19751 16164 19763 16167
rect 21082 16164 21088 16176
rect 19751 16136 20944 16164
rect 21043 16136 21088 16164
rect 19751 16133 19763 16136
rect 19705 16127 19763 16133
rect 8941 16099 8999 16105
rect 8168 16068 8340 16096
rect 8168 16056 8174 16068
rect 5736 16000 6040 16028
rect 6178 15988 6184 16040
rect 6236 16028 6242 16040
rect 6546 16028 6552 16040
rect 6236 16000 6552 16028
rect 6236 15988 6242 16000
rect 6546 15988 6552 16000
rect 6604 16028 6610 16040
rect 7009 16031 7067 16037
rect 7009 16028 7021 16031
rect 6604 16000 7021 16028
rect 6604 15988 6610 16000
rect 7009 15997 7021 16000
rect 7055 15997 7067 16031
rect 8202 16028 8208 16040
rect 8163 16000 8208 16028
rect 7009 15991 7067 15997
rect 8202 15988 8208 16000
rect 8260 15988 8266 16040
rect 8312 16037 8340 16068
rect 8941 16065 8953 16099
rect 8987 16065 8999 16099
rect 9208 16099 9266 16105
rect 9208 16096 9220 16099
rect 8941 16059 8999 16065
rect 9048 16068 9220 16096
rect 8297 16031 8355 16037
rect 8297 15997 8309 16031
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 8386 15988 8392 16040
rect 8444 16028 8450 16040
rect 9048 16028 9076 16068
rect 9208 16065 9220 16068
rect 9254 16096 9266 16099
rect 9582 16096 9588 16108
rect 9254 16068 9588 16096
rect 9254 16065 9266 16068
rect 9208 16059 9266 16065
rect 9582 16056 9588 16068
rect 9640 16056 9646 16108
rect 10962 16096 10968 16108
rect 10923 16068 10968 16096
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 11057 16099 11115 16105
rect 11057 16065 11069 16099
rect 11103 16096 11115 16099
rect 11330 16096 11336 16108
rect 11103 16068 11336 16096
rect 11103 16065 11115 16068
rect 11057 16059 11115 16065
rect 11330 16056 11336 16068
rect 11388 16056 11394 16108
rect 12529 16099 12587 16105
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 12802 16096 12808 16108
rect 12575 16068 12808 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 13170 16056 13176 16108
rect 13228 16096 13234 16108
rect 13357 16099 13415 16105
rect 13357 16096 13369 16099
rect 13228 16068 13369 16096
rect 13228 16056 13234 16068
rect 13357 16065 13369 16068
rect 13403 16065 13415 16099
rect 13357 16059 13415 16065
rect 13630 16056 13636 16108
rect 13688 16096 13694 16108
rect 14185 16099 14243 16105
rect 14185 16096 14197 16099
rect 13688 16068 14197 16096
rect 13688 16056 13694 16068
rect 14185 16065 14197 16068
rect 14231 16065 14243 16099
rect 14185 16059 14243 16065
rect 16669 16099 16727 16105
rect 16669 16065 16681 16099
rect 16715 16096 16727 16099
rect 16758 16096 16764 16108
rect 16715 16068 16764 16096
rect 16715 16065 16727 16068
rect 16669 16059 16727 16065
rect 16758 16056 16764 16068
rect 16816 16056 16822 16108
rect 17696 16068 20024 16096
rect 8444 16000 9076 16028
rect 8444 15988 8450 16000
rect 10870 15988 10876 16040
rect 10928 16028 10934 16040
rect 11149 16031 11207 16037
rect 11149 16028 11161 16031
rect 10928 16000 11161 16028
rect 10928 15988 10934 16000
rect 11149 15997 11161 16000
rect 11195 15997 11207 16031
rect 12710 16028 12716 16040
rect 12671 16000 12716 16028
rect 11149 15991 11207 15997
rect 12710 15988 12716 16000
rect 12768 15988 12774 16040
rect 13446 16028 13452 16040
rect 13407 16000 13452 16028
rect 13446 15988 13452 16000
rect 13504 15988 13510 16040
rect 13538 15988 13544 16040
rect 13596 16028 13602 16040
rect 14369 16031 14427 16037
rect 14369 16028 14381 16031
rect 13596 16000 14381 16028
rect 13596 15988 13602 16000
rect 14369 15997 14381 16000
rect 14415 15997 14427 16031
rect 14369 15991 14427 15997
rect 14829 16031 14887 16037
rect 14829 15997 14841 16031
rect 14875 15997 14887 16031
rect 14829 15991 14887 15997
rect 4856 15932 5028 15960
rect 4856 15920 4862 15932
rect 5902 15920 5908 15972
rect 5960 15960 5966 15972
rect 6454 15960 6460 15972
rect 5960 15932 6460 15960
rect 5960 15920 5966 15932
rect 6454 15920 6460 15932
rect 6512 15920 6518 15972
rect 6730 15920 6736 15972
rect 6788 15960 6794 15972
rect 6914 15960 6920 15972
rect 6788 15932 6920 15960
rect 6788 15920 6794 15932
rect 6914 15920 6920 15932
rect 6972 15920 6978 15972
rect 7374 15920 7380 15972
rect 7432 15960 7438 15972
rect 7745 15963 7803 15969
rect 7745 15960 7757 15963
rect 7432 15932 7757 15960
rect 7432 15920 7438 15932
rect 7745 15929 7757 15932
rect 7791 15929 7803 15963
rect 7745 15923 7803 15929
rect 8846 15920 8852 15972
rect 8904 15920 8910 15972
rect 13078 15960 13084 15972
rect 10152 15932 13084 15960
rect 6086 15892 6092 15904
rect 4724 15864 6092 15892
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 6549 15895 6607 15901
rect 6549 15861 6561 15895
rect 6595 15892 6607 15895
rect 6638 15892 6644 15904
rect 6595 15864 6644 15892
rect 6595 15861 6607 15864
rect 6549 15855 6607 15861
rect 6638 15852 6644 15864
rect 6696 15852 6702 15904
rect 8570 15892 8576 15904
rect 8531 15864 8576 15892
rect 8570 15852 8576 15864
rect 8628 15852 8634 15904
rect 8864 15892 8892 15920
rect 10152 15892 10180 15932
rect 13078 15920 13084 15932
rect 13136 15920 13142 15972
rect 14844 15960 14872 15991
rect 15102 15988 15108 16040
rect 15160 16028 15166 16040
rect 15565 16031 15623 16037
rect 15565 16028 15577 16031
rect 15160 16000 15577 16028
rect 15160 15988 15166 16000
rect 15565 15997 15577 16000
rect 15611 15997 15623 16031
rect 15565 15991 15623 15997
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 16028 15807 16031
rect 16022 16028 16028 16040
rect 15795 16000 16028 16028
rect 15795 15997 15807 16000
rect 15749 15991 15807 15997
rect 16022 15988 16028 16000
rect 16080 15988 16086 16040
rect 15120 15960 15148 15988
rect 14844 15932 15148 15960
rect 8864 15864 10180 15892
rect 10226 15852 10232 15904
rect 10284 15892 10290 15904
rect 10778 15892 10784 15904
rect 10284 15864 10784 15892
rect 10284 15852 10290 15864
rect 10778 15852 10784 15864
rect 10836 15892 10842 15904
rect 11330 15892 11336 15904
rect 10836 15864 11336 15892
rect 10836 15852 10842 15864
rect 11330 15852 11336 15864
rect 11388 15892 11394 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11388 15864 11529 15892
rect 11388 15852 11394 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11698 15892 11704 15904
rect 11659 15864 11704 15892
rect 11517 15855 11575 15861
rect 11698 15852 11704 15864
rect 11756 15852 11762 15904
rect 11882 15892 11888 15904
rect 11843 15864 11888 15892
rect 11882 15852 11888 15864
rect 11940 15852 11946 15904
rect 12158 15892 12164 15904
rect 12119 15864 12164 15892
rect 12158 15852 12164 15864
rect 12216 15852 12222 15904
rect 14642 15852 14648 15904
rect 14700 15892 14706 15904
rect 17696 15892 17724 16068
rect 19337 16031 19395 16037
rect 19337 15997 19349 16031
rect 19383 16028 19395 16031
rect 19794 16028 19800 16040
rect 19383 16000 19800 16028
rect 19383 15997 19395 16000
rect 19337 15991 19395 15997
rect 19794 15988 19800 16000
rect 19852 15988 19858 16040
rect 18322 15920 18328 15972
rect 18380 15960 18386 15972
rect 19610 15960 19616 15972
rect 18380 15932 19616 15960
rect 18380 15920 18386 15932
rect 19610 15920 19616 15932
rect 19668 15920 19674 15972
rect 19996 15960 20024 16068
rect 20162 16056 20168 16108
rect 20220 16096 20226 16108
rect 20717 16099 20775 16105
rect 20717 16096 20729 16099
rect 20220 16068 20729 16096
rect 20220 16056 20226 16068
rect 20717 16065 20729 16068
rect 20763 16065 20775 16099
rect 20717 16059 20775 16065
rect 20817 16099 20875 16105
rect 20817 16065 20829 16099
rect 20863 16065 20875 16099
rect 20916 16096 20944 16136
rect 21082 16124 21088 16136
rect 21140 16124 21146 16176
rect 20990 16096 20996 16108
rect 20916 16068 20996 16096
rect 20817 16059 20875 16065
rect 20073 16031 20131 16037
rect 20073 15997 20085 16031
rect 20119 16028 20131 16031
rect 20824 16028 20852 16059
rect 20990 16056 20996 16068
rect 21048 16056 21054 16108
rect 21100 16028 21128 16124
rect 21284 16105 21312 16204
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 20119 16000 20677 16028
rect 20824 16000 21128 16028
rect 20119 15997 20131 16000
rect 20073 15991 20131 15997
rect 20165 15963 20223 15969
rect 20165 15960 20177 15963
rect 19996 15932 20177 15960
rect 20165 15929 20177 15932
rect 20211 15929 20223 15963
rect 20346 15960 20352 15972
rect 20307 15932 20352 15960
rect 20165 15923 20223 15929
rect 14700 15864 17724 15892
rect 14700 15852 14706 15864
rect 17954 15852 17960 15904
rect 18012 15892 18018 15904
rect 18049 15895 18107 15901
rect 18049 15892 18061 15895
rect 18012 15864 18061 15892
rect 18012 15852 18018 15864
rect 18049 15861 18061 15864
rect 18095 15861 18107 15895
rect 18506 15892 18512 15904
rect 18467 15864 18512 15892
rect 18049 15855 18107 15861
rect 18506 15852 18512 15864
rect 18564 15852 18570 15904
rect 19518 15892 19524 15904
rect 19479 15864 19524 15892
rect 19518 15852 19524 15864
rect 19576 15852 19582 15904
rect 20180 15892 20208 15923
rect 20346 15920 20352 15932
rect 20404 15920 20410 15972
rect 20530 15892 20536 15904
rect 20180 15864 20536 15892
rect 20530 15852 20536 15864
rect 20588 15852 20594 15904
rect 20649 15892 20677 16000
rect 21910 15960 21916 15972
rect 21284 15932 21916 15960
rect 21284 15892 21312 15932
rect 21910 15920 21916 15932
rect 21968 15920 21974 15972
rect 21450 15892 21456 15904
rect 20649 15864 21312 15892
rect 21411 15864 21456 15892
rect 21450 15852 21456 15864
rect 21508 15852 21514 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 2222 15688 2228 15700
rect 2183 15660 2228 15688
rect 2222 15648 2228 15660
rect 2280 15648 2286 15700
rect 3234 15648 3240 15700
rect 3292 15688 3298 15700
rect 3973 15691 4031 15697
rect 3973 15688 3985 15691
rect 3292 15660 3985 15688
rect 3292 15648 3298 15660
rect 3620 15561 3648 15660
rect 3973 15657 3985 15660
rect 4019 15657 4031 15691
rect 3973 15651 4031 15657
rect 5445 15691 5503 15697
rect 5445 15657 5457 15691
rect 5491 15688 5503 15691
rect 5534 15688 5540 15700
rect 5491 15660 5540 15688
rect 5491 15657 5503 15660
rect 5445 15651 5503 15657
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 5626 15648 5632 15700
rect 5684 15688 5690 15700
rect 6178 15688 6184 15700
rect 5684 15660 6184 15688
rect 5684 15648 5690 15660
rect 6178 15648 6184 15660
rect 6236 15648 6242 15700
rect 8757 15691 8815 15697
rect 8757 15657 8769 15691
rect 8803 15688 8815 15691
rect 9122 15688 9128 15700
rect 8803 15660 9128 15688
rect 8803 15657 8815 15660
rect 8757 15651 8815 15657
rect 9122 15648 9128 15660
rect 9180 15648 9186 15700
rect 9401 15691 9459 15697
rect 9401 15657 9413 15691
rect 9447 15688 9459 15691
rect 9490 15688 9496 15700
rect 9447 15660 9496 15688
rect 9447 15657 9459 15660
rect 9401 15651 9459 15657
rect 4798 15580 4804 15632
rect 4856 15580 4862 15632
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 8941 15623 8999 15629
rect 8941 15620 8953 15623
rect 8720 15592 8953 15620
rect 8720 15580 8726 15592
rect 8941 15589 8953 15592
rect 8987 15589 8999 15623
rect 8941 15583 8999 15589
rect 3605 15555 3663 15561
rect 3605 15521 3617 15555
rect 3651 15521 3663 15555
rect 3605 15515 3663 15521
rect 4525 15555 4583 15561
rect 4525 15521 4537 15555
rect 4571 15552 4583 15555
rect 4816 15552 4844 15580
rect 7469 15555 7527 15561
rect 7469 15552 7481 15555
rect 4571 15524 4844 15552
rect 6748 15524 7481 15552
rect 4571 15521 4583 15524
rect 4525 15515 4583 15521
rect 1670 15484 1676 15496
rect 1631 15456 1676 15484
rect 1670 15444 1676 15456
rect 1728 15444 1734 15496
rect 2038 15484 2044 15496
rect 1999 15456 2044 15484
rect 2038 15444 2044 15456
rect 2096 15444 2102 15496
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4246 15484 4252 15496
rect 4203 15456 4252 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4246 15444 4252 15456
rect 4304 15444 4310 15496
rect 4614 15444 4620 15496
rect 4672 15484 4678 15496
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4672 15456 4813 15484
rect 4672 15444 4678 15456
rect 4801 15453 4813 15456
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 5810 15444 5816 15496
rect 5868 15484 5874 15496
rect 6270 15484 6276 15496
rect 5868 15456 6276 15484
rect 5868 15444 5874 15456
rect 6270 15444 6276 15456
rect 6328 15444 6334 15496
rect 6546 15444 6552 15496
rect 6604 15493 6610 15496
rect 6604 15484 6616 15493
rect 6748 15484 6776 15524
rect 7469 15521 7481 15524
rect 7515 15521 7527 15555
rect 7834 15552 7840 15564
rect 7469 15515 7527 15521
rect 7760 15524 7840 15552
rect 6604 15456 6776 15484
rect 6825 15487 6883 15493
rect 6604 15447 6616 15456
rect 6825 15453 6837 15487
rect 6871 15484 6883 15487
rect 7760 15484 7788 15524
rect 7834 15512 7840 15524
rect 7892 15512 7898 15564
rect 8205 15555 8263 15561
rect 8205 15521 8217 15555
rect 8251 15552 8263 15555
rect 8386 15552 8392 15564
rect 8251 15524 8392 15552
rect 8251 15521 8263 15524
rect 8205 15515 8263 15521
rect 8386 15512 8392 15524
rect 8444 15512 8450 15564
rect 9416 15552 9444 15651
rect 9490 15648 9496 15660
rect 9548 15648 9554 15700
rect 9582 15648 9588 15700
rect 9640 15648 9646 15700
rect 9766 15648 9772 15700
rect 9824 15688 9830 15700
rect 10413 15691 10471 15697
rect 10413 15688 10425 15691
rect 9824 15660 10425 15688
rect 9824 15648 9830 15660
rect 10413 15657 10425 15660
rect 10459 15657 10471 15691
rect 10413 15651 10471 15657
rect 12253 15691 12311 15697
rect 12253 15657 12265 15691
rect 12299 15688 12311 15691
rect 12342 15688 12348 15700
rect 12299 15660 12348 15688
rect 12299 15657 12311 15660
rect 12253 15651 12311 15657
rect 12342 15648 12348 15660
rect 12400 15648 12406 15700
rect 13170 15688 13176 15700
rect 13131 15660 13176 15688
rect 13170 15648 13176 15660
rect 13228 15648 13234 15700
rect 14461 15691 14519 15697
rect 14461 15657 14473 15691
rect 14507 15688 14519 15691
rect 14642 15688 14648 15700
rect 14507 15660 14648 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 14642 15648 14648 15660
rect 14700 15648 14706 15700
rect 15289 15691 15347 15697
rect 15289 15657 15301 15691
rect 15335 15688 15347 15691
rect 15378 15688 15384 15700
rect 15335 15660 15384 15688
rect 15335 15657 15347 15660
rect 15289 15651 15347 15657
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 16669 15691 16727 15697
rect 16669 15657 16681 15691
rect 16715 15688 16727 15691
rect 16758 15688 16764 15700
rect 16715 15660 16764 15688
rect 16715 15657 16727 15660
rect 16669 15651 16727 15657
rect 9600 15620 9628 15648
rect 12434 15620 12440 15632
rect 9600 15592 11008 15620
rect 9140 15524 9444 15552
rect 7926 15484 7932 15496
rect 6871 15456 7788 15484
rect 7887 15456 7932 15484
rect 6871 15453 6883 15456
rect 6825 15447 6883 15453
rect 6604 15444 6610 15447
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 9140 15493 9168 15524
rect 9582 15512 9588 15564
rect 9640 15552 9646 15564
rect 10980 15561 11008 15592
rect 11716 15592 12440 15620
rect 11716 15561 11744 15592
rect 12434 15580 12440 15592
rect 12492 15620 12498 15632
rect 13081 15623 13139 15629
rect 12492 15592 12572 15620
rect 12492 15580 12498 15592
rect 10137 15555 10195 15561
rect 10137 15552 10149 15555
rect 9640 15524 10149 15552
rect 9640 15512 9646 15524
rect 10137 15521 10149 15524
rect 10183 15521 10195 15555
rect 10137 15515 10195 15521
rect 10965 15555 11023 15561
rect 10965 15521 10977 15555
rect 11011 15521 11023 15555
rect 10965 15515 11023 15521
rect 11701 15555 11759 15561
rect 11701 15521 11713 15555
rect 11747 15521 11759 15555
rect 11701 15515 11759 15521
rect 11793 15555 11851 15561
rect 11793 15521 11805 15555
rect 11839 15552 11851 15555
rect 12250 15552 12256 15564
rect 11839 15524 12256 15552
rect 11839 15521 11851 15524
rect 11793 15515 11851 15521
rect 12250 15512 12256 15524
rect 12308 15512 12314 15564
rect 12544 15561 12572 15592
rect 13081 15589 13093 15623
rect 13127 15620 13139 15623
rect 13630 15620 13636 15632
rect 13127 15592 13636 15620
rect 13127 15589 13139 15592
rect 13081 15583 13139 15589
rect 13630 15580 13636 15592
rect 13688 15580 13694 15632
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15552 12587 15555
rect 13725 15555 13783 15561
rect 13725 15552 13737 15555
rect 12575 15524 13737 15552
rect 12575 15521 12587 15524
rect 12529 15515 12587 15521
rect 13725 15521 13737 15524
rect 13771 15521 13783 15555
rect 13725 15515 13783 15521
rect 14737 15555 14795 15561
rect 14737 15521 14749 15555
rect 14783 15552 14795 15555
rect 15102 15552 15108 15564
rect 14783 15524 15108 15552
rect 14783 15521 14795 15524
rect 14737 15515 14795 15521
rect 15102 15512 15108 15524
rect 15160 15512 15166 15564
rect 15286 15512 15292 15564
rect 15344 15552 15350 15564
rect 15473 15555 15531 15561
rect 15473 15552 15485 15555
rect 15344 15524 15485 15552
rect 15344 15512 15350 15524
rect 15473 15521 15485 15524
rect 15519 15521 15531 15555
rect 15473 15515 15531 15521
rect 9125 15487 9183 15493
rect 9125 15453 9137 15487
rect 9171 15453 9183 15487
rect 9125 15447 9183 15453
rect 9217 15487 9275 15493
rect 9217 15453 9229 15487
rect 9263 15484 9275 15487
rect 9858 15484 9864 15496
rect 9263 15456 9864 15484
rect 9263 15453 9275 15456
rect 9217 15447 9275 15453
rect 9858 15444 9864 15456
rect 9916 15444 9922 15496
rect 10502 15444 10508 15496
rect 10560 15484 10566 15496
rect 11885 15487 11943 15493
rect 10560 15456 11836 15484
rect 10560 15444 10566 15456
rect 3360 15419 3418 15425
rect 3360 15385 3372 15419
rect 3406 15416 3418 15419
rect 4632 15416 4660 15444
rect 3406 15388 4660 15416
rect 3406 15385 3418 15388
rect 3360 15379 3418 15385
rect 6454 15376 6460 15428
rect 6512 15416 6518 15428
rect 8389 15419 8447 15425
rect 6512 15388 6960 15416
rect 6512 15376 6518 15388
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 1854 15348 1860 15360
rect 1815 15320 1860 15348
rect 1854 15308 1860 15320
rect 1912 15308 1918 15360
rect 2682 15308 2688 15360
rect 2740 15348 2746 15360
rect 3789 15351 3847 15357
rect 3789 15348 3801 15351
rect 2740 15320 3801 15348
rect 2740 15308 2746 15320
rect 3789 15317 3801 15320
rect 3835 15317 3847 15351
rect 3789 15311 3847 15317
rect 4433 15351 4491 15357
rect 4433 15317 4445 15351
rect 4479 15348 4491 15351
rect 4706 15348 4712 15360
rect 4479 15320 4712 15348
rect 4479 15317 4491 15320
rect 4433 15311 4491 15317
rect 4706 15308 4712 15320
rect 4764 15308 4770 15360
rect 5074 15308 5080 15360
rect 5132 15348 5138 15360
rect 5534 15348 5540 15360
rect 5132 15320 5540 15348
rect 5132 15308 5138 15320
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 6932 15357 6960 15388
rect 8389 15385 8401 15419
rect 8435 15416 8447 15419
rect 11241 15419 11299 15425
rect 11241 15416 11253 15419
rect 8435 15388 9628 15416
rect 8435 15385 8447 15388
rect 8389 15379 8447 15385
rect 6917 15351 6975 15357
rect 6917 15317 6929 15351
rect 6963 15317 6975 15351
rect 7282 15348 7288 15360
rect 7243 15320 7288 15348
rect 6917 15311 6975 15317
rect 7282 15308 7288 15320
rect 7340 15308 7346 15360
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 7742 15348 7748 15360
rect 7432 15320 7477 15348
rect 7703 15320 7748 15348
rect 7432 15308 7438 15320
rect 7742 15308 7748 15320
rect 7800 15308 7806 15360
rect 8294 15348 8300 15360
rect 8255 15320 8300 15348
rect 8294 15308 8300 15320
rect 8352 15308 8358 15360
rect 9600 15357 9628 15388
rect 9968 15388 11253 15416
rect 9585 15351 9643 15357
rect 9585 15317 9597 15351
rect 9631 15317 9643 15351
rect 9585 15311 9643 15317
rect 9766 15308 9772 15360
rect 9824 15348 9830 15360
rect 9968 15357 9996 15388
rect 11241 15385 11253 15388
rect 11287 15385 11299 15419
rect 11808 15416 11836 15456
rect 11885 15453 11897 15487
rect 11931 15484 11943 15487
rect 12158 15484 12164 15496
rect 11931 15456 12164 15484
rect 11931 15453 11943 15456
rect 11885 15447 11943 15453
rect 12158 15444 12164 15456
rect 12216 15444 12222 15496
rect 14366 15484 14372 15496
rect 13464 15456 14372 15484
rect 13464 15416 13492 15456
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14918 15484 14924 15496
rect 14879 15456 14924 15484
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 15654 15444 15660 15496
rect 15712 15484 15718 15496
rect 16209 15487 16267 15493
rect 16209 15484 16221 15487
rect 15712 15456 16221 15484
rect 15712 15444 15718 15456
rect 16209 15453 16221 15456
rect 16255 15484 16267 15487
rect 16390 15484 16396 15496
rect 16255 15456 16396 15484
rect 16255 15453 16267 15456
rect 16209 15447 16267 15453
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16577 15487 16635 15493
rect 16577 15453 16589 15487
rect 16623 15484 16635 15487
rect 16684 15484 16712 15651
rect 16758 15648 16764 15660
rect 16816 15648 16822 15700
rect 17221 15691 17279 15697
rect 17221 15657 17233 15691
rect 17267 15688 17279 15691
rect 17402 15688 17408 15700
rect 17267 15660 17408 15688
rect 17267 15657 17279 15660
rect 17221 15651 17279 15657
rect 17402 15648 17408 15660
rect 17460 15648 17466 15700
rect 17494 15648 17500 15700
rect 17552 15688 17558 15700
rect 18966 15688 18972 15700
rect 17552 15660 18972 15688
rect 17552 15648 17558 15660
rect 18966 15648 18972 15660
rect 19024 15648 19030 15700
rect 19058 15648 19064 15700
rect 19116 15688 19122 15700
rect 19521 15691 19579 15697
rect 19116 15660 19161 15688
rect 19116 15648 19122 15660
rect 19521 15657 19533 15691
rect 19567 15688 19579 15691
rect 19978 15688 19984 15700
rect 19567 15660 19984 15688
rect 19567 15657 19579 15660
rect 19521 15651 19579 15657
rect 19978 15648 19984 15660
rect 20036 15648 20042 15700
rect 20162 15688 20168 15700
rect 20123 15660 20168 15688
rect 20162 15648 20168 15660
rect 20220 15648 20226 15700
rect 20254 15648 20260 15700
rect 20312 15688 20318 15700
rect 20349 15691 20407 15697
rect 20349 15688 20361 15691
rect 20312 15660 20361 15688
rect 20312 15648 20318 15660
rect 20349 15657 20361 15660
rect 20395 15657 20407 15691
rect 20349 15651 20407 15657
rect 20809 15691 20867 15697
rect 20809 15657 20821 15691
rect 20855 15688 20867 15691
rect 21266 15688 21272 15700
rect 20855 15660 21272 15688
rect 20855 15657 20867 15660
rect 20809 15651 20867 15657
rect 21266 15648 21272 15660
rect 21324 15648 21330 15700
rect 17313 15623 17371 15629
rect 17313 15589 17325 15623
rect 17359 15589 17371 15623
rect 17420 15620 17448 15648
rect 18693 15623 18751 15629
rect 17420 15592 17724 15620
rect 17313 15583 17371 15589
rect 17328 15552 17356 15583
rect 17402 15552 17408 15564
rect 17328 15524 17408 15552
rect 16623 15456 16712 15484
rect 16853 15487 16911 15493
rect 16623 15453 16635 15456
rect 16577 15447 16635 15453
rect 16853 15453 16865 15487
rect 16899 15484 16911 15487
rect 17328 15484 17356 15524
rect 17402 15512 17408 15524
rect 17460 15552 17466 15564
rect 17696 15552 17724 15592
rect 18693 15589 18705 15623
rect 18739 15620 18751 15623
rect 18739 15592 19656 15620
rect 18739 15589 18751 15592
rect 18693 15583 18751 15589
rect 19628 15564 19656 15592
rect 19886 15580 19892 15632
rect 19944 15620 19950 15632
rect 22370 15620 22376 15632
rect 19944 15592 22376 15620
rect 19944 15580 19950 15592
rect 22370 15580 22376 15592
rect 22428 15580 22434 15632
rect 17862 15552 17868 15564
rect 17460 15524 17632 15552
rect 17696 15524 17868 15552
rect 17460 15512 17466 15524
rect 17494 15484 17500 15496
rect 16899 15456 17356 15484
rect 17455 15456 17500 15484
rect 16899 15453 16911 15456
rect 16853 15447 16911 15453
rect 17494 15444 17500 15456
rect 17552 15444 17558 15496
rect 17604 15493 17632 15524
rect 17862 15512 17868 15524
rect 17920 15512 17926 15564
rect 18141 15555 18199 15561
rect 18141 15521 18153 15555
rect 18187 15552 18199 15555
rect 18414 15552 18420 15564
rect 18187 15524 18420 15552
rect 18187 15521 18199 15524
rect 18141 15515 18199 15521
rect 18414 15512 18420 15524
rect 18472 15512 18478 15564
rect 19610 15512 19616 15564
rect 19668 15512 19674 15564
rect 19794 15512 19800 15564
rect 19852 15552 19858 15564
rect 22002 15552 22008 15564
rect 19852 15524 22008 15552
rect 19852 15512 19858 15524
rect 22002 15512 22008 15524
rect 22060 15512 22066 15564
rect 17589 15487 17647 15493
rect 17589 15453 17601 15487
rect 17635 15453 17647 15487
rect 17589 15447 17647 15453
rect 17696 15456 17991 15484
rect 11808 15388 13492 15416
rect 13541 15419 13599 15425
rect 11241 15379 11299 15385
rect 13541 15385 13553 15419
rect 13587 15416 13599 15419
rect 14093 15419 14151 15425
rect 14093 15416 14105 15419
rect 13587 15388 14105 15416
rect 13587 15385 13599 15388
rect 13541 15379 13599 15385
rect 14093 15385 14105 15388
rect 14139 15385 14151 15419
rect 14093 15379 14151 15385
rect 14274 15376 14280 15428
rect 14332 15416 14338 15428
rect 15749 15419 15807 15425
rect 15749 15416 15761 15419
rect 14332 15388 15761 15416
rect 14332 15376 14338 15388
rect 15749 15385 15761 15388
rect 15795 15416 15807 15419
rect 16945 15419 17003 15425
rect 16945 15416 16957 15419
rect 15795 15388 16957 15416
rect 15795 15385 15807 15388
rect 15749 15379 15807 15385
rect 16945 15385 16957 15388
rect 16991 15416 17003 15419
rect 17696 15416 17724 15456
rect 16991 15388 17724 15416
rect 17963 15416 17991 15456
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18325 15487 18383 15493
rect 18325 15484 18337 15487
rect 18288 15456 18337 15484
rect 18288 15444 18294 15456
rect 18325 15453 18337 15456
rect 18371 15453 18383 15487
rect 18325 15447 18383 15453
rect 19334 15444 19340 15496
rect 19392 15484 19398 15496
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19392 15456 19993 15484
rect 19392 15444 19398 15456
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 20530 15484 20536 15496
rect 20491 15456 20536 15484
rect 19981 15447 20039 15453
rect 20530 15444 20536 15456
rect 20588 15444 20594 15496
rect 20625 15487 20683 15493
rect 20625 15453 20637 15487
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 19613 15419 19671 15425
rect 19613 15416 19625 15419
rect 17963 15388 19625 15416
rect 16991 15385 17003 15388
rect 16945 15379 17003 15385
rect 19613 15385 19625 15388
rect 19659 15416 19671 15419
rect 20640 15416 20668 15447
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 20901 15487 20959 15493
rect 20901 15484 20913 15487
rect 20772 15456 20913 15484
rect 20772 15444 20778 15456
rect 20901 15453 20913 15456
rect 20947 15453 20959 15487
rect 21266 15484 21272 15496
rect 21227 15456 21272 15484
rect 20901 15447 20959 15453
rect 21266 15444 21272 15456
rect 21324 15444 21330 15496
rect 19659 15388 20668 15416
rect 19659 15385 19671 15388
rect 19613 15379 19671 15385
rect 20990 15376 20996 15428
rect 21048 15416 21054 15428
rect 22186 15416 22192 15428
rect 21048 15388 22192 15416
rect 21048 15376 21054 15388
rect 22186 15376 22192 15388
rect 22244 15376 22250 15428
rect 9953 15351 10011 15357
rect 9953 15348 9965 15351
rect 9824 15320 9965 15348
rect 9824 15308 9830 15320
rect 9953 15317 9965 15320
rect 9999 15317 10011 15351
rect 9953 15311 10011 15317
rect 10042 15308 10048 15360
rect 10100 15348 10106 15360
rect 10100 15320 10145 15348
rect 10100 15308 10106 15320
rect 10318 15308 10324 15360
rect 10376 15348 10382 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 10376 15320 10793 15348
rect 10376 15308 10382 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10781 15311 10839 15317
rect 10870 15308 10876 15360
rect 10928 15348 10934 15360
rect 12618 15348 12624 15360
rect 10928 15320 10973 15348
rect 12579 15320 12624 15348
rect 10928 15308 10934 15320
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 12713 15351 12771 15357
rect 12713 15317 12725 15351
rect 12759 15348 12771 15351
rect 13354 15348 13360 15360
rect 12759 15320 13360 15348
rect 12759 15317 12771 15320
rect 12713 15311 12771 15317
rect 13354 15308 13360 15320
rect 13412 15308 13418 15360
rect 13633 15351 13691 15357
rect 13633 15317 13645 15351
rect 13679 15348 13691 15351
rect 14642 15348 14648 15360
rect 13679 15320 14648 15348
rect 13679 15317 13691 15320
rect 13633 15311 13691 15317
rect 14642 15308 14648 15320
rect 14700 15308 14706 15360
rect 14826 15348 14832 15360
rect 14787 15320 14832 15348
rect 14826 15308 14832 15320
rect 14884 15308 14890 15360
rect 15194 15308 15200 15360
rect 15252 15348 15258 15360
rect 15654 15348 15660 15360
rect 15252 15320 15660 15348
rect 15252 15308 15258 15320
rect 15654 15308 15660 15320
rect 15712 15308 15718 15360
rect 16114 15348 16120 15360
rect 16075 15320 16120 15348
rect 16114 15308 16120 15320
rect 16172 15308 16178 15360
rect 16298 15308 16304 15360
rect 16356 15348 16362 15360
rect 16393 15351 16451 15357
rect 16393 15348 16405 15351
rect 16356 15320 16405 15348
rect 16356 15308 16362 15320
rect 16393 15317 16405 15320
rect 16439 15317 16451 15351
rect 17770 15348 17776 15360
rect 17731 15320 17776 15348
rect 16393 15311 16451 15317
rect 17770 15308 17776 15320
rect 17828 15308 17834 15360
rect 17862 15308 17868 15360
rect 17920 15348 17926 15360
rect 18233 15351 18291 15357
rect 18233 15348 18245 15351
rect 17920 15320 18245 15348
rect 17920 15308 17926 15320
rect 18233 15317 18245 15320
rect 18279 15317 18291 15351
rect 18233 15311 18291 15317
rect 18690 15308 18696 15360
rect 18748 15348 18754 15360
rect 18785 15351 18843 15357
rect 18785 15348 18797 15351
rect 18748 15320 18797 15348
rect 18748 15308 18754 15320
rect 18785 15317 18797 15320
rect 18831 15317 18843 15351
rect 18785 15311 18843 15317
rect 19337 15351 19395 15357
rect 19337 15317 19349 15351
rect 19383 15348 19395 15351
rect 19889 15351 19947 15357
rect 19889 15348 19901 15351
rect 19383 15320 19901 15348
rect 19383 15317 19395 15320
rect 19337 15311 19395 15317
rect 19889 15317 19901 15320
rect 19935 15348 19947 15351
rect 20806 15348 20812 15360
rect 19935 15320 20812 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20806 15308 20812 15320
rect 20864 15308 20870 15360
rect 21082 15348 21088 15360
rect 21043 15320 21088 15348
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21450 15348 21456 15360
rect 21411 15320 21456 15348
rect 21450 15308 21456 15320
rect 21508 15308 21514 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 1857 15147 1915 15153
rect 1857 15113 1869 15147
rect 1903 15113 1915 15147
rect 1857 15107 1915 15113
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1872 15008 1900 15107
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 2409 15147 2467 15153
rect 2409 15144 2421 15147
rect 2096 15116 2421 15144
rect 2096 15104 2102 15116
rect 2409 15113 2421 15116
rect 2455 15113 2467 15147
rect 2409 15107 2467 15113
rect 2590 15104 2596 15156
rect 2648 15104 2654 15156
rect 2777 15147 2835 15153
rect 2777 15113 2789 15147
rect 2823 15144 2835 15147
rect 2958 15144 2964 15156
rect 2823 15116 2964 15144
rect 2823 15113 2835 15116
rect 2777 15107 2835 15113
rect 2958 15104 2964 15116
rect 3016 15104 3022 15156
rect 3973 15147 4031 15153
rect 3973 15113 3985 15147
rect 4019 15144 4031 15147
rect 4062 15144 4068 15156
rect 4019 15116 4068 15144
rect 4019 15113 4031 15116
rect 3973 15107 4031 15113
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 4433 15147 4491 15153
rect 4433 15113 4445 15147
rect 4479 15144 4491 15147
rect 5166 15144 5172 15156
rect 4479 15116 5172 15144
rect 4479 15113 4491 15116
rect 4433 15107 4491 15113
rect 5166 15104 5172 15116
rect 5224 15104 5230 15156
rect 6181 15147 6239 15153
rect 6181 15113 6193 15147
rect 6227 15144 6239 15147
rect 6546 15144 6552 15156
rect 6227 15116 6552 15144
rect 6227 15113 6239 15116
rect 6181 15107 6239 15113
rect 6546 15104 6552 15116
rect 6604 15104 6610 15156
rect 6733 15147 6791 15153
rect 6733 15113 6745 15147
rect 6779 15144 6791 15147
rect 7926 15144 7932 15156
rect 6779 15116 7932 15144
rect 6779 15113 6791 15116
rect 6733 15107 6791 15113
rect 2608 15076 2636 15104
rect 2056 15048 2636 15076
rect 2056 15017 2084 15048
rect 4246 15036 4252 15088
rect 4304 15076 4310 15088
rect 6748 15076 6776 15107
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8389 15147 8447 15153
rect 8389 15113 8401 15147
rect 8435 15113 8447 15147
rect 8389 15107 8447 15113
rect 8404 15076 8432 15107
rect 8478 15104 8484 15156
rect 8536 15144 8542 15156
rect 8536 15116 8581 15144
rect 8536 15104 8542 15116
rect 8754 15104 8760 15156
rect 8812 15144 8818 15156
rect 9953 15147 10011 15153
rect 8812 15116 9904 15144
rect 8812 15104 8818 15116
rect 9582 15076 9588 15088
rect 9640 15085 9646 15088
rect 4304 15048 6776 15076
rect 7024 15048 7420 15076
rect 8404 15048 9588 15076
rect 4304 15036 4310 15048
rect 1719 14980 1900 15008
rect 2041 15011 2099 15017
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 2041 14977 2053 15011
rect 2087 14977 2099 15011
rect 2314 15008 2320 15020
rect 2275 14980 2320 15008
rect 2041 14971 2099 14977
rect 1578 14900 1584 14952
rect 1636 14940 1642 14952
rect 2056 14940 2084 14971
rect 2314 14968 2320 14980
rect 2372 14968 2378 15020
rect 2590 15008 2596 15020
rect 2551 14980 2596 15008
rect 2590 14968 2596 14980
rect 2648 14968 2654 15020
rect 4816 15017 4844 15048
rect 3145 15011 3203 15017
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 3605 15011 3663 15017
rect 3605 15008 3617 15011
rect 3191 14980 3617 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3605 14977 3617 14980
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4801 15011 4859 15017
rect 4387 14980 4752 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 3234 14940 3240 14952
rect 1636 14912 2084 14940
rect 3195 14912 3240 14940
rect 1636 14900 1642 14912
rect 3234 14900 3240 14912
rect 3292 14900 3298 14952
rect 3421 14943 3479 14949
rect 3421 14909 3433 14943
rect 3467 14909 3479 14943
rect 4614 14940 4620 14952
rect 4575 14912 4620 14940
rect 3421 14903 3479 14909
rect 1394 14832 1400 14884
rect 1452 14872 1458 14884
rect 1452 14844 1624 14872
rect 1452 14832 1458 14844
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 1596 14804 1624 14844
rect 1670 14832 1676 14884
rect 1728 14872 1734 14884
rect 2133 14875 2191 14881
rect 2133 14872 2145 14875
rect 1728 14844 2145 14872
rect 1728 14832 1734 14844
rect 2133 14841 2145 14844
rect 2179 14841 2191 14875
rect 3436 14872 3464 14903
rect 4614 14900 4620 14912
rect 4672 14900 4678 14952
rect 4154 14872 4160 14884
rect 3436 14844 4160 14872
rect 2133 14835 2191 14841
rect 4154 14832 4160 14844
rect 4212 14872 4218 14884
rect 4632 14872 4660 14900
rect 4212 14844 4660 14872
rect 4724 14872 4752 14980
rect 4801 14977 4813 15011
rect 4847 14977 4859 15011
rect 4801 14971 4859 14977
rect 5068 15011 5126 15017
rect 5068 14977 5080 15011
rect 5114 15008 5126 15011
rect 6730 15008 6736 15020
rect 5114 14980 6736 15008
rect 5114 14977 5126 14980
rect 5068 14971 5126 14977
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 7024 15017 7052 15048
rect 6917 15011 6975 15017
rect 6917 14977 6929 15011
rect 6963 15008 6975 15011
rect 7009 15011 7067 15017
rect 7009 15008 7021 15011
rect 6963 14980 7021 15008
rect 6963 14977 6975 14980
rect 6917 14971 6975 14977
rect 7009 14977 7021 14980
rect 7055 14977 7067 15011
rect 7009 14971 7067 14977
rect 7098 14968 7104 15020
rect 7156 15008 7162 15020
rect 7265 15011 7323 15017
rect 7265 15008 7277 15011
rect 7156 14980 7277 15008
rect 7156 14968 7162 14980
rect 7265 14977 7277 14980
rect 7311 14977 7323 15011
rect 7392 15008 7420 15048
rect 9582 15036 9588 15048
rect 9640 15076 9652 15085
rect 9876 15076 9904 15116
rect 9953 15113 9965 15147
rect 9999 15144 10011 15147
rect 10042 15144 10048 15156
rect 9999 15116 10048 15144
rect 9999 15113 10011 15116
rect 9953 15107 10011 15113
rect 10042 15104 10048 15116
rect 10100 15104 10106 15156
rect 10321 15147 10379 15153
rect 10321 15144 10333 15147
rect 10152 15116 10333 15144
rect 10152 15076 10180 15116
rect 10321 15113 10333 15116
rect 10367 15144 10379 15147
rect 10410 15144 10416 15156
rect 10367 15116 10416 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 10410 15104 10416 15116
rect 10468 15104 10474 15156
rect 10594 15104 10600 15156
rect 10652 15144 10658 15156
rect 10652 15116 11560 15144
rect 10652 15104 10658 15116
rect 11054 15076 11060 15088
rect 9640 15048 9685 15076
rect 9876 15048 10180 15076
rect 10244 15048 11060 15076
rect 9640 15039 9652 15048
rect 9640 15036 9646 15039
rect 8662 15008 8668 15020
rect 7392 14980 8668 15008
rect 7265 14971 7323 14977
rect 8662 14968 8668 14980
rect 8720 14968 8726 15020
rect 10244 15008 10272 15048
rect 11054 15036 11060 15048
rect 11112 15036 11118 15088
rect 8864 14980 10272 15008
rect 10413 15011 10471 15017
rect 8018 14900 8024 14952
rect 8076 14940 8082 14952
rect 8864 14940 8892 14980
rect 10413 14977 10425 15011
rect 10459 15008 10471 15011
rect 10962 15008 10968 15020
rect 10459 14980 10968 15008
rect 10459 14977 10471 14980
rect 10413 14971 10471 14977
rect 9858 14940 9864 14952
rect 8076 14912 8892 14940
rect 9819 14912 9864 14940
rect 8076 14900 8082 14912
rect 9858 14900 9864 14912
rect 9916 14900 9922 14952
rect 10042 14900 10048 14952
rect 10100 14940 10106 14952
rect 10428 14940 10456 14971
rect 10962 14968 10968 14980
rect 11020 14968 11026 15020
rect 11532 14952 11560 15116
rect 12618 15104 12624 15156
rect 12676 15144 12682 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12676 15116 13001 15144
rect 12676 15104 12682 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 14001 15147 14059 15153
rect 14001 15144 14013 15147
rect 13412 15116 14013 15144
rect 13412 15104 13418 15116
rect 14001 15113 14013 15116
rect 14047 15113 14059 15147
rect 14001 15107 14059 15113
rect 14921 15147 14979 15153
rect 14921 15113 14933 15147
rect 14967 15144 14979 15147
rect 15381 15147 15439 15153
rect 15381 15144 15393 15147
rect 14967 15116 15393 15144
rect 14967 15113 14979 15116
rect 14921 15107 14979 15113
rect 15381 15113 15393 15116
rect 15427 15113 15439 15147
rect 15381 15107 15439 15113
rect 15841 15147 15899 15153
rect 15841 15113 15853 15147
rect 15887 15144 15899 15147
rect 16114 15144 16120 15156
rect 15887 15116 16120 15144
rect 15887 15113 15899 15116
rect 15841 15107 15899 15113
rect 11784 15079 11842 15085
rect 11784 15045 11796 15079
rect 11830 15076 11842 15079
rect 12710 15076 12716 15088
rect 11830 15048 12716 15076
rect 11830 15045 11842 15048
rect 11784 15039 11842 15045
rect 12710 15036 12716 15048
rect 12768 15076 12774 15088
rect 14016 15076 14044 15107
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 17586 15104 17592 15156
rect 17644 15144 17650 15156
rect 18874 15144 18880 15156
rect 17644 15116 18880 15144
rect 17644 15104 17650 15116
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 20441 15147 20499 15153
rect 20441 15113 20453 15147
rect 20487 15144 20499 15147
rect 20714 15144 20720 15156
rect 20487 15116 20720 15144
rect 20487 15113 20499 15116
rect 20441 15107 20499 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 15194 15076 15200 15088
rect 12768 15048 13492 15076
rect 14016 15048 15200 15076
rect 12768 15036 12774 15048
rect 13354 15008 13360 15020
rect 13315 14980 13360 15008
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13464 15008 13492 15048
rect 15194 15036 15200 15048
rect 15252 15036 15258 15088
rect 19334 15076 19340 15088
rect 15304 15048 19340 15076
rect 13464 14980 13584 15008
rect 10100 14912 10456 14940
rect 10597 14943 10655 14949
rect 10100 14900 10106 14912
rect 10597 14909 10609 14943
rect 10643 14909 10655 14943
rect 10597 14903 10655 14909
rect 10781 14943 10839 14949
rect 10781 14909 10793 14943
rect 10827 14940 10839 14943
rect 11514 14940 11520 14952
rect 10827 14912 10916 14940
rect 11427 14912 11520 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 4798 14872 4804 14884
rect 4724 14844 4804 14872
rect 4212 14832 4218 14844
rect 4798 14832 4804 14844
rect 4856 14832 4862 14884
rect 6086 14832 6092 14884
rect 6144 14872 6150 14884
rect 7006 14872 7012 14884
rect 6144 14844 7012 14872
rect 6144 14832 6150 14844
rect 7006 14832 7012 14844
rect 7064 14832 7070 14884
rect 10612 14816 10640 14903
rect 5994 14804 6000 14816
rect 1596 14776 6000 14804
rect 5994 14764 6000 14776
rect 6052 14804 6058 14816
rect 6365 14807 6423 14813
rect 6365 14804 6377 14807
rect 6052 14776 6377 14804
rect 6052 14764 6058 14776
rect 6365 14773 6377 14776
rect 6411 14773 6423 14807
rect 6638 14804 6644 14816
rect 6599 14776 6644 14804
rect 6365 14767 6423 14773
rect 6638 14764 6644 14776
rect 6696 14764 6702 14816
rect 7190 14764 7196 14816
rect 7248 14804 7254 14816
rect 10594 14804 10600 14816
rect 7248 14776 10600 14804
rect 7248 14764 7254 14776
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 10778 14764 10784 14816
rect 10836 14804 10842 14816
rect 10888 14804 10916 14912
rect 11514 14900 11520 14912
rect 11572 14900 11578 14952
rect 13262 14900 13268 14952
rect 13320 14940 13326 14952
rect 13556 14949 13584 14980
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13320 14912 13461 14940
rect 13320 14900 13326 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13541 14943 13599 14949
rect 13541 14909 13553 14943
rect 13587 14909 13599 14943
rect 14458 14940 14464 14952
rect 13541 14903 13599 14909
rect 14292 14912 14464 14940
rect 13464 14872 13492 14903
rect 14185 14875 14243 14881
rect 14185 14872 14197 14875
rect 13464 14844 14197 14872
rect 14185 14841 14197 14844
rect 14231 14841 14243 14875
rect 14185 14835 14243 14841
rect 10836 14776 10916 14804
rect 10836 14764 10842 14776
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11057 14807 11115 14813
rect 11057 14804 11069 14807
rect 11020 14776 11069 14804
rect 11020 14764 11026 14776
rect 11057 14773 11069 14776
rect 11103 14773 11115 14807
rect 11057 14767 11115 14773
rect 11333 14807 11391 14813
rect 11333 14773 11345 14807
rect 11379 14804 11391 14807
rect 11422 14804 11428 14816
rect 11379 14776 11428 14804
rect 11379 14773 11391 14776
rect 11333 14767 11391 14773
rect 11422 14764 11428 14776
rect 11480 14764 11486 14816
rect 12434 14764 12440 14816
rect 12492 14804 12498 14816
rect 12897 14807 12955 14813
rect 12897 14804 12909 14807
rect 12492 14776 12909 14804
rect 12492 14764 12498 14776
rect 12897 14773 12909 14776
rect 12943 14773 12955 14807
rect 12897 14767 12955 14773
rect 13354 14764 13360 14816
rect 13412 14804 13418 14816
rect 13722 14804 13728 14816
rect 13412 14776 13728 14804
rect 13412 14764 13418 14776
rect 13722 14764 13728 14776
rect 13780 14804 13786 14816
rect 13817 14807 13875 14813
rect 13817 14804 13829 14807
rect 13780 14776 13829 14804
rect 13780 14764 13786 14776
rect 13817 14773 13829 14776
rect 13863 14804 13875 14807
rect 14292 14804 14320 14912
rect 14458 14900 14464 14912
rect 14516 14900 14522 14952
rect 14734 14940 14740 14952
rect 14695 14912 14740 14940
rect 14734 14900 14740 14912
rect 14792 14900 14798 14952
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 15194 14940 15200 14952
rect 14875 14912 15200 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 15194 14900 15200 14912
rect 15252 14900 15258 14952
rect 15304 14881 15332 15048
rect 19334 15036 19340 15048
rect 19392 15036 19398 15088
rect 21085 15079 21143 15085
rect 21085 15076 21097 15079
rect 20548 15048 21097 15076
rect 15746 15008 15752 15020
rect 15707 14980 15752 15008
rect 15746 14968 15752 14980
rect 15804 14968 15810 15020
rect 17793 15011 17851 15017
rect 17793 14977 17805 15011
rect 17839 15008 17851 15011
rect 18230 15008 18236 15020
rect 17839 14980 18236 15008
rect 17839 14977 17851 14980
rect 17793 14971 17851 14977
rect 18230 14968 18236 14980
rect 18288 14968 18294 15020
rect 18414 15017 18420 15020
rect 18408 15008 18420 15017
rect 18375 14980 18420 15008
rect 18408 14971 18420 14980
rect 18472 15008 18478 15020
rect 18966 15008 18972 15020
rect 18472 14980 18972 15008
rect 18414 14968 18420 14971
rect 18472 14968 18478 14980
rect 18966 14968 18972 14980
rect 19024 14968 19030 15020
rect 19978 15008 19984 15020
rect 19939 14980 19984 15008
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20257 15011 20315 15017
rect 20257 15008 20269 15011
rect 20180 14980 20269 15008
rect 15930 14940 15936 14952
rect 15891 14912 15936 14940
rect 15930 14900 15936 14912
rect 15988 14900 15994 14952
rect 16390 14940 16396 14952
rect 16351 14912 16396 14940
rect 16390 14900 16396 14912
rect 16448 14900 16454 14952
rect 18049 14943 18107 14949
rect 18049 14909 18061 14943
rect 18095 14940 18107 14943
rect 18141 14943 18199 14949
rect 18141 14940 18153 14943
rect 18095 14912 18153 14940
rect 18095 14909 18107 14912
rect 18049 14903 18107 14909
rect 18141 14909 18153 14912
rect 18187 14909 18199 14943
rect 19794 14940 19800 14952
rect 19755 14912 19800 14940
rect 18141 14903 18199 14909
rect 15289 14875 15347 14881
rect 15289 14841 15301 14875
rect 15335 14841 15347 14875
rect 15289 14835 15347 14841
rect 14458 14804 14464 14816
rect 13863 14776 14320 14804
rect 14419 14776 14464 14804
rect 13863 14773 13875 14776
rect 13817 14767 13875 14773
rect 14458 14764 14464 14776
rect 14516 14804 14522 14816
rect 14826 14804 14832 14816
rect 14516 14776 14832 14804
rect 14516 14764 14522 14776
rect 14826 14764 14832 14776
rect 14884 14764 14890 14816
rect 16669 14807 16727 14813
rect 16669 14773 16681 14807
rect 16715 14804 16727 14807
rect 16942 14804 16948 14816
rect 16715 14776 16948 14804
rect 16715 14773 16727 14776
rect 16669 14767 16727 14773
rect 16942 14764 16948 14776
rect 17000 14764 17006 14816
rect 17402 14764 17408 14816
rect 17460 14804 17466 14816
rect 18064 14804 18092 14903
rect 19794 14900 19800 14912
rect 19852 14900 19858 14952
rect 20180 14881 20208 14980
rect 20257 14977 20269 14980
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20438 14968 20444 15020
rect 20496 15008 20502 15020
rect 20548 15017 20576 15048
rect 21085 15045 21097 15048
rect 21131 15045 21143 15079
rect 21085 15039 21143 15045
rect 20533 15011 20591 15017
rect 20533 15008 20545 15011
rect 20496 14980 20545 15008
rect 20496 14968 20502 14980
rect 20533 14977 20545 14980
rect 20579 14977 20591 15011
rect 20806 15008 20812 15020
rect 20719 14980 20812 15008
rect 20533 14971 20591 14977
rect 20806 14968 20812 14980
rect 20864 14968 20870 15020
rect 21174 14968 21180 15020
rect 21232 15008 21238 15020
rect 21269 15011 21327 15017
rect 21269 15008 21281 15011
rect 21232 14980 21281 15008
rect 21232 14968 21238 14980
rect 21269 14977 21281 14980
rect 21315 14977 21327 15011
rect 21269 14971 21327 14977
rect 20824 14940 20852 14968
rect 22738 14940 22744 14952
rect 20824 14912 22744 14940
rect 22738 14900 22744 14912
rect 22796 14900 22802 14952
rect 20165 14875 20223 14881
rect 20165 14841 20177 14875
rect 20211 14841 20223 14875
rect 20165 14835 20223 14841
rect 20717 14875 20775 14881
rect 20717 14841 20729 14875
rect 20763 14872 20775 14875
rect 21266 14872 21272 14884
rect 20763 14844 21272 14872
rect 20763 14841 20775 14844
rect 20717 14835 20775 14841
rect 21266 14832 21272 14844
rect 21324 14832 21330 14884
rect 17460 14776 18092 14804
rect 19521 14807 19579 14813
rect 17460 14764 17466 14776
rect 19521 14773 19533 14807
rect 19567 14804 19579 14807
rect 19886 14804 19892 14816
rect 19567 14776 19892 14804
rect 19567 14773 19579 14776
rect 19521 14767 19579 14773
rect 19886 14764 19892 14776
rect 19944 14764 19950 14816
rect 20990 14804 20996 14816
rect 20951 14776 20996 14804
rect 20990 14764 20996 14776
rect 21048 14764 21054 14816
rect 21450 14804 21456 14816
rect 21411 14776 21456 14804
rect 21450 14764 21456 14776
rect 21508 14764 21514 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 2777 14603 2835 14609
rect 2777 14569 2789 14603
rect 2823 14600 2835 14603
rect 3050 14600 3056 14612
rect 2823 14572 3056 14600
rect 2823 14569 2835 14572
rect 2777 14563 2835 14569
rect 3050 14560 3056 14572
rect 3108 14560 3114 14612
rect 3973 14603 4031 14609
rect 3973 14569 3985 14603
rect 4019 14600 4031 14603
rect 4522 14600 4528 14612
rect 4019 14572 4528 14600
rect 4019 14569 4031 14572
rect 3973 14563 4031 14569
rect 4522 14560 4528 14572
rect 4580 14560 4586 14612
rect 4798 14560 4804 14612
rect 4856 14600 4862 14612
rect 5169 14603 5227 14609
rect 5169 14600 5181 14603
rect 4856 14572 5181 14600
rect 4856 14560 4862 14572
rect 5169 14569 5181 14572
rect 5215 14600 5227 14603
rect 5258 14600 5264 14612
rect 5215 14572 5264 14600
rect 5215 14569 5227 14572
rect 5169 14563 5227 14569
rect 5258 14560 5264 14572
rect 5316 14560 5322 14612
rect 5718 14560 5724 14612
rect 5776 14600 5782 14612
rect 5997 14603 6055 14609
rect 5997 14600 6009 14603
rect 5776 14572 6009 14600
rect 5776 14560 5782 14572
rect 5997 14569 6009 14572
rect 6043 14569 6055 14603
rect 5997 14563 6055 14569
rect 6638 14560 6644 14612
rect 6696 14600 6702 14612
rect 9953 14603 10011 14609
rect 6696 14572 8432 14600
rect 6696 14560 6702 14572
rect 2958 14492 2964 14544
rect 3016 14532 3022 14544
rect 6822 14532 6828 14544
rect 3016 14504 6828 14532
rect 3016 14492 3022 14504
rect 6822 14492 6828 14504
rect 6880 14492 6886 14544
rect 7101 14535 7159 14541
rect 7101 14501 7113 14535
rect 7147 14532 7159 14535
rect 8202 14532 8208 14544
rect 7147 14504 8208 14532
rect 7147 14501 7159 14504
rect 7101 14495 7159 14501
rect 8202 14492 8208 14504
rect 8260 14492 8266 14544
rect 106 14424 112 14476
rect 164 14464 170 14476
rect 3421 14467 3479 14473
rect 164 14436 3372 14464
rect 164 14424 170 14436
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 1857 14399 1915 14405
rect 1857 14365 1869 14399
rect 1903 14396 1915 14399
rect 2222 14396 2228 14408
rect 1903 14368 2228 14396
rect 1903 14365 1915 14368
rect 1857 14359 1915 14365
rect 1688 14328 1716 14359
rect 2222 14356 2228 14368
rect 2280 14356 2286 14408
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2682 14396 2688 14408
rect 2639 14368 2688 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2332 14328 2360 14359
rect 2682 14356 2688 14368
rect 2740 14356 2746 14408
rect 3344 14396 3372 14436
rect 3421 14433 3433 14467
rect 3467 14464 3479 14467
rect 4154 14464 4160 14476
rect 3467 14436 4160 14464
rect 3467 14433 3479 14436
rect 3421 14427 3479 14433
rect 4154 14424 4160 14436
rect 4212 14424 4218 14476
rect 4709 14467 4767 14473
rect 4709 14433 4721 14467
rect 4755 14464 4767 14467
rect 5902 14464 5908 14476
rect 4755 14436 5908 14464
rect 4755 14433 4767 14436
rect 4709 14427 4767 14433
rect 5902 14424 5908 14436
rect 5960 14424 5966 14476
rect 6546 14464 6552 14476
rect 6507 14436 6552 14464
rect 6546 14424 6552 14436
rect 6604 14424 6610 14476
rect 6730 14424 6736 14476
rect 6788 14464 6794 14476
rect 7837 14467 7895 14473
rect 7837 14464 7849 14467
rect 6788 14436 7849 14464
rect 6788 14424 6794 14436
rect 7837 14433 7849 14436
rect 7883 14464 7895 14467
rect 8018 14464 8024 14476
rect 7883 14436 8024 14464
rect 7883 14433 7895 14436
rect 7837 14427 7895 14433
rect 8018 14424 8024 14436
rect 8076 14424 8082 14476
rect 8404 14464 8432 14572
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10870 14600 10876 14612
rect 9999 14572 10876 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10870 14560 10876 14572
rect 10928 14560 10934 14612
rect 11790 14600 11796 14612
rect 10980 14572 11796 14600
rect 8478 14492 8484 14544
rect 8536 14532 8542 14544
rect 10980 14532 11008 14572
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 11885 14603 11943 14609
rect 11885 14569 11897 14603
rect 11931 14600 11943 14603
rect 12158 14600 12164 14612
rect 11931 14572 12164 14600
rect 11931 14569 11943 14572
rect 11885 14563 11943 14569
rect 12158 14560 12164 14572
rect 12216 14560 12222 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12342 14600 12348 14612
rect 12299 14572 12348 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12342 14560 12348 14572
rect 12400 14600 12406 14612
rect 12618 14600 12624 14612
rect 12400 14572 12624 14600
rect 12400 14560 12406 14572
rect 12618 14560 12624 14572
rect 12676 14560 12682 14612
rect 13081 14603 13139 14609
rect 13081 14569 13093 14603
rect 13127 14600 13139 14603
rect 13446 14600 13452 14612
rect 13127 14572 13452 14600
rect 13127 14569 13139 14572
rect 13081 14563 13139 14569
rect 13446 14560 13452 14572
rect 13504 14560 13510 14612
rect 14093 14603 14151 14609
rect 14093 14569 14105 14603
rect 14139 14600 14151 14603
rect 15930 14600 15936 14612
rect 14139 14572 15936 14600
rect 14139 14569 14151 14572
rect 14093 14563 14151 14569
rect 8536 14504 11008 14532
rect 8536 14492 8542 14504
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 13265 14535 13323 14541
rect 13265 14532 13277 14535
rect 11572 14504 13277 14532
rect 11572 14492 11578 14504
rect 13265 14501 13277 14504
rect 13311 14501 13323 14535
rect 13265 14495 13323 14501
rect 8754 14464 8760 14476
rect 8404 14436 8760 14464
rect 8754 14424 8760 14436
rect 8812 14464 8818 14476
rect 9214 14464 9220 14476
rect 8812 14436 9220 14464
rect 8812 14424 8818 14436
rect 9214 14424 9220 14436
rect 9272 14424 9278 14476
rect 9401 14467 9459 14473
rect 9401 14433 9413 14467
rect 9447 14464 9459 14467
rect 9582 14464 9588 14476
rect 9447 14436 9588 14464
rect 9447 14433 9459 14436
rect 9401 14427 9459 14433
rect 9582 14424 9588 14436
rect 9640 14424 9646 14476
rect 10594 14464 10600 14476
rect 10555 14436 10600 14464
rect 10594 14424 10600 14436
rect 10652 14424 10658 14476
rect 11333 14467 11391 14473
rect 11333 14433 11345 14467
rect 11379 14433 11391 14467
rect 12434 14464 12440 14476
rect 12395 14436 12440 14464
rect 11333 14427 11391 14433
rect 3789 14399 3847 14405
rect 3789 14396 3801 14399
rect 3344 14368 3801 14396
rect 3789 14365 3801 14368
rect 3835 14396 3847 14399
rect 3878 14396 3884 14408
rect 3835 14368 3884 14396
rect 3835 14365 3847 14368
rect 3789 14359 3847 14365
rect 3878 14356 3884 14368
rect 3936 14356 3942 14408
rect 5077 14399 5135 14405
rect 5077 14365 5089 14399
rect 5123 14396 5135 14399
rect 5166 14396 5172 14408
rect 5123 14368 5172 14396
rect 5123 14365 5135 14368
rect 5077 14359 5135 14365
rect 5166 14356 5172 14368
rect 5224 14356 5230 14408
rect 5258 14356 5264 14408
rect 5316 14396 5322 14408
rect 5721 14399 5779 14405
rect 5721 14396 5733 14399
rect 5316 14368 5733 14396
rect 5316 14356 5322 14368
rect 5721 14365 5733 14368
rect 5767 14396 5779 14399
rect 6086 14396 6092 14408
rect 5767 14368 6092 14396
rect 5767 14365 5779 14368
rect 5721 14359 5779 14365
rect 6086 14356 6092 14368
rect 6144 14356 6150 14408
rect 6641 14399 6699 14405
rect 6641 14365 6653 14399
rect 6687 14396 6699 14399
rect 8110 14396 8116 14408
rect 6687 14368 8116 14396
rect 6687 14365 6699 14368
rect 6641 14359 6699 14365
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 8297 14399 8355 14405
rect 8297 14365 8309 14399
rect 8343 14396 8355 14399
rect 8386 14396 8392 14408
rect 8343 14368 8392 14396
rect 8343 14365 8355 14368
rect 8297 14359 8355 14365
rect 8386 14356 8392 14368
rect 8444 14356 8450 14408
rect 8481 14399 8539 14405
rect 8481 14365 8493 14399
rect 8527 14396 8539 14399
rect 9122 14396 9128 14408
rect 8527 14368 9128 14396
rect 8527 14365 8539 14368
rect 8481 14359 8539 14365
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9306 14356 9312 14408
rect 9364 14396 9370 14408
rect 10505 14399 10563 14405
rect 10505 14396 10517 14399
rect 9364 14368 10517 14396
rect 9364 14356 9370 14368
rect 10505 14365 10517 14368
rect 10551 14396 10563 14399
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10551 14368 10977 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11348 14396 11376 14427
rect 12434 14424 12440 14436
rect 12492 14424 12498 14476
rect 12618 14424 12624 14476
rect 12676 14464 12682 14476
rect 13280 14464 13308 14495
rect 13354 14492 13360 14544
rect 13412 14532 13418 14544
rect 13412 14504 13952 14532
rect 13412 14492 13418 14504
rect 13924 14464 13952 14504
rect 13998 14492 14004 14544
rect 14056 14532 14062 14544
rect 14108 14532 14136 14563
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 18230 14560 18236 14612
rect 18288 14600 18294 14612
rect 18877 14603 18935 14609
rect 18877 14600 18889 14603
rect 18288 14572 18889 14600
rect 18288 14560 18294 14572
rect 18877 14569 18889 14572
rect 18923 14569 18935 14603
rect 19978 14600 19984 14612
rect 19939 14572 19984 14600
rect 18877 14563 18935 14569
rect 14056 14504 14136 14532
rect 14056 14492 14062 14504
rect 14274 14464 14280 14476
rect 12676 14436 12721 14464
rect 13280 14436 13768 14464
rect 13924 14436 14280 14464
rect 12676 14424 12682 14436
rect 11204 14368 11376 14396
rect 11204 14356 11210 14368
rect 11422 14356 11428 14408
rect 11480 14396 11486 14408
rect 13446 14396 13452 14408
rect 11480 14368 13023 14396
rect 13407 14368 13452 14396
rect 11480 14356 11486 14368
rect 1688 14300 2176 14328
rect 2332 14300 4752 14328
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2038 14260 2044 14272
rect 1999 14232 2044 14260
rect 2038 14220 2044 14232
rect 2096 14220 2102 14272
rect 2148 14269 2176 14300
rect 2133 14263 2191 14269
rect 2133 14229 2145 14263
rect 2179 14229 2191 14263
rect 2406 14260 2412 14272
rect 2367 14232 2412 14260
rect 2133 14223 2191 14229
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 3142 14260 3148 14272
rect 3103 14232 3148 14260
rect 3142 14220 3148 14232
rect 3200 14220 3206 14272
rect 3237 14263 3295 14269
rect 3237 14229 3249 14263
rect 3283 14260 3295 14263
rect 3510 14260 3516 14272
rect 3283 14232 3516 14260
rect 3283 14229 3295 14232
rect 3237 14223 3295 14229
rect 3510 14220 3516 14232
rect 3568 14220 3574 14272
rect 4062 14260 4068 14272
rect 4023 14232 4068 14260
rect 4062 14220 4068 14232
rect 4120 14220 4126 14272
rect 4430 14260 4436 14272
rect 4391 14232 4436 14260
rect 4430 14220 4436 14232
rect 4488 14220 4494 14272
rect 4522 14220 4528 14272
rect 4580 14260 4586 14272
rect 4724 14260 4752 14300
rect 4890 14288 4896 14340
rect 4948 14328 4954 14340
rect 5905 14331 5963 14337
rect 4948 14300 5580 14328
rect 4948 14288 4954 14300
rect 5552 14272 5580 14300
rect 5905 14297 5917 14331
rect 5951 14328 5963 14331
rect 6730 14328 6736 14340
rect 5951 14300 6736 14328
rect 5951 14297 5963 14300
rect 5905 14291 5963 14297
rect 6730 14288 6736 14300
rect 6788 14288 6794 14340
rect 7834 14288 7840 14340
rect 7892 14328 7898 14340
rect 8573 14331 8631 14337
rect 8573 14328 8585 14331
rect 7892 14300 8585 14328
rect 7892 14288 7898 14300
rect 8573 14297 8585 14300
rect 8619 14297 8631 14331
rect 8573 14291 8631 14297
rect 9398 14288 9404 14340
rect 9456 14328 9462 14340
rect 9585 14331 9643 14337
rect 9585 14328 9597 14331
rect 9456 14300 9597 14328
rect 9456 14288 9462 14300
rect 9585 14297 9597 14300
rect 9631 14297 9643 14331
rect 12894 14328 12900 14340
rect 9585 14291 9643 14297
rect 10888 14300 12900 14328
rect 10888 14272 10916 14300
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 12995 14328 13023 14368
rect 13446 14356 13452 14368
rect 13504 14356 13510 14408
rect 13740 14405 13768 14436
rect 14274 14424 14280 14436
rect 14332 14424 14338 14476
rect 17494 14464 17500 14476
rect 17455 14436 17500 14464
rect 17494 14424 17500 14436
rect 17552 14424 17558 14476
rect 18892 14464 18920 14563
rect 19978 14560 19984 14572
rect 20036 14560 20042 14612
rect 20901 14603 20959 14609
rect 20901 14569 20913 14603
rect 20947 14600 20959 14603
rect 21082 14600 21088 14612
rect 20947 14572 21088 14600
rect 20947 14569 20959 14572
rect 20901 14563 20959 14569
rect 21082 14560 21088 14572
rect 21140 14560 21146 14612
rect 18966 14492 18972 14544
rect 19024 14532 19030 14544
rect 19150 14532 19156 14544
rect 19024 14504 19156 14532
rect 19024 14492 19030 14504
rect 19150 14492 19156 14504
rect 19208 14532 19214 14544
rect 19208 14504 20668 14532
rect 19208 14492 19214 14504
rect 19337 14467 19395 14473
rect 19337 14464 19349 14467
rect 18892 14436 19349 14464
rect 19337 14433 19349 14436
rect 19383 14433 19395 14467
rect 19337 14427 19395 14433
rect 19702 14424 19708 14476
rect 19760 14464 19766 14476
rect 20530 14464 20536 14476
rect 19760 14436 20536 14464
rect 19760 14424 19766 14436
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 20640 14473 20668 14504
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14433 20683 14467
rect 20625 14427 20683 14433
rect 20990 14424 20996 14476
rect 21048 14464 21054 14476
rect 21048 14436 21312 14464
rect 21048 14424 21054 14436
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14365 13783 14399
rect 15470 14396 15476 14408
rect 15431 14368 15476 14396
rect 13725 14359 13783 14365
rect 15470 14356 15476 14368
rect 15528 14356 15534 14408
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 16945 14399 17003 14405
rect 16945 14396 16957 14399
rect 16356 14368 16957 14396
rect 16356 14356 16362 14368
rect 16945 14365 16957 14368
rect 16991 14365 17003 14399
rect 16945 14359 17003 14365
rect 18782 14356 18788 14408
rect 18840 14396 18846 14408
rect 19426 14396 19432 14408
rect 18840 14368 19432 14396
rect 18840 14356 18846 14368
rect 19426 14356 19432 14368
rect 19484 14356 19490 14408
rect 19794 14356 19800 14408
rect 19852 14396 19858 14408
rect 21284 14405 21312 14436
rect 20441 14399 20499 14405
rect 20441 14396 20453 14399
rect 19852 14368 20453 14396
rect 19852 14356 19858 14368
rect 20441 14365 20453 14368
rect 20487 14365 20499 14399
rect 20441 14359 20499 14365
rect 21085 14399 21143 14405
rect 21085 14365 21097 14399
rect 21131 14365 21143 14399
rect 21085 14359 21143 14365
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 15286 14337 15292 14340
rect 15228 14331 15292 14337
rect 15228 14328 15240 14331
rect 12995 14300 14964 14328
rect 15199 14300 15240 14328
rect 5258 14260 5264 14272
rect 4580 14232 4625 14260
rect 4724 14232 5264 14260
rect 4580 14220 4586 14232
rect 5258 14220 5264 14232
rect 5316 14220 5322 14272
rect 5534 14260 5540 14272
rect 5495 14232 5540 14260
rect 5534 14220 5540 14232
rect 5592 14220 5598 14272
rect 6273 14263 6331 14269
rect 6273 14229 6285 14263
rect 6319 14260 6331 14263
rect 6546 14260 6552 14272
rect 6319 14232 6552 14260
rect 6319 14229 6331 14232
rect 6273 14223 6331 14229
rect 6546 14220 6552 14232
rect 6604 14220 6610 14272
rect 7190 14260 7196 14272
rect 7151 14232 7196 14260
rect 7190 14220 7196 14232
rect 7248 14220 7254 14272
rect 7282 14220 7288 14272
rect 7340 14260 7346 14272
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 7340 14232 7573 14260
rect 7340 14220 7346 14232
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 7653 14263 7711 14269
rect 7653 14229 7665 14263
rect 7699 14260 7711 14263
rect 7926 14260 7932 14272
rect 7699 14232 7932 14260
rect 7699 14229 7711 14232
rect 7653 14223 7711 14229
rect 7926 14220 7932 14232
rect 7984 14260 7990 14272
rect 8021 14263 8079 14269
rect 8021 14260 8033 14263
rect 7984 14232 8033 14260
rect 7984 14220 7990 14232
rect 8021 14229 8033 14232
rect 8067 14229 8079 14263
rect 8021 14223 8079 14229
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14260 9183 14263
rect 9214 14260 9220 14272
rect 9171 14232 9220 14260
rect 9171 14229 9183 14232
rect 9125 14223 9183 14229
rect 9214 14220 9220 14232
rect 9272 14260 9278 14272
rect 9490 14260 9496 14272
rect 9272 14232 9496 14260
rect 9272 14220 9278 14232
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 10042 14220 10048 14272
rect 10100 14260 10106 14272
rect 10413 14263 10471 14269
rect 10100 14232 10145 14260
rect 10100 14220 10106 14232
rect 10413 14229 10425 14263
rect 10459 14260 10471 14263
rect 10870 14260 10876 14272
rect 10459 14232 10876 14260
rect 10459 14229 10471 14232
rect 10413 14223 10471 14229
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11425 14263 11483 14269
rect 11425 14260 11437 14263
rect 11296 14232 11437 14260
rect 11296 14220 11302 14232
rect 11425 14229 11437 14232
rect 11471 14229 11483 14263
rect 11425 14223 11483 14229
rect 11517 14263 11575 14269
rect 11517 14229 11529 14263
rect 11563 14260 11575 14263
rect 11698 14260 11704 14272
rect 11563 14232 11704 14260
rect 11563 14229 11575 14232
rect 11517 14223 11575 14229
rect 11698 14220 11704 14232
rect 11756 14220 11762 14272
rect 11882 14220 11888 14272
rect 11940 14260 11946 14272
rect 11977 14263 12035 14269
rect 11977 14260 11989 14263
rect 11940 14232 11989 14260
rect 11940 14220 11946 14232
rect 11977 14229 11989 14232
rect 12023 14260 12035 14263
rect 12713 14263 12771 14269
rect 12713 14260 12725 14263
rect 12023 14232 12725 14260
rect 12023 14229 12035 14232
rect 11977 14223 12035 14229
rect 12713 14229 12725 14232
rect 12759 14260 12771 14263
rect 13354 14260 13360 14272
rect 12759 14232 13360 14260
rect 12759 14229 12771 14232
rect 12713 14223 12771 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13538 14260 13544 14272
rect 13499 14232 13544 14260
rect 13538 14220 13544 14232
rect 13596 14220 13602 14272
rect 13909 14263 13967 14269
rect 13909 14229 13921 14263
rect 13955 14260 13967 14263
rect 14826 14260 14832 14272
rect 13955 14232 14832 14260
rect 13955 14229 13967 14232
rect 13909 14223 13967 14229
rect 14826 14220 14832 14232
rect 14884 14220 14890 14272
rect 14936 14260 14964 14300
rect 15228 14297 15240 14300
rect 15274 14297 15292 14331
rect 15228 14291 15292 14297
rect 15286 14288 15292 14291
rect 15344 14328 15350 14340
rect 16700 14331 16758 14337
rect 15344 14300 15608 14328
rect 15344 14288 15350 14300
rect 15378 14260 15384 14272
rect 14936 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 15580 14269 15608 14300
rect 16700 14297 16712 14331
rect 16746 14328 16758 14331
rect 17764 14331 17822 14337
rect 16746 14300 16988 14328
rect 16746 14297 16758 14300
rect 16700 14291 16758 14297
rect 16960 14272 16988 14300
rect 17764 14297 17776 14331
rect 17810 14328 17822 14331
rect 17862 14328 17868 14340
rect 17810 14300 17868 14328
rect 17810 14297 17822 14300
rect 17764 14291 17822 14297
rect 17862 14288 17868 14300
rect 17920 14288 17926 14340
rect 19334 14288 19340 14340
rect 19392 14328 19398 14340
rect 19613 14331 19671 14337
rect 19613 14328 19625 14331
rect 19392 14300 19625 14328
rect 19392 14288 19398 14300
rect 19613 14297 19625 14300
rect 19659 14297 19671 14331
rect 19613 14291 19671 14297
rect 20162 14288 20168 14340
rect 20220 14328 20226 14340
rect 21100 14328 21128 14359
rect 20220 14300 21128 14328
rect 20220 14288 20226 14300
rect 15565 14263 15623 14269
rect 15565 14229 15577 14263
rect 15611 14260 15623 14263
rect 16114 14260 16120 14272
rect 15611 14232 16120 14260
rect 15611 14229 15623 14232
rect 15565 14223 15623 14229
rect 16114 14220 16120 14232
rect 16172 14220 16178 14272
rect 16942 14220 16948 14272
rect 17000 14220 17006 14272
rect 17129 14263 17187 14269
rect 17129 14229 17141 14263
rect 17175 14260 17187 14263
rect 17218 14260 17224 14272
rect 17175 14232 17224 14260
rect 17175 14229 17187 14232
rect 17129 14223 17187 14229
rect 17218 14220 17224 14232
rect 17276 14220 17282 14272
rect 17402 14260 17408 14272
rect 17363 14232 17408 14260
rect 17402 14220 17408 14232
rect 17460 14220 17466 14272
rect 18598 14220 18604 14272
rect 18656 14260 18662 14272
rect 18969 14263 19027 14269
rect 18969 14260 18981 14263
rect 18656 14232 18981 14260
rect 18656 14220 18662 14232
rect 18969 14229 18981 14232
rect 19015 14229 19027 14263
rect 19518 14260 19524 14272
rect 19479 14232 19524 14260
rect 18969 14223 19027 14229
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 19702 14220 19708 14272
rect 19760 14260 19766 14272
rect 20073 14263 20131 14269
rect 20073 14260 20085 14263
rect 19760 14232 20085 14260
rect 19760 14220 19766 14232
rect 20073 14229 20085 14232
rect 20119 14229 20131 14263
rect 20530 14260 20536 14272
rect 20491 14232 20536 14260
rect 20073 14223 20131 14229
rect 20530 14220 20536 14232
rect 20588 14220 20594 14272
rect 21450 14260 21456 14272
rect 21411 14232 21456 14260
rect 21450 14220 21456 14232
rect 21508 14220 21514 14272
rect 21818 14220 21824 14272
rect 21876 14260 21882 14272
rect 22462 14260 22468 14272
rect 21876 14232 22468 14260
rect 21876 14220 21882 14232
rect 22462 14220 22468 14232
rect 22520 14220 22526 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 2317 14059 2375 14065
rect 2317 14025 2329 14059
rect 2363 14056 2375 14059
rect 2590 14056 2596 14068
rect 2363 14028 2596 14056
rect 2363 14025 2375 14028
rect 2317 14019 2375 14025
rect 2590 14016 2596 14028
rect 2648 14016 2654 14068
rect 5258 14056 5264 14068
rect 2884 14028 5264 14056
rect 2406 13988 2412 14000
rect 1688 13960 2412 13988
rect 1688 13929 1716 13960
rect 2406 13948 2412 13960
rect 2464 13948 2470 14000
rect 2884 13988 2912 14028
rect 5258 14016 5264 14028
rect 5316 14016 5322 14068
rect 5902 14056 5908 14068
rect 5863 14028 5908 14056
rect 5902 14016 5908 14028
rect 5960 14056 5966 14068
rect 7098 14056 7104 14068
rect 5960 14028 7104 14056
rect 5960 14016 5966 14028
rect 7098 14016 7104 14028
rect 7156 14016 7162 14068
rect 7193 14059 7251 14065
rect 7193 14025 7205 14059
rect 7239 14056 7251 14059
rect 7745 14059 7803 14065
rect 7745 14056 7757 14059
rect 7239 14028 7757 14056
rect 7239 14025 7251 14028
rect 7193 14019 7251 14025
rect 7745 14025 7757 14028
rect 7791 14025 7803 14059
rect 7745 14019 7803 14025
rect 8294 14016 8300 14068
rect 8352 14056 8358 14068
rect 8757 14059 8815 14065
rect 8757 14056 8769 14059
rect 8352 14028 8769 14056
rect 8352 14016 8358 14028
rect 8757 14025 8769 14028
rect 8803 14025 8815 14059
rect 8757 14019 8815 14025
rect 9125 14059 9183 14065
rect 9125 14025 9137 14059
rect 9171 14056 9183 14059
rect 10042 14056 10048 14068
rect 9171 14028 10048 14056
rect 9171 14025 9183 14028
rect 9125 14019 9183 14025
rect 10042 14016 10048 14028
rect 10100 14016 10106 14068
rect 10318 14056 10324 14068
rect 10279 14028 10324 14056
rect 10318 14016 10324 14028
rect 10376 14016 10382 14068
rect 10870 14056 10876 14068
rect 10831 14028 10876 14056
rect 10870 14016 10876 14028
rect 10928 14016 10934 14068
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 11112 14028 11253 14056
rect 11112 14016 11118 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 11241 14019 11299 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11698 14056 11704 14068
rect 11563 14028 11704 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 4614 13988 4620 14000
rect 2516 13960 2912 13988
rect 3068 13960 4620 13988
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 2038 13920 2044 13932
rect 1999 13892 2044 13920
rect 1673 13883 1731 13889
rect 2038 13880 2044 13892
rect 2096 13880 2102 13932
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2516 13920 2544 13960
rect 2179 13892 2544 13920
rect 2593 13923 2651 13929
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2682 13920 2688 13932
rect 2639 13892 2688 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2682 13880 2688 13892
rect 2740 13880 2746 13932
rect 2969 13927 3027 13933
rect 2969 13893 2981 13927
rect 3015 13920 3027 13927
rect 3068 13920 3096 13960
rect 4614 13948 4620 13960
rect 4672 13948 4678 14000
rect 5994 13948 6000 14000
rect 6052 13988 6058 14000
rect 6089 13991 6147 13997
rect 6089 13988 6101 13991
rect 6052 13960 6101 13988
rect 6052 13948 6058 13960
rect 6089 13957 6101 13960
rect 6135 13988 6147 13991
rect 6638 13988 6644 14000
rect 6135 13960 6644 13988
rect 6135 13957 6147 13960
rect 6089 13951 6147 13957
rect 6638 13948 6644 13960
rect 6696 13988 6702 14000
rect 6733 13991 6791 13997
rect 6733 13988 6745 13991
rect 6696 13960 6745 13988
rect 6696 13948 6702 13960
rect 6733 13957 6745 13960
rect 6779 13957 6791 13991
rect 6733 13951 6791 13957
rect 6822 13948 6828 14000
rect 6880 13988 6886 14000
rect 8478 13988 8484 14000
rect 6880 13960 6925 13988
rect 8439 13960 8484 13988
rect 6880 13948 6886 13960
rect 8478 13948 8484 13960
rect 8536 13948 8542 14000
rect 8570 13948 8576 14000
rect 8628 13988 8634 14000
rect 9217 13991 9275 13997
rect 9217 13988 9229 13991
rect 8628 13960 9229 13988
rect 8628 13948 8634 13960
rect 9217 13957 9229 13960
rect 9263 13957 9275 13991
rect 9217 13951 9275 13957
rect 9953 13991 10011 13997
rect 9953 13957 9965 13991
rect 9999 13988 10011 13991
rect 10778 13988 10784 14000
rect 9999 13960 10784 13988
rect 9999 13957 10011 13960
rect 9953 13951 10011 13957
rect 10778 13948 10784 13960
rect 10836 13948 10842 14000
rect 3326 13929 3332 13932
rect 3320 13920 3332 13929
rect 3015 13893 3096 13920
rect 2969 13892 3096 13893
rect 3239 13892 3332 13920
rect 2969 13887 3027 13892
rect 2222 13812 2228 13864
rect 2280 13852 2286 13864
rect 3068 13861 3096 13892
rect 3320 13883 3332 13892
rect 3384 13920 3390 13932
rect 4781 13923 4839 13929
rect 4781 13920 4793 13923
rect 3384 13892 4108 13920
rect 3326 13880 3332 13883
rect 3384 13880 3390 13892
rect 4080 13864 4108 13892
rect 4448 13892 4793 13920
rect 3053 13855 3111 13861
rect 2280 13824 2452 13852
rect 2280 13812 2286 13824
rect 1854 13784 1860 13796
rect 1815 13756 1860 13784
rect 1854 13744 1860 13756
rect 1912 13744 1918 13796
rect 2424 13793 2452 13824
rect 3053 13821 3065 13855
rect 3099 13821 3111 13855
rect 3053 13815 3111 13821
rect 4062 13812 4068 13864
rect 4120 13812 4126 13864
rect 2409 13787 2467 13793
rect 2409 13753 2421 13787
rect 2455 13753 2467 13787
rect 2409 13747 2467 13753
rect 1486 13716 1492 13728
rect 1447 13688 1492 13716
rect 1486 13676 1492 13688
rect 1544 13676 1550 13728
rect 2682 13676 2688 13728
rect 2740 13716 2746 13728
rect 2777 13719 2835 13725
rect 2777 13716 2789 13719
rect 2740 13688 2789 13716
rect 2740 13676 2746 13688
rect 2777 13685 2789 13688
rect 2823 13685 2835 13719
rect 2777 13679 2835 13685
rect 4338 13676 4344 13728
rect 4396 13716 4402 13728
rect 4448 13725 4476 13892
rect 4781 13889 4793 13892
rect 4827 13889 4839 13923
rect 4781 13883 4839 13889
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 7653 13923 7711 13929
rect 7653 13920 7665 13923
rect 7064 13892 7665 13920
rect 7064 13880 7070 13892
rect 7653 13889 7665 13892
rect 7699 13889 7711 13923
rect 9306 13920 9312 13932
rect 7653 13883 7711 13889
rect 7760 13892 9312 13920
rect 4525 13855 4583 13861
rect 4525 13821 4537 13855
rect 4571 13821 4583 13855
rect 4525 13815 4583 13821
rect 4433 13719 4491 13725
rect 4433 13716 4445 13719
rect 4396 13688 4445 13716
rect 4396 13676 4402 13688
rect 4433 13685 4445 13688
rect 4479 13685 4491 13719
rect 4540 13716 4568 13815
rect 5902 13812 5908 13864
rect 5960 13852 5966 13864
rect 6454 13852 6460 13864
rect 5960 13824 6460 13852
rect 5960 13812 5966 13824
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13821 6607 13855
rect 7760 13852 7788 13892
rect 9306 13880 9312 13892
rect 9364 13880 9370 13932
rect 9490 13880 9496 13932
rect 9548 13920 9554 13932
rect 9861 13923 9919 13929
rect 9861 13920 9873 13923
rect 9548 13892 9873 13920
rect 9548 13880 9554 13892
rect 9861 13889 9873 13892
rect 9907 13889 9919 13923
rect 9861 13883 9919 13889
rect 6549 13815 6607 13821
rect 6757 13824 7788 13852
rect 7837 13855 7895 13861
rect 6362 13744 6368 13796
rect 6420 13784 6426 13796
rect 6564 13784 6592 13815
rect 6420 13756 6592 13784
rect 6420 13744 6426 13756
rect 4706 13716 4712 13728
rect 4540 13688 4712 13716
rect 4433 13679 4491 13685
rect 4706 13676 4712 13688
rect 4764 13676 4770 13728
rect 6546 13676 6552 13728
rect 6604 13716 6610 13728
rect 6757 13716 6785 13824
rect 7837 13821 7849 13855
rect 7883 13821 7895 13855
rect 7837 13815 7895 13821
rect 6822 13744 6828 13796
rect 6880 13784 6886 13796
rect 7852 13784 7880 13815
rect 8570 13812 8576 13864
rect 8628 13852 8634 13864
rect 8754 13852 8760 13864
rect 8628 13824 8760 13852
rect 8628 13812 8634 13824
rect 8754 13812 8760 13824
rect 8812 13812 8818 13864
rect 9401 13855 9459 13861
rect 9401 13821 9413 13855
rect 9447 13852 9459 13855
rect 9582 13852 9588 13864
rect 9447 13824 9588 13852
rect 9447 13821 9459 13824
rect 9401 13815 9459 13821
rect 9582 13812 9588 13824
rect 9640 13852 9646 13864
rect 9677 13855 9735 13861
rect 9677 13852 9689 13855
rect 9640 13824 9689 13852
rect 9640 13812 9646 13824
rect 9677 13821 9689 13824
rect 9723 13821 9735 13855
rect 10410 13852 10416 13864
rect 10371 13824 10416 13852
rect 9677 13815 9735 13821
rect 10410 13812 10416 13824
rect 10468 13812 10474 13864
rect 10686 13852 10692 13864
rect 10647 13824 10692 13852
rect 10686 13812 10692 13824
rect 10744 13812 10750 13864
rect 11146 13852 11152 13864
rect 11107 13824 11152 13852
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 11256 13852 11284 14019
rect 11698 14016 11704 14028
rect 11756 14016 11762 14068
rect 11790 14016 11796 14068
rect 11848 14056 11854 14068
rect 11974 14056 11980 14068
rect 11848 14028 11980 14056
rect 11848 14016 11854 14028
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12986 14016 12992 14068
rect 13044 14056 13050 14068
rect 13541 14059 13599 14065
rect 13541 14056 13553 14059
rect 13044 14028 13553 14056
rect 13044 14016 13050 14028
rect 13541 14025 13553 14028
rect 13587 14025 13599 14059
rect 15194 14056 15200 14068
rect 15155 14028 15200 14056
rect 13541 14019 13599 14025
rect 15194 14016 15200 14028
rect 15252 14016 15258 14068
rect 15470 14016 15476 14068
rect 15528 14056 15534 14068
rect 16025 14059 16083 14065
rect 16025 14056 16037 14059
rect 15528 14028 16037 14056
rect 15528 14016 15534 14028
rect 16025 14025 16037 14028
rect 16071 14025 16083 14059
rect 16025 14019 16083 14025
rect 17126 14016 17132 14068
rect 17184 14056 17190 14068
rect 17497 14059 17555 14065
rect 17497 14056 17509 14059
rect 17184 14028 17509 14056
rect 17184 14016 17190 14028
rect 17497 14025 17509 14028
rect 17543 14025 17555 14059
rect 17497 14019 17555 14025
rect 17957 14059 18015 14065
rect 17957 14025 17969 14059
rect 18003 14056 18015 14059
rect 18509 14059 18567 14065
rect 18509 14056 18521 14059
rect 18003 14028 18521 14056
rect 18003 14025 18015 14028
rect 17957 14019 18015 14025
rect 18509 14025 18521 14028
rect 18555 14025 18567 14059
rect 19334 14056 19340 14068
rect 19295 14028 19340 14056
rect 18509 14019 18567 14025
rect 19334 14016 19340 14028
rect 19392 14016 19398 14068
rect 19702 14056 19708 14068
rect 19663 14028 19708 14056
rect 19702 14016 19708 14028
rect 19760 14016 19766 14068
rect 20809 14059 20867 14065
rect 20809 14025 20821 14059
rect 20855 14025 20867 14059
rect 21082 14056 21088 14068
rect 21043 14028 21088 14056
rect 20809 14019 20867 14025
rect 12066 13948 12072 14000
rect 12124 13988 12130 14000
rect 12526 13988 12532 14000
rect 12124 13960 12532 13988
rect 12124 13948 12130 13960
rect 12526 13948 12532 13960
rect 12584 13988 12590 14000
rect 13357 13991 13415 13997
rect 13357 13988 13369 13991
rect 12584 13960 13369 13988
rect 12584 13948 12590 13960
rect 13357 13957 13369 13960
rect 13403 13957 13415 13991
rect 13357 13951 13415 13957
rect 13446 13948 13452 14000
rect 13504 13988 13510 14000
rect 15488 13988 15516 14016
rect 13504 13960 15516 13988
rect 13504 13948 13510 13960
rect 11330 13880 11336 13932
rect 11388 13920 11394 13932
rect 11790 13920 11796 13932
rect 11388 13892 11796 13920
rect 11388 13880 11394 13892
rect 11790 13880 11796 13892
rect 11848 13880 11854 13932
rect 13740 13929 13768 13960
rect 15654 13948 15660 14000
rect 15712 13988 15718 14000
rect 16393 13991 16451 13997
rect 16393 13988 16405 13991
rect 15712 13960 16405 13988
rect 15712 13948 15718 13960
rect 16393 13957 16405 13960
rect 16439 13988 16451 13991
rect 18414 13988 18420 14000
rect 16439 13960 18420 13988
rect 16439 13957 16451 13960
rect 16393 13951 16451 13957
rect 18414 13948 18420 13960
rect 18472 13948 18478 14000
rect 19518 13988 19524 14000
rect 18708 13960 19524 13988
rect 13998 13929 14004 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 11931 13892 12357 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 13725 13923 13783 13929
rect 13725 13889 13737 13923
rect 13771 13889 13783 13923
rect 13992 13920 14004 13929
rect 13959 13892 14004 13920
rect 13725 13883 13783 13889
rect 13992 13883 14004 13892
rect 13998 13880 14004 13883
rect 14056 13880 14062 13932
rect 15102 13880 15108 13932
rect 15160 13920 15166 13932
rect 15565 13923 15623 13929
rect 15565 13920 15577 13923
rect 15160 13892 15577 13920
rect 15160 13880 15166 13892
rect 15565 13889 15577 13892
rect 15611 13889 15623 13923
rect 15565 13883 15623 13889
rect 16209 13923 16267 13929
rect 16209 13889 16221 13923
rect 16255 13920 16267 13923
rect 16298 13920 16304 13932
rect 16255 13892 16304 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 17218 13920 17224 13932
rect 17179 13892 17224 13920
rect 17218 13880 17224 13892
rect 17276 13880 17282 13932
rect 18046 13920 18052 13932
rect 18007 13892 18052 13920
rect 18046 13880 18052 13892
rect 18104 13880 18110 13932
rect 11606 13852 11612 13864
rect 11256 13824 11612 13852
rect 11606 13812 11612 13824
rect 11664 13852 11670 13864
rect 11977 13855 12035 13861
rect 11977 13852 11989 13855
rect 11664 13824 11989 13852
rect 11664 13812 11670 13824
rect 11977 13821 11989 13824
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 12069 13855 12127 13861
rect 12069 13821 12081 13855
rect 12115 13821 12127 13855
rect 12986 13852 12992 13864
rect 12947 13824 12992 13852
rect 12069 13815 12127 13821
rect 6880 13756 7880 13784
rect 6880 13744 6886 13756
rect 7926 13744 7932 13796
rect 7984 13784 7990 13796
rect 8113 13787 8171 13793
rect 8113 13784 8125 13787
rect 7984 13756 8125 13784
rect 7984 13744 7990 13756
rect 8113 13753 8125 13756
rect 8159 13753 8171 13787
rect 8294 13784 8300 13796
rect 8255 13756 8300 13784
rect 8113 13747 8171 13753
rect 8294 13744 8300 13756
rect 8352 13744 8358 13796
rect 10134 13744 10140 13796
rect 10192 13784 10198 13796
rect 10192 13756 11652 13784
rect 10192 13744 10198 13756
rect 6604 13688 6785 13716
rect 6604 13676 6610 13688
rect 6914 13676 6920 13728
rect 6972 13716 6978 13728
rect 7285 13719 7343 13725
rect 7285 13716 7297 13719
rect 6972 13688 7297 13716
rect 6972 13676 6978 13688
rect 7285 13685 7297 13688
rect 7331 13685 7343 13719
rect 7285 13679 7343 13685
rect 7650 13676 7656 13728
rect 7708 13716 7714 13728
rect 8478 13716 8484 13728
rect 7708 13688 8484 13716
rect 7708 13676 7714 13688
rect 8478 13676 8484 13688
rect 8536 13716 8542 13728
rect 11514 13716 11520 13728
rect 8536 13688 11520 13716
rect 8536 13676 8542 13688
rect 11514 13676 11520 13688
rect 11572 13676 11578 13728
rect 11624 13716 11652 13756
rect 11790 13744 11796 13796
rect 11848 13784 11854 13796
rect 12084 13784 12112 13815
rect 12986 13812 12992 13824
rect 13044 13812 13050 13864
rect 13170 13852 13176 13864
rect 13131 13824 13176 13852
rect 13170 13812 13176 13824
rect 13228 13812 13234 13864
rect 14734 13812 14740 13864
rect 14792 13852 14798 13864
rect 15654 13852 15660 13864
rect 14792 13824 15148 13852
rect 15615 13824 15660 13852
rect 14792 13812 14798 13824
rect 15120 13793 15148 13824
rect 15654 13812 15660 13824
rect 15712 13812 15718 13864
rect 15841 13855 15899 13861
rect 15841 13821 15853 13855
rect 15887 13852 15899 13855
rect 15930 13852 15936 13864
rect 15887 13824 15936 13852
rect 15887 13821 15899 13824
rect 15841 13815 15899 13821
rect 15930 13812 15936 13824
rect 15988 13812 15994 13864
rect 16574 13812 16580 13864
rect 16632 13852 16638 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16632 13824 16681 13852
rect 16632 13812 16638 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 17126 13852 17132 13864
rect 17087 13824 17132 13852
rect 16669 13815 16727 13821
rect 17126 13812 17132 13824
rect 17184 13812 17190 13864
rect 17586 13852 17592 13864
rect 17236 13824 17592 13852
rect 17236 13796 17264 13824
rect 17586 13812 17592 13824
rect 17644 13812 17650 13864
rect 17862 13852 17868 13864
rect 17775 13824 17868 13852
rect 17862 13812 17868 13824
rect 17920 13852 17926 13864
rect 18708 13852 18736 13960
rect 19518 13948 19524 13960
rect 19576 13948 19582 14000
rect 19610 13948 19616 14000
rect 19668 13988 19674 14000
rect 19797 13991 19855 13997
rect 19797 13988 19809 13991
rect 19668 13960 19809 13988
rect 19668 13948 19674 13960
rect 19797 13957 19809 13960
rect 19843 13957 19855 13991
rect 20824 13988 20852 14019
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21174 13988 21180 14000
rect 20824 13960 21180 13988
rect 19797 13951 19855 13957
rect 21174 13948 21180 13960
rect 21232 13948 21238 14000
rect 18874 13920 18880 13932
rect 18835 13892 18880 13920
rect 18874 13880 18880 13892
rect 18932 13880 18938 13932
rect 20438 13920 20444 13932
rect 20399 13892 20444 13920
rect 20438 13880 20444 13892
rect 20496 13920 20502 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20496 13892 20637 13920
rect 20496 13880 20502 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20772 13892 20913 13920
rect 20772 13880 20778 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 21266 13920 21272 13932
rect 21227 13892 21272 13920
rect 20901 13883 20959 13889
rect 21266 13880 21272 13892
rect 21324 13880 21330 13932
rect 18966 13852 18972 13864
rect 17920 13824 18368 13852
rect 17920 13812 17926 13824
rect 15105 13787 15163 13793
rect 11848 13756 12112 13784
rect 12176 13756 12940 13784
rect 11848 13744 11854 13756
rect 12176 13716 12204 13756
rect 12618 13716 12624 13728
rect 11624 13688 12204 13716
rect 12579 13688 12624 13716
rect 12618 13676 12624 13688
rect 12676 13676 12682 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 12805 13719 12863 13725
rect 12805 13716 12817 13719
rect 12768 13688 12817 13716
rect 12768 13676 12774 13688
rect 12805 13685 12817 13688
rect 12851 13685 12863 13719
rect 12912 13716 12940 13756
rect 15105 13753 15117 13787
rect 15151 13753 15163 13787
rect 15105 13747 15163 13753
rect 17218 13744 17224 13796
rect 17276 13744 17282 13796
rect 14826 13716 14832 13728
rect 12912 13688 14832 13716
rect 12805 13679 12863 13685
rect 14826 13676 14832 13688
rect 14884 13676 14890 13728
rect 16206 13676 16212 13728
rect 16264 13716 16270 13728
rect 16666 13716 16672 13728
rect 16264 13688 16672 13716
rect 16264 13676 16270 13688
rect 16666 13676 16672 13688
rect 16724 13716 16730 13728
rect 16853 13719 16911 13725
rect 16853 13716 16865 13719
rect 16724 13688 16865 13716
rect 16724 13676 16730 13688
rect 16853 13685 16865 13688
rect 16899 13685 16911 13719
rect 18340 13716 18368 13824
rect 18432 13824 18736 13852
rect 18927 13824 18972 13852
rect 18432 13793 18460 13824
rect 18966 13812 18972 13824
rect 19024 13812 19030 13864
rect 19150 13852 19156 13864
rect 19111 13824 19156 13852
rect 19150 13812 19156 13824
rect 19208 13812 19214 13864
rect 19886 13812 19892 13864
rect 19944 13852 19950 13864
rect 19944 13824 19989 13852
rect 19944 13812 19950 13824
rect 20070 13812 20076 13864
rect 20128 13852 20134 13864
rect 20165 13855 20223 13861
rect 20165 13852 20177 13855
rect 20128 13824 20177 13852
rect 20128 13812 20134 13824
rect 20165 13821 20177 13824
rect 20211 13852 20223 13855
rect 20530 13852 20536 13864
rect 20211 13824 20536 13852
rect 20211 13821 20223 13824
rect 20165 13815 20223 13821
rect 20530 13812 20536 13824
rect 20588 13812 20594 13864
rect 18417 13787 18475 13793
rect 18417 13753 18429 13787
rect 18463 13753 18475 13787
rect 18417 13747 18475 13753
rect 19904 13716 19932 13812
rect 21450 13716 21456 13728
rect 18340 13688 19932 13716
rect 21411 13688 21456 13716
rect 16853 13679 16911 13685
rect 21450 13676 21456 13688
rect 21508 13676 21514 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 3326 13512 3332 13524
rect 2271 13484 3332 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 3326 13472 3332 13484
rect 3384 13472 3390 13524
rect 3418 13472 3424 13524
rect 3476 13512 3482 13524
rect 3878 13512 3884 13524
rect 3476 13484 3740 13512
rect 3839 13484 3884 13512
rect 3476 13472 3482 13484
rect 3712 13444 3740 13484
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4522 13472 4528 13524
rect 4580 13512 4586 13524
rect 4617 13515 4675 13521
rect 4617 13512 4629 13515
rect 4580 13484 4629 13512
rect 4580 13472 4586 13484
rect 4617 13481 4629 13484
rect 4663 13481 4675 13515
rect 4617 13475 4675 13481
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 6730 13512 6736 13524
rect 5040 13484 6736 13512
rect 5040 13472 5046 13484
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 7006 13512 7012 13524
rect 6967 13484 7012 13512
rect 7006 13472 7012 13484
rect 7064 13472 7070 13524
rect 7742 13512 7748 13524
rect 7116 13484 7748 13512
rect 6914 13444 6920 13456
rect 3712 13416 6040 13444
rect 4062 13376 4068 13388
rect 3528 13348 4068 13376
rect 1670 13308 1676 13320
rect 1631 13280 1676 13308
rect 1670 13268 1676 13280
rect 1728 13268 1734 13320
rect 2041 13311 2099 13317
rect 2041 13277 2053 13311
rect 2087 13308 2099 13311
rect 3528 13308 3556 13348
rect 4062 13336 4068 13348
rect 4120 13336 4126 13388
rect 4338 13336 4344 13388
rect 4396 13376 4402 13388
rect 5169 13379 5227 13385
rect 5169 13376 5181 13379
rect 4396 13348 5181 13376
rect 4396 13336 4402 13348
rect 5169 13345 5181 13348
rect 5215 13345 5227 13379
rect 5169 13339 5227 13345
rect 5718 13336 5724 13388
rect 5776 13376 5782 13388
rect 6012 13385 6040 13416
rect 6472 13416 6920 13444
rect 5905 13379 5963 13385
rect 5905 13376 5917 13379
rect 5776 13348 5917 13376
rect 5776 13336 5782 13348
rect 5905 13345 5917 13348
rect 5951 13345 5963 13379
rect 5905 13339 5963 13345
rect 5997 13379 6055 13385
rect 5997 13345 6009 13379
rect 6043 13376 6055 13379
rect 6362 13376 6368 13388
rect 6043 13348 6368 13376
rect 6043 13345 6055 13348
rect 5997 13339 6055 13345
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 2087 13280 3556 13308
rect 3605 13311 3663 13317
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 3605 13277 3617 13311
rect 3651 13308 3663 13311
rect 4706 13308 4712 13320
rect 3651 13280 4712 13308
rect 3651 13277 3663 13280
rect 3605 13271 3663 13277
rect 4706 13268 4712 13280
rect 4764 13268 4770 13320
rect 5077 13311 5135 13317
rect 5077 13277 5089 13311
rect 5123 13308 5135 13311
rect 6472 13308 6500 13416
rect 6914 13404 6920 13416
rect 6972 13404 6978 13456
rect 7116 13388 7144 13484
rect 7742 13472 7748 13484
rect 7800 13472 7806 13524
rect 8018 13472 8024 13524
rect 8076 13512 8082 13524
rect 9033 13515 9091 13521
rect 9033 13512 9045 13515
rect 8076 13484 9045 13512
rect 8076 13472 8082 13484
rect 9033 13481 9045 13484
rect 9079 13481 9091 13515
rect 11330 13512 11336 13524
rect 9033 13475 9091 13481
rect 9600 13484 11336 13512
rect 8481 13447 8539 13453
rect 8481 13413 8493 13447
rect 8527 13444 8539 13447
rect 9122 13444 9128 13456
rect 8527 13416 9128 13444
rect 8527 13413 8539 13416
rect 8481 13407 8539 13413
rect 9122 13404 9128 13416
rect 9180 13404 9186 13456
rect 7098 13376 7104 13388
rect 7011 13348 7104 13376
rect 7098 13336 7104 13348
rect 7156 13336 7162 13388
rect 5123 13280 6500 13308
rect 5123 13277 5135 13280
rect 5077 13271 5135 13277
rect 6546 13268 6552 13320
rect 6604 13308 6610 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 6604 13280 6653 13308
rect 6604 13268 6610 13280
rect 6641 13277 6653 13280
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 7190 13268 7196 13320
rect 7248 13308 7254 13320
rect 7357 13311 7415 13317
rect 7357 13308 7369 13311
rect 7248 13280 7369 13308
rect 7248 13268 7254 13280
rect 7357 13277 7369 13280
rect 7403 13277 7415 13311
rect 9600 13308 9628 13484
rect 11330 13472 11336 13484
rect 11388 13472 11394 13524
rect 11514 13472 11520 13524
rect 11572 13512 11578 13524
rect 15102 13512 15108 13524
rect 11572 13484 14780 13512
rect 15063 13484 15108 13512
rect 11572 13472 11578 13484
rect 13078 13404 13084 13456
rect 13136 13444 13142 13456
rect 13354 13444 13360 13456
rect 13136 13416 13360 13444
rect 13136 13404 13142 13416
rect 13354 13404 13360 13416
rect 13412 13404 13418 13456
rect 13541 13447 13599 13453
rect 13541 13413 13553 13447
rect 13587 13444 13599 13447
rect 13814 13444 13820 13456
rect 13587 13416 13820 13444
rect 13587 13413 13599 13416
rect 13541 13407 13599 13413
rect 13814 13404 13820 13416
rect 13872 13444 13878 13456
rect 14366 13444 14372 13456
rect 13872 13416 14372 13444
rect 13872 13404 13878 13416
rect 14366 13404 14372 13416
rect 14424 13404 14430 13456
rect 14752 13444 14780 13484
rect 15102 13472 15108 13484
rect 15160 13472 15166 13524
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15804 13484 16037 13512
rect 15804 13472 15810 13484
rect 16025 13481 16037 13484
rect 16071 13481 16083 13515
rect 18046 13512 18052 13524
rect 18007 13484 18052 13512
rect 16025 13475 16083 13481
rect 18046 13472 18052 13484
rect 18104 13472 18110 13524
rect 18414 13472 18420 13524
rect 18472 13512 18478 13524
rect 19429 13515 19487 13521
rect 19429 13512 19441 13515
rect 18472 13484 19441 13512
rect 18472 13472 18478 13484
rect 19429 13481 19441 13484
rect 19475 13481 19487 13515
rect 20714 13512 20720 13524
rect 20675 13484 20720 13512
rect 19429 13475 19487 13481
rect 20714 13472 20720 13484
rect 20772 13472 20778 13524
rect 20993 13515 21051 13521
rect 20993 13481 21005 13515
rect 21039 13512 21051 13515
rect 21266 13512 21272 13524
rect 21039 13484 21272 13512
rect 21039 13481 21051 13484
rect 20993 13475 21051 13481
rect 21266 13472 21272 13484
rect 21324 13472 21330 13524
rect 17037 13447 17095 13453
rect 17037 13444 17049 13447
rect 14752 13416 17049 13444
rect 17037 13413 17049 13416
rect 17083 13413 17095 13447
rect 17037 13407 17095 13413
rect 17957 13447 18015 13453
rect 17957 13413 17969 13447
rect 18003 13444 18015 13447
rect 18966 13444 18972 13456
rect 18003 13416 18972 13444
rect 18003 13413 18015 13416
rect 17957 13407 18015 13413
rect 9674 13336 9680 13388
rect 9732 13376 9738 13388
rect 11606 13376 11612 13388
rect 9732 13348 9777 13376
rect 11567 13348 11612 13376
rect 9732 13336 9738 13348
rect 11606 13336 11612 13348
rect 11664 13336 11670 13388
rect 14553 13379 14611 13385
rect 14553 13345 14565 13379
rect 14599 13376 14611 13379
rect 15286 13376 15292 13388
rect 14599 13348 15292 13376
rect 14599 13345 14611 13348
rect 14553 13339 14611 13345
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15841 13379 15899 13385
rect 15841 13345 15853 13379
rect 15887 13345 15899 13379
rect 15841 13339 15899 13345
rect 9950 13308 9956 13320
rect 7357 13271 7415 13277
rect 7484 13280 9628 13308
rect 9784 13280 9956 13308
rect 2314 13200 2320 13252
rect 2372 13240 2378 13252
rect 3326 13240 3332 13252
rect 3384 13249 3390 13252
rect 2372 13212 2774 13240
rect 3296 13212 3332 13240
rect 2372 13200 2378 13212
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1854 13172 1860 13184
rect 1815 13144 1860 13172
rect 1854 13132 1860 13144
rect 1912 13132 1918 13184
rect 2746 13172 2774 13212
rect 3326 13200 3332 13212
rect 3384 13203 3396 13249
rect 3973 13243 4031 13249
rect 3973 13240 3985 13243
rect 3436 13212 3985 13240
rect 3384 13200 3390 13203
rect 3142 13172 3148 13184
rect 2746 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13172 3206 13184
rect 3436 13172 3464 13212
rect 3973 13209 3985 13212
rect 4019 13209 4031 13243
rect 7484 13240 7512 13280
rect 3973 13203 4031 13209
rect 4080 13212 7512 13240
rect 3200 13144 3464 13172
rect 3200 13132 3206 13144
rect 3510 13132 3516 13184
rect 3568 13172 3574 13184
rect 4080 13172 4108 13212
rect 8202 13200 8208 13252
rect 8260 13240 8266 13252
rect 9125 13243 9183 13249
rect 9125 13240 9137 13243
rect 8260 13212 9137 13240
rect 8260 13200 8266 13212
rect 9125 13209 9137 13212
rect 9171 13209 9183 13243
rect 9490 13240 9496 13252
rect 9451 13212 9496 13240
rect 9125 13203 9183 13209
rect 9490 13200 9496 13212
rect 9548 13200 9554 13252
rect 4246 13172 4252 13184
rect 3568 13144 4108 13172
rect 4207 13144 4252 13172
rect 3568 13132 3574 13144
rect 4246 13132 4252 13144
rect 4304 13132 4310 13184
rect 4982 13172 4988 13184
rect 4943 13144 4988 13172
rect 4982 13132 4988 13144
rect 5040 13132 5046 13184
rect 5442 13172 5448 13184
rect 5403 13144 5448 13172
rect 5442 13132 5448 13144
rect 5500 13132 5506 13184
rect 5813 13175 5871 13181
rect 5813 13141 5825 13175
rect 5859 13172 5871 13175
rect 5994 13172 6000 13184
rect 5859 13144 6000 13172
rect 5859 13141 5871 13144
rect 5813 13135 5871 13141
rect 5994 13132 6000 13144
rect 6052 13132 6058 13184
rect 6549 13175 6607 13181
rect 6549 13141 6561 13175
rect 6595 13172 6607 13175
rect 7558 13172 7564 13184
rect 6595 13144 7564 13172
rect 6595 13141 6607 13144
rect 6549 13135 6607 13141
rect 7558 13132 7564 13144
rect 7616 13172 7622 13184
rect 7926 13172 7932 13184
rect 7616 13144 7932 13172
rect 7616 13132 7622 13144
rect 7926 13132 7932 13144
rect 7984 13132 7990 13184
rect 8662 13172 8668 13184
rect 8623 13144 8668 13172
rect 8662 13132 8668 13144
rect 8720 13132 8726 13184
rect 8754 13132 8760 13184
rect 8812 13172 8818 13184
rect 9784 13181 9812 13280
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10137 13311 10195 13317
rect 10137 13277 10149 13311
rect 10183 13308 10195 13311
rect 11624 13308 11652 13336
rect 11865 13311 11923 13317
rect 11865 13308 11877 13311
rect 10183 13280 11652 13308
rect 11716 13280 11877 13308
rect 10183 13277 10195 13280
rect 10137 13271 10195 13277
rect 10336 13184 10364 13280
rect 10404 13243 10462 13249
rect 10404 13209 10416 13243
rect 10450 13240 10462 13243
rect 10870 13240 10876 13252
rect 10450 13212 10876 13240
rect 10450 13209 10462 13212
rect 10404 13203 10462 13209
rect 10870 13200 10876 13212
rect 10928 13200 10934 13252
rect 9769 13175 9827 13181
rect 9769 13172 9781 13175
rect 8812 13144 9781 13172
rect 8812 13132 8818 13144
rect 9769 13141 9781 13144
rect 9815 13141 9827 13175
rect 9950 13172 9956 13184
rect 9911 13144 9956 13172
rect 9769 13135 9827 13141
rect 9950 13132 9956 13144
rect 10008 13132 10014 13184
rect 10318 13132 10324 13184
rect 10376 13132 10382 13184
rect 11054 13132 11060 13184
rect 11112 13172 11118 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11112 13144 11529 13172
rect 11112 13132 11118 13144
rect 11517 13141 11529 13144
rect 11563 13172 11575 13175
rect 11716 13172 11744 13280
rect 11865 13277 11877 13280
rect 11911 13277 11923 13311
rect 13725 13311 13783 13317
rect 13725 13308 13737 13311
rect 11865 13271 11923 13277
rect 11992 13280 13737 13308
rect 11992 13252 12020 13280
rect 13725 13277 13737 13280
rect 13771 13277 13783 13311
rect 13725 13271 13783 13277
rect 14645 13311 14703 13317
rect 14645 13277 14657 13311
rect 14691 13308 14703 13311
rect 15194 13308 15200 13320
rect 14691 13280 15200 13308
rect 14691 13277 14703 13280
rect 14645 13271 14703 13277
rect 15194 13268 15200 13280
rect 15252 13268 15258 13320
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 15657 13311 15715 13317
rect 15657 13308 15669 13311
rect 15528 13280 15669 13308
rect 15528 13268 15534 13280
rect 15657 13277 15669 13280
rect 15703 13277 15715 13311
rect 15856 13308 15884 13339
rect 16114 13336 16120 13388
rect 16172 13376 16178 13388
rect 16577 13379 16635 13385
rect 16577 13376 16589 13379
rect 16172 13348 16589 13376
rect 16172 13336 16178 13348
rect 16577 13345 16589 13348
rect 16623 13345 16635 13379
rect 16577 13339 16635 13345
rect 16206 13308 16212 13320
rect 15856 13280 16212 13308
rect 15657 13271 15715 13277
rect 16206 13268 16212 13280
rect 16264 13268 16270 13320
rect 16390 13308 16396 13320
rect 16351 13280 16396 13308
rect 16390 13268 16396 13280
rect 16448 13268 16454 13320
rect 17052 13308 17080 13407
rect 18966 13404 18972 13416
rect 19024 13404 19030 13456
rect 19337 13447 19395 13453
rect 19337 13413 19349 13447
rect 19383 13444 19395 13447
rect 19518 13444 19524 13456
rect 19383 13416 19524 13444
rect 19383 13413 19395 13416
rect 19337 13407 19395 13413
rect 19518 13404 19524 13416
rect 19576 13404 19582 13456
rect 19610 13404 19616 13456
rect 19668 13444 19674 13456
rect 22922 13444 22928 13456
rect 19668 13416 22928 13444
rect 19668 13404 19674 13416
rect 22922 13404 22928 13416
rect 22980 13404 22986 13456
rect 17405 13379 17463 13385
rect 17405 13345 17417 13379
rect 17451 13376 17463 13379
rect 18138 13376 18144 13388
rect 17451 13348 18144 13376
rect 17451 13345 17463 13348
rect 17405 13339 17463 13345
rect 18138 13336 18144 13348
rect 18196 13336 18202 13388
rect 18693 13379 18751 13385
rect 18693 13345 18705 13379
rect 18739 13376 18751 13379
rect 19058 13376 19064 13388
rect 18739 13348 19064 13376
rect 18739 13345 18751 13348
rect 18693 13339 18751 13345
rect 19058 13336 19064 13348
rect 19116 13336 19122 13388
rect 20364 13348 20852 13376
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17052 13280 17509 13308
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 17497 13271 17555 13277
rect 17604 13280 20177 13308
rect 11974 13200 11980 13252
rect 12032 13200 12038 13252
rect 12526 13200 12532 13252
rect 12584 13240 12590 13252
rect 12584 13212 13308 13240
rect 12584 13200 12590 13212
rect 12250 13172 12256 13184
rect 11563 13144 12256 13172
rect 11563 13141 11575 13144
rect 11517 13135 11575 13141
rect 12250 13132 12256 13144
rect 12308 13132 12314 13184
rect 12986 13172 12992 13184
rect 12947 13144 12992 13172
rect 12986 13132 12992 13144
rect 13044 13132 13050 13184
rect 13078 13132 13084 13184
rect 13136 13172 13142 13184
rect 13280 13172 13308 13212
rect 13354 13200 13360 13252
rect 13412 13240 13418 13252
rect 13814 13240 13820 13252
rect 13412 13212 13457 13240
rect 13775 13212 13820 13240
rect 13412 13200 13418 13212
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 14737 13243 14795 13249
rect 14737 13240 14749 13243
rect 14200 13212 14749 13240
rect 13722 13172 13728 13184
rect 13136 13144 13181 13172
rect 13280 13144 13728 13172
rect 13136 13132 13142 13144
rect 13722 13132 13728 13144
rect 13780 13172 13786 13184
rect 14200 13181 14228 13212
rect 14737 13209 14749 13212
rect 14783 13209 14795 13243
rect 15102 13240 15108 13252
rect 14737 13203 14795 13209
rect 14844 13212 15108 13240
rect 14185 13175 14243 13181
rect 14185 13172 14197 13175
rect 13780 13144 14197 13172
rect 13780 13132 13786 13144
rect 14185 13141 14197 13144
rect 14231 13141 14243 13175
rect 14185 13135 14243 13141
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 14844 13172 14872 13212
rect 15102 13200 15108 13212
rect 15160 13240 15166 13252
rect 15930 13240 15936 13252
rect 15160 13212 15936 13240
rect 15160 13200 15166 13212
rect 15930 13200 15936 13212
rect 15988 13240 15994 13252
rect 16485 13243 16543 13249
rect 16485 13240 16497 13243
rect 15988 13212 16497 13240
rect 15988 13200 15994 13212
rect 16485 13209 16497 13212
rect 16531 13209 16543 13243
rect 16485 13203 16543 13209
rect 17604 13184 17632 13280
rect 20165 13277 20177 13280
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 18877 13243 18935 13249
rect 18877 13240 18889 13243
rect 18432 13212 18889 13240
rect 18432 13184 18460 13212
rect 18877 13209 18889 13212
rect 18923 13209 18935 13243
rect 18877 13203 18935 13209
rect 19518 13200 19524 13252
rect 19576 13240 19582 13252
rect 20364 13240 20392 13348
rect 20530 13308 20536 13320
rect 20491 13280 20536 13308
rect 20530 13268 20536 13280
rect 20588 13268 20594 13320
rect 20824 13317 20852 13348
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 20855 13280 21097 13308
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21266 13308 21272 13320
rect 21227 13280 21272 13308
rect 21085 13271 21143 13277
rect 21266 13268 21272 13280
rect 21324 13268 21330 13320
rect 19576 13212 20392 13240
rect 20441 13243 20499 13249
rect 19576 13200 19582 13212
rect 20441 13209 20453 13243
rect 20487 13240 20499 13243
rect 21818 13240 21824 13252
rect 20487 13212 21824 13240
rect 20487 13209 20499 13212
rect 20441 13203 20499 13209
rect 21818 13200 21824 13212
rect 21876 13200 21882 13252
rect 14700 13144 14872 13172
rect 15197 13175 15255 13181
rect 14700 13132 14706 13144
rect 15197 13141 15209 13175
rect 15243 13172 15255 13175
rect 15286 13172 15292 13184
rect 15243 13144 15292 13172
rect 15243 13141 15255 13144
rect 15197 13135 15255 13141
rect 15286 13132 15292 13144
rect 15344 13132 15350 13184
rect 15562 13172 15568 13184
rect 15523 13144 15568 13172
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 16206 13132 16212 13184
rect 16264 13172 16270 13184
rect 16390 13172 16396 13184
rect 16264 13144 16396 13172
rect 16264 13132 16270 13144
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 16945 13175 17003 13181
rect 16945 13141 16957 13175
rect 16991 13172 17003 13175
rect 17586 13172 17592 13184
rect 16991 13144 17592 13172
rect 16991 13141 17003 13144
rect 16945 13135 17003 13141
rect 17586 13132 17592 13144
rect 17644 13132 17650 13184
rect 18414 13172 18420 13184
rect 18375 13144 18420 13172
rect 18414 13132 18420 13144
rect 18472 13132 18478 13184
rect 18506 13132 18512 13184
rect 18564 13172 18570 13184
rect 19886 13172 19892 13184
rect 18564 13144 18609 13172
rect 19847 13144 19892 13172
rect 18564 13132 18570 13144
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 20070 13172 20076 13184
rect 20031 13144 20076 13172
rect 20070 13132 20076 13144
rect 20128 13132 20134 13184
rect 21450 13172 21456 13184
rect 21411 13144 21456 13172
rect 21450 13132 21456 13144
rect 21508 13132 21514 13184
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 1670 12928 1676 12980
rect 1728 12968 1734 12980
rect 3421 12971 3479 12977
rect 3421 12968 3433 12971
rect 1728 12940 3433 12968
rect 1728 12928 1734 12940
rect 3421 12937 3433 12940
rect 3467 12937 3479 12971
rect 4430 12968 4436 12980
rect 4391 12940 4436 12968
rect 3421 12931 3479 12937
rect 4430 12928 4436 12940
rect 4488 12928 4494 12980
rect 4890 12928 4896 12980
rect 4948 12968 4954 12980
rect 4948 12940 5212 12968
rect 4948 12928 4954 12940
rect 1857 12903 1915 12909
rect 1857 12869 1869 12903
rect 1903 12900 1915 12903
rect 2038 12900 2044 12912
rect 1903 12872 2044 12900
rect 1903 12869 1915 12872
rect 1857 12863 1915 12869
rect 2038 12860 2044 12872
rect 2096 12860 2102 12912
rect 2774 12860 2780 12912
rect 2832 12900 2838 12912
rect 3510 12900 3516 12912
rect 2832 12872 3516 12900
rect 2832 12860 2838 12872
rect 3510 12860 3516 12872
rect 3568 12860 3574 12912
rect 1670 12832 1676 12844
rect 1631 12804 1676 12832
rect 1670 12792 1676 12804
rect 1728 12792 1734 12844
rect 1762 12792 1768 12844
rect 1820 12832 1826 12844
rect 2205 12835 2263 12841
rect 2205 12832 2217 12835
rect 1820 12804 2217 12832
rect 1820 12792 1826 12804
rect 2205 12801 2217 12804
rect 2251 12801 2263 12835
rect 2205 12795 2263 12801
rect 3234 12792 3240 12844
rect 3292 12832 3298 12844
rect 3605 12835 3663 12841
rect 3605 12832 3617 12835
rect 3292 12804 3617 12832
rect 3292 12792 3298 12804
rect 3605 12801 3617 12804
rect 3651 12801 3663 12835
rect 4062 12832 4068 12844
rect 4023 12804 4068 12832
rect 3605 12795 3663 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 4338 12792 4344 12844
rect 4396 12832 4402 12844
rect 4893 12835 4951 12841
rect 4893 12832 4905 12835
rect 4396 12804 4905 12832
rect 4396 12792 4402 12804
rect 4893 12801 4905 12804
rect 4939 12801 4951 12835
rect 4893 12795 4951 12801
rect 4985 12835 5043 12841
rect 4985 12801 4997 12835
rect 5031 12832 5043 12835
rect 5074 12832 5080 12844
rect 5031 12804 5080 12832
rect 5031 12801 5043 12804
rect 4985 12795 5043 12801
rect 5074 12792 5080 12804
rect 5132 12792 5138 12844
rect 5184 12832 5212 12940
rect 5442 12928 5448 12980
rect 5500 12968 5506 12980
rect 5905 12971 5963 12977
rect 5905 12968 5917 12971
rect 5500 12940 5917 12968
rect 5500 12928 5506 12940
rect 5905 12937 5917 12940
rect 5951 12937 5963 12971
rect 5905 12931 5963 12937
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6549 12971 6607 12977
rect 6549 12968 6561 12971
rect 6052 12940 6561 12968
rect 6052 12928 6058 12940
rect 6472 12912 6500 12940
rect 6549 12937 6561 12940
rect 6595 12937 6607 12971
rect 6549 12931 6607 12937
rect 7374 12928 7380 12980
rect 7432 12968 7438 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7432 12940 7665 12968
rect 7432 12928 7438 12940
rect 7653 12937 7665 12940
rect 7699 12937 7711 12971
rect 8018 12968 8024 12980
rect 7979 12940 8024 12968
rect 7653 12931 7711 12937
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 8113 12971 8171 12977
rect 8113 12937 8125 12971
rect 8159 12968 8171 12971
rect 8662 12968 8668 12980
rect 8159 12940 8668 12968
rect 8159 12937 8171 12940
rect 8113 12931 8171 12937
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 9766 12968 9772 12980
rect 8956 12940 9772 12968
rect 6454 12860 6460 12912
rect 6512 12860 6518 12912
rect 6730 12860 6736 12912
rect 6788 12900 6794 12912
rect 6788 12872 7696 12900
rect 6788 12860 6794 12872
rect 5813 12835 5871 12841
rect 5813 12832 5825 12835
rect 5184 12804 5825 12832
rect 5813 12801 5825 12804
rect 5859 12832 5871 12835
rect 7190 12832 7196 12844
rect 5859 12804 7052 12832
rect 7151 12804 7196 12832
rect 5859 12801 5871 12804
rect 5813 12795 5871 12801
rect 1949 12767 2007 12773
rect 1949 12733 1961 12767
rect 1995 12733 2007 12767
rect 3878 12764 3884 12776
rect 3839 12736 3884 12764
rect 1949 12727 2007 12733
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 1964 12628 1992 12727
rect 3878 12724 3884 12736
rect 3936 12724 3942 12776
rect 3973 12767 4031 12773
rect 3973 12733 3985 12767
rect 4019 12764 4031 12767
rect 5169 12767 5227 12773
rect 5169 12764 5181 12767
rect 4019 12736 4568 12764
rect 4019 12733 4031 12736
rect 3973 12727 4031 12733
rect 3326 12696 3332 12708
rect 3287 12668 3332 12696
rect 3326 12656 3332 12668
rect 3384 12656 3390 12708
rect 4540 12705 4568 12736
rect 4632 12736 5181 12764
rect 4525 12699 4583 12705
rect 4525 12665 4537 12699
rect 4571 12665 4583 12699
rect 4525 12659 4583 12665
rect 2222 12628 2228 12640
rect 1964 12600 2228 12628
rect 2222 12588 2228 12600
rect 2280 12628 2286 12640
rect 2682 12628 2688 12640
rect 2280 12600 2688 12628
rect 2280 12588 2286 12600
rect 2682 12588 2688 12600
rect 2740 12588 2746 12640
rect 3970 12588 3976 12640
rect 4028 12628 4034 12640
rect 4632 12628 4660 12736
rect 5169 12733 5181 12736
rect 5215 12764 5227 12767
rect 6089 12767 6147 12773
rect 6089 12764 6101 12767
rect 5215 12736 6101 12764
rect 5215 12733 5227 12736
rect 5169 12727 5227 12733
rect 6089 12733 6101 12736
rect 6135 12764 6147 12767
rect 6822 12764 6828 12776
rect 6135 12736 6828 12764
rect 6135 12733 6147 12736
rect 6089 12727 6147 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 4982 12656 4988 12708
rect 5040 12696 5046 12708
rect 5445 12699 5503 12705
rect 5445 12696 5457 12699
rect 5040 12668 5457 12696
rect 5040 12656 5046 12668
rect 5445 12665 5457 12668
rect 5491 12665 5503 12699
rect 5445 12659 5503 12665
rect 6454 12656 6460 12708
rect 6512 12696 6518 12708
rect 6914 12696 6920 12708
rect 6512 12668 6920 12696
rect 6512 12656 6518 12668
rect 6914 12656 6920 12668
rect 6972 12656 6978 12708
rect 7024 12696 7052 12804
rect 7190 12792 7196 12804
rect 7248 12792 7254 12844
rect 7668 12832 7696 12872
rect 7742 12860 7748 12912
rect 7800 12900 7806 12912
rect 8754 12900 8760 12912
rect 7800 12872 8760 12900
rect 7800 12860 7806 12872
rect 8754 12860 8760 12872
rect 8812 12860 8818 12912
rect 8956 12841 8984 12940
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 10042 12928 10048 12980
rect 10100 12968 10106 12980
rect 10413 12971 10471 12977
rect 10413 12968 10425 12971
rect 10100 12940 10425 12968
rect 10100 12928 10106 12940
rect 10413 12937 10425 12940
rect 10459 12968 10471 12971
rect 10873 12971 10931 12977
rect 10873 12968 10885 12971
rect 10459 12940 10885 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 10873 12937 10885 12940
rect 10919 12937 10931 12971
rect 10873 12931 10931 12937
rect 10962 12928 10968 12980
rect 11020 12968 11026 12980
rect 11020 12940 11100 12968
rect 11020 12928 11026 12940
rect 9030 12860 9036 12912
rect 9088 12900 9094 12912
rect 9493 12903 9551 12909
rect 9493 12900 9505 12903
rect 9088 12872 9505 12900
rect 9088 12860 9094 12872
rect 9493 12869 9505 12872
rect 9539 12900 9551 12903
rect 10134 12900 10140 12912
rect 9539 12872 10140 12900
rect 9539 12869 9551 12872
rect 9493 12863 9551 12869
rect 10134 12860 10140 12872
rect 10192 12860 10198 12912
rect 11072 12900 11100 12940
rect 11238 12928 11244 12980
rect 11296 12968 11302 12980
rect 11333 12971 11391 12977
rect 11333 12968 11345 12971
rect 11296 12940 11345 12968
rect 11296 12928 11302 12940
rect 11333 12937 11345 12940
rect 11379 12937 11391 12971
rect 11333 12931 11391 12937
rect 12253 12971 12311 12977
rect 12253 12937 12265 12971
rect 12299 12968 12311 12971
rect 12342 12968 12348 12980
rect 12299 12940 12348 12968
rect 12299 12937 12311 12940
rect 12253 12931 12311 12937
rect 12342 12928 12348 12940
rect 12400 12928 12406 12980
rect 12621 12971 12679 12977
rect 12621 12937 12633 12971
rect 12667 12968 12679 12971
rect 13262 12968 13268 12980
rect 12667 12940 13268 12968
rect 12667 12937 12679 12940
rect 12621 12931 12679 12937
rect 13262 12928 13268 12940
rect 13320 12928 13326 12980
rect 14093 12971 14151 12977
rect 14093 12937 14105 12971
rect 14139 12968 14151 12971
rect 14918 12968 14924 12980
rect 14139 12940 14924 12968
rect 14139 12937 14151 12940
rect 14093 12931 14151 12937
rect 14918 12928 14924 12940
rect 14976 12928 14982 12980
rect 15286 12968 15292 12980
rect 15247 12940 15292 12968
rect 15286 12928 15292 12940
rect 15344 12928 15350 12980
rect 15654 12928 15660 12980
rect 15712 12968 15718 12980
rect 15749 12971 15807 12977
rect 15749 12968 15761 12971
rect 15712 12940 15761 12968
rect 15712 12928 15718 12940
rect 15749 12937 15761 12940
rect 15795 12937 15807 12971
rect 15749 12931 15807 12937
rect 15930 12928 15936 12980
rect 15988 12968 15994 12980
rect 16025 12971 16083 12977
rect 16025 12968 16037 12971
rect 15988 12940 16037 12968
rect 15988 12928 15994 12940
rect 16025 12937 16037 12940
rect 16071 12937 16083 12971
rect 16025 12931 16083 12937
rect 16669 12971 16727 12977
rect 16669 12937 16681 12971
rect 16715 12937 16727 12971
rect 16669 12931 16727 12937
rect 12986 12909 12992 12912
rect 11517 12903 11575 12909
rect 11517 12900 11529 12903
rect 11072 12872 11529 12900
rect 11517 12869 11529 12872
rect 11563 12869 11575 12903
rect 12980 12900 12992 12909
rect 11517 12863 11575 12869
rect 11992 12872 12992 12900
rect 8941 12835 8999 12841
rect 8941 12832 8953 12835
rect 7668 12804 8953 12832
rect 8941 12801 8953 12804
rect 8987 12801 8999 12835
rect 9784 12832 9996 12836
rect 10965 12835 11023 12841
rect 10965 12832 10977 12835
rect 8941 12795 8999 12801
rect 9692 12808 10977 12832
rect 9692 12804 9812 12808
rect 9968 12804 10977 12808
rect 7282 12764 7288 12776
rect 7243 12736 7288 12764
rect 7282 12724 7288 12736
rect 7340 12724 7346 12776
rect 7374 12724 7380 12776
rect 7432 12764 7438 12776
rect 7432 12736 7477 12764
rect 7432 12724 7438 12736
rect 7558 12724 7564 12776
rect 7616 12764 7622 12776
rect 8202 12764 8208 12776
rect 7616 12736 8208 12764
rect 7616 12724 7622 12736
rect 8202 12724 8208 12736
rect 8260 12724 8266 12776
rect 8478 12724 8484 12776
rect 8536 12764 8542 12776
rect 9033 12767 9091 12773
rect 9033 12764 9045 12767
rect 8536 12736 9045 12764
rect 8536 12724 8542 12736
rect 9033 12733 9045 12736
rect 9079 12733 9091 12767
rect 9033 12727 9091 12733
rect 8846 12696 8852 12708
rect 7024 12668 8852 12696
rect 8846 12656 8852 12668
rect 8904 12656 8910 12708
rect 4028 12600 4660 12628
rect 4028 12588 4034 12600
rect 5534 12588 5540 12640
rect 5592 12628 5598 12640
rect 5810 12628 5816 12640
rect 5592 12600 5816 12628
rect 5592 12588 5598 12600
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 6546 12588 6552 12640
rect 6604 12628 6610 12640
rect 6641 12631 6699 12637
rect 6641 12628 6653 12631
rect 6604 12600 6653 12628
rect 6604 12588 6610 12600
rect 6641 12597 6653 12600
rect 6687 12597 6699 12631
rect 6822 12628 6828 12640
rect 6783 12600 6828 12628
rect 6641 12591 6699 12597
rect 6822 12588 6828 12600
rect 6880 12588 6886 12640
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 8573 12631 8631 12637
rect 8573 12628 8585 12631
rect 8536 12600 8585 12628
rect 8536 12588 8542 12600
rect 8573 12597 8585 12600
rect 8619 12597 8631 12631
rect 9048 12628 9076 12727
rect 9122 12724 9128 12776
rect 9180 12764 9186 12776
rect 9180 12736 9225 12764
rect 9180 12724 9186 12736
rect 9214 12656 9220 12708
rect 9272 12696 9278 12708
rect 9692 12696 9720 12804
rect 10965 12801 10977 12804
rect 11011 12801 11023 12835
rect 10965 12795 11023 12801
rect 9766 12724 9772 12776
rect 9824 12764 9830 12776
rect 10781 12767 10839 12773
rect 9824 12736 9869 12764
rect 9824 12724 9830 12736
rect 10781 12733 10793 12767
rect 10827 12764 10839 12767
rect 10870 12764 10876 12776
rect 10827 12736 10876 12764
rect 10827 12733 10839 12736
rect 10781 12727 10839 12733
rect 10870 12724 10876 12736
rect 10928 12764 10934 12776
rect 11698 12764 11704 12776
rect 10928 12736 11704 12764
rect 10928 12724 10934 12736
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11992 12773 12020 12872
rect 12980 12863 12992 12872
rect 12986 12860 12992 12863
rect 13044 12860 13050 12912
rect 15381 12903 15439 12909
rect 15381 12869 15393 12903
rect 15427 12900 15439 12903
rect 16684 12900 16712 12931
rect 17586 12928 17592 12980
rect 17644 12968 17650 12980
rect 19337 12971 19395 12977
rect 19337 12968 19349 12971
rect 17644 12940 19349 12968
rect 17644 12928 17650 12940
rect 19337 12937 19349 12940
rect 19383 12937 19395 12971
rect 21542 12968 21548 12980
rect 19337 12931 19395 12937
rect 20548 12940 21548 12968
rect 18138 12909 18144 12912
rect 15427 12872 16712 12900
rect 17037 12903 17095 12909
rect 15427 12869 15439 12872
rect 15381 12863 15439 12869
rect 17037 12869 17049 12903
rect 17083 12900 17095 12903
rect 17083 12872 17724 12900
rect 17083 12869 17095 12872
rect 17037 12863 17095 12869
rect 12526 12792 12532 12844
rect 12584 12792 12590 12844
rect 12713 12835 12771 12841
rect 12713 12801 12725 12835
rect 12759 12832 12771 12835
rect 13538 12832 13544 12844
rect 12759 12804 13544 12832
rect 12759 12801 12771 12804
rect 12713 12795 12771 12801
rect 13538 12792 13544 12804
rect 13596 12832 13602 12844
rect 13722 12832 13728 12844
rect 13596 12804 13728 12832
rect 13596 12792 13602 12804
rect 13722 12792 13728 12804
rect 13780 12792 13786 12844
rect 15470 12792 15476 12844
rect 15528 12832 15534 12844
rect 15930 12832 15936 12844
rect 15528 12804 15936 12832
rect 15528 12792 15534 12804
rect 15930 12792 15936 12804
rect 15988 12792 15994 12844
rect 16390 12792 16396 12844
rect 16448 12832 16454 12844
rect 16942 12832 16948 12844
rect 16448 12804 16948 12832
rect 16448 12792 16454 12804
rect 16942 12792 16948 12804
rect 17000 12832 17006 12844
rect 17586 12832 17592 12844
rect 17000 12804 17264 12832
rect 17547 12804 17592 12832
rect 17000 12792 17006 12804
rect 11977 12767 12035 12773
rect 11977 12733 11989 12767
rect 12023 12733 12035 12767
rect 12158 12764 12164 12776
rect 12119 12736 12164 12764
rect 11977 12727 12035 12733
rect 12158 12724 12164 12736
rect 12216 12724 12222 12776
rect 9272 12668 9720 12696
rect 9272 12656 9278 12668
rect 11238 12656 11244 12708
rect 11296 12696 11302 12708
rect 12544 12696 12572 12792
rect 15197 12767 15255 12773
rect 15197 12733 15209 12767
rect 15243 12764 15255 12767
rect 16114 12764 16120 12776
rect 15243 12736 16120 12764
rect 15243 12733 15255 12736
rect 15197 12727 15255 12733
rect 16114 12724 16120 12736
rect 16172 12724 16178 12776
rect 16206 12724 16212 12776
rect 16264 12764 16270 12776
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 16264 12736 16313 12764
rect 16264 12724 16270 12736
rect 16301 12733 16313 12736
rect 16347 12764 16359 12767
rect 17034 12764 17040 12776
rect 16347 12736 17040 12764
rect 16347 12733 16359 12736
rect 16301 12727 16359 12733
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 17236 12773 17264 12804
rect 17586 12792 17592 12804
rect 17644 12792 17650 12844
rect 17129 12767 17187 12773
rect 17129 12733 17141 12767
rect 17175 12733 17187 12767
rect 17129 12727 17187 12733
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12733 17279 12767
rect 17221 12727 17279 12733
rect 11296 12668 12572 12696
rect 11296 12656 11302 12668
rect 14274 12656 14280 12708
rect 14332 12696 14338 12708
rect 14553 12699 14611 12705
rect 14553 12696 14565 12699
rect 14332 12668 14565 12696
rect 14332 12656 14338 12668
rect 14553 12665 14565 12668
rect 14599 12665 14611 12699
rect 14553 12659 14611 12665
rect 15562 12656 15568 12708
rect 15620 12696 15626 12708
rect 16393 12699 16451 12705
rect 16393 12696 16405 12699
rect 15620 12668 16405 12696
rect 15620 12656 15626 12668
rect 16393 12665 16405 12668
rect 16439 12696 16451 12699
rect 17144 12696 17172 12727
rect 16439 12668 17172 12696
rect 17696 12696 17724 12872
rect 18132 12863 18144 12909
rect 18196 12900 18202 12912
rect 18196 12872 18232 12900
rect 18138 12860 18144 12863
rect 18196 12860 18202 12872
rect 18690 12860 18696 12912
rect 18748 12900 18754 12912
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 18748 12872 19809 12900
rect 18748 12860 18754 12872
rect 19797 12869 19809 12872
rect 19843 12869 19855 12903
rect 19797 12863 19855 12869
rect 17770 12792 17776 12844
rect 17828 12832 17834 12844
rect 17865 12835 17923 12841
rect 17865 12832 17877 12835
rect 17828 12804 17877 12832
rect 17828 12792 17834 12804
rect 17865 12801 17877 12804
rect 17911 12832 17923 12835
rect 18984 12832 19288 12836
rect 19521 12835 19579 12841
rect 19521 12832 19533 12835
rect 17911 12808 19533 12832
rect 17911 12804 19012 12808
rect 19260 12804 19533 12808
rect 17911 12801 17923 12804
rect 17865 12795 17923 12801
rect 19521 12801 19533 12804
rect 19567 12801 19579 12835
rect 19521 12795 19579 12801
rect 20548 12764 20576 12940
rect 21542 12928 21548 12940
rect 21600 12928 21606 12980
rect 20625 12903 20683 12909
rect 20625 12869 20637 12903
rect 20671 12900 20683 12903
rect 21634 12900 21640 12912
rect 20671 12872 21640 12900
rect 20671 12869 20683 12872
rect 20625 12863 20683 12869
rect 21634 12860 21640 12872
rect 21692 12860 21698 12912
rect 20809 12835 20867 12841
rect 20809 12801 20821 12835
rect 20855 12832 20867 12835
rect 21174 12832 21180 12844
rect 20855 12804 21180 12832
rect 20855 12801 20867 12804
rect 20809 12795 20867 12801
rect 21174 12792 21180 12804
rect 21232 12792 21238 12844
rect 21269 12835 21327 12841
rect 21269 12801 21281 12835
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 18892 12736 20576 12764
rect 17696 12668 17908 12696
rect 16439 12665 16451 12668
rect 16393 12659 16451 12665
rect 9585 12631 9643 12637
rect 9585 12628 9597 12631
rect 9048 12600 9597 12628
rect 8573 12591 8631 12597
rect 9585 12597 9597 12600
rect 9631 12597 9643 12631
rect 10042 12628 10048 12640
rect 10003 12600 10048 12628
rect 9585 12591 9643 12597
rect 10042 12588 10048 12600
rect 10100 12588 10106 12640
rect 10229 12631 10287 12637
rect 10229 12597 10241 12631
rect 10275 12628 10287 12631
rect 10502 12628 10508 12640
rect 10275 12600 10508 12628
rect 10275 12597 10287 12600
rect 10229 12591 10287 12597
rect 10502 12588 10508 12600
rect 10560 12588 10566 12640
rect 11790 12628 11796 12640
rect 11751 12600 11796 12628
rect 11790 12588 11796 12600
rect 11848 12588 11854 12640
rect 12618 12588 12624 12640
rect 12676 12628 12682 12640
rect 14185 12631 14243 12637
rect 14185 12628 14197 12631
rect 12676 12600 14197 12628
rect 12676 12588 12682 12600
rect 14185 12597 14197 12600
rect 14231 12597 14243 12631
rect 14458 12628 14464 12640
rect 14419 12600 14464 12628
rect 14185 12591 14243 12597
rect 14458 12588 14464 12600
rect 14516 12588 14522 12640
rect 14642 12588 14648 12640
rect 14700 12628 14706 12640
rect 14737 12631 14795 12637
rect 14737 12628 14749 12631
rect 14700 12600 14749 12628
rect 14700 12588 14706 12600
rect 14737 12597 14749 12600
rect 14783 12597 14795 12631
rect 14737 12591 14795 12597
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 16114 12628 16120 12640
rect 15068 12600 16120 12628
rect 15068 12588 15074 12600
rect 16114 12588 16120 12600
rect 16172 12588 16178 12640
rect 17770 12628 17776 12640
rect 17731 12600 17776 12628
rect 17770 12588 17776 12600
rect 17828 12588 17834 12640
rect 17880 12628 17908 12668
rect 18892 12628 18920 12736
rect 20714 12724 20720 12776
rect 20772 12764 20778 12776
rect 21284 12764 21312 12795
rect 20772 12736 21312 12764
rect 20772 12724 20778 12736
rect 18966 12656 18972 12708
rect 19024 12696 19030 12708
rect 19981 12699 20039 12705
rect 19981 12696 19993 12699
rect 19024 12668 19993 12696
rect 19024 12656 19030 12668
rect 19981 12665 19993 12668
rect 20027 12665 20039 12699
rect 19981 12659 20039 12665
rect 20441 12699 20499 12705
rect 20441 12665 20453 12699
rect 20487 12696 20499 12699
rect 21082 12696 21088 12708
rect 20487 12668 21088 12696
rect 20487 12665 20499 12668
rect 20441 12659 20499 12665
rect 21082 12656 21088 12668
rect 21140 12656 21146 12708
rect 21177 12699 21235 12705
rect 21177 12665 21189 12699
rect 21223 12696 21235 12699
rect 21358 12696 21364 12708
rect 21223 12668 21364 12696
rect 21223 12665 21235 12668
rect 21177 12659 21235 12665
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 17880 12600 18920 12628
rect 19058 12588 19064 12640
rect 19116 12628 19122 12640
rect 19245 12631 19303 12637
rect 19245 12628 19257 12631
rect 19116 12600 19257 12628
rect 19116 12588 19122 12600
rect 19245 12597 19257 12600
rect 19291 12597 19303 12631
rect 19702 12628 19708 12640
rect 19663 12600 19708 12628
rect 19245 12591 19303 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 20254 12628 20260 12640
rect 20215 12600 20260 12628
rect 20254 12588 20260 12600
rect 20312 12588 20318 12640
rect 20990 12628 20996 12640
rect 20951 12600 20996 12628
rect 20990 12588 20996 12600
rect 21048 12588 21054 12640
rect 21450 12628 21456 12640
rect 21411 12600 21456 12628
rect 21450 12588 21456 12600
rect 21508 12588 21514 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 1762 12424 1768 12436
rect 1627 12396 1768 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 1762 12384 1768 12396
rect 1820 12384 1826 12436
rect 2682 12384 2688 12436
rect 2740 12424 2746 12436
rect 3234 12424 3240 12436
rect 2740 12396 3004 12424
rect 3195 12396 3240 12424
rect 2740 12384 2746 12396
rect 2976 12297 3004 12396
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 3789 12427 3847 12433
rect 3789 12393 3801 12427
rect 3835 12424 3847 12427
rect 4062 12424 4068 12436
rect 3835 12396 4068 12424
rect 3835 12393 3847 12396
rect 3789 12387 3847 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 5350 12424 5356 12436
rect 5132 12396 5356 12424
rect 5132 12384 5138 12396
rect 5350 12384 5356 12396
rect 5408 12384 5414 12436
rect 7006 12424 7012 12436
rect 5460 12396 7012 12424
rect 3050 12316 3056 12368
rect 3108 12356 3114 12368
rect 3108 12328 4476 12356
rect 3108 12316 3114 12328
rect 2961 12291 3019 12297
rect 2961 12257 2973 12291
rect 3007 12257 3019 12291
rect 2961 12251 3019 12257
rect 3970 12248 3976 12300
rect 4028 12288 4034 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 4028 12260 4353 12288
rect 4028 12248 4034 12260
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4448 12288 4476 12328
rect 4614 12316 4620 12368
rect 4672 12356 4678 12368
rect 4709 12359 4767 12365
rect 4709 12356 4721 12359
rect 4672 12328 4721 12356
rect 4672 12316 4678 12328
rect 4709 12325 4721 12328
rect 4755 12356 4767 12359
rect 5460 12356 5488 12396
rect 7006 12384 7012 12396
rect 7064 12384 7070 12436
rect 7190 12424 7196 12436
rect 7151 12396 7196 12424
rect 7190 12384 7196 12396
rect 7248 12384 7254 12436
rect 7282 12384 7288 12436
rect 7340 12424 7346 12436
rect 8021 12427 8079 12433
rect 8021 12424 8033 12427
rect 7340 12396 8033 12424
rect 7340 12384 7346 12396
rect 8021 12393 8033 12396
rect 8067 12393 8079 12427
rect 8021 12387 8079 12393
rect 8110 12384 8116 12436
rect 8168 12424 8174 12436
rect 9214 12424 9220 12436
rect 8168 12396 9220 12424
rect 8168 12384 8174 12396
rect 9214 12384 9220 12396
rect 9272 12384 9278 12436
rect 10318 12384 10324 12436
rect 10376 12384 10382 12436
rect 11698 12384 11704 12436
rect 11756 12424 11762 12436
rect 11793 12427 11851 12433
rect 11793 12424 11805 12427
rect 11756 12396 11805 12424
rect 11756 12384 11762 12396
rect 11793 12393 11805 12396
rect 11839 12393 11851 12427
rect 11793 12387 11851 12393
rect 11885 12427 11943 12433
rect 11885 12393 11897 12427
rect 11931 12424 11943 12427
rect 12158 12424 12164 12436
rect 11931 12396 12164 12424
rect 11931 12393 11943 12396
rect 11885 12387 11943 12393
rect 8941 12359 8999 12365
rect 8941 12356 8953 12359
rect 4755 12328 5488 12356
rect 7760 12328 8953 12356
rect 4755 12325 4767 12328
rect 4709 12319 4767 12325
rect 4448 12260 5212 12288
rect 4341 12251 4399 12257
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 1360 12192 2820 12220
rect 1360 12180 1366 12192
rect 2406 12152 2412 12164
rect 1504 12124 2412 12152
rect 1504 12096 1532 12124
rect 2406 12112 2412 12124
rect 2464 12112 2470 12164
rect 2498 12112 2504 12164
rect 2556 12152 2562 12164
rect 2694 12155 2752 12161
rect 2694 12152 2706 12155
rect 2556 12124 2706 12152
rect 2556 12112 2562 12124
rect 2694 12121 2706 12124
rect 2740 12121 2752 12155
rect 2792 12152 2820 12192
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 3053 12223 3111 12229
rect 3053 12220 3065 12223
rect 2924 12192 3065 12220
rect 2924 12180 2930 12192
rect 3053 12189 3065 12192
rect 3099 12189 3111 12223
rect 3053 12183 3111 12189
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12220 3571 12223
rect 3878 12220 3884 12232
rect 3559 12192 3884 12220
rect 3559 12189 3571 12192
rect 3513 12183 3571 12189
rect 3878 12180 3884 12192
rect 3936 12180 3942 12232
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4246 12220 4252 12232
rect 4203 12192 4252 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4522 12152 4528 12164
rect 2792 12124 4528 12152
rect 2694 12115 2752 12121
rect 4522 12112 4528 12124
rect 4580 12112 4586 12164
rect 4982 12112 4988 12164
rect 5040 12152 5046 12164
rect 5077 12155 5135 12161
rect 5077 12152 5089 12155
rect 5040 12124 5089 12152
rect 5040 12112 5046 12124
rect 5077 12121 5089 12124
rect 5123 12121 5135 12155
rect 5184 12152 5212 12260
rect 5718 12248 5724 12300
rect 5776 12288 5782 12300
rect 5994 12288 6000 12300
rect 5776 12260 6000 12288
rect 5776 12248 5782 12260
rect 5994 12248 6000 12260
rect 6052 12248 6058 12300
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7760 12297 7788 12328
rect 7745 12291 7803 12297
rect 7745 12288 7757 12291
rect 7248 12260 7757 12288
rect 7248 12248 7254 12260
rect 7745 12257 7757 12260
rect 7791 12257 7803 12291
rect 8478 12288 8484 12300
rect 8439 12260 8484 12288
rect 7745 12251 7803 12257
rect 8478 12248 8484 12260
rect 8536 12248 8542 12300
rect 8588 12297 8616 12328
rect 8941 12325 8953 12328
rect 8987 12325 8999 12359
rect 8941 12319 8999 12325
rect 10336 12297 10364 12384
rect 11808 12356 11836 12387
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 13817 12427 13875 12433
rect 13817 12393 13829 12427
rect 13863 12424 13875 12427
rect 14366 12424 14372 12436
rect 13863 12396 14372 12424
rect 13863 12393 13875 12396
rect 13817 12387 13875 12393
rect 14366 12384 14372 12396
rect 14424 12384 14430 12436
rect 15746 12424 15752 12436
rect 14476 12396 15752 12424
rect 12066 12356 12072 12368
rect 11808 12328 12072 12356
rect 12066 12316 12072 12328
rect 12124 12316 12130 12368
rect 12250 12316 12256 12368
rect 12308 12356 12314 12368
rect 12805 12359 12863 12365
rect 12308 12328 12480 12356
rect 12308 12316 12314 12328
rect 8573 12291 8631 12297
rect 8573 12257 8585 12291
rect 8619 12257 8631 12291
rect 8573 12251 8631 12257
rect 10314 12291 10372 12297
rect 10314 12257 10326 12291
rect 10360 12257 10372 12291
rect 10314 12251 10372 12257
rect 10410 12248 10416 12300
rect 10468 12288 10474 12300
rect 10468 12260 10513 12288
rect 10468 12248 10474 12260
rect 11790 12248 11796 12300
rect 11848 12288 11854 12300
rect 12158 12288 12164 12300
rect 11848 12260 12164 12288
rect 11848 12248 11854 12260
rect 12158 12248 12164 12260
rect 12216 12248 12222 12300
rect 12452 12297 12480 12328
rect 12805 12325 12817 12359
rect 12851 12325 12863 12359
rect 12805 12319 12863 12325
rect 12437 12291 12495 12297
rect 12437 12257 12449 12291
rect 12483 12257 12495 12291
rect 12437 12251 12495 12257
rect 5902 12180 5908 12232
rect 5960 12220 5966 12232
rect 5960 12192 6224 12220
rect 5960 12180 5966 12192
rect 6196 12152 6224 12192
rect 6730 12180 6736 12232
rect 6788 12229 6794 12232
rect 6788 12220 6800 12229
rect 7009 12223 7067 12229
rect 6788 12192 6833 12220
rect 6788 12183 6800 12192
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7098 12220 7104 12232
rect 7055 12192 7104 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 6788 12180 6794 12183
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9824 12192 10180 12220
rect 9824 12180 9830 12192
rect 6822 12152 6828 12164
rect 5184 12124 6132 12152
rect 6196 12124 6828 12152
rect 5077 12115 5135 12121
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 1670 12044 1676 12096
rect 1728 12084 1734 12096
rect 3329 12087 3387 12093
rect 3329 12084 3341 12087
rect 1728 12056 3341 12084
rect 1728 12044 1734 12056
rect 3329 12053 3341 12056
rect 3375 12053 3387 12087
rect 3329 12047 3387 12053
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12084 4307 12087
rect 4614 12084 4620 12096
rect 4295 12056 4620 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 4890 12084 4896 12096
rect 4851 12056 4896 12084
rect 4890 12044 4896 12056
rect 4948 12044 4954 12096
rect 5350 12044 5356 12096
rect 5408 12084 5414 12096
rect 5445 12087 5503 12093
rect 5445 12084 5457 12087
rect 5408 12056 5457 12084
rect 5408 12044 5414 12056
rect 5445 12053 5457 12056
rect 5491 12053 5503 12087
rect 5445 12047 5503 12053
rect 5629 12087 5687 12093
rect 5629 12053 5641 12087
rect 5675 12084 5687 12087
rect 5994 12084 6000 12096
rect 5675 12056 6000 12084
rect 5675 12053 5687 12056
rect 5629 12047 5687 12053
rect 5994 12044 6000 12056
rect 6052 12044 6058 12096
rect 6104 12084 6132 12124
rect 6822 12112 6828 12124
rect 6880 12112 6886 12164
rect 7024 12124 8984 12152
rect 7024 12084 7052 12124
rect 6104 12056 7052 12084
rect 7374 12044 7380 12096
rect 7432 12084 7438 12096
rect 7561 12087 7619 12093
rect 7561 12084 7573 12087
rect 7432 12056 7573 12084
rect 7432 12044 7438 12056
rect 7561 12053 7573 12056
rect 7607 12053 7619 12087
rect 7561 12047 7619 12053
rect 7650 12044 7656 12096
rect 7708 12084 7714 12096
rect 8389 12087 8447 12093
rect 7708 12056 7753 12084
rect 7708 12044 7714 12056
rect 8389 12053 8401 12087
rect 8435 12084 8447 12087
rect 8846 12084 8852 12096
rect 8435 12056 8852 12084
rect 8435 12053 8447 12056
rect 8389 12047 8447 12053
rect 8846 12044 8852 12056
rect 8904 12044 8910 12096
rect 8956 12084 8984 12124
rect 9122 12112 9128 12164
rect 9180 12152 9186 12164
rect 10054 12155 10112 12161
rect 10054 12152 10066 12155
rect 9180 12124 10066 12152
rect 9180 12112 9186 12124
rect 10054 12121 10066 12124
rect 10100 12121 10112 12155
rect 10152 12152 10180 12192
rect 10502 12180 10508 12232
rect 10560 12180 10566 12232
rect 10962 12180 10968 12232
rect 11020 12220 11026 12232
rect 11882 12220 11888 12232
rect 11020 12192 11888 12220
rect 11020 12180 11026 12192
rect 11882 12180 11888 12192
rect 11940 12180 11946 12232
rect 12253 12223 12311 12229
rect 12253 12189 12265 12223
rect 12299 12220 12311 12223
rect 12526 12220 12532 12232
rect 12299 12192 12532 12220
rect 12299 12189 12311 12192
rect 12253 12183 12311 12189
rect 12526 12180 12532 12192
rect 12584 12180 12590 12232
rect 10520 12152 10548 12180
rect 10152 12124 10548 12152
rect 10680 12155 10738 12161
rect 10054 12115 10112 12121
rect 10680 12121 10692 12155
rect 10726 12152 10738 12155
rect 11146 12152 11152 12164
rect 10726 12124 11152 12152
rect 10726 12121 10738 12124
rect 10680 12115 10738 12121
rect 11146 12112 11152 12124
rect 11204 12112 11210 12164
rect 11606 12112 11612 12164
rect 11664 12152 11670 12164
rect 12820 12152 12848 12319
rect 12986 12316 12992 12368
rect 13044 12356 13050 12368
rect 13081 12359 13139 12365
rect 13081 12356 13093 12359
rect 13044 12328 13093 12356
rect 13044 12316 13050 12328
rect 13081 12325 13093 12328
rect 13127 12325 13139 12359
rect 13081 12319 13139 12325
rect 13630 12316 13636 12368
rect 13688 12356 13694 12368
rect 14476 12356 14504 12396
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 15838 12384 15844 12436
rect 15896 12424 15902 12436
rect 16390 12424 16396 12436
rect 15896 12396 16396 12424
rect 15896 12384 15902 12396
rect 16390 12384 16396 12396
rect 16448 12384 16454 12436
rect 16761 12427 16819 12433
rect 16761 12393 16773 12427
rect 16807 12424 16819 12427
rect 17218 12424 17224 12436
rect 16807 12396 17224 12424
rect 16807 12393 16819 12396
rect 16761 12387 16819 12393
rect 17218 12384 17224 12396
rect 17276 12384 17282 12436
rect 18874 12384 18880 12436
rect 18932 12424 18938 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18932 12396 19257 12424
rect 18932 12384 18938 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 20257 12427 20315 12433
rect 20257 12393 20269 12427
rect 20303 12424 20315 12427
rect 20530 12424 20536 12436
rect 20303 12396 20536 12424
rect 20303 12393 20315 12396
rect 20257 12387 20315 12393
rect 20530 12384 20536 12396
rect 20588 12384 20594 12436
rect 20622 12384 20628 12436
rect 20680 12384 20686 12436
rect 20993 12427 21051 12433
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21266 12424 21272 12436
rect 21039 12396 21272 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 13688 12328 14504 12356
rect 13688 12316 13694 12328
rect 16114 12316 16120 12368
rect 16172 12356 16178 12368
rect 17310 12356 17316 12368
rect 16172 12328 17316 12356
rect 16172 12316 16178 12328
rect 17310 12316 17316 12328
rect 17368 12316 17374 12368
rect 20640 12356 20668 12384
rect 20806 12356 20812 12368
rect 18708 12328 19932 12356
rect 20640 12328 20812 12356
rect 13722 12288 13728 12300
rect 13004 12260 13728 12288
rect 13004 12232 13032 12260
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 16574 12288 16580 12300
rect 16487 12260 16580 12288
rect 16574 12248 16580 12260
rect 16632 12288 16638 12300
rect 17034 12288 17040 12300
rect 16632 12260 17040 12288
rect 16632 12248 16638 12260
rect 17034 12248 17040 12260
rect 17092 12288 17098 12300
rect 17402 12288 17408 12300
rect 17092 12260 17408 12288
rect 17092 12248 17098 12260
rect 17402 12248 17408 12260
rect 17460 12248 17466 12300
rect 17678 12288 17684 12300
rect 17639 12260 17684 12288
rect 17678 12248 17684 12260
rect 17736 12248 17742 12300
rect 12986 12220 12992 12232
rect 12899 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 14366 12180 14372 12232
rect 14424 12220 14430 12232
rect 14553 12223 14611 12229
rect 14553 12220 14565 12223
rect 14424 12192 14565 12220
rect 14424 12180 14430 12192
rect 14553 12189 14565 12192
rect 14599 12189 14611 12223
rect 14553 12183 14611 12189
rect 14829 12223 14887 12229
rect 14829 12189 14841 12223
rect 14875 12220 14887 12223
rect 15378 12220 15384 12232
rect 14875 12192 15384 12220
rect 14875 12189 14887 12192
rect 14829 12183 14887 12189
rect 15378 12180 15384 12192
rect 15436 12220 15442 12232
rect 16298 12220 16304 12232
rect 15436 12192 16304 12220
rect 15436 12180 15442 12192
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 18708 12220 18736 12328
rect 19242 12288 19248 12300
rect 16448 12192 18736 12220
rect 19076 12260 19248 12288
rect 16448 12180 16454 12192
rect 11664 12124 12848 12152
rect 13357 12155 13415 12161
rect 11664 12112 11670 12124
rect 13357 12121 13369 12155
rect 13403 12152 13415 12155
rect 13403 12124 14596 12152
rect 13403 12121 13415 12124
rect 13357 12115 13415 12121
rect 9950 12084 9956 12096
rect 8956 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10502 12044 10508 12096
rect 10560 12084 10566 12096
rect 11238 12084 11244 12096
rect 10560 12056 11244 12084
rect 10560 12044 10566 12056
rect 11238 12044 11244 12056
rect 11296 12044 11302 12096
rect 12342 12084 12348 12096
rect 12303 12056 12348 12084
rect 12342 12044 12348 12056
rect 12400 12044 12406 12096
rect 13449 12087 13507 12093
rect 13449 12053 13461 12087
rect 13495 12084 13507 12087
rect 13538 12084 13544 12096
rect 13495 12056 13544 12084
rect 13495 12053 13507 12056
rect 13449 12047 13507 12053
rect 13538 12044 13544 12056
rect 13596 12044 13602 12096
rect 14090 12084 14096 12096
rect 14051 12056 14096 12084
rect 14090 12044 14096 12056
rect 14148 12044 14154 12096
rect 14369 12087 14427 12093
rect 14369 12053 14381 12087
rect 14415 12084 14427 12087
rect 14458 12084 14464 12096
rect 14415 12056 14464 12084
rect 14415 12053 14427 12056
rect 14369 12047 14427 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14568 12084 14596 12124
rect 14734 12112 14740 12164
rect 14792 12152 14798 12164
rect 15074 12155 15132 12161
rect 15074 12152 15086 12155
rect 14792 12124 15086 12152
rect 14792 12112 14798 12124
rect 15074 12121 15086 12124
rect 15120 12121 15132 12155
rect 15074 12115 15132 12121
rect 16666 12112 16672 12164
rect 16724 12112 16730 12164
rect 16758 12112 16764 12164
rect 16816 12112 16822 12164
rect 16942 12112 16948 12164
rect 17000 12152 17006 12164
rect 17678 12152 17684 12164
rect 17000 12124 17684 12152
rect 17000 12112 17006 12124
rect 17678 12112 17684 12124
rect 17736 12112 17742 12164
rect 17948 12155 18006 12161
rect 17948 12121 17960 12155
rect 17994 12152 18006 12155
rect 18230 12152 18236 12164
rect 17994 12124 18236 12152
rect 17994 12121 18006 12124
rect 17948 12115 18006 12121
rect 18230 12112 18236 12124
rect 18288 12112 18294 12164
rect 15286 12084 15292 12096
rect 14568 12056 15292 12084
rect 15286 12044 15292 12056
rect 15344 12084 15350 12096
rect 15654 12084 15660 12096
rect 15344 12056 15660 12084
rect 15344 12044 15350 12056
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16206 12084 16212 12096
rect 16167 12056 16212 12084
rect 16206 12044 16212 12056
rect 16264 12044 16270 12096
rect 16393 12087 16451 12093
rect 16393 12053 16405 12087
rect 16439 12084 16451 12087
rect 16684 12084 16712 12112
rect 16439 12056 16712 12084
rect 16776 12084 16804 12112
rect 17037 12087 17095 12093
rect 17037 12084 17049 12087
rect 16776 12056 17049 12084
rect 16439 12053 16451 12056
rect 16393 12047 16451 12053
rect 17037 12053 17049 12056
rect 17083 12053 17095 12087
rect 17218 12084 17224 12096
rect 17179 12056 17224 12084
rect 17037 12047 17095 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 17494 12084 17500 12096
rect 17455 12056 17500 12084
rect 17494 12044 17500 12056
rect 17552 12044 17558 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 19076 12093 19104 12260
rect 19242 12248 19248 12260
rect 19300 12288 19306 12300
rect 19797 12291 19855 12297
rect 19797 12288 19809 12291
rect 19300 12260 19809 12288
rect 19300 12248 19306 12260
rect 19797 12257 19809 12260
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 19610 12152 19616 12164
rect 19571 12124 19616 12152
rect 19610 12112 19616 12124
rect 19668 12112 19674 12164
rect 19702 12112 19708 12164
rect 19760 12152 19766 12164
rect 19904 12152 19932 12328
rect 20806 12316 20812 12328
rect 20864 12316 20870 12368
rect 19978 12248 19984 12300
rect 20036 12288 20042 12300
rect 21082 12288 21088 12300
rect 20036 12260 21088 12288
rect 20036 12248 20042 12260
rect 21082 12248 21088 12260
rect 21140 12248 21146 12300
rect 21542 12248 21548 12300
rect 21600 12288 21606 12300
rect 22186 12288 22192 12300
rect 21600 12260 22192 12288
rect 21600 12248 21606 12260
rect 22186 12248 22192 12260
rect 22244 12248 22250 12300
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20809 12223 20867 12229
rect 20809 12220 20821 12223
rect 20073 12183 20131 12189
rect 20272 12192 20821 12220
rect 19760 12124 19932 12152
rect 19760 12112 19766 12124
rect 19061 12087 19119 12093
rect 19061 12084 19073 12087
rect 18196 12056 19073 12084
rect 18196 12044 18202 12056
rect 19061 12053 19073 12056
rect 19107 12053 19119 12087
rect 19061 12047 19119 12053
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 20088 12084 20116 12183
rect 20272 12164 20300 12192
rect 20809 12189 20821 12192
rect 20855 12189 20867 12223
rect 21269 12223 21327 12229
rect 21269 12220 21281 12223
rect 20809 12183 20867 12189
rect 20916 12192 21281 12220
rect 20254 12112 20260 12164
rect 20312 12112 20318 12164
rect 20346 12112 20352 12164
rect 20404 12152 20410 12164
rect 20916 12152 20944 12192
rect 21269 12189 21281 12192
rect 21315 12189 21327 12223
rect 21269 12183 21327 12189
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21508 12192 21956 12220
rect 21508 12180 21514 12192
rect 20404 12124 20944 12152
rect 21177 12155 21235 12161
rect 20404 12112 20410 12124
rect 21177 12121 21189 12155
rect 21223 12152 21235 12155
rect 21542 12152 21548 12164
rect 21223 12124 21548 12152
rect 21223 12121 21235 12124
rect 21177 12115 21235 12121
rect 21542 12112 21548 12124
rect 21600 12112 21606 12164
rect 20530 12084 20536 12096
rect 19208 12056 20116 12084
rect 20491 12056 20536 12084
rect 19208 12044 19214 12056
rect 20530 12044 20536 12056
rect 20588 12044 20594 12096
rect 20717 12087 20775 12093
rect 20717 12053 20729 12087
rect 20763 12084 20775 12087
rect 21082 12084 21088 12096
rect 20763 12056 21088 12084
rect 20763 12053 20775 12056
rect 20717 12047 20775 12053
rect 21082 12044 21088 12056
rect 21140 12044 21146 12096
rect 21450 12084 21456 12096
rect 21411 12056 21456 12084
rect 21450 12044 21456 12056
rect 21508 12044 21514 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2777 11883 2835 11889
rect 2777 11880 2789 11883
rect 1728 11852 2789 11880
rect 1728 11840 1734 11852
rect 2777 11849 2789 11852
rect 2823 11849 2835 11883
rect 3050 11880 3056 11892
rect 2777 11843 2835 11849
rect 2976 11852 3056 11880
rect 2976 11812 3004 11852
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 3145 11883 3203 11889
rect 3145 11849 3157 11883
rect 3191 11880 3203 11883
rect 3605 11883 3663 11889
rect 3605 11880 3617 11883
rect 3191 11852 3617 11880
rect 3191 11849 3203 11852
rect 3145 11843 3203 11849
rect 3605 11849 3617 11852
rect 3651 11849 3663 11883
rect 3605 11843 3663 11849
rect 4154 11840 4160 11892
rect 4212 11880 4218 11892
rect 4433 11883 4491 11889
rect 4433 11880 4445 11883
rect 4212 11852 4445 11880
rect 4212 11840 4218 11852
rect 4433 11849 4445 11852
rect 4479 11849 4491 11883
rect 4433 11843 4491 11849
rect 5258 11840 5264 11892
rect 5316 11880 5322 11892
rect 5445 11883 5503 11889
rect 5445 11880 5457 11883
rect 5316 11852 5457 11880
rect 5316 11840 5322 11852
rect 5445 11849 5457 11852
rect 5491 11849 5503 11883
rect 7282 11880 7288 11892
rect 5445 11843 5503 11849
rect 5644 11852 6224 11880
rect 2240 11784 3004 11812
rect 3068 11784 5304 11812
rect 1854 11704 1860 11756
rect 1912 11744 1918 11756
rect 1912 11716 2075 11744
rect 1912 11704 1918 11716
rect 1949 11679 2007 11685
rect 1949 11645 1961 11679
rect 1995 11645 2007 11679
rect 2047 11676 2075 11716
rect 2130 11704 2136 11756
rect 2188 11744 2194 11756
rect 2240 11753 2268 11784
rect 2225 11747 2283 11753
rect 2225 11744 2237 11747
rect 2188 11716 2237 11744
rect 2188 11704 2194 11716
rect 2225 11713 2237 11716
rect 2271 11713 2283 11747
rect 2225 11707 2283 11713
rect 2409 11747 2467 11753
rect 2409 11713 2421 11747
rect 2455 11744 2467 11747
rect 3068 11744 3096 11784
rect 5276 11756 5304 11784
rect 3973 11747 4031 11753
rect 2455 11716 3096 11744
rect 3160 11716 3924 11744
rect 2455 11713 2467 11716
rect 2409 11707 2467 11713
rect 2424 11676 2452 11707
rect 2047 11648 2452 11676
rect 2593 11679 2651 11685
rect 1949 11639 2007 11645
rect 2593 11645 2605 11679
rect 2639 11676 2651 11679
rect 3160 11676 3188 11716
rect 2639 11648 3188 11676
rect 3237 11679 3295 11685
rect 2639 11645 2651 11648
rect 2593 11639 2651 11645
rect 3237 11645 3249 11679
rect 3283 11645 3295 11679
rect 3237 11639 3295 11645
rect 1964 11540 1992 11639
rect 2406 11540 2412 11552
rect 1964 11512 2412 11540
rect 2406 11500 2412 11512
rect 2464 11500 2470 11552
rect 3252 11540 3280 11639
rect 3326 11636 3332 11688
rect 3384 11676 3390 11688
rect 3384 11648 3429 11676
rect 3384 11636 3390 11648
rect 3896 11608 3924 11716
rect 3973 11713 3985 11747
rect 4019 11744 4031 11747
rect 4246 11744 4252 11756
rect 4019 11716 4252 11744
rect 4019 11713 4031 11716
rect 3973 11707 4031 11713
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4614 11744 4620 11756
rect 4575 11716 4620 11744
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 5258 11704 5264 11756
rect 5316 11704 5322 11756
rect 5644 11744 5672 11852
rect 5902 11812 5908 11824
rect 5863 11784 5908 11812
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 5810 11744 5816 11756
rect 5460 11716 5672 11744
rect 5771 11716 5816 11744
rect 4062 11676 4068 11688
rect 4023 11648 4068 11676
rect 4062 11636 4068 11648
rect 4120 11636 4126 11688
rect 4154 11636 4160 11688
rect 4212 11676 4218 11688
rect 4212 11648 4257 11676
rect 4212 11636 4218 11648
rect 4982 11636 4988 11688
rect 5040 11676 5046 11688
rect 5077 11679 5135 11685
rect 5077 11676 5089 11679
rect 5040 11648 5089 11676
rect 5040 11636 5046 11648
rect 5077 11645 5089 11648
rect 5123 11676 5135 11679
rect 5460 11676 5488 11716
rect 5810 11704 5816 11716
rect 5868 11704 5874 11756
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6196 11744 6224 11852
rect 6886 11852 7288 11880
rect 6362 11772 6368 11824
rect 6420 11812 6426 11824
rect 6730 11812 6736 11824
rect 6420 11784 6736 11812
rect 6420 11772 6426 11784
rect 6730 11772 6736 11784
rect 6788 11812 6794 11824
rect 6886 11812 6914 11852
rect 7282 11840 7288 11852
rect 7340 11840 7346 11892
rect 7650 11840 7656 11892
rect 7708 11880 7714 11892
rect 8021 11883 8079 11889
rect 8021 11880 8033 11883
rect 7708 11852 8033 11880
rect 7708 11840 7714 11852
rect 8021 11849 8033 11852
rect 8067 11849 8079 11883
rect 8846 11880 8852 11892
rect 8807 11852 8852 11880
rect 8021 11843 8079 11849
rect 8846 11840 8852 11852
rect 8904 11840 8910 11892
rect 10318 11880 10324 11892
rect 8956 11852 10180 11880
rect 10279 11852 10324 11880
rect 6788 11784 6914 11812
rect 6788 11772 6794 11784
rect 7098 11772 7104 11824
rect 7156 11812 7162 11824
rect 7156 11784 7788 11812
rect 7156 11772 7162 11784
rect 6638 11744 6644 11756
rect 6052 11716 6132 11744
rect 6196 11716 6644 11744
rect 6052 11704 6058 11716
rect 5123 11648 5488 11676
rect 5123 11645 5135 11648
rect 5077 11639 5135 11645
rect 5534 11636 5540 11688
rect 5592 11676 5598 11688
rect 5902 11676 5908 11688
rect 5592 11648 5908 11676
rect 5592 11636 5598 11648
rect 5902 11636 5908 11648
rect 5960 11636 5966 11688
rect 6104 11685 6132 11716
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 7190 11704 7196 11756
rect 7248 11744 7254 11756
rect 7760 11753 7788 11784
rect 8662 11772 8668 11824
rect 8720 11772 8726 11824
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 8956 11812 8984 11852
rect 8812 11784 8984 11812
rect 9309 11815 9367 11821
rect 8812 11772 8818 11784
rect 9309 11781 9321 11815
rect 9355 11812 9367 11815
rect 9953 11815 10011 11821
rect 9953 11812 9965 11815
rect 9355 11784 9965 11812
rect 9355 11781 9367 11784
rect 9309 11775 9367 11781
rect 9953 11781 9965 11784
rect 9999 11812 10011 11815
rect 10042 11812 10048 11824
rect 9999 11784 10048 11812
rect 9999 11781 10011 11784
rect 9953 11775 10011 11781
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10152 11812 10180 11852
rect 10318 11840 10324 11852
rect 10376 11840 10382 11892
rect 11333 11883 11391 11889
rect 11333 11849 11345 11883
rect 11379 11880 11391 11883
rect 11885 11883 11943 11889
rect 11885 11880 11897 11883
rect 11379 11852 11897 11880
rect 11379 11849 11391 11852
rect 11333 11843 11391 11849
rect 11885 11849 11897 11852
rect 11931 11849 11943 11883
rect 11885 11843 11943 11849
rect 12253 11883 12311 11889
rect 12253 11849 12265 11883
rect 12299 11880 12311 11883
rect 12342 11880 12348 11892
rect 12299 11852 12348 11880
rect 12299 11849 12311 11852
rect 12253 11843 12311 11849
rect 12342 11840 12348 11852
rect 12400 11840 12406 11892
rect 12437 11883 12495 11889
rect 12437 11849 12449 11883
rect 12483 11880 12495 11883
rect 12802 11880 12808 11892
rect 12483 11852 12808 11880
rect 12483 11849 12495 11852
rect 12437 11843 12495 11849
rect 10873 11815 10931 11821
rect 10873 11812 10885 11815
rect 10152 11784 10885 11812
rect 10873 11781 10885 11784
rect 10919 11812 10931 11815
rect 10919 11784 12204 11812
rect 10919 11781 10931 11784
rect 10873 11775 10931 11781
rect 7478 11747 7536 11753
rect 7478 11744 7490 11747
rect 7248 11716 7490 11744
rect 7248 11704 7254 11716
rect 7478 11713 7490 11716
rect 7524 11713 7536 11747
rect 7478 11707 7536 11713
rect 7745 11747 7803 11753
rect 7745 11713 7757 11747
rect 7791 11713 7803 11747
rect 7745 11707 7803 11713
rect 7929 11747 7987 11753
rect 7929 11713 7941 11747
rect 7975 11744 7987 11747
rect 8386 11744 8392 11756
rect 7975 11716 8392 11744
rect 7975 11713 7987 11716
rect 7929 11707 7987 11713
rect 8386 11704 8392 11716
rect 8444 11704 8450 11756
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11744 8539 11747
rect 8680 11744 8708 11772
rect 9030 11744 9036 11756
rect 8527 11716 9036 11744
rect 8527 11713 8539 11716
rect 8481 11707 8539 11713
rect 9030 11704 9036 11716
rect 9088 11704 9094 11756
rect 9217 11747 9275 11753
rect 9217 11713 9229 11747
rect 9263 11744 9275 11747
rect 9263 11716 9674 11744
rect 9263 11713 9275 11716
rect 9217 11707 9275 11713
rect 6089 11679 6147 11685
rect 6089 11645 6101 11679
rect 6135 11645 6147 11679
rect 6089 11639 6147 11645
rect 8665 11679 8723 11685
rect 8665 11645 8677 11679
rect 8711 11676 8723 11679
rect 9122 11676 9128 11688
rect 8711 11648 9128 11676
rect 8711 11645 8723 11648
rect 8665 11639 8723 11645
rect 9122 11636 9128 11648
rect 9180 11676 9186 11688
rect 9401 11679 9459 11685
rect 9401 11676 9413 11679
rect 9180 11648 9413 11676
rect 9180 11636 9186 11648
rect 9401 11645 9413 11648
rect 9447 11645 9459 11679
rect 9646 11676 9674 11716
rect 10410 11704 10416 11756
rect 10468 11744 10474 11756
rect 10505 11747 10563 11753
rect 10505 11744 10517 11747
rect 10468 11716 10517 11744
rect 10468 11704 10474 11716
rect 10505 11713 10517 11716
rect 10551 11713 10563 11747
rect 10965 11747 11023 11753
rect 10965 11744 10977 11747
rect 10505 11707 10563 11713
rect 10704 11716 10977 11744
rect 9769 11679 9827 11685
rect 9769 11676 9781 11679
rect 9646 11648 9781 11676
rect 9401 11639 9459 11645
rect 9769 11645 9781 11648
rect 9815 11676 9827 11679
rect 10226 11676 10232 11688
rect 9815 11648 10232 11676
rect 9815 11645 9827 11648
rect 9769 11639 9827 11645
rect 10226 11636 10232 11648
rect 10284 11676 10290 11688
rect 10704 11676 10732 11716
rect 10965 11713 10977 11716
rect 11011 11744 11023 11747
rect 11882 11744 11888 11756
rect 11011 11716 11376 11744
rect 11011 11713 11023 11716
rect 10965 11707 11023 11713
rect 10284 11648 10732 11676
rect 10781 11679 10839 11685
rect 10284 11636 10290 11648
rect 10781 11645 10793 11679
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 10796 11608 10824 11639
rect 11146 11608 11152 11620
rect 3896 11580 6877 11608
rect 4522 11540 4528 11552
rect 3252 11512 4528 11540
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 4706 11540 4712 11552
rect 4667 11512 4712 11540
rect 4706 11500 4712 11512
rect 4764 11500 4770 11552
rect 5074 11500 5080 11552
rect 5132 11540 5138 11552
rect 5169 11543 5227 11549
rect 5169 11540 5181 11543
rect 5132 11512 5181 11540
rect 5132 11500 5138 11512
rect 5169 11509 5181 11512
rect 5215 11509 5227 11543
rect 6362 11540 6368 11552
rect 6323 11512 6368 11540
rect 5169 11503 5227 11509
rect 6362 11500 6368 11512
rect 6420 11500 6426 11552
rect 6849 11540 6877 11580
rect 7760 11580 10732 11608
rect 10796 11580 11152 11608
rect 7760 11540 7788 11580
rect 10134 11540 10140 11552
rect 6849 11512 7788 11540
rect 10095 11512 10140 11540
rect 10134 11500 10140 11512
rect 10192 11500 10198 11552
rect 10704 11540 10732 11580
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 11348 11608 11376 11716
rect 11624 11716 11888 11744
rect 11624 11685 11652 11716
rect 11882 11704 11888 11716
rect 11940 11744 11946 11756
rect 12066 11744 12072 11756
rect 11940 11716 12072 11744
rect 11940 11704 11946 11716
rect 12066 11704 12072 11716
rect 12124 11704 12130 11756
rect 11609 11679 11667 11685
rect 11609 11645 11621 11679
rect 11655 11645 11667 11679
rect 11609 11639 11667 11645
rect 11698 11636 11704 11688
rect 11756 11676 11762 11688
rect 11793 11679 11851 11685
rect 11793 11676 11805 11679
rect 11756 11648 11805 11676
rect 11756 11636 11762 11648
rect 11793 11645 11805 11648
rect 11839 11645 11851 11679
rect 12176 11676 12204 11784
rect 12342 11704 12348 11756
rect 12400 11744 12406 11756
rect 12452 11744 12480 11843
rect 12802 11840 12808 11852
rect 12860 11840 12866 11892
rect 15194 11840 15200 11892
rect 15252 11880 15258 11892
rect 15289 11883 15347 11889
rect 15289 11880 15301 11883
rect 15252 11852 15301 11880
rect 15252 11840 15258 11852
rect 15289 11849 15301 11852
rect 15335 11849 15347 11883
rect 15289 11843 15347 11849
rect 15746 11840 15752 11892
rect 15804 11880 15810 11892
rect 18049 11883 18107 11889
rect 15804 11852 17724 11880
rect 15804 11840 15810 11852
rect 12621 11815 12679 11821
rect 12621 11781 12633 11815
rect 12667 11812 12679 11815
rect 15930 11812 15936 11824
rect 12667 11784 15936 11812
rect 12667 11781 12679 11784
rect 12621 11775 12679 11781
rect 12400 11716 12480 11744
rect 12400 11704 12406 11716
rect 12636 11676 12664 11775
rect 15930 11772 15936 11784
rect 15988 11772 15994 11824
rect 16298 11772 16304 11824
rect 16356 11812 16362 11824
rect 16393 11815 16451 11821
rect 16393 11812 16405 11815
rect 16356 11784 16405 11812
rect 16356 11772 16362 11784
rect 16393 11781 16405 11784
rect 16439 11781 16451 11815
rect 17586 11812 17592 11824
rect 16393 11775 16451 11781
rect 16684 11784 17592 11812
rect 16684 11756 16712 11784
rect 17586 11772 17592 11784
rect 17644 11772 17650 11824
rect 17696 11812 17724 11852
rect 18049 11849 18061 11883
rect 18095 11880 18107 11883
rect 18230 11880 18236 11892
rect 18095 11852 18236 11880
rect 18095 11849 18107 11852
rect 18049 11843 18107 11849
rect 18230 11840 18236 11852
rect 18288 11840 18294 11892
rect 18506 11840 18512 11892
rect 18564 11880 18570 11892
rect 18969 11883 19027 11889
rect 18969 11880 18981 11883
rect 18564 11852 18981 11880
rect 18564 11840 18570 11852
rect 18969 11849 18981 11852
rect 19015 11849 19027 11883
rect 19334 11880 19340 11892
rect 19295 11852 19340 11880
rect 18969 11843 19027 11849
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19797 11883 19855 11889
rect 19797 11880 19809 11883
rect 19576 11852 19809 11880
rect 19576 11840 19582 11852
rect 19797 11849 19809 11852
rect 19843 11849 19855 11883
rect 20346 11880 20352 11892
rect 20307 11852 20352 11880
rect 19797 11843 19855 11849
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 20622 11880 20628 11892
rect 20583 11852 20628 11880
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 21450 11812 21456 11824
rect 17696 11784 21456 11812
rect 21450 11772 21456 11784
rect 21508 11772 21514 11824
rect 12802 11704 12808 11756
rect 12860 11744 12866 11756
rect 13265 11747 13323 11753
rect 13265 11744 13277 11747
rect 12860 11716 13277 11744
rect 12860 11704 12866 11716
rect 13265 11713 13277 11716
rect 13311 11713 13323 11747
rect 13265 11707 13323 11713
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11744 13415 11747
rect 13538 11744 13544 11756
rect 13403 11716 13544 11744
rect 13403 11713 13415 11716
rect 13357 11707 13415 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 14918 11744 14924 11756
rect 14976 11753 14982 11756
rect 14976 11747 14999 11753
rect 14851 11716 14924 11744
rect 14918 11704 14924 11716
rect 14987 11744 14999 11747
rect 15102 11744 15108 11756
rect 14987 11716 15108 11744
rect 14987 11713 14999 11716
rect 14976 11707 14999 11713
rect 14976 11704 14982 11707
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15197 11747 15255 11753
rect 15197 11713 15209 11747
rect 15243 11744 15255 11747
rect 15378 11744 15384 11756
rect 15243 11716 15384 11744
rect 15243 11713 15255 11716
rect 15197 11707 15255 11713
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15654 11744 15660 11756
rect 15615 11716 15660 11744
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11744 15807 11747
rect 16482 11744 16488 11756
rect 15795 11716 16488 11744
rect 15795 11713 15807 11716
rect 15749 11707 15807 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 16936 11747 16994 11753
rect 16724 11716 16817 11744
rect 16724 11704 16730 11716
rect 16936 11713 16948 11747
rect 16982 11744 16994 11747
rect 17954 11744 17960 11756
rect 16982 11716 17960 11744
rect 16982 11713 16994 11716
rect 16936 11707 16994 11713
rect 17954 11704 17960 11716
rect 18012 11704 18018 11756
rect 18506 11744 18512 11756
rect 18467 11716 18512 11744
rect 18506 11704 18512 11716
rect 18564 11704 18570 11756
rect 19429 11747 19487 11753
rect 19429 11713 19441 11747
rect 19475 11744 19487 11747
rect 19794 11744 19800 11756
rect 19475 11716 19800 11744
rect 19475 11713 19487 11716
rect 19429 11707 19487 11713
rect 19794 11704 19800 11716
rect 19852 11704 19858 11756
rect 20165 11747 20223 11753
rect 20165 11713 20177 11747
rect 20211 11744 20223 11747
rect 20346 11744 20352 11756
rect 20211 11716 20352 11744
rect 20211 11713 20223 11716
rect 20165 11707 20223 11713
rect 20346 11704 20352 11716
rect 20404 11704 20410 11756
rect 20438 11704 20444 11756
rect 20496 11744 20502 11756
rect 21269 11747 21327 11753
rect 20496 11716 20541 11744
rect 20496 11704 20502 11716
rect 21269 11713 21281 11747
rect 21315 11744 21327 11747
rect 21928 11744 21956 12192
rect 21315 11716 21956 11744
rect 21315 11713 21327 11716
rect 21269 11707 21327 11713
rect 12176 11648 12664 11676
rect 13173 11679 13231 11685
rect 11793 11639 11851 11645
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 12342 11608 12348 11620
rect 11348 11580 12348 11608
rect 12342 11568 12348 11580
rect 12400 11568 12406 11620
rect 13188 11608 13216 11639
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 15838 11676 15844 11688
rect 13504 11648 13952 11676
rect 15799 11648 15844 11676
rect 13504 11636 13510 11648
rect 13630 11608 13636 11620
rect 12452 11580 13032 11608
rect 13188 11580 13636 11608
rect 12452 11540 12480 11580
rect 12802 11540 12808 11552
rect 10704 11512 12480 11540
rect 12763 11512 12808 11540
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13004 11540 13032 11580
rect 13630 11568 13636 11580
rect 13688 11608 13694 11620
rect 13817 11611 13875 11617
rect 13817 11608 13829 11611
rect 13688 11580 13829 11608
rect 13688 11568 13694 11580
rect 13817 11577 13829 11580
rect 13863 11577 13875 11611
rect 13817 11571 13875 11577
rect 13538 11540 13544 11552
rect 13004 11512 13544 11540
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 13722 11540 13728 11552
rect 13683 11512 13728 11540
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 13924 11540 13952 11648
rect 15838 11636 15844 11648
rect 15896 11636 15902 11688
rect 18230 11676 18236 11688
rect 18191 11648 18236 11676
rect 18230 11636 18236 11648
rect 18288 11636 18294 11688
rect 18414 11676 18420 11688
rect 18375 11648 18420 11676
rect 18414 11636 18420 11648
rect 18472 11636 18478 11688
rect 19150 11676 19156 11688
rect 18892 11648 19156 11676
rect 18892 11617 18920 11648
rect 19150 11636 19156 11648
rect 19208 11636 19214 11688
rect 19242 11636 19248 11688
rect 19300 11676 19306 11688
rect 19521 11679 19579 11685
rect 19521 11676 19533 11679
rect 19300 11648 19533 11676
rect 19300 11636 19306 11648
rect 19521 11645 19533 11648
rect 19567 11645 19579 11679
rect 21542 11676 21548 11688
rect 21503 11648 21548 11676
rect 19521 11639 19579 11645
rect 21542 11636 21548 11648
rect 21600 11636 21606 11688
rect 18877 11611 18935 11617
rect 18877 11577 18889 11611
rect 18923 11577 18935 11611
rect 20622 11608 20628 11620
rect 18877 11571 18935 11577
rect 19812 11580 20628 11608
rect 16209 11543 16267 11549
rect 16209 11540 16221 11543
rect 13924 11512 16221 11540
rect 16209 11509 16221 11512
rect 16255 11509 16267 11543
rect 16209 11503 16267 11509
rect 17402 11500 17408 11552
rect 17460 11540 17466 11552
rect 19812 11540 19840 11580
rect 20622 11568 20628 11580
rect 20680 11568 20686 11620
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 22738 11608 22744 11620
rect 20864 11580 22744 11608
rect 20864 11568 20870 11580
rect 22738 11568 22744 11580
rect 22796 11568 22802 11620
rect 17460 11512 19840 11540
rect 17460 11500 17466 11512
rect 19886 11500 19892 11552
rect 19944 11540 19950 11552
rect 19981 11543 20039 11549
rect 19981 11540 19993 11543
rect 19944 11512 19993 11540
rect 19944 11500 19950 11512
rect 19981 11509 19993 11512
rect 20027 11509 20039 11543
rect 19981 11503 20039 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2133 11339 2191 11345
rect 2133 11305 2145 11339
rect 2179 11336 2191 11339
rect 2866 11336 2872 11348
rect 2179 11308 2872 11336
rect 2179 11305 2191 11308
rect 2133 11299 2191 11305
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3605 11339 3663 11345
rect 3605 11305 3617 11339
rect 3651 11336 3663 11339
rect 3970 11336 3976 11348
rect 3651 11308 3976 11336
rect 3651 11305 3663 11308
rect 3605 11299 3663 11305
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 4120 11308 4169 11336
rect 4120 11296 4126 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 8573 11339 8631 11345
rect 8573 11336 8585 11339
rect 4157 11299 4215 11305
rect 5920 11308 8585 11336
rect 1762 11268 1768 11280
rect 1504 11240 1768 11268
rect 1504 11209 1532 11240
rect 1762 11228 1768 11240
rect 1820 11228 1826 11280
rect 5810 11268 5816 11280
rect 5771 11240 5816 11268
rect 5810 11228 5816 11240
rect 5868 11228 5874 11280
rect 1489 11203 1547 11209
rect 1489 11169 1501 11203
rect 1535 11169 1547 11203
rect 1670 11200 1676 11212
rect 1631 11172 1676 11200
rect 1489 11163 1547 11169
rect 1670 11160 1676 11172
rect 1728 11160 1734 11212
rect 2222 11200 2228 11212
rect 2183 11172 2228 11200
rect 2222 11160 2228 11172
rect 2280 11160 2286 11212
rect 4062 11160 4068 11212
rect 4120 11200 4126 11212
rect 4706 11200 4712 11212
rect 4120 11172 4712 11200
rect 4120 11160 4126 11172
rect 4706 11160 4712 11172
rect 4764 11160 4770 11212
rect 4801 11203 4859 11209
rect 4801 11169 4813 11203
rect 4847 11200 4859 11203
rect 4890 11200 4896 11212
rect 4847 11172 4896 11200
rect 4847 11169 4859 11172
rect 4801 11163 4859 11169
rect 4890 11160 4896 11172
rect 4948 11160 4954 11212
rect 5169 11203 5227 11209
rect 5169 11169 5181 11203
rect 5215 11169 5227 11203
rect 5169 11163 5227 11169
rect 3786 11132 3792 11144
rect 3747 11104 3792 11132
rect 3786 11092 3792 11104
rect 3844 11092 3850 11144
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11132 4675 11135
rect 4982 11132 4988 11144
rect 4663 11104 4988 11132
rect 4663 11101 4675 11104
rect 4617 11095 4675 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5184 11132 5212 11163
rect 5258 11160 5264 11212
rect 5316 11200 5322 11212
rect 5920 11200 5948 11308
rect 8573 11305 8585 11308
rect 8619 11305 8631 11339
rect 8573 11299 8631 11305
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9125 11339 9183 11345
rect 9125 11336 9137 11339
rect 8720 11308 9137 11336
rect 8720 11296 8726 11308
rect 9125 11305 9137 11308
rect 9171 11305 9183 11339
rect 9858 11336 9864 11348
rect 9771 11308 9864 11336
rect 9125 11299 9183 11305
rect 9858 11296 9864 11308
rect 9916 11336 9922 11348
rect 11238 11336 11244 11348
rect 9916 11308 11244 11336
rect 9916 11296 9922 11308
rect 11238 11296 11244 11308
rect 11296 11296 11302 11348
rect 11698 11336 11704 11348
rect 11659 11308 11704 11336
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12342 11296 12348 11348
rect 12400 11336 12406 11348
rect 12529 11339 12587 11345
rect 12529 11336 12541 11339
rect 12400 11308 12541 11336
rect 12400 11296 12406 11308
rect 12529 11305 12541 11308
rect 12575 11305 12587 11339
rect 12529 11299 12587 11305
rect 12802 11296 12808 11348
rect 12860 11336 12866 11348
rect 13170 11336 13176 11348
rect 12860 11308 13176 11336
rect 12860 11296 12866 11308
rect 13170 11296 13176 11308
rect 13228 11296 13234 11348
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 15010 11336 15016 11348
rect 13596 11308 15016 11336
rect 13596 11296 13602 11308
rect 15010 11296 15016 11308
rect 15068 11296 15074 11348
rect 15194 11296 15200 11348
rect 15252 11336 15258 11348
rect 15473 11339 15531 11345
rect 15473 11336 15485 11339
rect 15252 11308 15485 11336
rect 15252 11296 15258 11308
rect 15473 11305 15485 11308
rect 15519 11336 15531 11339
rect 16114 11336 16120 11348
rect 15519 11308 16120 11336
rect 15519 11305 15531 11308
rect 15473 11299 15531 11305
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 16666 11336 16672 11348
rect 16316 11308 16672 11336
rect 9950 11268 9956 11280
rect 9911 11240 9956 11268
rect 9950 11228 9956 11240
rect 10008 11228 10014 11280
rect 10594 11228 10600 11280
rect 10652 11268 10658 11280
rect 10778 11268 10784 11280
rect 10652 11240 10784 11268
rect 10652 11228 10658 11240
rect 10778 11228 10784 11240
rect 10836 11228 10842 11280
rect 10873 11271 10931 11277
rect 10873 11237 10885 11271
rect 10919 11268 10931 11271
rect 10919 11240 12112 11268
rect 10919 11237 10931 11240
rect 10873 11231 10931 11237
rect 5316 11172 5948 11200
rect 5316 11160 5322 11172
rect 5994 11160 6000 11212
rect 6052 11160 6058 11212
rect 6362 11200 6368 11212
rect 6323 11172 6368 11200
rect 6362 11160 6368 11172
rect 6420 11160 6426 11212
rect 7742 11160 7748 11212
rect 7800 11200 7806 11212
rect 10042 11200 10048 11212
rect 7800 11172 10048 11200
rect 7800 11160 7806 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 10321 11203 10379 11209
rect 10321 11169 10333 11203
rect 10367 11200 10379 11203
rect 11146 11200 11152 11212
rect 10367 11172 11152 11200
rect 10367 11169 10379 11172
rect 10321 11163 10379 11169
rect 11146 11160 11152 11172
rect 11204 11160 11210 11212
rect 11882 11200 11888 11212
rect 11843 11172 11888 11200
rect 11882 11160 11888 11172
rect 11940 11160 11946 11212
rect 12084 11209 12112 11240
rect 12250 11228 12256 11280
rect 12308 11268 12314 11280
rect 12621 11271 12679 11277
rect 12621 11268 12633 11271
rect 12308 11240 12633 11268
rect 12308 11228 12314 11240
rect 12621 11237 12633 11240
rect 12667 11237 12679 11271
rect 12621 11231 12679 11237
rect 12989 11271 13047 11277
rect 12989 11237 13001 11271
rect 13035 11268 13047 11271
rect 13354 11268 13360 11280
rect 13035 11240 13360 11268
rect 13035 11237 13047 11240
rect 12989 11231 13047 11237
rect 13354 11228 13360 11240
rect 13412 11228 13418 11280
rect 14093 11271 14151 11277
rect 14093 11268 14105 11271
rect 13464 11240 14105 11268
rect 13464 11209 13492 11240
rect 14093 11237 14105 11240
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 14366 11228 14372 11280
rect 14424 11268 14430 11280
rect 14734 11268 14740 11280
rect 14424 11240 14740 11268
rect 14424 11228 14430 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 15286 11228 15292 11280
rect 15344 11268 15350 11280
rect 15565 11271 15623 11277
rect 15565 11268 15577 11271
rect 15344 11240 15577 11268
rect 15344 11228 15350 11240
rect 15565 11237 15577 11240
rect 15611 11237 15623 11271
rect 15565 11231 15623 11237
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 16316 11268 16344 11308
rect 16666 11296 16672 11308
rect 16724 11296 16730 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18509 11339 18567 11345
rect 18509 11336 18521 11339
rect 18472 11308 18521 11336
rect 18472 11296 18478 11308
rect 18509 11305 18521 11308
rect 18555 11305 18567 11339
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 18509 11299 18567 11305
rect 19260 11308 19533 11336
rect 15896 11240 16344 11268
rect 15896 11228 15902 11240
rect 12069 11203 12127 11209
rect 12069 11169 12081 11203
rect 12115 11169 12127 11203
rect 13449 11203 13507 11209
rect 12069 11163 12127 11169
rect 12728 11172 13308 11200
rect 5810 11132 5816 11144
rect 5184 11104 5816 11132
rect 5810 11092 5816 11104
rect 5868 11092 5874 11144
rect 6012 11132 6040 11160
rect 6012 11104 6224 11132
rect 2492 11067 2550 11073
rect 2492 11033 2504 11067
rect 2538 11064 2550 11067
rect 3418 11064 3424 11076
rect 2538 11036 3424 11064
rect 2538 11033 2550 11036
rect 2492 11027 2550 11033
rect 3418 11024 3424 11036
rect 3476 11024 3482 11076
rect 4154 11024 4160 11076
rect 4212 11064 4218 11076
rect 4525 11067 4583 11073
rect 4525 11064 4537 11067
rect 4212 11036 4537 11064
rect 4212 11024 4218 11036
rect 4525 11033 4537 11036
rect 4571 11064 4583 11067
rect 5074 11064 5080 11076
rect 4571 11036 5080 11064
rect 4571 11033 4583 11036
rect 4525 11027 4583 11033
rect 5074 11024 5080 11036
rect 5132 11024 5138 11076
rect 5353 11067 5411 11073
rect 5353 11033 5365 11067
rect 5399 11064 5411 11067
rect 6196 11064 6224 11104
rect 6270 11092 6276 11144
rect 6328 11132 6334 11144
rect 6730 11132 6736 11144
rect 6328 11104 6373 11132
rect 6691 11104 6736 11132
rect 6328 11092 6334 11104
rect 6730 11092 6736 11104
rect 6788 11092 6794 11144
rect 8481 11135 8539 11141
rect 8481 11101 8493 11135
rect 8527 11132 8539 11135
rect 9214 11132 9220 11144
rect 8527 11104 9220 11132
rect 8527 11101 8539 11104
rect 8481 11095 8539 11101
rect 9214 11092 9220 11104
rect 9272 11132 9278 11144
rect 9401 11135 9459 11141
rect 9401 11132 9413 11135
rect 9272 11104 9413 11132
rect 9272 11092 9278 11104
rect 9401 11101 9413 11104
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 9677 11135 9735 11141
rect 9677 11101 9689 11135
rect 9723 11132 9735 11135
rect 10505 11135 10563 11141
rect 10505 11132 10517 11135
rect 9723 11104 10517 11132
rect 9723 11101 9735 11104
rect 9677 11095 9735 11101
rect 10505 11101 10517 11104
rect 10551 11132 10563 11135
rect 10962 11132 10968 11144
rect 10551 11104 10968 11132
rect 10551 11101 10563 11104
rect 10505 11095 10563 11101
rect 10962 11092 10968 11104
rect 11020 11092 11026 11144
rect 12728 11132 12756 11172
rect 11348 11104 12756 11132
rect 12805 11135 12863 11141
rect 6978 11067 7036 11073
rect 6978 11064 6990 11067
rect 5399 11036 5672 11064
rect 5399 11033 5411 11036
rect 5353 11027 5411 11033
rect 5644 11008 5672 11036
rect 5736 11036 6040 11064
rect 6196 11036 6990 11064
rect 1762 10956 1768 11008
rect 1820 10996 1826 11008
rect 1820 10968 1865 10996
rect 1820 10956 1826 10968
rect 2958 10956 2964 11008
rect 3016 10996 3022 11008
rect 3973 10999 4031 11005
rect 3973 10996 3985 10999
rect 3016 10968 3985 10996
rect 3016 10956 3022 10968
rect 3973 10965 3985 10968
rect 4019 10965 4031 10999
rect 5258 10996 5264 11008
rect 5219 10968 5264 10996
rect 3973 10959 4031 10965
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5626 10956 5632 11008
rect 5684 10956 5690 11008
rect 5736 11005 5764 11036
rect 5721 10999 5779 11005
rect 5721 10965 5733 10999
rect 5767 10965 5779 10999
rect 6012 10996 6040 11036
rect 6978 11033 6990 11036
rect 7024 11033 7036 11067
rect 6978 11027 7036 11033
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 8297 11067 8355 11073
rect 8297 11064 8309 11067
rect 7432 11036 8309 11064
rect 7432 11024 7438 11036
rect 8297 11033 8309 11036
rect 8343 11033 8355 11067
rect 8297 11027 8355 11033
rect 9033 11067 9091 11073
rect 9033 11033 9045 11067
rect 9079 11064 9091 11067
rect 9122 11064 9128 11076
rect 9079 11036 9128 11064
rect 9079 11033 9091 11036
rect 9033 11027 9091 11033
rect 9122 11024 9128 11036
rect 9180 11064 9186 11076
rect 9180 11036 9904 11064
rect 9180 11024 9186 11036
rect 6181 10999 6239 11005
rect 6181 10996 6193 10999
rect 6012 10968 6193 10996
rect 5721 10959 5779 10965
rect 6181 10965 6193 10968
rect 6227 10965 6239 10999
rect 8110 10996 8116 11008
rect 8071 10968 8116 10996
rect 6181 10959 6239 10965
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 8478 10956 8484 11008
rect 8536 10996 8542 11008
rect 9306 10996 9312 11008
rect 8536 10968 9312 10996
rect 8536 10956 8542 10968
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 9876 10996 9904 11036
rect 9950 11024 9956 11076
rect 10008 11064 10014 11076
rect 11348 11073 11376 11104
rect 12805 11101 12817 11135
rect 12851 11132 12863 11135
rect 12986 11132 12992 11144
rect 12851 11104 12992 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 12986 11092 12992 11104
rect 13044 11092 13050 11144
rect 11333 11067 11391 11073
rect 11333 11064 11345 11067
rect 10008 11036 11345 11064
rect 10008 11024 10014 11036
rect 11333 11033 11345 11036
rect 11379 11033 11391 11067
rect 11790 11064 11796 11076
rect 11333 11027 11391 11033
rect 11624 11036 11796 11064
rect 10413 10999 10471 11005
rect 10413 10996 10425 10999
rect 9876 10968 10425 10996
rect 10413 10965 10425 10968
rect 10459 10996 10471 10999
rect 10594 10996 10600 11008
rect 10459 10968 10600 10996
rect 10459 10965 10471 10968
rect 10413 10959 10471 10965
rect 10594 10956 10600 10968
rect 10652 10956 10658 11008
rect 11238 10996 11244 11008
rect 11151 10968 11244 10996
rect 11238 10956 11244 10968
rect 11296 10996 11302 11008
rect 11624 10996 11652 11036
rect 11790 11024 11796 11036
rect 11848 11024 11854 11076
rect 11882 11024 11888 11076
rect 11940 11064 11946 11076
rect 12161 11067 12219 11073
rect 12161 11064 12173 11067
rect 11940 11036 12173 11064
rect 11940 11024 11946 11036
rect 12161 11033 12173 11036
rect 12207 11064 12219 11067
rect 12618 11064 12624 11076
rect 12207 11036 12624 11064
rect 12207 11033 12219 11036
rect 12161 11027 12219 11033
rect 12618 11024 12624 11036
rect 12676 11024 12682 11076
rect 11296 10968 11652 10996
rect 13004 10996 13032 11092
rect 13280 11064 13308 11172
rect 13449 11169 13461 11203
rect 13495 11169 13507 11203
rect 13449 11163 13507 11169
rect 13538 11160 13544 11212
rect 13596 11200 13602 11212
rect 13814 11200 13820 11212
rect 13596 11172 13641 11200
rect 13775 11172 13820 11200
rect 13596 11160 13602 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 13906 11160 13912 11212
rect 13964 11200 13970 11212
rect 14645 11203 14703 11209
rect 14645 11200 14657 11203
rect 13964 11172 14657 11200
rect 13964 11160 13970 11172
rect 14645 11169 14657 11172
rect 14691 11169 14703 11203
rect 14645 11163 14703 11169
rect 14918 11160 14924 11212
rect 14976 11200 14982 11212
rect 15746 11200 15752 11212
rect 14976 11172 15752 11200
rect 14976 11160 14982 11172
rect 15746 11160 15752 11172
rect 15804 11160 15810 11212
rect 16316 11209 16344 11240
rect 17681 11271 17739 11277
rect 17681 11237 17693 11271
rect 17727 11237 17739 11271
rect 17681 11231 17739 11237
rect 16301 11203 16359 11209
rect 16301 11169 16313 11203
rect 16347 11169 16359 11203
rect 17696 11200 17724 11231
rect 17954 11200 17960 11212
rect 17696 11172 17960 11200
rect 16301 11163 16359 11169
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 19260 11200 19288 11308
rect 19521 11305 19533 11308
rect 19567 11336 19579 11339
rect 20162 11336 20168 11348
rect 19567 11308 20168 11336
rect 19567 11305 19579 11308
rect 19521 11299 19579 11305
rect 20162 11296 20168 11308
rect 20220 11296 20226 11348
rect 20346 11336 20352 11348
rect 20307 11308 20352 11336
rect 20346 11296 20352 11308
rect 20404 11296 20410 11348
rect 20622 11296 20628 11348
rect 20680 11336 20686 11348
rect 20993 11339 21051 11345
rect 20993 11336 21005 11339
rect 20680 11308 21005 11336
rect 20680 11296 20686 11308
rect 20993 11305 21005 11308
rect 21039 11305 21051 11339
rect 20993 11299 21051 11305
rect 21361 11339 21419 11345
rect 21361 11305 21373 11339
rect 21407 11336 21419 11339
rect 21450 11336 21456 11348
rect 21407 11308 21456 11336
rect 21407 11305 21419 11308
rect 21361 11299 21419 11305
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 19337 11271 19395 11277
rect 19337 11237 19349 11271
rect 19383 11268 19395 11271
rect 19702 11268 19708 11280
rect 19383 11240 19708 11268
rect 19383 11237 19395 11240
rect 19337 11231 19395 11237
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 20254 11268 20260 11280
rect 20215 11240 20260 11268
rect 20254 11228 20260 11240
rect 20312 11228 20318 11280
rect 20806 11268 20812 11280
rect 20767 11240 20812 11268
rect 20806 11228 20812 11240
rect 20864 11228 20870 11280
rect 19518 11200 19524 11212
rect 19260 11172 19524 11200
rect 19518 11160 19524 11172
rect 19576 11160 19582 11212
rect 20162 11160 20168 11212
rect 20220 11200 20226 11212
rect 20220 11172 20576 11200
rect 20220 11160 20226 11172
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11132 13415 11135
rect 13722 11132 13728 11144
rect 13403 11104 13728 11132
rect 13403 11101 13415 11104
rect 13357 11095 13415 11101
rect 13722 11092 13728 11104
rect 13780 11092 13786 11144
rect 13832 11132 13860 11160
rect 14553 11135 14611 11141
rect 14553 11132 14565 11135
rect 13832 11104 14565 11132
rect 14553 11101 14565 11104
rect 14599 11101 14611 11135
rect 15194 11132 15200 11144
rect 15155 11104 15200 11132
rect 14553 11095 14611 11101
rect 15194 11092 15200 11104
rect 15252 11132 15258 11144
rect 16114 11132 16120 11144
rect 15252 11128 15792 11132
rect 15856 11128 16120 11132
rect 15252 11104 16120 11128
rect 15252 11092 15258 11104
rect 15764 11100 15884 11104
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17770 11132 17776 11144
rect 17552 11104 17776 11132
rect 17552 11092 17558 11104
rect 17770 11092 17776 11104
rect 17828 11132 17834 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 17828 11104 18613 11132
rect 17828 11092 17834 11104
rect 18601 11101 18613 11104
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 20548 11141 20576 11172
rect 19705 11135 19763 11141
rect 19705 11132 19717 11135
rect 19392 11104 19717 11132
rect 19392 11092 19398 11104
rect 19705 11101 19717 11104
rect 19751 11101 19763 11135
rect 19705 11095 19763 11101
rect 20073 11135 20131 11141
rect 20073 11101 20085 11135
rect 20119 11132 20131 11135
rect 20533 11135 20591 11141
rect 20119 11104 20484 11132
rect 20119 11101 20131 11104
rect 20073 11095 20131 11101
rect 14461 11067 14519 11073
rect 13280 11036 14412 11064
rect 13906 10996 13912 11008
rect 13004 10968 13912 10996
rect 11296 10956 11302 10968
rect 13906 10956 13912 10968
rect 13964 10956 13970 11008
rect 14384 10996 14412 11036
rect 14461 11033 14473 11067
rect 14507 11064 14519 11067
rect 15010 11064 15016 11076
rect 14507 11036 15016 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 15010 11024 15016 11036
rect 15068 11024 15074 11076
rect 16390 11064 16396 11076
rect 15212 11036 16396 11064
rect 15212 10996 15240 11036
rect 16390 11024 16396 11036
rect 16448 11024 16454 11076
rect 16568 11067 16626 11073
rect 16568 11033 16580 11067
rect 16614 11064 16626 11067
rect 16942 11064 16948 11076
rect 16614 11036 16948 11064
rect 16614 11033 16626 11036
rect 16568 11027 16626 11033
rect 16942 11024 16948 11036
rect 17000 11024 17006 11076
rect 17310 11024 17316 11076
rect 17368 11064 17374 11076
rect 18141 11067 18199 11073
rect 18141 11064 18153 11067
rect 17368 11036 18153 11064
rect 17368 11024 17374 11036
rect 18141 11033 18153 11036
rect 18187 11033 18199 11067
rect 18141 11027 18199 11033
rect 19061 11067 19119 11073
rect 19061 11033 19073 11067
rect 19107 11064 19119 11067
rect 20346 11064 20352 11076
rect 19107 11036 20352 11064
rect 19107 11033 19119 11036
rect 19061 11027 19119 11033
rect 20346 11024 20352 11036
rect 20404 11024 20410 11076
rect 20456 11064 20484 11104
rect 20533 11101 20545 11135
rect 20579 11101 20591 11135
rect 20533 11095 20591 11101
rect 20625 11135 20683 11141
rect 20625 11101 20637 11135
rect 20671 11132 20683 11135
rect 20898 11132 20904 11144
rect 20671 11104 20904 11132
rect 20671 11101 20683 11104
rect 20625 11095 20683 11101
rect 20898 11092 20904 11104
rect 20956 11092 20962 11144
rect 21450 11132 21456 11144
rect 21411 11104 21456 11132
rect 21450 11092 21456 11104
rect 21508 11092 21514 11144
rect 21082 11064 21088 11076
rect 20456 11036 20852 11064
rect 21043 11036 21088 11064
rect 20824 11008 20852 11036
rect 21082 11024 21088 11036
rect 21140 11024 21146 11076
rect 14384 10968 15240 10996
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 15654 10996 15660 11008
rect 15344 10968 15660 10996
rect 15344 10956 15350 10968
rect 15654 10956 15660 10968
rect 15712 10956 15718 11008
rect 15746 10956 15752 11008
rect 15804 10996 15810 11008
rect 15804 10968 15849 10996
rect 15804 10956 15810 10968
rect 15930 10956 15936 11008
rect 15988 10996 15994 11008
rect 18046 10996 18052 11008
rect 15988 10968 16033 10996
rect 18007 10968 18052 10996
rect 15988 10956 15994 10968
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 18782 10996 18788 11008
rect 18743 10968 18788 10996
rect 18782 10956 18788 10968
rect 18840 10956 18846 11008
rect 19610 10956 19616 11008
rect 19668 10996 19674 11008
rect 19889 10999 19947 11005
rect 19889 10996 19901 10999
rect 19668 10968 19901 10996
rect 19668 10956 19674 10968
rect 19889 10965 19901 10968
rect 19935 10996 19947 10999
rect 20622 10996 20628 11008
rect 19935 10968 20628 10996
rect 19935 10965 19947 10968
rect 19889 10959 19947 10965
rect 20622 10956 20628 10968
rect 20680 10956 20686 11008
rect 20806 10956 20812 11008
rect 20864 10956 20870 11008
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 382 10752 388 10804
rect 440 10792 446 10804
rect 3142 10792 3148 10804
rect 440 10764 3148 10792
rect 440 10752 446 10764
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 3789 10795 3847 10801
rect 3789 10761 3801 10795
rect 3835 10792 3847 10795
rect 4062 10792 4068 10804
rect 3835 10764 4068 10792
rect 3835 10761 3847 10764
rect 3789 10755 3847 10761
rect 4062 10752 4068 10764
rect 4120 10752 4126 10804
rect 4157 10795 4215 10801
rect 4157 10761 4169 10795
rect 4203 10792 4215 10795
rect 5445 10795 5503 10801
rect 5445 10792 5457 10795
rect 4203 10764 5457 10792
rect 4203 10761 4215 10764
rect 4157 10755 4215 10761
rect 5445 10761 5457 10764
rect 5491 10761 5503 10795
rect 5445 10755 5503 10761
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 5997 10795 6055 10801
rect 5997 10792 6009 10795
rect 5684 10764 6009 10792
rect 5684 10752 5690 10764
rect 5997 10761 6009 10764
rect 6043 10761 6055 10795
rect 5997 10755 6055 10761
rect 6095 10764 6684 10792
rect 1486 10724 1492 10736
rect 1447 10696 1492 10724
rect 1486 10684 1492 10696
rect 1544 10684 1550 10736
rect 2222 10724 2228 10736
rect 1780 10696 2228 10724
rect 1780 10665 1808 10696
rect 2222 10684 2228 10696
rect 2280 10684 2286 10736
rect 2682 10684 2688 10736
rect 2740 10724 2746 10736
rect 3237 10727 3295 10733
rect 3237 10724 3249 10727
rect 2740 10696 3249 10724
rect 2740 10684 2746 10696
rect 3237 10693 3249 10696
rect 3283 10724 3295 10727
rect 3697 10727 3755 10733
rect 3697 10724 3709 10727
rect 3283 10696 3709 10724
rect 3283 10693 3295 10696
rect 3237 10687 3295 10693
rect 3697 10693 3709 10696
rect 3743 10693 3755 10727
rect 3697 10687 3755 10693
rect 3970 10684 3976 10736
rect 4028 10724 4034 10736
rect 4028 10696 4752 10724
rect 4028 10684 4034 10696
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10625 1823 10659
rect 1765 10619 1823 10625
rect 1854 10616 1860 10668
rect 1912 10656 1918 10668
rect 2032 10659 2090 10665
rect 2032 10656 2044 10659
rect 1912 10628 2044 10656
rect 1912 10616 1918 10628
rect 2032 10625 2044 10628
rect 2078 10656 2090 10659
rect 2078 10628 3740 10656
rect 2078 10625 2090 10628
rect 2032 10619 2090 10625
rect 3605 10591 3663 10597
rect 3605 10557 3617 10591
rect 3651 10557 3663 10591
rect 3712 10588 3740 10628
rect 3988 10588 4016 10684
rect 4338 10616 4344 10668
rect 4396 10656 4402 10668
rect 4617 10659 4675 10665
rect 4617 10656 4629 10659
rect 4396 10628 4629 10656
rect 4396 10616 4402 10628
rect 4617 10625 4629 10628
rect 4663 10625 4675 10659
rect 4724 10656 4752 10696
rect 4982 10684 4988 10736
rect 5040 10724 5046 10736
rect 5040 10696 5764 10724
rect 5040 10684 5046 10696
rect 5736 10656 5764 10696
rect 5810 10684 5816 10736
rect 5868 10724 5874 10736
rect 6095 10724 6123 10764
rect 5868 10696 6123 10724
rect 6656 10724 6684 10764
rect 7282 10752 7288 10804
rect 7340 10792 7346 10804
rect 7377 10795 7435 10801
rect 7377 10792 7389 10795
rect 7340 10764 7389 10792
rect 7340 10752 7346 10764
rect 7377 10761 7389 10764
rect 7423 10761 7435 10795
rect 7377 10755 7435 10761
rect 7653 10795 7711 10801
rect 7653 10761 7665 10795
rect 7699 10792 7711 10795
rect 7742 10792 7748 10804
rect 7699 10764 7748 10792
rect 7699 10761 7711 10764
rect 7653 10755 7711 10761
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 8018 10752 8024 10804
rect 8076 10792 8082 10804
rect 8205 10795 8263 10801
rect 8205 10792 8217 10795
rect 8076 10764 8217 10792
rect 8076 10752 8082 10764
rect 8205 10761 8217 10764
rect 8251 10761 8263 10795
rect 8205 10755 8263 10761
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 8941 10795 8999 10801
rect 8941 10792 8953 10795
rect 8343 10764 8953 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 8941 10761 8953 10764
rect 8987 10792 8999 10795
rect 10226 10792 10232 10804
rect 8987 10764 10232 10792
rect 8987 10761 8999 10764
rect 8941 10755 8999 10761
rect 7190 10724 7196 10736
rect 6656 10696 7196 10724
rect 5868 10684 5874 10696
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 4724 10628 5672 10656
rect 5736 10628 6745 10656
rect 4617 10619 4675 10625
rect 4706 10588 4712 10600
rect 3712 10560 4016 10588
rect 4667 10560 4712 10588
rect 3605 10551 3663 10557
rect 1581 10455 1639 10461
rect 1581 10421 1593 10455
rect 1627 10452 1639 10455
rect 1946 10452 1952 10464
rect 1627 10424 1952 10452
rect 1627 10421 1639 10424
rect 1581 10415 1639 10421
rect 1946 10412 1952 10424
rect 2004 10412 2010 10464
rect 2498 10412 2504 10464
rect 2556 10452 2562 10464
rect 3145 10455 3203 10461
rect 3145 10452 3157 10455
rect 2556 10424 3157 10452
rect 2556 10412 2562 10424
rect 3145 10421 3157 10424
rect 3191 10452 3203 10455
rect 3326 10452 3332 10464
rect 3191 10424 3332 10452
rect 3191 10421 3203 10424
rect 3145 10415 3203 10421
rect 3326 10412 3332 10424
rect 3384 10412 3390 10464
rect 3620 10452 3648 10551
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 4890 10588 4896 10600
rect 4851 10560 4896 10588
rect 4890 10548 4896 10560
rect 4948 10548 4954 10600
rect 5166 10548 5172 10600
rect 5224 10588 5230 10600
rect 5644 10597 5672 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 6932 10597 6960 10696
rect 7190 10684 7196 10696
rect 7248 10684 7254 10736
rect 8220 10656 8248 10755
rect 10226 10752 10232 10764
rect 10284 10792 10290 10804
rect 10284 10764 11100 10792
rect 10284 10752 10290 10764
rect 8570 10684 8576 10736
rect 8628 10724 8634 10736
rect 9769 10727 9827 10733
rect 9769 10724 9781 10727
rect 8628 10696 9781 10724
rect 8628 10684 8634 10696
rect 9769 10693 9781 10696
rect 9815 10693 9827 10727
rect 10318 10724 10324 10736
rect 9769 10687 9827 10693
rect 9968 10696 10324 10724
rect 9968 10665 9996 10696
rect 10318 10684 10324 10696
rect 10376 10684 10382 10736
rect 11072 10724 11100 10764
rect 11146 10752 11152 10804
rect 11204 10792 11210 10804
rect 11333 10795 11391 10801
rect 11333 10792 11345 10795
rect 11204 10764 11345 10792
rect 11204 10752 11210 10764
rect 11333 10761 11345 10764
rect 11379 10761 11391 10795
rect 11333 10755 11391 10761
rect 11701 10795 11759 10801
rect 11701 10761 11713 10795
rect 11747 10792 11759 10795
rect 11882 10792 11888 10804
rect 11747 10764 11888 10792
rect 11747 10761 11759 10764
rect 11701 10755 11759 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 12345 10795 12403 10801
rect 12345 10792 12357 10795
rect 12124 10764 12357 10792
rect 12124 10752 12130 10764
rect 12345 10761 12357 10764
rect 12391 10761 12403 10795
rect 12345 10755 12403 10761
rect 12529 10795 12587 10801
rect 12529 10761 12541 10795
rect 12575 10792 12587 10795
rect 14461 10795 14519 10801
rect 12575 10764 13308 10792
rect 12575 10761 12587 10764
rect 12529 10755 12587 10761
rect 12986 10724 12992 10736
rect 11072 10696 12992 10724
rect 12986 10684 12992 10696
rect 13044 10684 13050 10736
rect 13280 10724 13308 10764
rect 14461 10761 14473 10795
rect 14507 10792 14519 10795
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 14507 10764 14841 10792
rect 14507 10761 14519 10764
rect 14461 10755 14519 10761
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 15197 10795 15255 10801
rect 15197 10761 15209 10795
rect 15243 10792 15255 10795
rect 15657 10795 15715 10801
rect 15657 10792 15669 10795
rect 15243 10764 15669 10792
rect 15243 10761 15255 10764
rect 15197 10755 15255 10761
rect 15657 10761 15669 10764
rect 15703 10761 15715 10795
rect 15657 10755 15715 10761
rect 15930 10752 15936 10804
rect 15988 10792 15994 10804
rect 16025 10795 16083 10801
rect 16025 10792 16037 10795
rect 15988 10764 16037 10792
rect 15988 10752 15994 10764
rect 16025 10761 16037 10764
rect 16071 10761 16083 10795
rect 16025 10755 16083 10761
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 17037 10795 17095 10801
rect 17037 10792 17049 10795
rect 16172 10764 17049 10792
rect 16172 10752 16178 10764
rect 17037 10761 17049 10764
rect 17083 10761 17095 10795
rect 17037 10755 17095 10761
rect 17405 10795 17463 10801
rect 17405 10761 17417 10795
rect 17451 10792 17463 10795
rect 17773 10795 17831 10801
rect 17773 10792 17785 10795
rect 17451 10764 17785 10792
rect 17451 10761 17463 10764
rect 17405 10755 17463 10761
rect 17773 10761 17785 10764
rect 17819 10761 17831 10795
rect 17773 10755 17831 10761
rect 18046 10752 18052 10804
rect 18104 10792 18110 10804
rect 18233 10795 18291 10801
rect 18233 10792 18245 10795
rect 18104 10764 18245 10792
rect 18104 10752 18110 10764
rect 18233 10761 18245 10764
rect 18279 10761 18291 10795
rect 18233 10755 18291 10761
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10792 18383 10795
rect 18506 10792 18512 10804
rect 18371 10764 18512 10792
rect 18371 10761 18383 10764
rect 18325 10755 18383 10761
rect 18506 10752 18512 10764
rect 18564 10752 18570 10804
rect 18785 10795 18843 10801
rect 18785 10761 18797 10795
rect 18831 10792 18843 10795
rect 19153 10795 19211 10801
rect 19153 10792 19165 10795
rect 18831 10764 19165 10792
rect 18831 10761 18843 10764
rect 18785 10755 18843 10761
rect 19153 10761 19165 10764
rect 19199 10761 19211 10795
rect 19518 10792 19524 10804
rect 19479 10764 19524 10792
rect 19153 10755 19211 10761
rect 19518 10752 19524 10764
rect 19576 10752 19582 10804
rect 19981 10795 20039 10801
rect 19981 10761 19993 10795
rect 20027 10761 20039 10795
rect 20346 10792 20352 10804
rect 20307 10764 20352 10792
rect 19981 10755 20039 10761
rect 13538 10724 13544 10736
rect 13280 10696 13544 10724
rect 13538 10684 13544 10696
rect 13596 10684 13602 10736
rect 13722 10733 13728 10736
rect 13664 10727 13728 10733
rect 13664 10693 13676 10727
rect 13710 10693 13728 10727
rect 13664 10687 13728 10693
rect 13722 10684 13728 10687
rect 13780 10684 13786 10736
rect 15286 10684 15292 10736
rect 15344 10724 15350 10736
rect 15562 10724 15568 10736
rect 15344 10696 15568 10724
rect 15344 10684 15350 10696
rect 15562 10684 15568 10696
rect 15620 10684 15626 10736
rect 15746 10684 15752 10736
rect 15804 10724 15810 10736
rect 16945 10727 17003 10733
rect 16945 10724 16957 10727
rect 15804 10696 16957 10724
rect 15804 10684 15810 10696
rect 16945 10693 16957 10696
rect 16991 10693 17003 10727
rect 16945 10687 17003 10693
rect 18693 10727 18751 10733
rect 18693 10693 18705 10727
rect 18739 10724 18751 10727
rect 19996 10724 20024 10755
rect 20346 10752 20352 10764
rect 20404 10752 20410 10804
rect 20441 10795 20499 10801
rect 20441 10761 20453 10795
rect 20487 10792 20499 10795
rect 20622 10792 20628 10804
rect 20487 10764 20628 10792
rect 20487 10761 20499 10764
rect 20441 10755 20499 10761
rect 20622 10752 20628 10764
rect 20680 10752 20686 10804
rect 18739 10696 20024 10724
rect 18739 10693 18751 10696
rect 18693 10687 18751 10693
rect 8665 10659 8723 10665
rect 8665 10656 8677 10659
rect 8220 10628 8677 10656
rect 8665 10625 8677 10628
rect 8711 10625 8723 10659
rect 8665 10619 8723 10625
rect 9401 10659 9459 10665
rect 9401 10625 9413 10659
rect 9447 10625 9459 10659
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9401 10619 9459 10625
rect 9646 10628 9965 10656
rect 5537 10591 5595 10597
rect 5537 10588 5549 10591
rect 5224 10560 5549 10588
rect 5224 10548 5230 10560
rect 5537 10557 5549 10560
rect 5583 10557 5595 10591
rect 5537 10551 5595 10557
rect 5629 10591 5687 10597
rect 5629 10557 5641 10591
rect 5675 10557 5687 10591
rect 5629 10551 5687 10557
rect 6825 10591 6883 10597
rect 6825 10557 6837 10591
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10557 6975 10591
rect 6917 10551 6975 10557
rect 4246 10520 4252 10532
rect 4207 10492 4252 10520
rect 4246 10480 4252 10492
rect 4304 10480 4310 10532
rect 4522 10480 4528 10532
rect 4580 10520 4586 10532
rect 5077 10523 5135 10529
rect 5077 10520 5089 10523
rect 4580 10492 5089 10520
rect 4580 10480 4586 10492
rect 5077 10489 5089 10492
rect 5123 10489 5135 10523
rect 5077 10483 5135 10489
rect 5994 10480 6000 10532
rect 6052 10520 6058 10532
rect 6365 10523 6423 10529
rect 6365 10520 6377 10523
rect 6052 10492 6377 10520
rect 6052 10480 6058 10492
rect 6365 10489 6377 10492
rect 6411 10489 6423 10523
rect 6840 10520 6868 10551
rect 7190 10548 7196 10600
rect 7248 10588 7254 10600
rect 7834 10588 7840 10600
rect 7248 10560 7840 10588
rect 7248 10548 7254 10560
rect 7834 10548 7840 10560
rect 7892 10548 7898 10600
rect 8110 10548 8116 10600
rect 8168 10588 8174 10600
rect 8389 10591 8447 10597
rect 8389 10588 8401 10591
rect 8168 10560 8401 10588
rect 8168 10548 8174 10560
rect 8389 10557 8401 10560
rect 8435 10557 8447 10591
rect 8389 10551 8447 10557
rect 7285 10523 7343 10529
rect 7285 10520 7297 10523
rect 6840 10492 7297 10520
rect 6365 10483 6423 10489
rect 7285 10489 7297 10492
rect 7331 10520 7343 10523
rect 7466 10520 7472 10532
rect 7331 10492 7472 10520
rect 7331 10489 7343 10492
rect 7285 10483 7343 10489
rect 7466 10480 7472 10492
rect 7524 10520 7530 10532
rect 8018 10520 8024 10532
rect 7524 10492 8024 10520
rect 7524 10480 7530 10492
rect 8018 10480 8024 10492
rect 8076 10480 8082 10532
rect 8680 10520 8708 10619
rect 9125 10591 9183 10597
rect 9125 10557 9137 10591
rect 9171 10588 9183 10591
rect 9214 10588 9220 10600
rect 9171 10560 9220 10588
rect 9171 10557 9183 10560
rect 9125 10551 9183 10557
rect 9214 10548 9220 10560
rect 9272 10548 9278 10600
rect 9416 10588 9444 10619
rect 9646 10600 9674 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10220 10659 10278 10665
rect 10220 10625 10232 10659
rect 10266 10656 10278 10659
rect 10502 10656 10508 10668
rect 10266 10628 10508 10656
rect 10266 10625 10278 10628
rect 10220 10619 10278 10625
rect 10502 10616 10508 10628
rect 10560 10616 10566 10668
rect 10594 10616 10600 10668
rect 10652 10656 10658 10668
rect 11885 10659 11943 10665
rect 11885 10656 11897 10659
rect 10652 10628 11897 10656
rect 10652 10616 10658 10628
rect 11885 10625 11897 10628
rect 11931 10656 11943 10659
rect 12526 10656 12532 10668
rect 11931 10628 12532 10656
rect 11931 10625 11943 10628
rect 11885 10619 11943 10625
rect 12526 10616 12532 10628
rect 12584 10616 12590 10668
rect 13262 10656 13268 10668
rect 12912 10628 13268 10656
rect 9646 10588 9680 10600
rect 9416 10560 9680 10588
rect 9674 10548 9680 10560
rect 9732 10548 9738 10600
rect 10962 10548 10968 10600
rect 11020 10588 11026 10600
rect 12802 10588 12808 10600
rect 11020 10560 12808 10588
rect 11020 10548 11026 10560
rect 12802 10548 12808 10560
rect 12860 10548 12866 10600
rect 9858 10520 9864 10532
rect 8680 10492 9864 10520
rect 9858 10480 9864 10492
rect 9916 10480 9922 10532
rect 11882 10480 11888 10532
rect 11940 10520 11946 10532
rect 12912 10520 12940 10628
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 14366 10616 14372 10668
rect 14424 10656 14430 10668
rect 17862 10656 17868 10668
rect 14424 10628 14469 10656
rect 17823 10628 17868 10656
rect 14424 10616 14430 10628
rect 17862 10616 17868 10628
rect 17920 10616 17926 10668
rect 19720 10628 20576 10656
rect 19720 10600 19748 10628
rect 13906 10588 13912 10600
rect 13867 10560 13912 10588
rect 13906 10548 13912 10560
rect 13964 10548 13970 10600
rect 13998 10548 14004 10600
rect 14056 10588 14062 10600
rect 14553 10591 14611 10597
rect 14553 10588 14565 10591
rect 14056 10560 14565 10588
rect 14056 10548 14062 10560
rect 14553 10557 14565 10560
rect 14599 10557 14611 10591
rect 14553 10551 14611 10557
rect 14918 10548 14924 10600
rect 14976 10588 14982 10600
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14976 10560 15301 10588
rect 14976 10548 14982 10560
rect 15289 10557 15301 10560
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 15378 10548 15384 10600
rect 15436 10588 15442 10600
rect 16117 10591 16175 10597
rect 16117 10588 16129 10591
rect 15436 10560 15481 10588
rect 16040 10560 16129 10588
rect 15436 10548 15442 10560
rect 16040 10532 16068 10560
rect 16117 10557 16129 10560
rect 16163 10557 16175 10591
rect 16117 10551 16175 10557
rect 16209 10591 16267 10597
rect 16209 10557 16221 10591
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 16853 10591 16911 10597
rect 16853 10557 16865 10591
rect 16899 10557 16911 10591
rect 16853 10551 16911 10557
rect 11940 10492 12940 10520
rect 11940 10480 11946 10492
rect 16022 10480 16028 10532
rect 16080 10480 16086 10532
rect 4890 10452 4896 10464
rect 3620 10424 4896 10452
rect 4890 10412 4896 10424
rect 4948 10412 4954 10464
rect 5258 10412 5264 10464
rect 5316 10452 5322 10464
rect 5626 10452 5632 10464
rect 5316 10424 5632 10452
rect 5316 10412 5322 10424
rect 5626 10412 5632 10424
rect 5684 10412 5690 10464
rect 7834 10452 7840 10464
rect 7795 10424 7840 10452
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 9122 10412 9128 10464
rect 9180 10452 9186 10464
rect 9217 10455 9275 10461
rect 9217 10452 9229 10455
rect 9180 10424 9229 10452
rect 9180 10412 9186 10424
rect 9217 10421 9229 10424
rect 9263 10421 9275 10455
rect 9217 10415 9275 10421
rect 9677 10455 9735 10461
rect 9677 10421 9689 10455
rect 9723 10452 9735 10455
rect 10318 10452 10324 10464
rect 9723 10424 10324 10452
rect 9723 10421 9735 10424
rect 9677 10415 9735 10421
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 12066 10452 12072 10464
rect 12027 10424 12072 10452
rect 12066 10412 12072 10424
rect 12124 10412 12130 10464
rect 12158 10412 12164 10464
rect 12216 10452 12222 10464
rect 12216 10424 12261 10452
rect 12216 10412 12222 10424
rect 13262 10412 13268 10464
rect 13320 10452 13326 10464
rect 14001 10455 14059 10461
rect 14001 10452 14013 10455
rect 13320 10424 14013 10452
rect 13320 10412 13326 10424
rect 14001 10421 14013 10424
rect 14047 10421 14059 10455
rect 14001 10415 14059 10421
rect 15102 10412 15108 10464
rect 15160 10452 15166 10464
rect 16224 10452 16252 10551
rect 16868 10520 16896 10551
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17589 10591 17647 10597
rect 17589 10588 17601 10591
rect 17000 10560 17601 10588
rect 17000 10548 17006 10560
rect 17589 10557 17601 10560
rect 17635 10557 17647 10591
rect 17589 10551 17647 10557
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18877 10591 18935 10597
rect 18877 10588 18889 10591
rect 18012 10560 18889 10588
rect 18012 10548 18018 10560
rect 18877 10557 18889 10560
rect 18923 10557 18935 10591
rect 18877 10551 18935 10557
rect 18966 10548 18972 10600
rect 19024 10588 19030 10600
rect 19613 10591 19671 10597
rect 19613 10588 19625 10591
rect 19024 10560 19625 10588
rect 19024 10548 19030 10560
rect 19613 10557 19625 10560
rect 19659 10557 19671 10591
rect 19613 10551 19671 10557
rect 19702 10548 19708 10600
rect 19760 10588 19766 10600
rect 20548 10597 20576 10628
rect 20898 10616 20904 10668
rect 20956 10656 20962 10668
rect 21177 10659 21235 10665
rect 21177 10656 21189 10659
rect 20956 10628 21189 10656
rect 20956 10616 20962 10628
rect 21177 10625 21189 10628
rect 21223 10625 21235 10659
rect 21177 10619 21235 10625
rect 21269 10659 21327 10665
rect 21269 10625 21281 10659
rect 21315 10656 21327 10659
rect 22186 10656 22192 10668
rect 21315 10628 22192 10656
rect 21315 10625 21327 10628
rect 21269 10619 21327 10625
rect 22186 10616 22192 10628
rect 22244 10656 22250 10668
rect 22554 10656 22560 10668
rect 22244 10628 22560 10656
rect 22244 10616 22250 10628
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 20533 10591 20591 10597
rect 19760 10560 19805 10588
rect 19760 10548 19766 10560
rect 20533 10557 20545 10591
rect 20579 10557 20591 10591
rect 20533 10551 20591 10557
rect 21453 10591 21511 10597
rect 21453 10557 21465 10591
rect 21499 10588 21511 10591
rect 21542 10588 21548 10600
rect 21499 10560 21548 10588
rect 21499 10557 21511 10560
rect 21453 10551 21511 10557
rect 21542 10548 21548 10560
rect 21600 10548 21606 10600
rect 18230 10520 18236 10532
rect 16868 10492 18236 10520
rect 18230 10480 18236 10492
rect 18288 10480 18294 10532
rect 19628 10492 21312 10520
rect 19628 10464 19656 10492
rect 21284 10464 21312 10492
rect 15160 10424 16252 10452
rect 15160 10412 15166 10424
rect 19610 10412 19616 10464
rect 19668 10412 19674 10464
rect 20714 10412 20720 10464
rect 20772 10452 20778 10464
rect 20809 10455 20867 10461
rect 20809 10452 20821 10455
rect 20772 10424 20821 10452
rect 20772 10412 20778 10424
rect 20809 10421 20821 10424
rect 20855 10421 20867 10455
rect 20809 10415 20867 10421
rect 21266 10412 21272 10464
rect 21324 10412 21330 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1762 10208 1768 10260
rect 1820 10248 1826 10260
rect 1857 10251 1915 10257
rect 1857 10248 1869 10251
rect 1820 10220 1869 10248
rect 1820 10208 1826 10220
rect 1857 10217 1869 10220
rect 1903 10217 1915 10251
rect 3970 10248 3976 10260
rect 3931 10220 3976 10248
rect 1857 10211 1915 10217
rect 3970 10208 3976 10220
rect 4028 10208 4034 10260
rect 4982 10248 4988 10260
rect 4080 10220 4988 10248
rect 4080 10189 4108 10220
rect 4982 10208 4988 10220
rect 5040 10208 5046 10260
rect 5166 10248 5172 10260
rect 5127 10220 5172 10248
rect 5166 10208 5172 10220
rect 5224 10208 5230 10260
rect 5258 10208 5264 10260
rect 5316 10248 5322 10260
rect 5316 10220 6500 10248
rect 5316 10208 5322 10220
rect 4065 10183 4123 10189
rect 4065 10180 4077 10183
rect 3160 10152 4077 10180
rect 2498 10112 2504 10124
rect 2459 10084 2504 10112
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 3160 10056 3188 10152
rect 4065 10149 4077 10152
rect 4111 10149 4123 10183
rect 4065 10143 4123 10149
rect 4706 10140 4712 10192
rect 4764 10180 4770 10192
rect 5442 10180 5448 10192
rect 4764 10152 5448 10180
rect 4764 10140 4770 10152
rect 5442 10140 5448 10152
rect 5500 10180 5506 10192
rect 6365 10183 6423 10189
rect 6365 10180 6377 10183
rect 5500 10152 6377 10180
rect 5500 10140 5506 10152
rect 6365 10149 6377 10152
rect 6411 10149 6423 10183
rect 6472 10180 6500 10220
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 9122 10248 9128 10260
rect 6972 10220 9128 10248
rect 6972 10208 6978 10220
rect 7374 10180 7380 10192
rect 6472 10152 7380 10180
rect 6365 10143 6423 10149
rect 7374 10140 7380 10152
rect 7432 10140 7438 10192
rect 3329 10115 3387 10121
rect 3329 10081 3341 10115
rect 3375 10112 3387 10115
rect 3418 10112 3424 10124
rect 3375 10084 3424 10112
rect 3375 10081 3387 10084
rect 3329 10075 3387 10081
rect 3418 10072 3424 10084
rect 3476 10072 3482 10124
rect 4617 10115 4675 10121
rect 3528 10084 4384 10112
rect 1489 10047 1547 10053
rect 1489 10013 1501 10047
rect 1535 10044 1547 10047
rect 2774 10044 2780 10056
rect 1535 10016 2780 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 2774 10004 2780 10016
rect 2832 10004 2838 10056
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 1670 9976 1676 9988
rect 1631 9948 1676 9976
rect 1670 9936 1676 9948
rect 1728 9936 1734 9988
rect 2222 9908 2228 9920
rect 2183 9880 2228 9908
rect 2222 9868 2228 9880
rect 2280 9868 2286 9920
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 2682 9908 2688 9920
rect 2372 9880 2417 9908
rect 2643 9880 2688 9908
rect 2372 9868 2378 9880
rect 2682 9868 2688 9880
rect 2740 9868 2746 9920
rect 2774 9868 2780 9920
rect 2832 9908 2838 9920
rect 2958 9908 2964 9920
rect 2832 9880 2964 9908
rect 2832 9868 2838 9880
rect 2958 9868 2964 9880
rect 3016 9908 3022 9920
rect 3053 9911 3111 9917
rect 3053 9908 3065 9911
rect 3016 9880 3065 9908
rect 3016 9868 3022 9880
rect 3053 9877 3065 9880
rect 3099 9877 3111 9911
rect 3053 9871 3111 9877
rect 3326 9868 3332 9920
rect 3384 9908 3390 9920
rect 3528 9917 3556 10084
rect 3786 10044 3792 10056
rect 3747 10016 3792 10044
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 4246 10044 4252 10056
rect 4207 10016 4252 10044
rect 4246 10004 4252 10016
rect 4304 10004 4310 10056
rect 4356 10044 4384 10084
rect 4617 10081 4629 10115
rect 4663 10112 4675 10115
rect 4890 10112 4896 10124
rect 4663 10084 4896 10112
rect 4663 10081 4675 10084
rect 4617 10075 4675 10081
rect 4890 10072 4896 10084
rect 4948 10112 4954 10124
rect 5994 10112 6000 10124
rect 4948 10084 6000 10112
rect 4948 10072 4954 10084
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6181 10115 6239 10121
rect 6181 10081 6193 10115
rect 6227 10112 6239 10115
rect 7098 10112 7104 10124
rect 6227 10084 7104 10112
rect 6227 10081 6239 10084
rect 6181 10075 6239 10081
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 8404 10121 8432 10220
rect 8864 10192 8892 10220
rect 9122 10208 9128 10220
rect 9180 10208 9186 10260
rect 10502 10248 10508 10260
rect 10463 10220 10508 10248
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 10778 10208 10784 10260
rect 10836 10248 10842 10260
rect 11885 10251 11943 10257
rect 11885 10248 11897 10251
rect 10836 10220 11897 10248
rect 10836 10208 10842 10220
rect 11885 10217 11897 10220
rect 11931 10217 11943 10251
rect 11885 10211 11943 10217
rect 11974 10208 11980 10260
rect 12032 10248 12038 10260
rect 12069 10251 12127 10257
rect 12069 10248 12081 10251
rect 12032 10220 12081 10248
rect 12032 10208 12038 10220
rect 12069 10217 12081 10220
rect 12115 10217 12127 10251
rect 13630 10248 13636 10260
rect 12069 10211 12127 10217
rect 12176 10220 13636 10248
rect 8846 10140 8852 10192
rect 8904 10140 8910 10192
rect 10594 10180 10600 10192
rect 10555 10152 10600 10180
rect 10594 10140 10600 10152
rect 10652 10140 10658 10192
rect 11790 10180 11796 10192
rect 11703 10152 11796 10180
rect 11790 10140 11796 10152
rect 11848 10180 11854 10192
rect 12176 10180 12204 10220
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 14093 10251 14151 10257
rect 14093 10217 14105 10251
rect 14139 10248 14151 10251
rect 14366 10248 14372 10260
rect 14139 10220 14372 10248
rect 14139 10217 14151 10220
rect 14093 10211 14151 10217
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14918 10248 14924 10260
rect 14879 10220 14924 10248
rect 14918 10208 14924 10220
rect 14976 10208 14982 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 15930 10248 15936 10260
rect 15804 10220 15936 10248
rect 15804 10208 15810 10220
rect 15930 10208 15936 10220
rect 15988 10248 15994 10260
rect 16114 10248 16120 10260
rect 15988 10220 16120 10248
rect 15988 10208 15994 10220
rect 16114 10208 16120 10220
rect 16172 10208 16178 10260
rect 17310 10248 17316 10260
rect 17271 10220 17316 10248
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 18877 10251 18935 10257
rect 18877 10248 18889 10251
rect 17512 10220 18889 10248
rect 11848 10152 12204 10180
rect 11848 10140 11854 10152
rect 13814 10140 13820 10192
rect 13872 10180 13878 10192
rect 13909 10183 13967 10189
rect 13909 10180 13921 10183
rect 13872 10152 13921 10180
rect 13872 10140 13878 10152
rect 13909 10149 13921 10152
rect 13955 10180 13967 10183
rect 14182 10180 14188 10192
rect 13955 10152 14188 10180
rect 13955 10149 13967 10152
rect 13909 10143 13967 10149
rect 14182 10140 14188 10152
rect 14240 10180 14246 10192
rect 14550 10180 14556 10192
rect 14240 10152 14556 10180
rect 14240 10140 14246 10152
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 15378 10180 15384 10192
rect 14660 10152 15384 10180
rect 8389 10115 8447 10121
rect 8389 10081 8401 10115
rect 8435 10081 8447 10115
rect 8389 10075 8447 10081
rect 9125 10115 9183 10121
rect 9125 10081 9137 10115
rect 9171 10081 9183 10115
rect 9125 10075 9183 10081
rect 5445 10047 5503 10053
rect 5445 10044 5457 10047
rect 4356 10016 5457 10044
rect 5445 10013 5457 10016
rect 5491 10013 5503 10047
rect 6638 10044 6644 10056
rect 6599 10016 6644 10044
rect 5445 10007 5503 10013
rect 6638 10004 6644 10016
rect 6696 10004 6702 10056
rect 6914 10044 6920 10056
rect 6875 10016 6920 10044
rect 6914 10004 6920 10016
rect 6972 10004 6978 10056
rect 8110 10004 8116 10056
rect 8168 10053 8174 10056
rect 8168 10044 8180 10053
rect 8168 10016 8213 10044
rect 8168 10007 8180 10016
rect 8168 10004 8174 10007
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 9033 10047 9091 10053
rect 9033 10044 9045 10047
rect 8352 10016 9045 10044
rect 8352 10004 8358 10016
rect 9033 10013 9045 10016
rect 9079 10013 9091 10047
rect 9131 10044 9159 10075
rect 10134 10072 10140 10124
rect 10192 10112 10198 10124
rect 11149 10115 11207 10121
rect 11149 10112 11161 10115
rect 10192 10084 11161 10112
rect 10192 10072 10198 10084
rect 11149 10081 11161 10084
rect 11195 10081 11207 10115
rect 12250 10112 12256 10124
rect 12211 10084 12256 10112
rect 11149 10075 11207 10081
rect 12250 10072 12256 10084
rect 12308 10072 12314 10124
rect 13354 10072 13360 10124
rect 13412 10112 13418 10124
rect 13630 10112 13636 10124
rect 13412 10084 13636 10112
rect 13412 10072 13418 10084
rect 13630 10072 13636 10084
rect 13688 10072 13694 10124
rect 13722 10072 13728 10124
rect 13780 10112 13786 10124
rect 14660 10121 14688 10152
rect 15378 10140 15384 10152
rect 15436 10140 15442 10192
rect 16942 10180 16948 10192
rect 16776 10152 16948 10180
rect 14645 10115 14703 10121
rect 14645 10112 14657 10115
rect 13780 10084 14657 10112
rect 13780 10072 13786 10084
rect 14645 10081 14657 10084
rect 14691 10081 14703 10115
rect 15102 10112 15108 10124
rect 15015 10084 15108 10112
rect 14645 10075 14703 10081
rect 15102 10072 15108 10084
rect 15160 10112 15166 10124
rect 15473 10115 15531 10121
rect 15473 10112 15485 10115
rect 15160 10084 15485 10112
rect 15160 10072 15166 10084
rect 15473 10081 15485 10084
rect 15519 10081 15531 10115
rect 15930 10112 15936 10124
rect 15843 10084 15936 10112
rect 15473 10075 15531 10081
rect 15930 10072 15936 10084
rect 15988 10112 15994 10124
rect 16206 10112 16212 10124
rect 15988 10084 16212 10112
rect 15988 10072 15994 10084
rect 16206 10072 16212 10084
rect 16264 10072 16270 10124
rect 16776 10121 16804 10152
rect 16942 10140 16948 10152
rect 17000 10180 17006 10192
rect 17512 10180 17540 10220
rect 18877 10217 18889 10220
rect 18923 10248 18935 10251
rect 19702 10248 19708 10260
rect 18923 10220 19708 10248
rect 18923 10217 18935 10220
rect 18877 10211 18935 10217
rect 19702 10208 19708 10220
rect 19760 10208 19766 10260
rect 20530 10208 20536 10260
rect 20588 10248 20594 10260
rect 20588 10220 21220 10248
rect 20588 10208 20594 10220
rect 18966 10180 18972 10192
rect 17000 10152 17540 10180
rect 18927 10152 18972 10180
rect 17000 10140 17006 10152
rect 18966 10140 18972 10152
rect 19024 10140 19030 10192
rect 19245 10183 19303 10189
rect 19245 10149 19257 10183
rect 19291 10180 19303 10183
rect 19794 10180 19800 10192
rect 19291 10152 19800 10180
rect 19291 10149 19303 10152
rect 19245 10143 19303 10149
rect 19794 10140 19800 10152
rect 19852 10140 19858 10192
rect 20990 10180 20996 10192
rect 20951 10152 20996 10180
rect 20990 10140 20996 10152
rect 21048 10140 21054 10192
rect 16761 10115 16819 10121
rect 16761 10081 16773 10115
rect 16807 10081 16819 10115
rect 17494 10112 17500 10124
rect 17455 10084 17500 10112
rect 16761 10075 16819 10081
rect 17494 10072 17500 10084
rect 17552 10072 17558 10124
rect 18782 10072 18788 10124
rect 18840 10112 18846 10124
rect 19702 10112 19708 10124
rect 18840 10084 19708 10112
rect 18840 10072 18846 10084
rect 19702 10072 19708 10084
rect 19760 10072 19766 10124
rect 20901 10115 20959 10121
rect 20901 10081 20913 10115
rect 20947 10112 20959 10115
rect 21082 10112 21088 10124
rect 20947 10084 21088 10112
rect 20947 10081 20959 10084
rect 20901 10075 20959 10081
rect 21082 10072 21088 10084
rect 21140 10072 21146 10124
rect 9674 10044 9680 10056
rect 9131 10016 9680 10044
rect 9033 10007 9091 10013
rect 3602 9936 3608 9988
rect 3660 9976 3666 9988
rect 3660 9948 5304 9976
rect 3660 9936 3666 9948
rect 3513 9911 3571 9917
rect 3513 9908 3525 9911
rect 3384 9880 3525 9908
rect 3384 9868 3390 9880
rect 3513 9877 3525 9880
rect 3559 9877 3571 9911
rect 3513 9871 3571 9877
rect 4062 9868 4068 9920
rect 4120 9908 4126 9920
rect 4522 9908 4528 9920
rect 4120 9880 4528 9908
rect 4120 9868 4126 9880
rect 4522 9868 4528 9880
rect 4580 9868 4586 9920
rect 4706 9908 4712 9920
rect 4667 9880 4712 9908
rect 4706 9868 4712 9880
rect 4764 9868 4770 9920
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9908 4859 9911
rect 5166 9908 5172 9920
rect 4847 9880 5172 9908
rect 4847 9877 4859 9880
rect 4801 9871 4859 9877
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 5276 9917 5304 9948
rect 5350 9936 5356 9988
rect 5408 9976 5414 9988
rect 5997 9979 6055 9985
rect 5997 9976 6009 9979
rect 5408 9948 6009 9976
rect 5408 9936 5414 9948
rect 5997 9945 6009 9948
rect 6043 9976 6055 9979
rect 7374 9976 7380 9988
rect 6043 9948 7380 9976
rect 6043 9945 6055 9948
rect 5997 9939 6055 9945
rect 7374 9936 7380 9948
rect 7432 9936 7438 9988
rect 8386 9936 8392 9988
rect 8444 9976 8450 9988
rect 8665 9979 8723 9985
rect 8665 9976 8677 9979
rect 8444 9948 8677 9976
rect 8444 9936 8450 9948
rect 8665 9945 8677 9948
rect 8711 9945 8723 9979
rect 8665 9939 8723 9945
rect 5261 9911 5319 9917
rect 5261 9877 5273 9911
rect 5307 9877 5319 9911
rect 5534 9908 5540 9920
rect 5495 9880 5540 9908
rect 5261 9871 5319 9877
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5902 9908 5908 9920
rect 5863 9880 5908 9908
rect 5902 9868 5908 9880
rect 5960 9868 5966 9920
rect 6638 9868 6644 9920
rect 6696 9908 6702 9920
rect 6733 9911 6791 9917
rect 6733 9908 6745 9911
rect 6696 9880 6745 9908
rect 6696 9868 6702 9880
rect 6733 9877 6745 9880
rect 6779 9877 6791 9911
rect 6733 9871 6791 9877
rect 7009 9911 7067 9917
rect 7009 9877 7021 9911
rect 7055 9908 7067 9911
rect 7098 9908 7104 9920
rect 7055 9880 7104 9908
rect 7055 9877 7067 9880
rect 7009 9871 7067 9877
rect 7098 9868 7104 9880
rect 7156 9908 7162 9920
rect 7926 9908 7932 9920
rect 7156 9880 7932 9908
rect 7156 9868 7162 9880
rect 7926 9868 7932 9880
rect 7984 9868 7990 9920
rect 8570 9908 8576 9920
rect 8483 9880 8576 9908
rect 8570 9868 8576 9880
rect 8628 9908 8634 9920
rect 8938 9908 8944 9920
rect 8628 9880 8944 9908
rect 8628 9868 8634 9880
rect 8938 9868 8944 9880
rect 8996 9868 9002 9920
rect 9048 9908 9076 10007
rect 9674 10004 9680 10016
rect 9732 10004 9738 10056
rect 9858 10004 9864 10056
rect 9916 10044 9922 10056
rect 12520 10047 12578 10053
rect 9916 10016 12480 10044
rect 9916 10004 9922 10016
rect 9122 9936 9128 9988
rect 9180 9976 9186 9988
rect 9370 9979 9428 9985
rect 9370 9976 9382 9979
rect 9180 9948 9382 9976
rect 9180 9936 9186 9948
rect 9370 9945 9382 9948
rect 9416 9945 9428 9979
rect 10870 9976 10876 9988
rect 9370 9939 9428 9945
rect 9692 9948 10876 9976
rect 9692 9920 9720 9948
rect 10870 9936 10876 9948
rect 10928 9936 10934 9988
rect 10965 9979 11023 9985
rect 10965 9945 10977 9979
rect 11011 9976 11023 9979
rect 11425 9979 11483 9985
rect 11425 9976 11437 9979
rect 11011 9948 11437 9976
rect 11011 9945 11023 9948
rect 10965 9939 11023 9945
rect 11425 9945 11437 9948
rect 11471 9945 11483 9979
rect 12452 9976 12480 10016
rect 12520 10013 12532 10047
rect 12566 10044 12578 10047
rect 13538 10044 13544 10056
rect 12566 10016 13544 10044
rect 12566 10013 12578 10016
rect 12520 10007 12578 10013
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 15120 10044 15148 10072
rect 14056 10016 15148 10044
rect 14056 10004 14062 10016
rect 15378 10004 15384 10056
rect 15436 10044 15442 10056
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 15436 10016 16129 10044
rect 15436 10004 15442 10016
rect 16117 10013 16129 10016
rect 16163 10013 16175 10047
rect 16390 10044 16396 10056
rect 16117 10007 16175 10013
rect 16224 10016 16396 10044
rect 16224 9988 16252 10016
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 16853 10047 16911 10053
rect 16853 10013 16865 10047
rect 16899 10044 16911 10047
rect 16942 10044 16948 10056
rect 16899 10016 16948 10044
rect 16899 10013 16911 10016
rect 16853 10007 16911 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17512 10044 17540 10072
rect 21192 10056 21220 10220
rect 18046 10044 18052 10056
rect 17512 10016 18052 10044
rect 18046 10004 18052 10016
rect 18104 10004 18110 10056
rect 19426 10044 19432 10056
rect 19387 10016 19432 10044
rect 19426 10004 19432 10016
rect 19484 10004 19490 10056
rect 21174 10044 21180 10056
rect 21135 10016 21180 10044
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21450 10044 21456 10056
rect 21411 10016 21456 10044
rect 21450 10004 21456 10016
rect 21508 10004 21514 10056
rect 15746 9976 15752 9988
rect 12452 9948 15752 9976
rect 11425 9939 11483 9945
rect 15746 9936 15752 9948
rect 15804 9936 15810 9988
rect 16206 9936 16212 9988
rect 16264 9936 16270 9988
rect 16298 9936 16304 9988
rect 16356 9976 16362 9988
rect 17764 9979 17822 9985
rect 16356 9948 16988 9976
rect 16356 9936 16362 9948
rect 9582 9908 9588 9920
rect 9048 9880 9588 9908
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9674 9868 9680 9920
rect 9732 9868 9738 9920
rect 10042 9868 10048 9920
rect 10100 9908 10106 9920
rect 10778 9908 10784 9920
rect 10100 9880 10784 9908
rect 10100 9868 10106 9880
rect 10778 9868 10784 9880
rect 10836 9868 10842 9920
rect 11054 9908 11060 9920
rect 10967 9880 11060 9908
rect 11054 9868 11060 9880
rect 11112 9908 11118 9920
rect 11790 9908 11796 9920
rect 11112 9880 11796 9908
rect 11112 9868 11118 9880
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 13170 9868 13176 9920
rect 13228 9908 13234 9920
rect 13633 9911 13691 9917
rect 13633 9908 13645 9911
rect 13228 9880 13645 9908
rect 13228 9868 13234 9880
rect 13633 9877 13645 9880
rect 13679 9877 13691 9911
rect 13633 9871 13691 9877
rect 14182 9868 14188 9920
rect 14240 9908 14246 9920
rect 14461 9911 14519 9917
rect 14461 9908 14473 9911
rect 14240 9880 14473 9908
rect 14240 9868 14246 9880
rect 14461 9877 14473 9880
rect 14507 9877 14519 9911
rect 14461 9871 14519 9877
rect 14550 9868 14556 9920
rect 14608 9908 14614 9920
rect 14608 9880 14653 9908
rect 14608 9868 14614 9880
rect 14918 9868 14924 9920
rect 14976 9908 14982 9920
rect 15286 9908 15292 9920
rect 14976 9880 15292 9908
rect 14976 9868 14982 9880
rect 15286 9868 15292 9880
rect 15344 9868 15350 9920
rect 15381 9911 15439 9917
rect 15381 9877 15393 9911
rect 15427 9908 15439 9911
rect 15562 9908 15568 9920
rect 15427 9880 15568 9908
rect 15427 9877 15439 9880
rect 15381 9871 15439 9877
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 15654 9868 15660 9920
rect 15712 9908 15718 9920
rect 16025 9911 16083 9917
rect 16025 9908 16037 9911
rect 15712 9880 16037 9908
rect 15712 9868 15718 9880
rect 16025 9877 16037 9880
rect 16071 9877 16083 9911
rect 16025 9871 16083 9877
rect 16390 9868 16396 9920
rect 16448 9908 16454 9920
rect 16960 9917 16988 9948
rect 17764 9945 17776 9979
rect 17810 9976 17822 9979
rect 17810 9948 18276 9976
rect 17810 9945 17822 9948
rect 17764 9939 17822 9945
rect 18248 9920 18276 9948
rect 20530 9936 20536 9988
rect 20588 9976 20594 9988
rect 20634 9979 20692 9985
rect 20634 9976 20646 9979
rect 20588 9948 20646 9976
rect 20588 9936 20594 9948
rect 20634 9945 20646 9948
rect 20680 9945 20692 9979
rect 20634 9939 20692 9945
rect 20806 9936 20812 9988
rect 20864 9976 20870 9988
rect 20864 9948 21956 9976
rect 20864 9936 20870 9948
rect 16485 9911 16543 9917
rect 16485 9908 16497 9911
rect 16448 9880 16497 9908
rect 16448 9868 16454 9880
rect 16485 9877 16497 9880
rect 16531 9877 16543 9911
rect 16485 9871 16543 9877
rect 16945 9911 17003 9917
rect 16945 9877 16957 9911
rect 16991 9877 17003 9911
rect 16945 9871 17003 9877
rect 18230 9868 18236 9920
rect 18288 9908 18294 9920
rect 19521 9911 19579 9917
rect 19521 9908 19533 9911
rect 18288 9880 19533 9908
rect 18288 9868 18294 9880
rect 19521 9877 19533 9880
rect 19567 9877 19579 9911
rect 19521 9871 19579 9877
rect 20346 9868 20352 9920
rect 20404 9908 20410 9920
rect 21361 9911 21419 9917
rect 21361 9908 21373 9911
rect 20404 9880 21373 9908
rect 20404 9868 20410 9880
rect 21361 9877 21373 9880
rect 21407 9877 21419 9911
rect 21361 9871 21419 9877
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 2133 9707 2191 9713
rect 2133 9673 2145 9707
rect 2179 9704 2191 9707
rect 2314 9704 2320 9716
rect 2179 9676 2320 9704
rect 2179 9673 2191 9676
rect 2133 9667 2191 9673
rect 2314 9664 2320 9676
rect 2372 9664 2378 9716
rect 2593 9707 2651 9713
rect 2593 9673 2605 9707
rect 2639 9704 2651 9707
rect 2682 9704 2688 9716
rect 2639 9676 2688 9704
rect 2639 9673 2651 9676
rect 2593 9667 2651 9673
rect 2682 9664 2688 9676
rect 2740 9664 2746 9716
rect 2958 9664 2964 9716
rect 3016 9704 3022 9716
rect 3786 9704 3792 9716
rect 3016 9676 3792 9704
rect 3016 9664 3022 9676
rect 3786 9664 3792 9676
rect 3844 9664 3850 9716
rect 4065 9707 4123 9713
rect 4065 9673 4077 9707
rect 4111 9704 4123 9707
rect 4338 9704 4344 9716
rect 4111 9676 4344 9704
rect 4111 9673 4123 9676
rect 4065 9667 4123 9673
rect 4338 9664 4344 9676
rect 4396 9664 4402 9716
rect 4525 9707 4583 9713
rect 4525 9673 4537 9707
rect 4571 9704 4583 9707
rect 4706 9704 4712 9716
rect 4571 9676 4712 9704
rect 4571 9673 4583 9676
rect 4525 9667 4583 9673
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 4890 9704 4896 9716
rect 4851 9676 4896 9704
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 4982 9664 4988 9716
rect 5040 9704 5046 9716
rect 5350 9704 5356 9716
rect 5040 9676 5356 9704
rect 5040 9664 5046 9676
rect 5350 9664 5356 9676
rect 5408 9664 5414 9716
rect 5810 9704 5816 9716
rect 5771 9676 5816 9704
rect 5810 9664 5816 9676
rect 5868 9664 5874 9716
rect 5902 9664 5908 9716
rect 5960 9704 5966 9716
rect 6733 9707 6791 9713
rect 6733 9704 6745 9707
rect 5960 9676 6745 9704
rect 5960 9664 5966 9676
rect 6733 9673 6745 9676
rect 6779 9673 6791 9707
rect 6733 9667 6791 9673
rect 7377 9707 7435 9713
rect 7377 9673 7389 9707
rect 7423 9704 7435 9707
rect 7834 9704 7840 9716
rect 7423 9676 7840 9704
rect 7423 9673 7435 9676
rect 7377 9667 7435 9673
rect 7834 9664 7840 9676
rect 7892 9664 7898 9716
rect 9490 9704 9496 9716
rect 8128 9676 9496 9704
rect 1302 9596 1308 9648
rect 1360 9636 1366 9648
rect 1360 9608 1624 9636
rect 1360 9596 1366 9608
rect 1489 9571 1547 9577
rect 1489 9537 1501 9571
rect 1535 9537 1547 9571
rect 1596 9568 1624 9608
rect 1670 9596 1676 9648
rect 1728 9636 1734 9648
rect 3694 9636 3700 9648
rect 1728 9608 3700 9636
rect 1728 9596 1734 9608
rect 3694 9596 3700 9608
rect 3752 9596 3758 9648
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 3804 9608 6561 9636
rect 1765 9571 1823 9577
rect 1765 9568 1777 9571
rect 1596 9540 1777 9568
rect 1489 9531 1547 9537
rect 1765 9537 1777 9540
rect 1811 9537 1823 9571
rect 1765 9531 1823 9537
rect 2501 9571 2559 9577
rect 2501 9537 2513 9571
rect 2547 9568 2559 9571
rect 2866 9568 2872 9580
rect 2547 9540 2872 9568
rect 2547 9537 2559 9540
rect 2501 9531 2559 9537
rect 842 9460 848 9512
rect 900 9500 906 9512
rect 1026 9500 1032 9512
rect 900 9472 1032 9500
rect 900 9460 906 9472
rect 1026 9460 1032 9472
rect 1084 9500 1090 9512
rect 1504 9500 1532 9531
rect 2866 9528 2872 9540
rect 2924 9528 2930 9580
rect 3804 9577 3832 9608
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 8128 9636 8156 9676
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 10410 9704 10416 9716
rect 9876 9676 10416 9704
rect 6549 9599 6607 9605
rect 7760 9608 8156 9636
rect 8205 9639 8263 9645
rect 3789 9571 3847 9577
rect 3789 9568 3801 9571
rect 2976 9540 3801 9568
rect 1084 9472 1532 9500
rect 1084 9460 1090 9472
rect 1854 9460 1860 9512
rect 1912 9500 1918 9512
rect 2682 9500 2688 9512
rect 1912 9472 2688 9500
rect 1912 9460 1918 9472
rect 2682 9460 2688 9472
rect 2740 9460 2746 9512
rect 1946 9432 1952 9444
rect 1907 9404 1952 9432
rect 1946 9392 1952 9404
rect 2004 9432 2010 9444
rect 2314 9432 2320 9444
rect 2004 9404 2320 9432
rect 2004 9392 2010 9404
rect 2314 9392 2320 9404
rect 2372 9392 2378 9444
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 2976 9432 3004 9540
rect 3789 9537 3801 9540
rect 3835 9537 3847 9571
rect 3789 9531 3847 9537
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4246 9568 4252 9580
rect 4203 9540 4252 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4246 9528 4252 9540
rect 4304 9568 4310 9580
rect 4430 9568 4436 9580
rect 4304 9540 4436 9568
rect 4304 9528 4310 9540
rect 4430 9528 4436 9540
rect 4488 9528 4494 9580
rect 4540 9540 5304 9568
rect 4540 9500 4568 9540
rect 2464 9404 3004 9432
rect 3335 9472 4568 9500
rect 2464 9392 2470 9404
rect 1394 9324 1400 9376
rect 1452 9364 1458 9376
rect 1581 9367 1639 9373
rect 1581 9364 1593 9367
rect 1452 9336 1593 9364
rect 1452 9324 1458 9336
rect 1581 9333 1593 9336
rect 1627 9364 1639 9367
rect 2130 9364 2136 9376
rect 1627 9336 2136 9364
rect 1627 9333 1639 9336
rect 1581 9327 1639 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3335 9364 3363 9472
rect 4706 9460 4712 9512
rect 4764 9500 4770 9512
rect 4985 9503 5043 9509
rect 4985 9500 4997 9503
rect 4764 9472 4997 9500
rect 4764 9460 4770 9472
rect 4985 9469 4997 9472
rect 5031 9469 5043 9503
rect 4985 9463 5043 9469
rect 5074 9460 5080 9512
rect 5132 9500 5138 9512
rect 5276 9500 5304 9540
rect 5442 9528 5448 9580
rect 5500 9568 5506 9580
rect 5721 9571 5779 9577
rect 5721 9568 5733 9571
rect 5500 9540 5733 9568
rect 5500 9528 5506 9540
rect 5721 9537 5733 9540
rect 5767 9537 5779 9571
rect 5721 9531 5779 9537
rect 5828 9540 6040 9568
rect 5828 9500 5856 9540
rect 5132 9472 5177 9500
rect 5276 9472 5856 9500
rect 5905 9503 5963 9509
rect 5132 9460 5138 9472
rect 5905 9469 5917 9503
rect 5951 9469 5963 9503
rect 6012 9500 6040 9540
rect 6454 9528 6460 9580
rect 6512 9568 6518 9580
rect 7760 9568 7788 9608
rect 8205 9605 8217 9639
rect 8251 9636 8263 9639
rect 8386 9636 8392 9648
rect 8251 9608 8392 9636
rect 8251 9605 8263 9608
rect 8205 9599 8263 9605
rect 8386 9596 8392 9608
rect 8444 9636 8450 9648
rect 9876 9636 9904 9676
rect 10410 9664 10416 9676
rect 10468 9664 10474 9716
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10689 9707 10747 9713
rect 10689 9704 10701 9707
rect 10652 9676 10701 9704
rect 10652 9664 10658 9676
rect 10689 9673 10701 9676
rect 10735 9673 10747 9707
rect 10689 9667 10747 9673
rect 11974 9664 11980 9716
rect 12032 9704 12038 9716
rect 12710 9704 12716 9716
rect 12032 9676 12716 9704
rect 12032 9664 12038 9676
rect 12710 9664 12716 9676
rect 12768 9664 12774 9716
rect 14550 9704 14556 9716
rect 12820 9676 13584 9704
rect 14511 9676 14556 9704
rect 8444 9608 9904 9636
rect 8444 9596 8450 9608
rect 9950 9596 9956 9648
rect 10008 9636 10014 9648
rect 12820 9636 12848 9676
rect 10008 9608 12848 9636
rect 13357 9639 13415 9645
rect 10008 9596 10014 9608
rect 13357 9605 13369 9639
rect 13403 9636 13415 9639
rect 13556 9636 13584 9676
rect 14550 9664 14556 9676
rect 14608 9664 14614 9716
rect 15010 9704 15016 9716
rect 14971 9676 15016 9704
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 15378 9704 15384 9716
rect 15339 9676 15384 9704
rect 15378 9664 15384 9676
rect 15436 9664 15442 9716
rect 15654 9704 15660 9716
rect 15615 9676 15660 9704
rect 15654 9664 15660 9676
rect 15712 9664 15718 9716
rect 16206 9664 16212 9716
rect 16264 9704 16270 9716
rect 16761 9707 16819 9713
rect 16264 9676 16574 9704
rect 16264 9664 16270 9676
rect 16546 9648 16574 9676
rect 16761 9673 16773 9707
rect 16807 9704 16819 9707
rect 16942 9704 16948 9716
rect 16807 9676 16948 9704
rect 16807 9673 16819 9676
rect 16761 9667 16819 9673
rect 16942 9664 16948 9676
rect 17000 9664 17006 9716
rect 17589 9707 17647 9713
rect 17589 9673 17601 9707
rect 17635 9704 17647 9707
rect 17862 9704 17868 9716
rect 17635 9676 17868 9704
rect 17635 9673 17647 9676
rect 17589 9667 17647 9673
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 19518 9664 19524 9716
rect 19576 9664 19582 9716
rect 20530 9664 20536 9716
rect 20588 9704 20594 9716
rect 20625 9707 20683 9713
rect 20625 9704 20637 9707
rect 20588 9676 20637 9704
rect 20588 9664 20594 9676
rect 20625 9673 20637 9676
rect 20671 9673 20683 9707
rect 20625 9667 20683 9673
rect 20717 9707 20775 9713
rect 20717 9673 20729 9707
rect 20763 9704 20775 9707
rect 21928 9704 21956 9948
rect 20763 9676 21956 9704
rect 20763 9673 20775 9676
rect 20717 9667 20775 9673
rect 13403 9608 13492 9636
rect 13556 9608 15323 9636
rect 13403 9605 13415 9608
rect 13357 9599 13415 9605
rect 6512 9540 7788 9568
rect 8297 9571 8355 9577
rect 6512 9528 6518 9540
rect 8297 9537 8309 9571
rect 8343 9568 8355 9571
rect 8846 9568 8852 9580
rect 8343 9540 8708 9568
rect 8807 9540 8852 9568
rect 8343 9537 8355 9540
rect 8297 9531 8355 9537
rect 6914 9500 6920 9512
rect 6012 9472 6920 9500
rect 5905 9463 5963 9469
rect 3694 9392 3700 9444
rect 3752 9392 3758 9444
rect 4430 9392 4436 9444
rect 4488 9432 4494 9444
rect 4488 9404 5120 9432
rect 4488 9392 4494 9404
rect 3292 9336 3363 9364
rect 3559 9367 3617 9373
rect 3292 9324 3298 9336
rect 3559 9333 3571 9367
rect 3605 9364 3617 9367
rect 3712 9364 3740 9392
rect 4246 9364 4252 9376
rect 3605 9336 4252 9364
rect 3605 9333 3617 9336
rect 3559 9327 3617 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4341 9367 4399 9373
rect 4341 9333 4353 9367
rect 4387 9364 4399 9367
rect 4890 9364 4896 9376
rect 4387 9336 4896 9364
rect 4387 9333 4399 9336
rect 4341 9327 4399 9333
rect 4890 9324 4896 9336
rect 4948 9324 4954 9376
rect 5092 9364 5120 9404
rect 5166 9392 5172 9444
rect 5224 9432 5230 9444
rect 5353 9435 5411 9441
rect 5353 9432 5365 9435
rect 5224 9404 5365 9432
rect 5224 9392 5230 9404
rect 5353 9401 5365 9404
rect 5399 9401 5411 9435
rect 5353 9395 5411 9401
rect 5718 9392 5724 9444
rect 5776 9432 5782 9444
rect 5920 9432 5948 9463
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7466 9500 7472 9512
rect 7427 9472 7472 9500
rect 7466 9460 7472 9472
rect 7524 9460 7530 9512
rect 7653 9503 7711 9509
rect 7653 9469 7665 9503
rect 7699 9500 7711 9503
rect 7926 9500 7932 9512
rect 7699 9472 7932 9500
rect 7699 9469 7711 9472
rect 7653 9463 7711 9469
rect 7926 9460 7932 9472
rect 7984 9460 7990 9512
rect 8110 9460 8116 9512
rect 8168 9500 8174 9512
rect 8389 9503 8447 9509
rect 8389 9500 8401 9503
rect 8168 9472 8401 9500
rect 8168 9460 8174 9472
rect 8389 9469 8401 9472
rect 8435 9469 8447 9503
rect 8389 9463 8447 9469
rect 5776 9404 5948 9432
rect 5776 9392 5782 9404
rect 5994 9392 6000 9444
rect 6052 9432 6058 9444
rect 6365 9435 6423 9441
rect 6365 9432 6377 9435
rect 6052 9404 6377 9432
rect 6052 9392 6058 9404
rect 6365 9401 6377 9404
rect 6411 9401 6423 9435
rect 8294 9432 8300 9444
rect 6365 9395 6423 9401
rect 6932 9404 8300 9432
rect 6932 9364 6960 9404
rect 8294 9392 8300 9404
rect 8352 9392 8358 9444
rect 8680 9376 8708 9540
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 9116 9571 9174 9577
rect 9116 9537 9128 9571
rect 9162 9568 9174 9571
rect 10134 9568 10140 9580
rect 9162 9540 10140 9568
rect 9162 9537 9174 9540
rect 9116 9531 9174 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 11333 9571 11391 9577
rect 11333 9537 11345 9571
rect 11379 9568 11391 9571
rect 12250 9568 12256 9580
rect 11379 9540 12256 9568
rect 11379 9537 11391 9540
rect 11333 9531 11391 9537
rect 12250 9528 12256 9540
rect 12308 9528 12314 9580
rect 12641 9571 12699 9577
rect 12641 9537 12653 9571
rect 12687 9568 12699 9571
rect 12687 9540 13216 9568
rect 12687 9537 12699 9540
rect 12641 9531 12699 9537
rect 13188 9512 13216 9540
rect 13262 9528 13268 9580
rect 13320 9568 13326 9580
rect 13464 9568 13492 9608
rect 13538 9568 13544 9580
rect 13320 9540 13365 9568
rect 13464 9540 13544 9568
rect 13320 9528 13326 9540
rect 13538 9528 13544 9540
rect 13596 9528 13602 9580
rect 13630 9528 13636 9580
rect 13688 9568 13694 9580
rect 14185 9571 14243 9577
rect 14185 9568 14197 9571
rect 13688 9540 14197 9568
rect 13688 9528 13694 9540
rect 14185 9537 14197 9540
rect 14231 9537 14243 9571
rect 14185 9531 14243 9537
rect 10410 9500 10416 9512
rect 10371 9472 10416 9500
rect 10410 9460 10416 9472
rect 10468 9460 10474 9512
rect 10594 9500 10600 9512
rect 10555 9472 10600 9500
rect 10594 9460 10600 9472
rect 10652 9460 10658 9512
rect 12897 9503 12955 9509
rect 12897 9469 12909 9503
rect 12943 9469 12955 9503
rect 13170 9500 13176 9512
rect 13131 9472 13176 9500
rect 12897 9463 12955 9469
rect 9858 9392 9864 9444
rect 9916 9432 9922 9444
rect 9916 9404 11560 9432
rect 9916 9392 9922 9404
rect 5092 9336 6960 9364
rect 7006 9324 7012 9376
rect 7064 9364 7070 9376
rect 7834 9364 7840 9376
rect 7064 9336 7109 9364
rect 7795 9336 7840 9364
rect 7064 9324 7070 9336
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8662 9364 8668 9376
rect 8623 9336 8668 9364
rect 8662 9324 8668 9336
rect 8720 9324 8726 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 10229 9367 10287 9373
rect 10229 9364 10241 9367
rect 9180 9336 10241 9364
rect 9180 9324 9186 9336
rect 10229 9333 10241 9336
rect 10275 9364 10287 9367
rect 10410 9364 10416 9376
rect 10275 9336 10416 9364
rect 10275 9333 10287 9336
rect 10229 9327 10287 9333
rect 10410 9324 10416 9336
rect 10468 9324 10474 9376
rect 10778 9324 10784 9376
rect 10836 9364 10842 9376
rect 11057 9367 11115 9373
rect 11057 9364 11069 9367
rect 10836 9336 11069 9364
rect 10836 9324 10842 9336
rect 11057 9333 11069 9336
rect 11103 9333 11115 9367
rect 11057 9327 11115 9333
rect 11146 9324 11152 9376
rect 11204 9364 11210 9376
rect 11532 9373 11560 9404
rect 11517 9367 11575 9373
rect 11204 9336 11249 9364
rect 11204 9324 11210 9336
rect 11517 9333 11529 9367
rect 11563 9333 11575 9367
rect 11517 9327 11575 9333
rect 12250 9324 12256 9376
rect 12308 9364 12314 9376
rect 12912 9364 12940 9463
rect 13170 9460 13176 9472
rect 13228 9460 13234 9512
rect 13998 9500 14004 9512
rect 13959 9472 14004 9500
rect 13998 9460 14004 9472
rect 14056 9460 14062 9512
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9500 14151 9503
rect 15010 9500 15016 9512
rect 14139 9472 15016 9500
rect 14139 9469 14151 9472
rect 14093 9463 14151 9469
rect 12986 9392 12992 9444
rect 13044 9432 13050 9444
rect 14108 9432 14136 9463
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 13044 9404 14136 9432
rect 13044 9392 13050 9404
rect 14550 9392 14556 9444
rect 14608 9432 14614 9444
rect 14826 9432 14832 9444
rect 14608 9404 14832 9432
rect 14608 9392 14614 9404
rect 14826 9392 14832 9404
rect 14884 9432 14890 9444
rect 15197 9435 15255 9441
rect 15197 9432 15209 9435
rect 14884 9404 15209 9432
rect 14884 9392 14890 9404
rect 15197 9401 15209 9404
rect 15243 9401 15255 9435
rect 15295 9432 15323 9608
rect 15470 9596 15476 9648
rect 15528 9636 15534 9648
rect 16298 9636 16304 9648
rect 15528 9608 16304 9636
rect 15528 9596 15534 9608
rect 16298 9596 16304 9608
rect 16356 9636 16362 9648
rect 16393 9639 16451 9645
rect 16393 9636 16405 9639
rect 16356 9608 16405 9636
rect 16356 9596 16362 9608
rect 16393 9605 16405 9608
rect 16439 9605 16451 9639
rect 16393 9599 16451 9605
rect 16482 9596 16488 9648
rect 16540 9636 16574 9648
rect 16540 9608 17264 9636
rect 16540 9596 16546 9608
rect 16206 9568 16212 9580
rect 16167 9540 16212 9568
rect 16206 9528 16212 9540
rect 16264 9568 16270 9580
rect 17129 9571 17187 9577
rect 17129 9568 17141 9571
rect 16264 9540 17141 9568
rect 16264 9528 16270 9540
rect 17129 9537 17141 9540
rect 17175 9537 17187 9571
rect 17236 9568 17264 9608
rect 17310 9596 17316 9648
rect 17368 9636 17374 9648
rect 18049 9639 18107 9645
rect 18049 9636 18061 9639
rect 17368 9608 18061 9636
rect 17368 9596 17374 9608
rect 18049 9605 18061 9608
rect 18095 9605 18107 9639
rect 19536 9636 19564 9664
rect 20346 9636 20352 9648
rect 18049 9599 18107 9605
rect 18616 9608 20352 9636
rect 17236 9540 17540 9568
rect 17129 9531 17187 9537
rect 15654 9460 15660 9512
rect 15712 9500 15718 9512
rect 16025 9503 16083 9509
rect 16025 9500 16037 9503
rect 15712 9472 16037 9500
rect 15712 9460 15718 9472
rect 16025 9469 16037 9472
rect 16071 9469 16083 9503
rect 17218 9500 17224 9512
rect 17179 9472 17224 9500
rect 16025 9463 16083 9469
rect 17218 9460 17224 9472
rect 17276 9460 17282 9512
rect 17405 9503 17463 9509
rect 17405 9469 17417 9503
rect 17451 9469 17463 9503
rect 17512 9500 17540 9540
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 18616 9577 18644 9608
rect 20346 9596 20352 9608
rect 20404 9596 20410 9648
rect 20640 9636 20668 9667
rect 20640 9608 21312 9636
rect 17957 9571 18015 9577
rect 17957 9568 17969 9571
rect 17736 9540 17969 9568
rect 17736 9528 17742 9540
rect 17957 9537 17969 9540
rect 18003 9537 18015 9571
rect 18417 9571 18475 9577
rect 18417 9568 18429 9571
rect 17957 9531 18015 9537
rect 18064 9540 18429 9568
rect 18064 9500 18092 9540
rect 18417 9537 18429 9540
rect 18463 9537 18475 9571
rect 18417 9531 18475 9537
rect 18601 9571 18659 9577
rect 18601 9537 18613 9571
rect 18647 9537 18659 9571
rect 18601 9531 18659 9537
rect 18690 9528 18696 9580
rect 18748 9568 18754 9580
rect 19058 9568 19064 9580
rect 18748 9540 19064 9568
rect 18748 9528 18754 9540
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19518 9577 19524 9580
rect 19512 9568 19524 9577
rect 19479 9540 19524 9568
rect 19512 9531 19524 9540
rect 19518 9528 19524 9531
rect 19576 9528 19582 9580
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 21085 9571 21143 9577
rect 21085 9568 21097 9571
rect 20036 9540 21097 9568
rect 20036 9528 20042 9540
rect 21085 9537 21097 9540
rect 21131 9537 21143 9571
rect 21085 9531 21143 9537
rect 18230 9500 18236 9512
rect 17512 9472 18092 9500
rect 18191 9472 18236 9500
rect 17405 9463 17463 9469
rect 17310 9432 17316 9444
rect 15295 9404 17316 9432
rect 15197 9395 15255 9401
rect 17310 9392 17316 9404
rect 17368 9392 17374 9444
rect 17420 9432 17448 9463
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18782 9460 18788 9512
rect 18840 9500 18846 9512
rect 19245 9503 19303 9509
rect 19245 9500 19257 9503
rect 18840 9472 19257 9500
rect 18840 9460 18846 9472
rect 19245 9469 19257 9472
rect 19291 9469 19303 9503
rect 19245 9463 19303 9469
rect 20714 9460 20720 9512
rect 20772 9500 20778 9512
rect 21284 9509 21312 9608
rect 21177 9503 21235 9509
rect 21177 9500 21189 9503
rect 20772 9472 21189 9500
rect 20772 9460 20778 9472
rect 21177 9469 21189 9472
rect 21223 9469 21235 9503
rect 21177 9463 21235 9469
rect 21269 9503 21327 9509
rect 21269 9469 21281 9503
rect 21315 9469 21327 9503
rect 21269 9463 21327 9469
rect 18248 9432 18276 9460
rect 17420 9404 18276 9432
rect 18877 9435 18935 9441
rect 18877 9401 18889 9435
rect 18923 9432 18935 9435
rect 19150 9432 19156 9444
rect 18923 9404 19156 9432
rect 18923 9401 18935 9404
rect 18877 9395 18935 9401
rect 19150 9392 19156 9404
rect 19208 9392 19214 9444
rect 12308 9336 12940 9364
rect 12308 9324 12314 9336
rect 13354 9324 13360 9376
rect 13412 9364 13418 9376
rect 13725 9367 13783 9373
rect 13725 9364 13737 9367
rect 13412 9336 13737 9364
rect 13412 9324 13418 9336
rect 13725 9333 13737 9336
rect 13771 9333 13783 9367
rect 14642 9364 14648 9376
rect 14603 9336 14648 9364
rect 13725 9327 13783 9333
rect 14642 9324 14648 9336
rect 14700 9324 14706 9376
rect 14918 9364 14924 9376
rect 14879 9336 14924 9364
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15746 9364 15752 9376
rect 15707 9336 15752 9364
rect 15746 9324 15752 9336
rect 15804 9324 15810 9376
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17678 9364 17684 9376
rect 17276 9336 17684 9364
rect 17276 9324 17282 9336
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 18785 9367 18843 9373
rect 18785 9333 18797 9367
rect 18831 9364 18843 9367
rect 20162 9364 20168 9376
rect 18831 9336 20168 9364
rect 18831 9333 18843 9336
rect 18785 9327 18843 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1949 9163 2007 9169
rect 1949 9129 1961 9163
rect 1995 9129 2007 9163
rect 1949 9123 2007 9129
rect 2041 9163 2099 9169
rect 2041 9129 2053 9163
rect 2087 9160 2099 9163
rect 2222 9160 2228 9172
rect 2087 9132 2228 9160
rect 2087 9129 2099 9132
rect 2041 9123 2099 9129
rect 1964 9092 1992 9123
rect 2222 9120 2228 9132
rect 2280 9120 2286 9172
rect 2406 9120 2412 9172
rect 2464 9160 2470 9172
rect 2866 9160 2872 9172
rect 2464 9132 2774 9160
rect 2827 9132 2872 9160
rect 2464 9120 2470 9132
rect 2498 9092 2504 9104
rect 1964 9064 2504 9092
rect 2498 9052 2504 9064
rect 2556 9052 2562 9104
rect 2746 9092 2774 9132
rect 2866 9120 2872 9132
rect 2924 9120 2930 9172
rect 3789 9163 3847 9169
rect 3789 9129 3801 9163
rect 3835 9160 3847 9163
rect 3878 9160 3884 9172
rect 3835 9132 3884 9160
rect 3835 9129 3847 9132
rect 3789 9123 3847 9129
rect 3878 9120 3884 9132
rect 3936 9120 3942 9172
rect 4062 9120 4068 9172
rect 4120 9120 4126 9172
rect 4706 9120 4712 9172
rect 4764 9160 4770 9172
rect 4764 9132 7420 9160
rect 4764 9120 4770 9132
rect 2746 9064 3556 9092
rect 3528 9036 3556 9064
rect 2682 9024 2688 9036
rect 2643 8996 2688 9024
rect 2682 8984 2688 8996
rect 2740 8984 2746 9036
rect 3329 9027 3387 9033
rect 3329 8993 3341 9027
rect 3375 9024 3387 9027
rect 3418 9024 3424 9036
rect 3375 8996 3424 9024
rect 3375 8993 3387 8996
rect 3329 8987 3387 8993
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 3510 8984 3516 9036
rect 3568 9024 3574 9036
rect 4080 9024 4108 9120
rect 4249 9095 4307 9101
rect 4249 9061 4261 9095
rect 4295 9092 4307 9095
rect 4338 9092 4344 9104
rect 4295 9064 4344 9092
rect 4295 9061 4307 9064
rect 4249 9055 4307 9061
rect 4338 9052 4344 9064
rect 4396 9052 4402 9104
rect 6914 9052 6920 9104
rect 6972 9092 6978 9104
rect 7285 9095 7343 9101
rect 7285 9092 7297 9095
rect 6972 9064 7297 9092
rect 6972 9052 6978 9064
rect 7285 9061 7297 9064
rect 7331 9061 7343 9095
rect 7392 9092 7420 9132
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 7561 9163 7619 9169
rect 7561 9160 7573 9163
rect 7524 9132 7573 9160
rect 7524 9120 7530 9132
rect 7561 9129 7573 9132
rect 7607 9129 7619 9163
rect 7561 9123 7619 9129
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 9125 9163 9183 9169
rect 9125 9160 9137 9163
rect 7800 9132 9137 9160
rect 7800 9120 7806 9132
rect 9125 9129 9137 9132
rect 9171 9129 9183 9163
rect 9125 9123 9183 9129
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9401 9163 9459 9169
rect 9401 9160 9413 9163
rect 9364 9132 9413 9160
rect 9364 9120 9370 9132
rect 9401 9129 9413 9132
rect 9447 9129 9459 9163
rect 9401 9123 9459 9129
rect 10321 9163 10379 9169
rect 10321 9129 10333 9163
rect 10367 9160 10379 9163
rect 10594 9160 10600 9172
rect 10367 9132 10600 9160
rect 10367 9129 10379 9132
rect 10321 9123 10379 9129
rect 10594 9120 10600 9132
rect 10652 9120 10658 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 11790 9160 11796 9172
rect 10928 9132 11796 9160
rect 10928 9120 10934 9132
rect 11790 9120 11796 9132
rect 11848 9120 11854 9172
rect 11974 9160 11980 9172
rect 11935 9132 11980 9160
rect 11974 9120 11980 9132
rect 12032 9120 12038 9172
rect 12805 9163 12863 9169
rect 12805 9129 12817 9163
rect 12851 9160 12863 9163
rect 12894 9160 12900 9172
rect 12851 9132 12900 9160
rect 12851 9129 12863 9132
rect 12805 9123 12863 9129
rect 12894 9120 12900 9132
rect 12952 9160 12958 9172
rect 13538 9160 13544 9172
rect 12952 9132 13544 9160
rect 12952 9120 12958 9132
rect 13538 9120 13544 9132
rect 13596 9160 13602 9172
rect 14366 9160 14372 9172
rect 13596 9132 14372 9160
rect 13596 9120 13602 9132
rect 14366 9120 14372 9132
rect 14424 9120 14430 9172
rect 15102 9120 15108 9172
rect 15160 9160 15166 9172
rect 16577 9163 16635 9169
rect 15160 9132 16068 9160
rect 15160 9120 15166 9132
rect 8478 9092 8484 9104
rect 7392 9064 8484 9092
rect 7285 9055 7343 9061
rect 7300 9024 7328 9055
rect 8478 9052 8484 9064
rect 8536 9052 8542 9104
rect 8662 9052 8668 9104
rect 8720 9092 8726 9104
rect 8720 9064 11468 9092
rect 8720 9052 8726 9064
rect 3568 8996 3661 9024
rect 4080 8996 4476 9024
rect 7300 8996 8064 9024
rect 3568 8984 3574 8996
rect 4448 8968 4476 8996
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1486 8956 1492 8968
rect 1443 8928 1492 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1486 8916 1492 8928
rect 1544 8916 1550 8968
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 1765 8959 1823 8965
rect 1765 8956 1777 8959
rect 1636 8928 1777 8956
rect 1636 8916 1642 8928
rect 1765 8925 1777 8928
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 2774 8916 2780 8968
rect 2832 8956 2838 8968
rect 3973 8959 4031 8965
rect 3973 8956 3985 8959
rect 2832 8928 3985 8956
rect 2832 8916 2838 8928
rect 3973 8925 3985 8928
rect 4019 8925 4031 8959
rect 3973 8919 4031 8925
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 4338 8956 4344 8968
rect 4120 8928 4165 8956
rect 4299 8928 4344 8956
rect 4120 8916 4126 8928
rect 4338 8916 4344 8928
rect 4396 8916 4402 8968
rect 4430 8916 4436 8968
rect 4488 8916 4494 8968
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 4540 8928 5825 8956
rect 2866 8848 2872 8900
rect 2924 8888 2930 8900
rect 2924 8860 4108 8888
rect 2924 8848 2930 8860
rect 4080 8832 4108 8860
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2406 8820 2412 8832
rect 2367 8792 2412 8820
rect 2406 8780 2412 8792
rect 2464 8780 2470 8832
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 3234 8820 3240 8832
rect 2556 8792 2601 8820
rect 3195 8792 3240 8820
rect 2556 8780 2562 8792
rect 3234 8780 3240 8792
rect 3292 8780 3298 8832
rect 4062 8780 4068 8832
rect 4120 8780 4126 8832
rect 4338 8780 4344 8832
rect 4396 8820 4402 8832
rect 4540 8820 4568 8928
rect 5813 8925 5825 8928
rect 5859 8956 5871 8959
rect 6638 8956 6644 8968
rect 5859 8928 6644 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 6638 8916 6644 8928
rect 6696 8916 6702 8968
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8956 7527 8959
rect 7742 8956 7748 8968
rect 7515 8928 7748 8956
rect 7515 8925 7527 8928
rect 7469 8919 7527 8925
rect 7742 8916 7748 8928
rect 7800 8916 7806 8968
rect 7926 8956 7932 8968
rect 7852 8928 7932 8956
rect 4608 8891 4666 8897
rect 4608 8857 4620 8891
rect 4654 8888 4666 8891
rect 5626 8888 5632 8900
rect 4654 8860 5632 8888
rect 4654 8857 4666 8860
rect 4608 8851 4666 8857
rect 5626 8848 5632 8860
rect 5684 8888 5690 8900
rect 5684 8860 5856 8888
rect 5684 8848 5690 8860
rect 5718 8820 5724 8832
rect 4396 8792 4568 8820
rect 5679 8792 5724 8820
rect 4396 8780 4402 8792
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 5828 8820 5856 8860
rect 5902 8848 5908 8900
rect 5960 8888 5966 8900
rect 6080 8891 6138 8897
rect 6080 8888 6092 8891
rect 5960 8860 6092 8888
rect 5960 8848 5966 8860
rect 6080 8857 6092 8860
rect 6126 8888 6138 8891
rect 7852 8888 7880 8928
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8036 8956 8064 8996
rect 8110 8984 8116 9036
rect 8168 9024 8174 9036
rect 8386 9024 8392 9036
rect 8168 8996 8213 9024
rect 8347 8996 8392 9024
rect 8168 8984 8174 8996
rect 8386 8984 8392 8996
rect 8444 8984 8450 9036
rect 9769 9027 9827 9033
rect 8680 8996 9536 9024
rect 8680 8956 8708 8996
rect 8036 8928 8708 8956
rect 8757 8959 8815 8965
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 9030 8956 9036 8968
rect 8803 8928 9036 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 9030 8916 9036 8928
rect 9088 8916 9094 8968
rect 9508 8956 9536 8996
rect 9769 8993 9781 9027
rect 9815 9024 9827 9027
rect 10134 9024 10140 9036
rect 9815 8996 10140 9024
rect 9815 8993 9827 8996
rect 9769 8987 9827 8993
rect 10134 8984 10140 8996
rect 10192 8984 10198 9036
rect 10502 9024 10508 9036
rect 10463 8996 10508 9024
rect 10502 8984 10508 8996
rect 10560 8984 10566 9036
rect 10612 8996 10916 9024
rect 10612 8956 10640 8996
rect 10778 8956 10784 8968
rect 9508 8928 10640 8956
rect 10739 8928 10784 8956
rect 10778 8916 10784 8928
rect 10836 8916 10842 8968
rect 10888 8956 10916 8996
rect 11146 8984 11152 9036
rect 11204 9024 11210 9036
rect 11333 9027 11391 9033
rect 11333 9024 11345 9027
rect 11204 8996 11345 9024
rect 11204 8984 11210 8996
rect 11333 8993 11345 8996
rect 11379 8993 11391 9027
rect 11440 9024 11468 9064
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 12069 9095 12127 9101
rect 12069 9092 12081 9095
rect 11664 9064 12081 9092
rect 11664 9052 11670 9064
rect 12069 9061 12081 9064
rect 12115 9061 12127 9095
rect 12986 9092 12992 9104
rect 12069 9055 12127 9061
rect 12176 9064 12992 9092
rect 12176 9024 12204 9064
rect 12986 9052 12992 9064
rect 13044 9052 13050 9104
rect 11440 8996 12204 9024
rect 11333 8987 11391 8993
rect 12802 8984 12808 9036
rect 12860 9024 12866 9036
rect 13909 9027 13967 9033
rect 12860 8996 13860 9024
rect 12860 8984 12866 8996
rect 11514 8956 11520 8968
rect 10888 8928 11520 8956
rect 11514 8916 11520 8928
rect 11572 8916 11578 8968
rect 12434 8956 12440 8968
rect 11624 8928 12440 8956
rect 9582 8888 9588 8900
rect 6126 8860 7880 8888
rect 7944 8860 9588 8888
rect 6126 8857 6138 8860
rect 6080 8851 6138 8857
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 5828 8792 7205 8820
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 7282 8780 7288 8832
rect 7340 8820 7346 8832
rect 7944 8829 7972 8860
rect 9582 8848 9588 8860
rect 9640 8848 9646 8900
rect 10318 8848 10324 8900
rect 10376 8888 10382 8900
rect 11624 8888 11652 8928
rect 12434 8916 12440 8928
rect 12492 8916 12498 8968
rect 12989 8959 13047 8965
rect 12989 8925 13001 8959
rect 13035 8956 13047 8959
rect 13170 8956 13176 8968
rect 13035 8928 13176 8956
rect 13035 8925 13047 8928
rect 12989 8919 13047 8925
rect 13170 8916 13176 8928
rect 13228 8916 13234 8968
rect 13832 8956 13860 8996
rect 13909 8993 13921 9027
rect 13955 9024 13967 9027
rect 14182 9024 14188 9036
rect 13955 8996 14188 9024
rect 13955 8993 13967 8996
rect 13909 8987 13967 8993
rect 14182 8984 14188 8996
rect 14240 8984 14246 9036
rect 15562 9024 15568 9036
rect 15396 8996 15568 9024
rect 14826 8956 14832 8968
rect 13832 8928 14832 8956
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 15217 8959 15275 8965
rect 15217 8925 15229 8959
rect 15263 8956 15275 8959
rect 15396 8956 15424 8996
rect 15562 8984 15568 8996
rect 15620 9024 15626 9036
rect 15933 9027 15991 9033
rect 15933 9024 15945 9027
rect 15620 8996 15945 9024
rect 15620 8984 15626 8996
rect 15933 8993 15945 8996
rect 15979 8993 15991 9027
rect 15933 8987 15991 8993
rect 15263 8928 15424 8956
rect 15473 8959 15531 8965
rect 15263 8925 15275 8928
rect 15217 8919 15275 8925
rect 15473 8925 15485 8959
rect 15519 8925 15531 8959
rect 15473 8919 15531 8925
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 15838 8956 15844 8968
rect 15795 8928 15844 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 10376 8860 11652 8888
rect 10376 8848 10382 8860
rect 11790 8848 11796 8900
rect 11848 8888 11854 8900
rect 13630 8888 13636 8900
rect 11848 8860 13636 8888
rect 11848 8848 11854 8860
rect 13630 8848 13636 8860
rect 13688 8848 13694 8900
rect 14016 8860 14504 8888
rect 7929 8823 7987 8829
rect 7929 8820 7941 8823
rect 7340 8792 7941 8820
rect 7340 8780 7346 8792
rect 7929 8789 7941 8792
rect 7975 8789 7987 8823
rect 7929 8783 7987 8789
rect 8021 8823 8079 8829
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8110 8820 8116 8832
rect 8067 8792 8116 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8386 8780 8392 8832
rect 8444 8820 8450 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 8444 8792 8585 8820
rect 8444 8780 8450 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 8662 8780 8668 8832
rect 8720 8820 8726 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8720 8792 8953 8820
rect 8720 8780 8726 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 8941 8783 8999 8789
rect 9306 8780 9312 8832
rect 9364 8820 9370 8832
rect 9861 8823 9919 8829
rect 9861 8820 9873 8823
rect 9364 8792 9873 8820
rect 9364 8780 9370 8792
rect 9861 8789 9873 8792
rect 9907 8789 9919 8823
rect 9861 8783 9919 8789
rect 9953 8823 10011 8829
rect 9953 8789 9965 8823
rect 9999 8820 10011 8823
rect 10410 8820 10416 8832
rect 9999 8792 10416 8820
rect 9999 8789 10011 8792
rect 9953 8783 10011 8789
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10686 8820 10692 8832
rect 10647 8792 10692 8820
rect 10686 8780 10692 8792
rect 10744 8780 10750 8832
rect 10962 8780 10968 8832
rect 11020 8820 11026 8832
rect 11149 8823 11207 8829
rect 11149 8820 11161 8823
rect 11020 8792 11161 8820
rect 11020 8780 11026 8792
rect 11149 8789 11161 8792
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 11238 8780 11244 8832
rect 11296 8820 11302 8832
rect 11517 8823 11575 8829
rect 11517 8820 11529 8823
rect 11296 8792 11529 8820
rect 11296 8780 11302 8792
rect 11517 8789 11529 8792
rect 11563 8789 11575 8823
rect 11517 8783 11575 8789
rect 11609 8823 11667 8829
rect 11609 8789 11621 8823
rect 11655 8820 11667 8823
rect 11698 8820 11704 8832
rect 11655 8792 11704 8820
rect 11655 8789 11667 8792
rect 11609 8783 11667 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12526 8820 12532 8832
rect 12487 8792 12532 8820
rect 12526 8780 12532 8792
rect 12584 8780 12590 8832
rect 13078 8820 13084 8832
rect 13039 8792 13084 8820
rect 13078 8780 13084 8792
rect 13136 8780 13142 8832
rect 13357 8823 13415 8829
rect 13357 8789 13369 8823
rect 13403 8820 13415 8823
rect 13446 8820 13452 8832
rect 13403 8792 13452 8820
rect 13403 8789 13415 8792
rect 13357 8783 13415 8789
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 14016 8820 14044 8860
rect 14476 8832 14504 8860
rect 13587 8792 14044 8820
rect 14093 8823 14151 8829
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 14093 8789 14105 8823
rect 14139 8820 14151 8823
rect 14366 8820 14372 8832
rect 14139 8792 14372 8820
rect 14139 8789 14151 8792
rect 14093 8783 14151 8789
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14458 8780 14464 8832
rect 14516 8780 14522 8832
rect 15010 8780 15016 8832
rect 15068 8820 15074 8832
rect 15488 8820 15516 8919
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16040 8956 16068 9132
rect 16577 9129 16589 9163
rect 16623 9160 16635 9163
rect 17126 9160 17132 9172
rect 16623 9132 17132 9160
rect 16623 9129 16635 9132
rect 16577 9123 16635 9129
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17310 9120 17316 9172
rect 17368 9160 17374 9172
rect 17589 9163 17647 9169
rect 17589 9160 17601 9163
rect 17368 9132 17601 9160
rect 17368 9120 17374 9132
rect 17589 9129 17601 9132
rect 17635 9129 17647 9163
rect 17589 9123 17647 9129
rect 19518 9120 19524 9172
rect 19576 9160 19582 9172
rect 20714 9160 20720 9172
rect 19576 9132 20208 9160
rect 20675 9132 20720 9160
rect 19576 9120 19582 9132
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 17770 9092 17776 9104
rect 17092 9064 17776 9092
rect 17092 9052 17098 9064
rect 17770 9052 17776 9064
rect 17828 9052 17834 9104
rect 18690 9092 18696 9104
rect 17972 9064 18696 9092
rect 16206 8984 16212 9036
rect 16264 9024 16270 9036
rect 16482 9024 16488 9036
rect 16264 8996 16488 9024
rect 16264 8984 16270 8996
rect 16482 8984 16488 8996
rect 16540 8984 16546 9036
rect 17218 9024 17224 9036
rect 17179 8996 17224 9024
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 17972 9024 18000 9064
rect 18690 9052 18696 9064
rect 18748 9092 18754 9104
rect 18966 9092 18972 9104
rect 18748 9064 18972 9092
rect 18748 9052 18754 9064
rect 18966 9052 18972 9064
rect 19024 9052 19030 9104
rect 20180 9092 20208 9132
rect 20714 9120 20720 9132
rect 20772 9120 20778 9172
rect 20625 9095 20683 9101
rect 20625 9092 20637 9095
rect 20180 9064 20637 9092
rect 20625 9061 20637 9064
rect 20671 9061 20683 9095
rect 20625 9055 20683 9061
rect 17880 8996 18000 9024
rect 18509 9027 18567 9033
rect 17880 8965 17908 8996
rect 18509 8993 18521 9027
rect 18555 8993 18567 9027
rect 18509 8987 18567 8993
rect 17129 8959 17187 8965
rect 17129 8956 17141 8959
rect 16040 8928 17141 8956
rect 17129 8925 17141 8928
rect 17175 8925 17187 8959
rect 17129 8919 17187 8925
rect 17865 8959 17923 8965
rect 17865 8925 17877 8959
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 17957 8959 18015 8965
rect 17957 8925 17969 8959
rect 18003 8956 18015 8959
rect 18046 8956 18052 8968
rect 18003 8928 18052 8956
rect 18003 8925 18015 8928
rect 17957 8919 18015 8925
rect 18046 8916 18052 8928
rect 18104 8916 18110 8968
rect 18524 8956 18552 8987
rect 18782 8984 18788 9036
rect 18840 9024 18846 9036
rect 19245 9027 19303 9033
rect 19245 9024 19257 9027
rect 18840 8996 19257 9024
rect 18840 8984 18846 8996
rect 19245 8993 19257 8996
rect 19291 8993 19303 9027
rect 20640 9024 20668 9055
rect 21269 9027 21327 9033
rect 21269 9024 21281 9027
rect 20640 8996 21281 9024
rect 19245 8987 19303 8993
rect 21269 8993 21281 8996
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 19886 8956 19892 8968
rect 18524 8928 19892 8956
rect 19886 8916 19892 8928
rect 19944 8916 19950 8968
rect 20622 8916 20628 8968
rect 20680 8956 20686 8968
rect 21177 8959 21235 8965
rect 21177 8956 21189 8959
rect 20680 8928 21189 8956
rect 20680 8916 20686 8928
rect 21177 8925 21189 8928
rect 21223 8925 21235 8959
rect 21177 8919 21235 8925
rect 16209 8891 16267 8897
rect 16209 8857 16221 8891
rect 16255 8888 16267 8891
rect 16255 8860 16712 8888
rect 16255 8857 16267 8860
rect 16209 8851 16267 8857
rect 15565 8823 15623 8829
rect 15565 8820 15577 8823
rect 15068 8792 15577 8820
rect 15068 8780 15074 8792
rect 15565 8789 15577 8792
rect 15611 8789 15623 8823
rect 16114 8820 16120 8832
rect 16075 8792 16120 8820
rect 15565 8783 15623 8789
rect 16114 8780 16120 8792
rect 16172 8780 16178 8832
rect 16684 8829 16712 8860
rect 17586 8848 17592 8900
rect 17644 8888 17650 8900
rect 18693 8891 18751 8897
rect 18693 8888 18705 8891
rect 17644 8860 18705 8888
rect 17644 8848 17650 8860
rect 18693 8857 18705 8860
rect 18739 8857 18751 8891
rect 18693 8851 18751 8857
rect 19512 8891 19570 8897
rect 19512 8857 19524 8891
rect 19558 8888 19570 8891
rect 19794 8888 19800 8900
rect 19558 8860 19800 8888
rect 19558 8857 19570 8860
rect 19512 8851 19570 8857
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 16669 8823 16727 8829
rect 16669 8789 16681 8823
rect 16715 8789 16727 8823
rect 17034 8820 17040 8832
rect 16995 8792 17040 8820
rect 16669 8783 16727 8789
rect 17034 8780 17040 8792
rect 17092 8780 17098 8832
rect 17494 8780 17500 8832
rect 17552 8820 17558 8832
rect 17681 8823 17739 8829
rect 17681 8820 17693 8823
rect 17552 8792 17693 8820
rect 17552 8780 17558 8792
rect 17681 8789 17693 8792
rect 17727 8789 17739 8823
rect 17681 8783 17739 8789
rect 18141 8823 18199 8829
rect 18141 8789 18153 8823
rect 18187 8820 18199 8823
rect 18414 8820 18420 8832
rect 18187 8792 18420 8820
rect 18187 8789 18199 8792
rect 18141 8783 18199 8789
rect 18414 8780 18420 8792
rect 18472 8780 18478 8832
rect 18601 8823 18659 8829
rect 18601 8789 18613 8823
rect 18647 8820 18659 8823
rect 18966 8820 18972 8832
rect 18647 8792 18972 8820
rect 18647 8789 18659 8792
rect 18601 8783 18659 8789
rect 18966 8780 18972 8792
rect 19024 8780 19030 8832
rect 19061 8823 19119 8829
rect 19061 8789 19073 8823
rect 19107 8820 19119 8823
rect 19702 8820 19708 8832
rect 19107 8792 19708 8820
rect 19107 8789 19119 8792
rect 19061 8783 19119 8789
rect 19702 8780 19708 8792
rect 19760 8780 19766 8832
rect 21082 8820 21088 8832
rect 21043 8792 21088 8820
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 2498 8616 2504 8628
rect 2271 8588 2504 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 4982 8616 4988 8628
rect 2746 8588 4988 8616
rect 1857 8551 1915 8557
rect 1857 8517 1869 8551
rect 1903 8548 1915 8551
rect 2746 8548 2774 8588
rect 4982 8576 4988 8588
rect 5040 8576 5046 8628
rect 5166 8616 5172 8628
rect 5127 8588 5172 8616
rect 5166 8576 5172 8588
rect 5224 8576 5230 8628
rect 5258 8576 5264 8628
rect 5316 8576 5322 8628
rect 5810 8576 5816 8628
rect 5868 8616 5874 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 5868 8588 6561 8616
rect 5868 8576 5874 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 6917 8619 6975 8625
rect 6917 8585 6929 8619
rect 6963 8616 6975 8619
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 6963 8588 7389 8616
rect 6963 8585 6975 8588
rect 6917 8579 6975 8585
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7834 8616 7840 8628
rect 7795 8588 7840 8616
rect 7377 8579 7435 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8941 8619 8999 8625
rect 8941 8585 8953 8619
rect 8987 8616 8999 8619
rect 9401 8619 9459 8625
rect 9401 8616 9413 8619
rect 8987 8588 9413 8616
rect 8987 8585 8999 8588
rect 8941 8579 8999 8585
rect 9401 8585 9413 8588
rect 9447 8585 9459 8619
rect 9401 8579 9459 8585
rect 9769 8619 9827 8625
rect 9769 8585 9781 8619
rect 9815 8585 9827 8619
rect 9950 8616 9956 8628
rect 9911 8588 9956 8616
rect 9769 8579 9827 8585
rect 4056 8551 4114 8557
rect 4056 8548 4068 8551
rect 1903 8520 2774 8548
rect 3712 8520 4068 8548
rect 1903 8517 1915 8520
rect 1857 8511 1915 8517
rect 1946 8440 1952 8492
rect 2004 8480 2010 8492
rect 2573 8483 2631 8489
rect 2573 8480 2585 8483
rect 2004 8452 2585 8480
rect 2004 8440 2010 8452
rect 2573 8449 2585 8452
rect 2619 8449 2631 8483
rect 2573 8443 2631 8449
rect 1670 8412 1676 8424
rect 1631 8384 1676 8412
rect 1670 8372 1676 8384
rect 1728 8372 1734 8424
rect 1765 8415 1823 8421
rect 1765 8381 1777 8415
rect 1811 8412 1823 8415
rect 2222 8412 2228 8424
rect 1811 8384 2228 8412
rect 1811 8381 1823 8384
rect 1765 8375 1823 8381
rect 2222 8372 2228 8384
rect 2280 8372 2286 8424
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8381 2375 8415
rect 2317 8375 2375 8381
rect 2332 8276 2360 8375
rect 3712 8353 3740 8520
rect 4056 8517 4068 8520
rect 4102 8548 4114 8551
rect 5276 8548 5304 8576
rect 5902 8548 5908 8560
rect 4102 8520 5304 8548
rect 5552 8520 5908 8548
rect 4102 8517 4114 8520
rect 4056 8511 4114 8517
rect 4338 8480 4344 8492
rect 3804 8452 4344 8480
rect 3804 8421 3832 8452
rect 4338 8440 4344 8452
rect 4396 8440 4402 8492
rect 5258 8480 5264 8492
rect 5219 8452 5264 8480
rect 5258 8440 5264 8452
rect 5316 8440 5322 8492
rect 5552 8421 5580 8520
rect 5902 8508 5908 8520
rect 5960 8508 5966 8560
rect 8294 8508 8300 8560
rect 8352 8548 8358 8560
rect 9490 8548 9496 8560
rect 8352 8520 9496 8548
rect 8352 8508 8358 8520
rect 9490 8508 9496 8520
rect 9548 8508 9554 8560
rect 5813 8483 5871 8489
rect 5813 8449 5825 8483
rect 5859 8480 5871 8483
rect 6086 8480 6092 8492
rect 5859 8452 6092 8480
rect 5859 8449 5871 8452
rect 5813 8443 5871 8449
rect 6086 8440 6092 8452
rect 6144 8440 6150 8492
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 7745 8483 7803 8489
rect 7745 8480 7757 8483
rect 6420 8452 7135 8480
rect 6420 8440 6426 8452
rect 3789 8415 3847 8421
rect 3789 8381 3801 8415
rect 3835 8381 3847 8415
rect 3789 8375 3847 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8381 5595 8415
rect 5721 8415 5779 8421
rect 5721 8412 5733 8415
rect 5537 8375 5595 8381
rect 5644 8384 5733 8412
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8313 3755 8347
rect 3697 8307 3755 8313
rect 3804 8276 3832 8375
rect 2332 8248 3832 8276
rect 3970 8236 3976 8288
rect 4028 8276 4034 8288
rect 5644 8276 5672 8384
rect 5721 8381 5733 8384
rect 5767 8412 5779 8415
rect 6454 8412 6460 8424
rect 5767 8384 6460 8412
rect 5767 8381 5779 8384
rect 5721 8375 5779 8381
rect 6454 8372 6460 8384
rect 6512 8372 6518 8424
rect 6730 8372 6736 8424
rect 6788 8412 6794 8424
rect 7107 8421 7135 8452
rect 7280 8452 7757 8480
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 6788 8384 7021 8412
rect 6788 8372 6794 8384
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7009 8375 7067 8381
rect 7101 8415 7159 8421
rect 7101 8381 7113 8415
rect 7147 8381 7159 8415
rect 7101 8375 7159 8381
rect 6546 8304 6552 8356
rect 6604 8344 6610 8356
rect 7280 8344 7308 8452
rect 7745 8449 7757 8452
rect 7791 8449 7803 8483
rect 7745 8443 7803 8449
rect 7834 8440 7840 8492
rect 7892 8480 7898 8492
rect 8018 8480 8024 8492
rect 7892 8452 8024 8480
rect 7892 8440 7898 8452
rect 8018 8440 8024 8452
rect 8076 8440 8082 8492
rect 8573 8484 8631 8489
rect 8573 8483 8708 8484
rect 8573 8449 8585 8483
rect 8619 8480 8708 8483
rect 9398 8480 9404 8492
rect 8619 8456 9404 8480
rect 8619 8449 8631 8456
rect 8680 8452 9404 8456
rect 8573 8443 8631 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9784 8480 9812 8579
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10686 8616 10692 8628
rect 10060 8588 10692 8616
rect 10060 8480 10088 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 10870 8616 10876 8628
rect 10831 8588 10876 8616
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 11333 8619 11391 8625
rect 11333 8616 11345 8619
rect 11296 8588 11345 8616
rect 11296 8576 11302 8588
rect 11333 8585 11345 8588
rect 11379 8585 11391 8619
rect 11333 8579 11391 8585
rect 11517 8619 11575 8625
rect 11517 8585 11529 8619
rect 11563 8585 11575 8619
rect 12802 8616 12808 8628
rect 11517 8579 11575 8585
rect 11808 8588 12808 8616
rect 10594 8508 10600 8560
rect 10652 8548 10658 8560
rect 10965 8551 11023 8557
rect 10965 8548 10977 8551
rect 10652 8520 10977 8548
rect 10652 8508 10658 8520
rect 10965 8517 10977 8520
rect 11011 8517 11023 8551
rect 10965 8511 11023 8517
rect 11146 8508 11152 8560
rect 11204 8548 11210 8560
rect 11532 8548 11560 8579
rect 11204 8520 11560 8548
rect 11204 8508 11210 8520
rect 10410 8480 10416 8492
rect 9784 8452 10088 8480
rect 10371 8452 10416 8480
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 11808 8480 11836 8588
rect 12802 8576 12808 8588
rect 12860 8576 12866 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13817 8619 13875 8625
rect 13817 8616 13829 8619
rect 13403 8588 13829 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13817 8585 13829 8588
rect 13863 8585 13875 8619
rect 14182 8616 14188 8628
rect 14143 8588 14188 8616
rect 13817 8579 13875 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 14645 8619 14703 8625
rect 14645 8585 14657 8619
rect 14691 8585 14703 8619
rect 14645 8579 14703 8585
rect 12250 8508 12256 8560
rect 12308 8548 12314 8560
rect 13449 8551 13507 8557
rect 12308 8520 12940 8548
rect 12308 8508 12314 8520
rect 12912 8489 12940 8520
rect 13449 8517 13461 8551
rect 13495 8548 13507 8551
rect 13722 8548 13728 8560
rect 13495 8520 13728 8548
rect 13495 8517 13507 8520
rect 13449 8511 13507 8517
rect 13722 8508 13728 8520
rect 13780 8508 13786 8560
rect 14660 8548 14688 8579
rect 14826 8576 14832 8628
rect 14884 8616 14890 8628
rect 15470 8616 15476 8628
rect 14884 8588 15476 8616
rect 14884 8576 14890 8588
rect 15470 8576 15476 8588
rect 15528 8576 15534 8628
rect 16114 8576 16120 8628
rect 16172 8616 16178 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16172 8588 16681 8616
rect 16172 8576 16178 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 17034 8576 17040 8628
rect 17092 8616 17098 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17092 8588 17509 8616
rect 17092 8576 17098 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17954 8576 17960 8628
rect 18012 8616 18018 8628
rect 18601 8619 18659 8625
rect 18601 8616 18613 8619
rect 18012 8588 18613 8616
rect 18012 8576 18018 8588
rect 18601 8585 18613 8588
rect 18647 8585 18659 8619
rect 18601 8579 18659 8585
rect 19242 8576 19248 8628
rect 19300 8616 19306 8628
rect 19978 8616 19984 8628
rect 19300 8588 19656 8616
rect 19939 8588 19984 8616
rect 19300 8576 19306 8588
rect 13832 8520 14688 8548
rect 15280 8551 15338 8557
rect 12641 8483 12699 8489
rect 12641 8480 12653 8483
rect 10704 8452 11836 8480
rect 11900 8452 12653 8480
rect 7926 8412 7932 8424
rect 7887 8384 7932 8412
rect 7926 8372 7932 8384
rect 7984 8372 7990 8424
rect 8389 8415 8447 8421
rect 8389 8381 8401 8415
rect 8435 8381 8447 8415
rect 8389 8375 8447 8381
rect 6604 8316 7308 8344
rect 6604 8304 6610 8316
rect 7374 8304 7380 8356
rect 7432 8344 7438 8356
rect 8018 8344 8024 8356
rect 7432 8316 8024 8344
rect 7432 8304 7438 8316
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 8294 8304 8300 8356
rect 8352 8344 8358 8356
rect 8404 8344 8432 8375
rect 8478 8372 8484 8424
rect 8536 8412 8542 8424
rect 9122 8412 9128 8424
rect 8536 8384 8581 8412
rect 9083 8384 9128 8412
rect 8536 8372 8542 8384
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9306 8412 9312 8424
rect 9267 8384 9312 8412
rect 9306 8372 9312 8384
rect 9364 8372 9370 8424
rect 10042 8412 10048 8424
rect 10003 8384 10048 8412
rect 10042 8372 10048 8384
rect 10100 8412 10106 8424
rect 10704 8412 10732 8452
rect 10100 8384 10732 8412
rect 10781 8415 10839 8421
rect 10100 8372 10106 8384
rect 10781 8381 10793 8415
rect 10827 8412 10839 8415
rect 11900 8412 11928 8452
rect 12641 8449 12653 8452
rect 12687 8480 12699 8483
rect 12897 8483 12955 8489
rect 12687 8452 12848 8480
rect 12687 8449 12699 8452
rect 12641 8443 12699 8449
rect 10827 8384 11928 8412
rect 12820 8412 12848 8452
rect 12897 8449 12909 8483
rect 12943 8449 12955 8483
rect 13832 8480 13860 8520
rect 15280 8517 15292 8551
rect 15326 8548 15338 8551
rect 15930 8548 15936 8560
rect 15326 8520 15936 8548
rect 15326 8517 15338 8520
rect 15280 8511 15338 8517
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 16758 8508 16764 8560
rect 16816 8548 16822 8560
rect 17129 8551 17187 8557
rect 17129 8548 17141 8551
rect 16816 8520 17141 8548
rect 16816 8508 16822 8520
rect 17129 8517 17141 8520
rect 17175 8517 17187 8551
rect 17129 8511 17187 8517
rect 18506 8508 18512 8560
rect 18564 8548 18570 8560
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 18564 8520 18705 8548
rect 18564 8508 18570 8520
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 19518 8548 19524 8560
rect 18693 8511 18751 8517
rect 19352 8520 19524 8548
rect 12897 8443 12955 8449
rect 12995 8452 13860 8480
rect 14277 8483 14335 8489
rect 12995 8412 13023 8452
rect 14277 8449 14289 8483
rect 14323 8480 14335 8483
rect 14829 8483 14887 8489
rect 14323 8452 14504 8480
rect 14323 8449 14335 8452
rect 14277 8443 14335 8449
rect 13538 8412 13544 8424
rect 12820 8384 13023 8412
rect 13499 8384 13544 8412
rect 10827 8381 10839 8384
rect 10781 8375 10839 8381
rect 11164 8356 11192 8384
rect 13538 8372 13544 8384
rect 13596 8372 13602 8424
rect 14366 8412 14372 8424
rect 14327 8384 14372 8412
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 14476 8412 14504 8452
rect 14829 8449 14841 8483
rect 14875 8449 14887 8483
rect 17034 8480 17040 8492
rect 14829 8443 14887 8449
rect 16408 8452 16896 8480
rect 16995 8452 17040 8480
rect 14550 8412 14556 8424
rect 14476 8384 14556 8412
rect 14550 8372 14556 8384
rect 14608 8372 14614 8424
rect 14844 8412 14872 8443
rect 15010 8412 15016 8424
rect 14752 8384 14872 8412
rect 14923 8384 15016 8412
rect 10134 8344 10140 8356
rect 8352 8316 10140 8344
rect 8352 8304 8358 8316
rect 10134 8304 10140 8316
rect 10192 8304 10198 8356
rect 10318 8344 10324 8356
rect 10279 8316 10324 8344
rect 10318 8304 10324 8316
rect 10376 8344 10382 8356
rect 10376 8316 10824 8344
rect 10376 8304 10382 8316
rect 4028 8248 5672 8276
rect 4028 8236 4034 8248
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 6012 8285 6224 8294
rect 6012 8279 6239 8285
rect 6012 8276 6193 8279
rect 5776 8266 6193 8276
rect 5776 8248 6040 8266
rect 5776 8236 5782 8248
rect 6181 8245 6193 8266
rect 6227 8245 6239 8279
rect 6181 8239 6239 8245
rect 6457 8279 6515 8285
rect 6457 8245 6469 8279
rect 6503 8276 6515 8279
rect 7190 8276 7196 8288
rect 6503 8248 7196 8276
rect 6503 8245 6515 8248
rect 6457 8239 6515 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7466 8236 7472 8288
rect 7524 8276 7530 8288
rect 10686 8276 10692 8288
rect 7524 8248 10692 8276
rect 7524 8236 7530 8248
rect 10686 8236 10692 8248
rect 10744 8236 10750 8288
rect 10796 8276 10824 8316
rect 10870 8304 10876 8356
rect 10928 8344 10934 8356
rect 11054 8344 11060 8356
rect 10928 8316 11060 8344
rect 10928 8304 10934 8316
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 11146 8304 11152 8356
rect 11204 8304 11210 8356
rect 13262 8304 13268 8356
rect 13320 8344 13326 8356
rect 13446 8344 13452 8356
rect 13320 8316 13452 8344
rect 13320 8304 13326 8316
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 14384 8344 14412 8372
rect 14752 8344 14780 8384
rect 15010 8372 15016 8384
rect 15068 8372 15074 8424
rect 14384 8316 14780 8344
rect 14826 8304 14832 8356
rect 14884 8344 14890 8356
rect 15028 8344 15056 8372
rect 16408 8353 16436 8452
rect 16868 8424 16896 8452
rect 17034 8440 17040 8452
rect 17092 8440 17098 8492
rect 17310 8440 17316 8492
rect 17368 8480 17374 8492
rect 17865 8483 17923 8489
rect 17865 8480 17877 8483
rect 17368 8452 17877 8480
rect 17368 8440 17374 8452
rect 17865 8449 17877 8452
rect 17911 8449 17923 8483
rect 17865 8443 17923 8449
rect 17957 8483 18015 8489
rect 17957 8449 17969 8483
rect 18003 8480 18015 8483
rect 18230 8480 18236 8492
rect 18003 8452 18236 8480
rect 18003 8449 18015 8452
rect 17957 8443 18015 8449
rect 18230 8440 18236 8452
rect 18288 8440 18294 8492
rect 16850 8412 16856 8424
rect 16763 8384 16856 8412
rect 16850 8372 16856 8384
rect 16908 8412 16914 8424
rect 17218 8412 17224 8424
rect 16908 8384 17224 8412
rect 16908 8372 16914 8384
rect 17218 8372 17224 8384
rect 17276 8372 17282 8424
rect 18049 8415 18107 8421
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18506 8412 18512 8424
rect 18467 8384 18512 8412
rect 18049 8375 18107 8381
rect 14884 8316 15056 8344
rect 16393 8347 16451 8353
rect 14884 8304 14890 8316
rect 16393 8313 16405 8347
rect 16439 8313 16451 8347
rect 18064 8344 18092 8375
rect 18506 8372 18512 8384
rect 18564 8372 18570 8424
rect 19352 8421 19380 8520
rect 19518 8508 19524 8520
rect 19576 8508 19582 8560
rect 19628 8548 19656 8588
rect 19978 8576 19984 8588
rect 20036 8576 20042 8628
rect 20947 8619 21005 8625
rect 20947 8616 20959 8619
rect 20088 8588 20959 8616
rect 20088 8548 20116 8588
rect 20947 8585 20959 8588
rect 20993 8585 21005 8619
rect 20947 8579 21005 8585
rect 19628 8520 20116 8548
rect 20533 8551 20591 8557
rect 20533 8517 20545 8551
rect 20579 8548 20591 8551
rect 20714 8548 20720 8560
rect 20579 8520 20720 8548
rect 20579 8517 20591 8520
rect 20533 8511 20591 8517
rect 20714 8508 20720 8520
rect 20772 8508 20778 8560
rect 19610 8480 19616 8492
rect 19571 8452 19616 8480
rect 19610 8440 19616 8452
rect 19668 8440 19674 8492
rect 20346 8440 20352 8492
rect 20404 8480 20410 8492
rect 21266 8480 21272 8492
rect 20404 8452 21272 8480
rect 20404 8440 20410 8452
rect 21266 8440 21272 8452
rect 21324 8440 21330 8492
rect 19337 8415 19395 8421
rect 19337 8381 19349 8415
rect 19383 8381 19395 8415
rect 19518 8412 19524 8424
rect 19479 8384 19524 8412
rect 19337 8375 19395 8381
rect 19518 8372 19524 8384
rect 19576 8372 19582 8424
rect 20162 8372 20168 8424
rect 20220 8412 20226 8424
rect 20257 8415 20315 8421
rect 20257 8412 20269 8415
rect 20220 8384 20269 8412
rect 20220 8372 20226 8384
rect 20257 8381 20269 8384
rect 20303 8381 20315 8415
rect 20714 8412 20720 8424
rect 20675 8384 20720 8412
rect 20257 8375 20315 8381
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 16393 8307 16451 8313
rect 17880 8316 18092 8344
rect 19061 8347 19119 8353
rect 11330 8276 11336 8288
rect 10796 8248 11336 8276
rect 11330 8236 11336 8248
rect 11388 8236 11394 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 12526 8276 12532 8288
rect 11848 8248 12532 8276
rect 11848 8236 11854 8248
rect 12526 8236 12532 8248
rect 12584 8236 12590 8288
rect 12618 8236 12624 8288
rect 12676 8276 12682 8288
rect 12989 8279 13047 8285
rect 12989 8276 13001 8279
rect 12676 8248 13001 8276
rect 12676 8236 12682 8248
rect 12989 8245 13001 8248
rect 13035 8245 13047 8279
rect 12989 8239 13047 8245
rect 13170 8236 13176 8288
rect 13228 8276 13234 8288
rect 15378 8276 15384 8288
rect 13228 8248 15384 8276
rect 13228 8236 13234 8248
rect 15378 8236 15384 8248
rect 15436 8236 15442 8288
rect 15930 8236 15936 8288
rect 15988 8276 15994 8288
rect 17880 8276 17908 8316
rect 19061 8313 19073 8347
rect 19107 8344 19119 8347
rect 20070 8344 20076 8356
rect 19107 8316 20076 8344
rect 19107 8313 19119 8316
rect 19061 8307 19119 8313
rect 20070 8304 20076 8316
rect 20128 8304 20134 8356
rect 15988 8248 17908 8276
rect 15988 8236 15994 8248
rect 18966 8236 18972 8288
rect 19024 8276 19030 8288
rect 20441 8279 20499 8285
rect 20441 8276 20453 8279
rect 19024 8248 20453 8276
rect 19024 8236 19030 8248
rect 20441 8245 20453 8248
rect 20487 8245 20499 8279
rect 20441 8239 20499 8245
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 1946 8072 1952 8084
rect 1811 8044 1952 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 1946 8032 1952 8044
rect 2004 8032 2010 8084
rect 2406 8032 2412 8084
rect 2464 8072 2470 8084
rect 3789 8075 3847 8081
rect 3789 8072 3801 8075
rect 2464 8044 3801 8072
rect 2464 8032 2470 8044
rect 3789 8041 3801 8044
rect 3835 8041 3847 8075
rect 5442 8072 5448 8084
rect 5403 8044 5448 8072
rect 3789 8035 3847 8041
rect 5442 8032 5448 8044
rect 5500 8032 5506 8084
rect 7650 8072 7656 8084
rect 5552 8044 6868 8072
rect 3234 7964 3240 8016
rect 3292 8004 3298 8016
rect 4617 8007 4675 8013
rect 4617 8004 4629 8007
rect 3292 7976 4629 8004
rect 3292 7964 3298 7976
rect 4617 7973 4629 7976
rect 4663 7973 4675 8007
rect 4617 7967 4675 7973
rect 4890 7964 4896 8016
rect 4948 8004 4954 8016
rect 5552 8004 5580 8044
rect 4948 7976 5580 8004
rect 4948 7964 4954 7976
rect 5626 7964 5632 8016
rect 5684 8004 5690 8016
rect 6362 8004 6368 8016
rect 5684 7976 6368 8004
rect 5684 7964 5690 7976
rect 3605 7939 3663 7945
rect 3605 7905 3617 7939
rect 3651 7936 3663 7939
rect 3970 7936 3976 7948
rect 3651 7908 3976 7936
rect 3651 7905 3663 7908
rect 3605 7899 3663 7905
rect 3970 7896 3976 7908
rect 4028 7896 4034 7948
rect 4246 7896 4252 7948
rect 4304 7936 4310 7948
rect 4341 7939 4399 7945
rect 4341 7936 4353 7939
rect 4304 7908 4353 7936
rect 4304 7896 4310 7908
rect 4341 7905 4353 7908
rect 4387 7905 4399 7939
rect 5166 7936 5172 7948
rect 5127 7908 5172 7936
rect 4341 7899 4399 7905
rect 5166 7896 5172 7908
rect 5224 7896 5230 7948
rect 5718 7896 5724 7948
rect 5776 7936 5782 7948
rect 6012 7945 6040 7976
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 6840 7945 6868 8044
rect 7116 8044 7656 8072
rect 5905 7939 5963 7945
rect 5905 7936 5917 7939
rect 5776 7908 5917 7936
rect 5776 7896 5782 7908
rect 5905 7905 5917 7908
rect 5951 7905 5963 7939
rect 5905 7899 5963 7905
rect 5997 7939 6055 7945
rect 5997 7905 6009 7939
rect 6043 7905 6055 7939
rect 5997 7899 6055 7905
rect 6825 7939 6883 7945
rect 6825 7905 6837 7939
rect 6871 7905 6883 7939
rect 7116 7936 7144 8044
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 8662 8072 8668 8084
rect 7760 8044 8668 8072
rect 7374 7964 7380 8016
rect 7432 8004 7438 8016
rect 7760 8004 7788 8044
rect 8662 8032 8668 8044
rect 8720 8032 8726 8084
rect 8757 8075 8815 8081
rect 8757 8041 8769 8075
rect 8803 8072 8815 8075
rect 9306 8072 9312 8084
rect 8803 8044 9312 8072
rect 8803 8041 8815 8044
rect 8757 8035 8815 8041
rect 9306 8032 9312 8044
rect 9364 8032 9370 8084
rect 10134 8032 10140 8084
rect 10192 8072 10198 8084
rect 10321 8075 10379 8081
rect 10321 8072 10333 8075
rect 10192 8044 10333 8072
rect 10192 8032 10198 8044
rect 10321 8041 10333 8044
rect 10367 8041 10379 8075
rect 10321 8035 10379 8041
rect 10689 8075 10747 8081
rect 10689 8041 10701 8075
rect 10735 8072 10747 8075
rect 10778 8072 10784 8084
rect 10735 8044 10784 8072
rect 10735 8041 10747 8044
rect 10689 8035 10747 8041
rect 10778 8032 10784 8044
rect 10836 8032 10842 8084
rect 10870 8032 10876 8084
rect 10928 8072 10934 8084
rect 11606 8072 11612 8084
rect 10928 8044 11612 8072
rect 10928 8032 10934 8044
rect 8570 8004 8576 8016
rect 7432 7976 7788 8004
rect 8137 7976 8576 8004
rect 7432 7964 7438 7976
rect 7285 7939 7343 7945
rect 7285 7936 7297 7939
rect 7116 7908 7297 7936
rect 6825 7899 6883 7905
rect 7285 7905 7297 7908
rect 7331 7905 7343 7939
rect 7285 7899 7343 7905
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7936 7527 7939
rect 8137 7936 8165 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 7515 7908 8165 7936
rect 8205 7939 8263 7945
rect 7515 7905 7527 7908
rect 7469 7899 7527 7905
rect 8205 7905 8217 7939
rect 8251 7936 8263 7939
rect 8294 7936 8300 7948
rect 8251 7908 8300 7936
rect 8251 7905 8263 7908
rect 8205 7899 8263 7905
rect 8294 7896 8300 7908
rect 8352 7896 8358 7948
rect 10980 7945 11008 8044
rect 11606 8032 11612 8044
rect 11664 8032 11670 8084
rect 12434 8072 12440 8084
rect 12395 8044 12440 8072
rect 12434 8032 12440 8044
rect 12492 8072 12498 8084
rect 12710 8072 12716 8084
rect 12492 8044 12716 8072
rect 12492 8032 12498 8044
rect 12710 8032 12716 8044
rect 12768 8032 12774 8084
rect 12802 8032 12808 8084
rect 12860 8072 12866 8084
rect 12860 8044 13685 8072
rect 12860 8032 12866 8044
rect 10965 7939 11023 7945
rect 10965 7905 10977 7939
rect 11011 7905 11023 7939
rect 12526 7936 12532 7948
rect 10965 7899 11023 7905
rect 12176 7908 12532 7936
rect 14 7828 20 7880
rect 72 7868 78 7880
rect 1026 7868 1032 7880
rect 72 7840 1032 7868
rect 72 7828 78 7840
rect 1026 7828 1032 7840
rect 1084 7868 1090 7880
rect 1489 7871 1547 7877
rect 1489 7868 1501 7871
rect 1084 7840 1501 7868
rect 1084 7828 1090 7840
rect 1489 7837 1501 7840
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 1578 7828 1584 7880
rect 1636 7868 1642 7880
rect 2878 7871 2936 7877
rect 2878 7868 2890 7871
rect 1636 7840 2890 7868
rect 1636 7828 1642 7840
rect 2878 7837 2890 7840
rect 2924 7837 2936 7871
rect 2878 7831 2936 7837
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 3237 7871 3295 7877
rect 3237 7837 3249 7871
rect 3283 7868 3295 7871
rect 3510 7868 3516 7880
rect 3283 7840 3516 7868
rect 3283 7837 3295 7840
rect 3237 7831 3295 7837
rect 1670 7800 1676 7812
rect 1631 7772 1676 7800
rect 1670 7760 1676 7772
rect 1728 7760 1734 7812
rect 3160 7800 3188 7831
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4154 7868 4160 7880
rect 4115 7840 4160 7868
rect 4154 7828 4160 7840
rect 4212 7828 4218 7880
rect 5258 7828 5264 7880
rect 5316 7868 5322 7880
rect 5316 7840 6316 7868
rect 5316 7828 5322 7840
rect 3694 7800 3700 7812
rect 3160 7772 3700 7800
rect 3694 7760 3700 7772
rect 3752 7760 3758 7812
rect 4985 7803 5043 7809
rect 4985 7769 4997 7803
rect 5031 7800 5043 7803
rect 5994 7800 6000 7812
rect 5031 7772 6000 7800
rect 5031 7769 5043 7772
rect 4985 7763 5043 7769
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 3421 7735 3479 7741
rect 3421 7701 3433 7735
rect 3467 7732 3479 7735
rect 4062 7732 4068 7744
rect 3467 7704 4068 7732
rect 3467 7701 3479 7704
rect 3421 7695 3479 7701
rect 4062 7692 4068 7704
rect 4120 7692 4126 7744
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4338 7732 4344 7744
rect 4295 7704 4344 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4338 7692 4344 7704
rect 4396 7692 4402 7744
rect 5074 7692 5080 7744
rect 5132 7732 5138 7744
rect 5132 7704 5177 7732
rect 5132 7692 5138 7704
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 6288 7741 6316 7840
rect 6638 7828 6644 7880
rect 6696 7868 6702 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6696 7840 6745 7868
rect 6696 7828 6702 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 8941 7871 8999 7877
rect 7708 7840 8708 7868
rect 7708 7828 7714 7840
rect 6822 7760 6828 7812
rect 6880 7800 6886 7812
rect 8389 7803 8447 7809
rect 8389 7800 8401 7803
rect 6880 7772 7512 7800
rect 6880 7760 6886 7772
rect 7484 7744 7512 7772
rect 7944 7772 8401 7800
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 5776 7704 5825 7732
rect 5776 7692 5782 7704
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 5813 7695 5871 7701
rect 6273 7735 6331 7741
rect 6273 7701 6285 7735
rect 6319 7701 6331 7735
rect 6273 7695 6331 7701
rect 6641 7735 6699 7741
rect 6641 7701 6653 7735
rect 6687 7732 6699 7735
rect 7374 7732 7380 7744
rect 6687 7704 7380 7732
rect 6687 7701 6699 7704
rect 6641 7695 6699 7701
rect 7374 7692 7380 7704
rect 7432 7692 7438 7744
rect 7466 7692 7472 7744
rect 7524 7732 7530 7744
rect 7944 7741 7972 7772
rect 8389 7769 8401 7772
rect 8435 7769 8447 7803
rect 8680 7800 8708 7840
rect 8941 7837 8953 7871
rect 8987 7868 8999 7871
rect 9030 7868 9036 7880
rect 8987 7840 9036 7868
rect 8987 7837 8999 7840
rect 8941 7831 8999 7837
rect 9030 7828 9036 7840
rect 9088 7868 9094 7880
rect 10980 7868 11008 7899
rect 11238 7877 11244 7880
rect 9088 7840 11008 7868
rect 9088 7828 9094 7840
rect 11232 7831 11244 7877
rect 11296 7868 11302 7880
rect 12176 7868 12204 7908
rect 12526 7896 12532 7908
rect 12584 7936 12590 7948
rect 12989 7939 13047 7945
rect 12989 7936 13001 7939
rect 12584 7908 13001 7936
rect 12584 7896 12590 7908
rect 12989 7905 13001 7908
rect 13035 7936 13047 7939
rect 13538 7936 13544 7948
rect 13035 7908 13544 7936
rect 13035 7905 13047 7908
rect 12989 7899 13047 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 12802 7868 12808 7880
rect 11296 7840 12204 7868
rect 12763 7840 12808 7868
rect 11238 7828 11244 7831
rect 11296 7828 11302 7840
rect 12802 7828 12808 7840
rect 12860 7868 12866 7880
rect 13265 7871 13323 7877
rect 13265 7868 13277 7871
rect 12860 7840 13277 7868
rect 12860 7828 12866 7840
rect 13265 7837 13277 7840
rect 13311 7837 13323 7871
rect 13657 7868 13685 8044
rect 13722 8032 13728 8084
rect 13780 8072 13786 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13780 8044 14105 8072
rect 13780 8032 13786 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14093 8035 14151 8041
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 15010 8072 15016 8084
rect 14608 8044 15016 8072
rect 14608 8032 14614 8044
rect 15010 8032 15016 8044
rect 15068 8032 15074 8084
rect 15562 8072 15568 8084
rect 15523 8044 15568 8072
rect 15562 8032 15568 8044
rect 15620 8032 15626 8084
rect 15838 8032 15844 8084
rect 15896 8072 15902 8084
rect 18046 8072 18052 8084
rect 15896 8044 16988 8072
rect 15896 8032 15902 8044
rect 14458 7964 14464 8016
rect 14516 8004 14522 8016
rect 14826 8004 14832 8016
rect 14516 7976 14832 8004
rect 14516 7964 14522 7976
rect 14826 7964 14832 7976
rect 14884 7964 14890 8016
rect 15473 8007 15531 8013
rect 15473 7973 15485 8007
rect 15519 7973 15531 8007
rect 15473 7967 15531 7973
rect 13906 7896 13912 7948
rect 13964 7936 13970 7948
rect 14366 7936 14372 7948
rect 13964 7908 14372 7936
rect 13964 7896 13970 7908
rect 14366 7896 14372 7908
rect 14424 7936 14430 7948
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14424 7908 14657 7936
rect 14424 7896 14430 7908
rect 14645 7905 14657 7908
rect 14691 7905 14703 7939
rect 15488 7936 15516 7967
rect 15838 7936 15844 7948
rect 15488 7908 15844 7936
rect 14645 7899 14703 7905
rect 15838 7896 15844 7908
rect 15896 7896 15902 7948
rect 16960 7945 16988 8044
rect 17696 8044 18052 8072
rect 17589 8007 17647 8013
rect 17589 7973 17601 8007
rect 17635 7973 17647 8007
rect 17589 7967 17647 7973
rect 16945 7939 17003 7945
rect 16945 7905 16957 7939
rect 16991 7905 17003 7939
rect 16945 7899 17003 7905
rect 17221 7939 17279 7945
rect 17221 7905 17233 7939
rect 17267 7936 17279 7939
rect 17310 7936 17316 7948
rect 17267 7908 17316 7936
rect 17267 7905 17279 7908
rect 17221 7899 17279 7905
rect 17310 7896 17316 7908
rect 17368 7896 17374 7948
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 13657 7840 14473 7868
rect 13265 7831 13323 7837
rect 14461 7837 14473 7840
rect 14507 7868 14519 7871
rect 15105 7871 15163 7877
rect 15105 7868 15117 7871
rect 14507 7840 15117 7868
rect 14507 7837 14519 7840
rect 14461 7831 14519 7837
rect 15105 7837 15117 7840
rect 15151 7837 15163 7871
rect 15105 7831 15163 7837
rect 15289 7871 15347 7877
rect 15289 7837 15301 7871
rect 15335 7837 15347 7871
rect 15289 7831 15347 7837
rect 9186 7803 9244 7809
rect 9186 7800 9198 7803
rect 8680 7772 9198 7800
rect 8389 7763 8447 7769
rect 9186 7769 9198 7772
rect 9232 7800 9244 7803
rect 9582 7800 9588 7812
rect 9232 7772 9588 7800
rect 9232 7769 9244 7772
rect 9186 7763 9244 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 9858 7760 9864 7812
rect 9916 7800 9922 7812
rect 10134 7800 10140 7812
rect 9916 7772 10140 7800
rect 9916 7760 9922 7772
rect 10134 7760 10140 7772
rect 10192 7760 10198 7812
rect 10505 7803 10563 7809
rect 10505 7769 10517 7803
rect 10551 7800 10563 7803
rect 10686 7800 10692 7812
rect 10551 7772 10692 7800
rect 10551 7769 10563 7772
rect 10505 7763 10563 7769
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 12250 7760 12256 7812
rect 12308 7800 12314 7812
rect 12618 7800 12624 7812
rect 12308 7772 12624 7800
rect 12308 7760 12314 7772
rect 12618 7760 12624 7772
rect 12676 7760 12682 7812
rect 13078 7760 13084 7812
rect 13136 7760 13142 7812
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13725 7803 13783 7809
rect 13725 7800 13737 7803
rect 13228 7772 13273 7800
rect 13464 7772 13737 7800
rect 13228 7760 13234 7772
rect 7561 7735 7619 7741
rect 7561 7732 7573 7735
rect 7524 7704 7573 7732
rect 7524 7692 7530 7704
rect 7561 7701 7573 7704
rect 7607 7701 7619 7735
rect 7561 7695 7619 7701
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7701 7987 7735
rect 8294 7732 8300 7744
rect 8255 7704 8300 7732
rect 7929 7695 7987 7701
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8570 7692 8576 7744
rect 8628 7732 8634 7744
rect 9306 7732 9312 7744
rect 8628 7704 9312 7732
rect 8628 7692 8634 7704
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 10410 7732 10416 7744
rect 9548 7704 10416 7732
rect 9548 7692 9554 7704
rect 10410 7692 10416 7704
rect 10468 7692 10474 7744
rect 10870 7732 10876 7744
rect 10831 7704 10876 7732
rect 10870 7692 10876 7704
rect 10928 7732 10934 7744
rect 11882 7732 11888 7744
rect 10928 7704 11888 7732
rect 10928 7692 10934 7704
rect 11882 7692 11888 7704
rect 11940 7692 11946 7744
rect 12342 7732 12348 7744
rect 12303 7704 12348 7732
rect 12342 7692 12348 7704
rect 12400 7692 12406 7744
rect 13096 7732 13124 7760
rect 13464 7732 13492 7772
rect 13725 7769 13737 7772
rect 13771 7769 13783 7803
rect 13725 7763 13783 7769
rect 13096 7704 13492 7732
rect 13538 7692 13544 7744
rect 13596 7732 13602 7744
rect 13633 7735 13691 7741
rect 13633 7732 13645 7735
rect 13596 7704 13645 7732
rect 13596 7692 13602 7704
rect 13633 7701 13645 7704
rect 13679 7701 13691 7735
rect 13633 7695 13691 7701
rect 14553 7735 14611 7741
rect 14553 7701 14565 7735
rect 14599 7732 14611 7735
rect 14826 7732 14832 7744
rect 14599 7704 14832 7732
rect 14599 7701 14611 7704
rect 14553 7695 14611 7701
rect 14826 7692 14832 7704
rect 14884 7732 14890 7744
rect 14921 7735 14979 7741
rect 14921 7732 14933 7735
rect 14884 7704 14933 7732
rect 14884 7692 14890 7704
rect 14921 7701 14933 7704
rect 14967 7701 14979 7735
rect 15120 7732 15148 7831
rect 15304 7800 15332 7831
rect 15378 7828 15384 7880
rect 15436 7868 15442 7880
rect 16206 7868 16212 7880
rect 15436 7840 16212 7868
rect 15436 7828 15442 7840
rect 16206 7828 16212 7840
rect 16264 7828 16270 7880
rect 16678 7871 16736 7877
rect 16678 7837 16690 7871
rect 16724 7868 16736 7871
rect 16850 7868 16856 7880
rect 16724 7840 16856 7868
rect 16724 7837 16736 7840
rect 16678 7831 16736 7837
rect 16850 7828 16856 7840
rect 16908 7828 16914 7880
rect 17402 7868 17408 7880
rect 17363 7840 17408 7868
rect 17402 7828 17408 7840
rect 17460 7828 17466 7880
rect 17604 7868 17632 7967
rect 17696 7945 17724 8044
rect 18046 8032 18052 8044
rect 18104 8032 18110 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19981 8075 20039 8081
rect 19981 8072 19993 8075
rect 19576 8044 19993 8072
rect 19576 8032 19582 8044
rect 19981 8041 19993 8044
rect 20027 8041 20039 8075
rect 21358 8072 21364 8084
rect 21319 8044 21364 8072
rect 19981 8035 20039 8041
rect 21358 8032 21364 8044
rect 21416 8032 21422 8084
rect 19061 8007 19119 8013
rect 19061 7973 19073 8007
rect 19107 8004 19119 8007
rect 19794 8004 19800 8016
rect 19107 7976 19800 8004
rect 19107 7973 19119 7976
rect 19061 7967 19119 7973
rect 19444 7945 19472 7976
rect 19794 7964 19800 7976
rect 19852 7964 19858 8016
rect 17681 7939 17739 7945
rect 17681 7905 17693 7939
rect 17727 7905 17739 7939
rect 17681 7899 17739 7905
rect 19429 7939 19487 7945
rect 19429 7905 19441 7939
rect 19475 7905 19487 7939
rect 19429 7899 19487 7905
rect 19521 7939 19579 7945
rect 19521 7905 19533 7939
rect 19567 7936 19579 7939
rect 19702 7936 19708 7948
rect 19567 7908 19708 7936
rect 19567 7905 19579 7908
rect 19521 7899 19579 7905
rect 19702 7896 19708 7908
rect 19760 7896 19766 7948
rect 19886 7896 19892 7948
rect 19944 7936 19950 7948
rect 20165 7939 20223 7945
rect 20165 7936 20177 7939
rect 19944 7908 20177 7936
rect 19944 7896 19950 7908
rect 20165 7905 20177 7908
rect 20211 7936 20223 7939
rect 21358 7936 21364 7948
rect 20211 7908 21364 7936
rect 20211 7905 20223 7908
rect 20165 7899 20223 7905
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 19978 7868 19984 7880
rect 17604 7840 19984 7868
rect 19978 7828 19984 7840
rect 20036 7828 20042 7880
rect 20441 7871 20499 7877
rect 20441 7868 20453 7871
rect 20088 7840 20453 7868
rect 15746 7800 15752 7812
rect 15304 7772 15752 7800
rect 15746 7760 15752 7772
rect 15804 7800 15810 7812
rect 16942 7800 16948 7812
rect 15804 7772 16948 7800
rect 15804 7760 15810 7772
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 17948 7803 18006 7809
rect 17948 7769 17960 7803
rect 17994 7800 18006 7803
rect 18506 7800 18512 7812
rect 17994 7772 18512 7800
rect 17994 7769 18006 7772
rect 17948 7763 18006 7769
rect 18506 7760 18512 7772
rect 18564 7800 18570 7812
rect 18966 7800 18972 7812
rect 18564 7772 18972 7800
rect 18564 7760 18570 7772
rect 18966 7760 18972 7772
rect 19024 7800 19030 7812
rect 20088 7800 20116 7840
rect 20441 7837 20453 7840
rect 20487 7837 20499 7871
rect 20441 7831 20499 7837
rect 20530 7828 20536 7880
rect 20588 7868 20594 7880
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 20588 7840 21465 7868
rect 20588 7828 20594 7840
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21453 7831 21511 7837
rect 19024 7772 20116 7800
rect 19024 7760 19030 7772
rect 20714 7760 20720 7812
rect 20772 7800 20778 7812
rect 21085 7803 21143 7809
rect 21085 7800 21097 7803
rect 20772 7772 21097 7800
rect 20772 7760 20778 7772
rect 21085 7769 21097 7772
rect 21131 7769 21143 7803
rect 21085 7763 21143 7769
rect 15470 7732 15476 7744
rect 15120 7704 15476 7732
rect 14921 7695 14979 7701
rect 15470 7692 15476 7704
rect 15528 7692 15534 7744
rect 16206 7692 16212 7744
rect 16264 7732 16270 7744
rect 18230 7732 18236 7744
rect 16264 7704 18236 7732
rect 16264 7692 16270 7704
rect 18230 7692 18236 7704
rect 18288 7692 18294 7744
rect 19150 7692 19156 7744
rect 19208 7732 19214 7744
rect 19613 7735 19671 7741
rect 19613 7732 19625 7735
rect 19208 7704 19625 7732
rect 19208 7692 19214 7704
rect 19613 7701 19625 7704
rect 19659 7701 19671 7735
rect 19613 7695 19671 7701
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 750 7488 756 7540
rect 808 7528 814 7540
rect 2958 7528 2964 7540
rect 808 7500 2964 7528
rect 808 7488 814 7500
rect 2958 7488 2964 7500
rect 3016 7488 3022 7540
rect 5166 7528 5172 7540
rect 3160 7500 5172 7528
rect 1486 7460 1492 7472
rect 1447 7432 1492 7460
rect 1486 7420 1492 7432
rect 1544 7420 1550 7472
rect 2958 7352 2964 7404
rect 3016 7401 3022 7404
rect 3016 7392 3028 7401
rect 3160 7392 3188 7500
rect 5166 7488 5172 7500
rect 5224 7528 5230 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 5224 7500 5365 7528
rect 5224 7488 5230 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5859 7500 6377 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 6733 7531 6791 7537
rect 6733 7497 6745 7531
rect 6779 7528 6791 7531
rect 7282 7528 7288 7540
rect 6779 7500 7288 7528
rect 6779 7497 6791 7500
rect 6733 7491 6791 7497
rect 7282 7488 7288 7500
rect 7340 7488 7346 7540
rect 7650 7528 7656 7540
rect 7611 7500 7656 7528
rect 7650 7488 7656 7500
rect 7708 7488 7714 7540
rect 8386 7488 8392 7540
rect 8444 7488 8450 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8536 7500 9137 7528
rect 8536 7488 8542 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9125 7491 9183 7497
rect 9585 7531 9643 7537
rect 9585 7497 9597 7531
rect 9631 7528 9643 7531
rect 10045 7531 10103 7537
rect 10045 7528 10057 7531
rect 9631 7500 10057 7528
rect 9631 7497 9643 7500
rect 9585 7491 9643 7497
rect 10045 7497 10057 7500
rect 10091 7528 10103 7531
rect 10226 7528 10232 7540
rect 10091 7500 10232 7528
rect 10091 7497 10103 7500
rect 10045 7491 10103 7497
rect 10226 7488 10232 7500
rect 10284 7488 10290 7540
rect 10873 7531 10931 7537
rect 10873 7497 10885 7531
rect 10919 7528 10931 7531
rect 11609 7531 11667 7537
rect 11609 7528 11621 7531
rect 10919 7500 11621 7528
rect 10919 7497 10931 7500
rect 10873 7491 10931 7497
rect 11609 7497 11621 7500
rect 11655 7497 11667 7531
rect 11974 7528 11980 7540
rect 11935 7500 11980 7528
rect 11609 7491 11667 7497
rect 11974 7488 11980 7500
rect 12032 7488 12038 7540
rect 12069 7531 12127 7537
rect 12069 7497 12081 7531
rect 12115 7528 12127 7531
rect 12250 7528 12256 7540
rect 12115 7500 12256 7528
rect 12115 7497 12127 7500
rect 12069 7491 12127 7497
rect 12250 7488 12256 7500
rect 12308 7488 12314 7540
rect 12710 7528 12716 7540
rect 12671 7500 12716 7528
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7528 12863 7531
rect 13078 7528 13084 7540
rect 12851 7500 13084 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 13078 7488 13084 7500
rect 13136 7488 13142 7540
rect 13170 7488 13176 7540
rect 13228 7528 13234 7540
rect 13265 7531 13323 7537
rect 13265 7528 13277 7531
rect 13228 7500 13277 7528
rect 13228 7488 13234 7500
rect 13265 7497 13277 7500
rect 13311 7497 13323 7531
rect 13630 7528 13636 7540
rect 13591 7500 13636 7528
rect 13265 7491 13323 7497
rect 13630 7488 13636 7500
rect 13688 7488 13694 7540
rect 13725 7531 13783 7537
rect 13725 7497 13737 7531
rect 13771 7528 13783 7531
rect 13814 7528 13820 7540
rect 13771 7500 13820 7528
rect 13771 7497 13783 7500
rect 13725 7491 13783 7497
rect 5905 7463 5963 7469
rect 5905 7429 5917 7463
rect 5951 7460 5963 7463
rect 6178 7460 6184 7472
rect 5951 7432 6184 7460
rect 5951 7429 5963 7432
rect 5905 7423 5963 7429
rect 6178 7420 6184 7432
rect 6236 7420 6242 7472
rect 6454 7420 6460 7472
rect 6512 7460 6518 7472
rect 6638 7460 6644 7472
rect 6512 7432 6644 7460
rect 6512 7420 6518 7432
rect 6638 7420 6644 7432
rect 6696 7420 6702 7472
rect 6822 7460 6828 7472
rect 6783 7432 6828 7460
rect 6822 7420 6828 7432
rect 6880 7420 6886 7472
rect 8404 7460 8432 7488
rect 7576 7432 9076 7460
rect 3016 7364 3188 7392
rect 3237 7395 3295 7401
rect 3016 7355 3028 7364
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3694 7392 3700 7404
rect 3283 7364 3700 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3016 7352 3022 7355
rect 3694 7352 3700 7364
rect 3752 7352 3758 7404
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 3973 7395 4031 7401
rect 3973 7392 3985 7395
rect 3927 7364 3985 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 3973 7361 3985 7364
rect 4019 7392 4031 7395
rect 4062 7392 4068 7404
rect 4019 7364 4068 7392
rect 4019 7361 4031 7364
rect 3973 7355 4031 7361
rect 4062 7352 4068 7364
rect 4120 7352 4126 7404
rect 4246 7401 4252 7404
rect 4240 7392 4252 7401
rect 4207 7364 4252 7392
rect 4240 7355 4252 7364
rect 4246 7352 4252 7355
rect 4304 7352 4310 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5166 7352 5172 7404
rect 5224 7392 5230 7404
rect 5981 7392 6123 7396
rect 5224 7368 6123 7392
rect 5224 7364 6009 7368
rect 5224 7352 5230 7364
rect 3326 7284 3332 7336
rect 3384 7324 3390 7336
rect 3384 7296 3429 7324
rect 3384 7284 3390 7296
rect 3602 7284 3608 7336
rect 3660 7284 3666 7336
rect 1673 7259 1731 7265
rect 1673 7225 1685 7259
rect 1719 7256 1731 7259
rect 1719 7228 2360 7256
rect 1719 7225 1731 7228
rect 1673 7219 1731 7225
rect 1578 7148 1584 7200
rect 1636 7188 1642 7200
rect 1857 7191 1915 7197
rect 1857 7188 1869 7191
rect 1636 7160 1869 7188
rect 1636 7148 1642 7160
rect 1857 7157 1869 7160
rect 1903 7157 1915 7191
rect 2332 7188 2360 7228
rect 3620 7188 3648 7284
rect 3712 7197 3740 7352
rect 5000 7324 5028 7352
rect 5997 7327 6055 7333
rect 5000 7296 5856 7324
rect 4982 7216 4988 7268
rect 5040 7256 5046 7268
rect 5445 7259 5503 7265
rect 5445 7256 5457 7259
rect 5040 7228 5457 7256
rect 5040 7216 5046 7228
rect 5445 7225 5457 7228
rect 5491 7225 5503 7259
rect 5828 7256 5856 7296
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6095 7324 6123 7368
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 7466 7392 7472 7404
rect 7331 7364 7472 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 7466 7352 7472 7364
rect 7524 7352 7530 7404
rect 7576 7401 7604 7432
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 8386 7352 8392 7404
rect 8444 7392 8450 7404
rect 9048 7401 9076 7432
rect 9306 7420 9312 7472
rect 9364 7460 9370 7472
rect 9493 7463 9551 7469
rect 9493 7460 9505 7463
rect 9364 7432 9505 7460
rect 9364 7420 9370 7432
rect 9493 7429 9505 7432
rect 9539 7460 9551 7463
rect 10594 7460 10600 7472
rect 9539 7432 10600 7460
rect 9539 7429 9551 7432
rect 9493 7423 9551 7429
rect 10594 7420 10600 7432
rect 10652 7420 10658 7472
rect 12728 7460 12756 7488
rect 12728 7432 13124 7460
rect 13096 7404 13124 7432
rect 8766 7395 8824 7401
rect 8766 7392 8778 7395
rect 8444 7364 8778 7392
rect 8444 7352 8450 7364
rect 8766 7361 8778 7364
rect 8812 7361 8824 7395
rect 8766 7355 8824 7361
rect 9033 7395 9091 7401
rect 9033 7361 9045 7395
rect 9079 7392 9091 7395
rect 9122 7392 9128 7404
rect 9079 7364 9128 7392
rect 9079 7361 9091 7364
rect 9033 7355 9091 7361
rect 9122 7352 9128 7364
rect 9180 7352 9186 7404
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7392 11023 7395
rect 12894 7392 12900 7404
rect 11011 7364 12664 7392
rect 11011 7361 11023 7364
rect 10965 7355 11023 7361
rect 6043 7296 6123 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6638 7284 6644 7336
rect 6696 7324 6702 7336
rect 6917 7327 6975 7333
rect 6917 7324 6929 7327
rect 6696 7296 6929 7324
rect 6696 7284 6702 7296
rect 6917 7293 6929 7296
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9640 7296 9689 7324
rect 9640 7284 9646 7296
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 10226 7324 10232 7336
rect 10187 7296 10232 7324
rect 9677 7287 9735 7293
rect 10226 7284 10232 7296
rect 10284 7284 10290 7336
rect 10781 7327 10839 7333
rect 10781 7293 10793 7327
rect 10827 7324 10839 7327
rect 11790 7324 11796 7336
rect 10827 7296 11796 7324
rect 10827 7293 10839 7296
rect 10781 7287 10839 7293
rect 11790 7284 11796 7296
rect 11848 7284 11854 7336
rect 12253 7327 12311 7333
rect 12253 7293 12265 7327
rect 12299 7324 12311 7327
rect 12342 7324 12348 7336
rect 12299 7296 12348 7324
rect 12299 7293 12311 7296
rect 12253 7287 12311 7293
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12526 7324 12532 7336
rect 12487 7296 12532 7324
rect 12526 7284 12532 7296
rect 12584 7284 12590 7336
rect 5828 7228 7788 7256
rect 5445 7219 5503 7225
rect 2332 7160 3648 7188
rect 3697 7191 3755 7197
rect 1857 7151 1915 7157
rect 3697 7157 3709 7191
rect 3743 7188 3755 7191
rect 3970 7188 3976 7200
rect 3743 7160 3976 7188
rect 3743 7157 3755 7160
rect 3697 7151 3755 7157
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 6914 7188 6920 7200
rect 4396 7160 6920 7188
rect 4396 7148 4402 7160
rect 6914 7148 6920 7160
rect 6972 7148 6978 7200
rect 7377 7191 7435 7197
rect 7377 7157 7389 7191
rect 7423 7188 7435 7191
rect 7650 7188 7656 7200
rect 7423 7160 7656 7188
rect 7423 7157 7435 7160
rect 7377 7151 7435 7157
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 7760 7188 7788 7228
rect 10870 7216 10876 7268
rect 10928 7256 10934 7268
rect 10928 7228 12572 7256
rect 10928 7216 10934 7228
rect 12544 7200 12572 7228
rect 9306 7188 9312 7200
rect 7760 7160 9312 7188
rect 9306 7148 9312 7160
rect 9364 7148 9370 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10594 7188 10600 7200
rect 10192 7160 10600 7188
rect 10192 7148 10198 7160
rect 10594 7148 10600 7160
rect 10652 7148 10658 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11204 7160 11345 7188
rect 11204 7148 11210 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11333 7151 11391 7157
rect 12526 7148 12532 7200
rect 12584 7148 12590 7200
rect 12636 7188 12664 7364
rect 12728 7364 12900 7392
rect 12728 7268 12756 7364
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 13078 7352 13084 7404
rect 13136 7352 13142 7404
rect 13630 7352 13636 7404
rect 13688 7392 13694 7404
rect 13740 7392 13768 7491
rect 13814 7488 13820 7500
rect 13872 7528 13878 7540
rect 14093 7531 14151 7537
rect 14093 7528 14105 7531
rect 13872 7500 14105 7528
rect 13872 7488 13878 7500
rect 14093 7497 14105 7500
rect 14139 7497 14151 7531
rect 14093 7491 14151 7497
rect 15102 7488 15108 7540
rect 15160 7528 15166 7540
rect 15565 7531 15623 7537
rect 15565 7528 15577 7531
rect 15160 7500 15577 7528
rect 15160 7488 15166 7500
rect 15565 7497 15577 7500
rect 15611 7497 15623 7531
rect 16022 7528 16028 7540
rect 15983 7500 16028 7528
rect 15565 7491 15623 7497
rect 16022 7488 16028 7500
rect 16080 7488 16086 7540
rect 16298 7488 16304 7540
rect 16356 7528 16362 7540
rect 16356 7500 16436 7528
rect 16356 7488 16362 7500
rect 15378 7460 15384 7472
rect 13688 7364 13768 7392
rect 14108 7432 15384 7460
rect 13688 7352 13694 7364
rect 13354 7284 13360 7336
rect 13412 7284 13418 7336
rect 13906 7324 13912 7336
rect 13867 7296 13912 7324
rect 13906 7284 13912 7296
rect 13964 7284 13970 7336
rect 12710 7216 12716 7268
rect 12768 7216 12774 7268
rect 13372 7200 13400 7284
rect 13722 7216 13728 7268
rect 13780 7256 13786 7268
rect 14108 7256 14136 7432
rect 14458 7392 14464 7404
rect 14419 7364 14464 7392
rect 14458 7352 14464 7364
rect 14516 7352 14522 7404
rect 14553 7395 14611 7401
rect 14553 7361 14565 7395
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 14274 7256 14280 7268
rect 13780 7228 14136 7256
rect 14187 7228 14280 7256
rect 13780 7216 13786 7228
rect 14274 7216 14280 7228
rect 14332 7256 14338 7268
rect 14568 7256 14596 7355
rect 14826 7352 14832 7404
rect 14884 7352 14890 7404
rect 15194 7392 15200 7404
rect 15155 7364 15200 7392
rect 15194 7352 15200 7364
rect 15252 7352 15258 7404
rect 14332 7228 14596 7256
rect 14332 7216 14338 7228
rect 12986 7188 12992 7200
rect 12636 7160 12992 7188
rect 12986 7148 12992 7160
rect 13044 7148 13050 7200
rect 13170 7188 13176 7200
rect 13131 7160 13176 7188
rect 13170 7148 13176 7160
rect 13228 7148 13234 7200
rect 13354 7148 13360 7200
rect 13412 7148 13418 7200
rect 14734 7188 14740 7200
rect 14695 7160 14740 7188
rect 14734 7148 14740 7160
rect 14792 7148 14798 7200
rect 14844 7188 14872 7352
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7293 15071 7327
rect 15013 7287 15071 7293
rect 15105 7327 15163 7333
rect 15105 7293 15117 7327
rect 15151 7324 15163 7327
rect 15295 7324 15323 7432
rect 15378 7420 15384 7432
rect 15436 7420 15442 7472
rect 15746 7392 15752 7404
rect 15707 7364 15752 7392
rect 15746 7352 15752 7364
rect 15804 7352 15810 7404
rect 16206 7352 16212 7404
rect 16264 7392 16270 7404
rect 16408 7392 16436 7500
rect 17034 7488 17040 7540
rect 17092 7528 17098 7540
rect 17221 7531 17279 7537
rect 17221 7528 17233 7531
rect 17092 7500 17233 7528
rect 17092 7488 17098 7500
rect 17221 7497 17233 7500
rect 17267 7497 17279 7531
rect 17221 7491 17279 7497
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18325 7531 18383 7537
rect 18325 7528 18337 7531
rect 18012 7500 18337 7528
rect 18012 7488 18018 7500
rect 18325 7497 18337 7500
rect 18371 7497 18383 7531
rect 18325 7491 18383 7497
rect 18785 7531 18843 7537
rect 18785 7497 18797 7531
rect 18831 7528 18843 7531
rect 19150 7528 19156 7540
rect 18831 7500 19156 7528
rect 18831 7497 18843 7500
rect 18785 7491 18843 7497
rect 19150 7488 19156 7500
rect 19208 7488 19214 7540
rect 19242 7488 19248 7540
rect 19300 7528 19306 7540
rect 19300 7500 19345 7528
rect 19300 7488 19306 7500
rect 19610 7488 19616 7540
rect 19668 7528 19674 7540
rect 19705 7531 19763 7537
rect 19705 7528 19717 7531
rect 19668 7500 19717 7528
rect 19668 7488 19674 7500
rect 19705 7497 19717 7500
rect 19751 7497 19763 7531
rect 19705 7491 19763 7497
rect 20070 7488 20076 7540
rect 20128 7528 20134 7540
rect 20165 7531 20223 7537
rect 20165 7528 20177 7531
rect 20128 7500 20177 7528
rect 20128 7488 20134 7500
rect 20165 7497 20177 7500
rect 20211 7497 20223 7531
rect 20806 7528 20812 7540
rect 20767 7500 20812 7528
rect 20165 7491 20223 7497
rect 20806 7488 20812 7500
rect 20864 7488 20870 7540
rect 20898 7488 20904 7540
rect 20956 7488 20962 7540
rect 21082 7488 21088 7540
rect 21140 7528 21146 7540
rect 21269 7531 21327 7537
rect 21269 7528 21281 7531
rect 21140 7500 21281 7528
rect 21140 7488 21146 7500
rect 21269 7497 21281 7500
rect 21315 7497 21327 7531
rect 21269 7491 21327 7497
rect 21358 7488 21364 7540
rect 21416 7528 21422 7540
rect 21416 7500 21461 7528
rect 21416 7488 21422 7500
rect 16574 7420 16580 7472
rect 16632 7460 16638 7472
rect 16632 7432 17632 7460
rect 16632 7420 16638 7432
rect 17604 7404 17632 7432
rect 17770 7420 17776 7472
rect 17828 7460 17834 7472
rect 19058 7460 19064 7472
rect 17828 7432 19064 7460
rect 17828 7420 17834 7432
rect 19058 7420 19064 7432
rect 19116 7460 19122 7472
rect 20530 7460 20536 7472
rect 19116 7432 20536 7460
rect 19116 7420 19122 7432
rect 20530 7420 20536 7432
rect 20588 7420 20594 7472
rect 20916 7460 20944 7488
rect 20732 7432 20944 7460
rect 16485 7395 16543 7401
rect 16485 7392 16497 7395
rect 16264 7364 16309 7392
rect 16408 7364 16497 7392
rect 16264 7352 16270 7364
rect 16485 7361 16497 7364
rect 16531 7361 16543 7395
rect 16666 7392 16672 7404
rect 16627 7364 16672 7392
rect 16485 7355 16543 7361
rect 16666 7352 16672 7364
rect 16724 7352 16730 7404
rect 16945 7395 17003 7401
rect 16945 7361 16957 7395
rect 16991 7392 17003 7395
rect 17218 7392 17224 7404
rect 16991 7364 17224 7392
rect 16991 7361 17003 7364
rect 16945 7355 17003 7361
rect 17218 7352 17224 7364
rect 17276 7352 17282 7404
rect 17586 7392 17592 7404
rect 17547 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7352 17650 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 18417 7395 18475 7401
rect 17727 7364 18184 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 15151 7296 15323 7324
rect 15151 7293 15163 7296
rect 15105 7287 15163 7293
rect 15028 7256 15056 7287
rect 15930 7284 15936 7336
rect 15988 7324 15994 7336
rect 17773 7327 17831 7333
rect 17773 7324 17785 7327
rect 15988 7296 17785 7324
rect 15988 7284 15994 7296
rect 17773 7293 17785 7296
rect 17819 7293 17831 7327
rect 17773 7287 17831 7293
rect 15948 7256 15976 7284
rect 15028 7228 15976 7256
rect 16206 7216 16212 7268
rect 16264 7216 16270 7268
rect 16853 7259 16911 7265
rect 16853 7225 16865 7259
rect 16899 7256 16911 7259
rect 17310 7256 17316 7268
rect 16899 7228 17316 7256
rect 16899 7225 16911 7228
rect 16853 7219 16911 7225
rect 17310 7216 17316 7228
rect 17368 7216 17374 7268
rect 17402 7216 17408 7268
rect 17460 7256 17466 7268
rect 18156 7256 18184 7364
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 18506 7392 18512 7404
rect 18463 7364 18512 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 18506 7352 18512 7364
rect 18564 7352 18570 7404
rect 20070 7392 20076 7404
rect 20031 7364 20076 7392
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 18233 7327 18291 7333
rect 18233 7293 18245 7327
rect 18279 7324 18291 7327
rect 18966 7324 18972 7336
rect 18279 7296 18972 7324
rect 18279 7293 18291 7296
rect 18233 7287 18291 7293
rect 18966 7284 18972 7296
rect 19024 7284 19030 7336
rect 19058 7284 19064 7336
rect 19116 7324 19122 7336
rect 19153 7327 19211 7333
rect 19153 7324 19165 7327
rect 19116 7296 19165 7324
rect 19116 7284 19122 7296
rect 19153 7293 19165 7296
rect 19199 7293 19211 7327
rect 19153 7287 19211 7293
rect 19794 7284 19800 7336
rect 19852 7324 19858 7336
rect 20257 7327 20315 7333
rect 20257 7324 20269 7327
rect 19852 7296 20269 7324
rect 19852 7284 19858 7296
rect 20257 7293 20269 7296
rect 20303 7324 20315 7327
rect 20625 7327 20683 7333
rect 20625 7324 20637 7327
rect 20303 7296 20637 7324
rect 20303 7293 20315 7296
rect 20257 7287 20315 7293
rect 20625 7293 20637 7296
rect 20671 7293 20683 7327
rect 20625 7287 20683 7293
rect 19702 7256 19708 7268
rect 17460 7228 19708 7256
rect 17460 7216 17466 7228
rect 19702 7216 19708 7228
rect 19760 7256 19766 7268
rect 20732 7256 20760 7432
rect 20898 7392 20904 7404
rect 20859 7364 20904 7392
rect 20898 7352 20904 7364
rect 20956 7352 20962 7404
rect 21542 7392 21548 7404
rect 21503 7364 21548 7392
rect 21542 7352 21548 7364
rect 21600 7352 21606 7404
rect 19760 7228 20760 7256
rect 19760 7216 19766 7228
rect 15102 7188 15108 7200
rect 14844 7160 15108 7188
rect 15102 7148 15108 7160
rect 15160 7148 15166 7200
rect 15930 7188 15936 7200
rect 15891 7160 15936 7188
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16224 7188 16252 7216
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 16224 7160 16313 7188
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 16482 7148 16488 7200
rect 16540 7188 16546 7200
rect 16574 7188 16580 7200
rect 16540 7160 16580 7188
rect 16540 7148 16546 7160
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 17129 7191 17187 7197
rect 17129 7157 17141 7191
rect 17175 7188 17187 7191
rect 17862 7188 17868 7200
rect 17175 7160 17868 7188
rect 17175 7157 17187 7160
rect 17129 7151 17187 7157
rect 17862 7148 17868 7160
rect 17920 7148 17926 7200
rect 19610 7188 19616 7200
rect 19571 7160 19616 7188
rect 19610 7148 19616 7160
rect 19668 7148 19674 7200
rect 19978 7148 19984 7200
rect 20036 7188 20042 7200
rect 20806 7188 20812 7200
rect 20036 7160 20812 7188
rect 20036 7148 20042 7160
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 21726 7148 21732 7200
rect 21784 7188 21790 7200
rect 22002 7188 22008 7200
rect 21784 7160 22008 7188
rect 21784 7148 21790 7160
rect 22002 7148 22008 7160
rect 22060 7148 22066 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 22002 7012 22008 7064
rect 22060 7052 22066 7064
rect 22370 7052 22376 7064
rect 22060 7024 22376 7052
rect 22060 7012 22066 7024
rect 22370 7012 22376 7024
rect 22428 7012 22434 7064
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4120 6956 7236 6984
rect 4120 6944 4126 6956
rect 2869 6919 2927 6925
rect 2869 6916 2881 6919
rect 2332 6888 2881 6916
rect 1026 6808 1032 6860
rect 1084 6848 1090 6860
rect 1084 6820 1808 6848
rect 1084 6808 1090 6820
rect 1302 6740 1308 6792
rect 1360 6780 1366 6792
rect 1780 6789 1808 6820
rect 1946 6808 1952 6860
rect 2004 6848 2010 6860
rect 2332 6857 2360 6888
rect 2869 6885 2881 6888
rect 2915 6885 2927 6919
rect 4890 6916 4896 6928
rect 2869 6879 2927 6885
rect 2976 6888 4896 6916
rect 2133 6851 2191 6857
rect 2133 6848 2145 6851
rect 2004 6820 2145 6848
rect 2004 6808 2010 6820
rect 2133 6817 2145 6820
rect 2179 6817 2191 6851
rect 2133 6811 2191 6817
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6817 2375 6851
rect 2317 6811 2375 6817
rect 2590 6808 2596 6860
rect 2648 6848 2654 6860
rect 2976 6848 3004 6888
rect 4890 6876 4896 6888
rect 4948 6876 4954 6928
rect 3510 6848 3516 6860
rect 2648 6820 3004 6848
rect 3471 6820 3516 6848
rect 2648 6808 2654 6820
rect 3510 6808 3516 6820
rect 3568 6808 3574 6860
rect 5736 6857 5764 6956
rect 7098 6916 7104 6928
rect 7059 6888 7104 6916
rect 7098 6876 7104 6888
rect 7156 6876 7162 6928
rect 7208 6916 7236 6956
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 8202 6984 8208 6996
rect 7340 6956 8208 6984
rect 7340 6944 7346 6956
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8294 6944 8300 6996
rect 8352 6984 8358 6996
rect 8941 6987 8999 6993
rect 8941 6984 8953 6987
rect 8352 6956 8953 6984
rect 8352 6944 8358 6956
rect 8941 6953 8953 6956
rect 8987 6953 8999 6987
rect 8941 6947 8999 6953
rect 9398 6944 9404 6996
rect 9456 6984 9462 6996
rect 11974 6984 11980 6996
rect 9456 6956 10088 6984
rect 9456 6944 9462 6956
rect 7650 6916 7656 6928
rect 7208 6888 7656 6916
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 8220 6888 8800 6916
rect 3881 6851 3939 6857
rect 3881 6817 3893 6851
rect 3927 6848 3939 6851
rect 5721 6851 5779 6857
rect 3927 6820 5672 6848
rect 3927 6817 3939 6820
rect 3881 6811 3939 6817
rect 1489 6783 1547 6789
rect 1489 6780 1501 6783
rect 1360 6752 1501 6780
rect 1360 6740 1366 6752
rect 1489 6749 1501 6752
rect 1535 6749 1547 6783
rect 1489 6743 1547 6749
rect 1765 6783 1823 6789
rect 1765 6749 1777 6783
rect 1811 6749 1823 6783
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 1765 6743 1823 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3970 6780 3976 6792
rect 3931 6752 3976 6780
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4062 6740 4068 6792
rect 4120 6780 4126 6792
rect 4246 6780 4252 6792
rect 4120 6752 4252 6780
rect 4120 6740 4126 6752
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4522 6780 4528 6792
rect 4483 6752 4528 6780
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 4890 6740 4896 6792
rect 4948 6780 4954 6792
rect 5166 6780 5172 6792
rect 4948 6752 5172 6780
rect 4948 6740 4954 6752
rect 5166 6740 5172 6752
rect 5224 6740 5230 6792
rect 5442 6780 5448 6792
rect 5403 6752 5448 6780
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 2038 6712 2044 6724
rect 1719 6684 2044 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 2038 6672 2044 6684
rect 2096 6672 2102 6724
rect 3329 6715 3387 6721
rect 3329 6681 3341 6715
rect 3375 6712 3387 6715
rect 4982 6712 4988 6724
rect 3375 6684 4988 6712
rect 3375 6681 3387 6684
rect 3329 6675 3387 6681
rect 4982 6672 4988 6684
rect 5040 6672 5046 6724
rect 5644 6712 5672 6820
rect 5721 6817 5733 6851
rect 5767 6817 5779 6851
rect 5721 6811 5779 6817
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 8220 6857 8248 6888
rect 7745 6851 7803 6857
rect 7745 6848 7757 6851
rect 6788 6820 7757 6848
rect 6788 6808 6794 6820
rect 7745 6817 7757 6820
rect 7791 6817 7803 6851
rect 7745 6811 7803 6817
rect 8205 6851 8263 6857
rect 8205 6817 8217 6851
rect 8251 6817 8263 6851
rect 8205 6811 8263 6817
rect 8294 6808 8300 6860
rect 8352 6848 8358 6860
rect 8662 6848 8668 6860
rect 8352 6820 8668 6848
rect 8352 6808 8358 6820
rect 8662 6808 8668 6820
rect 8720 6808 8726 6860
rect 8772 6848 8800 6888
rect 9324 6888 9628 6916
rect 9324 6848 9352 6888
rect 9490 6848 9496 6860
rect 8772 6820 9352 6848
rect 9451 6820 9496 6848
rect 9490 6808 9496 6820
rect 9548 6808 9554 6860
rect 9600 6848 9628 6888
rect 10060 6848 10088 6956
rect 10888 6956 11980 6984
rect 10594 6876 10600 6928
rect 10652 6916 10658 6928
rect 10888 6916 10916 6956
rect 11974 6944 11980 6956
rect 12032 6944 12038 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 13081 6987 13139 6993
rect 13081 6984 13093 6987
rect 13044 6956 13093 6984
rect 13044 6944 13050 6956
rect 13081 6953 13093 6956
rect 13127 6953 13139 6987
rect 13081 6947 13139 6953
rect 14369 6987 14427 6993
rect 14369 6953 14381 6987
rect 14415 6984 14427 6987
rect 15654 6984 15660 6996
rect 14415 6956 15660 6984
rect 14415 6953 14427 6956
rect 14369 6947 14427 6953
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 15746 6944 15752 6996
rect 15804 6984 15810 6996
rect 18046 6984 18052 6996
rect 15804 6956 18052 6984
rect 15804 6944 15810 6956
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18230 6944 18236 6996
rect 18288 6984 18294 6996
rect 20901 6987 20959 6993
rect 18288 6956 19288 6984
rect 18288 6944 18294 6956
rect 19260 6928 19288 6956
rect 20901 6953 20913 6987
rect 20947 6984 20959 6987
rect 21542 6984 21548 6996
rect 20947 6956 21548 6984
rect 20947 6953 20959 6956
rect 20901 6947 20959 6953
rect 21542 6944 21548 6956
rect 21600 6944 21606 6996
rect 10652 6888 10916 6916
rect 10652 6876 10658 6888
rect 10413 6851 10471 6857
rect 9600 6820 9904 6848
rect 10060 6820 10364 6848
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5977 6783 6035 6789
rect 5977 6780 5989 6783
rect 5868 6752 5989 6780
rect 5868 6740 5874 6752
rect 5977 6749 5989 6752
rect 6023 6749 6035 6783
rect 7561 6783 7619 6789
rect 7561 6780 7573 6783
rect 5977 6743 6035 6749
rect 6095 6752 7573 6780
rect 6095 6712 6123 6752
rect 7561 6749 7573 6752
rect 7607 6780 7619 6783
rect 8110 6780 8116 6792
rect 7607 6752 8116 6780
rect 7607 6749 7619 6752
rect 7561 6743 7619 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 8478 6740 8484 6792
rect 8536 6780 8542 6792
rect 9214 6780 9220 6792
rect 8536 6752 9220 6780
rect 8536 6740 8542 6752
rect 9214 6740 9220 6752
rect 9272 6740 9278 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9876 6780 9904 6820
rect 10042 6780 10048 6792
rect 9364 6752 9409 6780
rect 9876 6752 10048 6780
rect 9364 6740 9370 6752
rect 10042 6740 10048 6752
rect 10100 6740 10106 6792
rect 10137 6783 10195 6789
rect 10137 6749 10149 6783
rect 10183 6780 10195 6783
rect 10226 6780 10232 6792
rect 10183 6752 10232 6780
rect 10183 6749 10195 6752
rect 10137 6743 10195 6749
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10336 6780 10364 6820
rect 10413 6817 10425 6851
rect 10459 6848 10471 6851
rect 10888 6848 10916 6888
rect 15930 6876 15936 6928
rect 15988 6916 15994 6928
rect 16482 6916 16488 6928
rect 15988 6888 16488 6916
rect 15988 6876 15994 6888
rect 16482 6876 16488 6888
rect 16540 6876 16546 6928
rect 16761 6919 16819 6925
rect 16761 6885 16773 6919
rect 16807 6885 16819 6919
rect 16761 6879 16819 6885
rect 10459 6820 10916 6848
rect 10965 6851 11023 6857
rect 10459 6817 10471 6820
rect 10413 6811 10471 6817
rect 10965 6817 10977 6851
rect 11011 6848 11023 6851
rect 11054 6848 11060 6860
rect 11011 6820 11060 6848
rect 11011 6817 11023 6820
rect 10965 6811 11023 6817
rect 11054 6808 11060 6820
rect 11112 6808 11118 6860
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 11609 6851 11667 6857
rect 11609 6848 11621 6851
rect 11296 6820 11621 6848
rect 11296 6808 11302 6820
rect 11609 6817 11621 6820
rect 11655 6817 11667 6851
rect 13538 6848 13544 6860
rect 13499 6820 13544 6848
rect 11609 6811 11667 6817
rect 13538 6808 13544 6820
rect 13596 6808 13602 6860
rect 13633 6851 13691 6857
rect 13633 6817 13645 6851
rect 13679 6817 13691 6851
rect 14458 6848 14464 6860
rect 14419 6820 14464 6848
rect 13633 6811 13691 6817
rect 11149 6783 11207 6789
rect 11149 6780 11161 6783
rect 10336 6752 11161 6780
rect 11149 6749 11161 6752
rect 11195 6749 11207 6783
rect 12434 6780 12440 6792
rect 11149 6743 11207 6749
rect 11440 6752 12440 6780
rect 5644 6684 6123 6712
rect 6546 6672 6552 6724
rect 6604 6712 6610 6724
rect 10597 6715 10655 6721
rect 10597 6712 10609 6715
rect 6604 6684 10609 6712
rect 6604 6672 6610 6684
rect 10597 6681 10609 6684
rect 10643 6712 10655 6715
rect 11238 6712 11244 6724
rect 10643 6684 11244 6712
rect 10643 6681 10655 6684
rect 10597 6675 10655 6681
rect 11238 6672 11244 6684
rect 11296 6672 11302 6724
rect 1854 6604 1860 6656
rect 1912 6644 1918 6656
rect 1949 6647 2007 6653
rect 1949 6644 1961 6647
rect 1912 6616 1961 6644
rect 1912 6604 1918 6616
rect 1949 6613 1961 6616
rect 1995 6613 2007 6647
rect 1949 6607 2007 6613
rect 2130 6604 2136 6656
rect 2188 6644 2194 6656
rect 2409 6647 2467 6653
rect 2409 6644 2421 6647
rect 2188 6616 2421 6644
rect 2188 6604 2194 6616
rect 2409 6613 2421 6616
rect 2455 6613 2467 6647
rect 2409 6607 2467 6613
rect 2774 6604 2780 6656
rect 2832 6644 2838 6656
rect 4154 6644 4160 6656
rect 2832 6616 2877 6644
rect 4115 6616 4160 6644
rect 2832 6604 2838 6616
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4706 6604 4712 6656
rect 4764 6644 4770 6656
rect 5353 6647 5411 6653
rect 5353 6644 5365 6647
rect 4764 6616 5365 6644
rect 4764 6604 4770 6616
rect 5353 6613 5365 6616
rect 5399 6613 5411 6647
rect 5626 6644 5632 6656
rect 5587 6616 5632 6644
rect 5353 6607 5411 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5902 6604 5908 6656
rect 5960 6644 5966 6656
rect 7193 6647 7251 6653
rect 7193 6644 7205 6647
rect 5960 6616 7205 6644
rect 5960 6604 5966 6616
rect 7193 6613 7205 6616
rect 7239 6613 7251 6647
rect 7193 6607 7251 6613
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 7524 6616 7665 6644
rect 7524 6604 7530 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 7926 6604 7932 6656
rect 7984 6644 7990 6656
rect 8389 6647 8447 6653
rect 8389 6644 8401 6647
rect 7984 6616 8401 6644
rect 7984 6604 7990 6616
rect 8389 6613 8401 6616
rect 8435 6613 8447 6647
rect 8389 6607 8447 6613
rect 8757 6647 8815 6653
rect 8757 6613 8769 6647
rect 8803 6644 8815 6647
rect 9214 6644 9220 6656
rect 8803 6616 9220 6644
rect 8803 6613 8815 6616
rect 8757 6607 8815 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 9401 6647 9459 6653
rect 9401 6644 9413 6647
rect 9364 6616 9413 6644
rect 9364 6604 9370 6616
rect 9401 6613 9413 6616
rect 9447 6613 9459 6647
rect 9766 6644 9772 6656
rect 9727 6616 9772 6644
rect 9401 6607 9459 6613
rect 9766 6604 9772 6616
rect 9824 6604 9830 6656
rect 10134 6604 10140 6656
rect 10192 6644 10198 6656
rect 10229 6647 10287 6653
rect 10229 6644 10241 6647
rect 10192 6616 10241 6644
rect 10192 6604 10198 6616
rect 10229 6613 10241 6616
rect 10275 6613 10287 6647
rect 10229 6607 10287 6613
rect 10870 6604 10876 6656
rect 10928 6644 10934 6656
rect 11057 6647 11115 6653
rect 11057 6644 11069 6647
rect 10928 6616 11069 6644
rect 10928 6604 10934 6616
rect 11057 6613 11069 6616
rect 11103 6644 11115 6647
rect 11440 6644 11468 6752
rect 12434 6740 12440 6752
rect 12492 6740 12498 6792
rect 13170 6740 13176 6792
rect 13228 6780 13234 6792
rect 13449 6783 13507 6789
rect 13449 6780 13461 6783
rect 13228 6752 13461 6780
rect 13228 6740 13234 6752
rect 13449 6749 13461 6752
rect 13495 6749 13507 6783
rect 13449 6743 13507 6749
rect 11876 6715 11934 6721
rect 11876 6681 11888 6715
rect 11922 6712 11934 6715
rect 12066 6712 12072 6724
rect 11922 6684 12072 6712
rect 11922 6681 11934 6684
rect 11876 6675 11934 6681
rect 12066 6672 12072 6684
rect 12124 6712 12130 6724
rect 13648 6712 13676 6811
rect 14458 6808 14464 6820
rect 14516 6808 14522 6860
rect 16209 6851 16267 6857
rect 16209 6817 16221 6851
rect 16255 6817 16267 6851
rect 16776 6848 16804 6879
rect 17218 6876 17224 6928
rect 17276 6916 17282 6928
rect 18138 6916 18144 6928
rect 17276 6888 18144 6916
rect 17276 6876 17282 6888
rect 16942 6848 16948 6860
rect 16776 6820 16948 6848
rect 16209 6811 16267 6817
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6780 14243 6783
rect 15930 6780 15936 6792
rect 14231 6752 15936 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 15930 6740 15936 6752
rect 15988 6740 15994 6792
rect 16114 6740 16120 6792
rect 16172 6780 16178 6792
rect 16224 6780 16252 6811
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17126 6808 17132 6860
rect 17184 6848 17190 6860
rect 17512 6857 17540 6888
rect 18138 6876 18144 6888
rect 18196 6876 18202 6928
rect 18693 6919 18751 6925
rect 18693 6885 18705 6919
rect 18739 6885 18751 6919
rect 18693 6879 18751 6885
rect 17313 6851 17371 6857
rect 17313 6848 17325 6851
rect 17184 6820 17325 6848
rect 17184 6808 17190 6820
rect 17313 6817 17325 6820
rect 17359 6817 17371 6851
rect 17313 6811 17371 6817
rect 17497 6851 17555 6857
rect 17497 6817 17509 6851
rect 17543 6817 17555 6851
rect 18230 6848 18236 6860
rect 17497 6811 17555 6817
rect 17604 6820 18236 6848
rect 17604 6780 17632 6820
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 18414 6808 18420 6860
rect 18472 6848 18478 6860
rect 18708 6848 18736 6879
rect 19242 6876 19248 6928
rect 19300 6876 19306 6928
rect 18472 6820 18644 6848
rect 18708 6820 19656 6848
rect 18472 6808 18478 6820
rect 16172 6752 17632 6780
rect 16172 6740 16178 6752
rect 17954 6740 17960 6792
rect 18012 6780 18018 6792
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 18012 6752 18153 6780
rect 18012 6740 18018 6752
rect 18141 6749 18153 6752
rect 18187 6749 18199 6783
rect 18506 6780 18512 6792
rect 18467 6752 18512 6780
rect 18141 6743 18199 6749
rect 18506 6740 18512 6752
rect 18564 6740 18570 6792
rect 18616 6780 18644 6820
rect 18874 6780 18880 6792
rect 18616 6752 18880 6780
rect 18874 6740 18880 6752
rect 18932 6780 18938 6792
rect 18932 6752 19104 6780
rect 18932 6740 18938 6752
rect 12124 6684 13676 6712
rect 12124 6672 12130 6684
rect 13722 6672 13728 6724
rect 13780 6712 13786 6724
rect 14728 6715 14786 6721
rect 13780 6684 14688 6712
rect 13780 6672 13786 6684
rect 11103 6616 11468 6644
rect 11517 6647 11575 6653
rect 11103 6613 11115 6616
rect 11057 6607 11115 6613
rect 11517 6613 11529 6647
rect 11563 6644 11575 6647
rect 11698 6644 11704 6656
rect 11563 6616 11704 6644
rect 11563 6613 11575 6616
rect 11517 6607 11575 6613
rect 11698 6604 11704 6616
rect 11756 6604 11762 6656
rect 11790 6604 11796 6656
rect 11848 6644 11854 6656
rect 12342 6644 12348 6656
rect 11848 6616 12348 6644
rect 11848 6604 11854 6616
rect 12342 6604 12348 6616
rect 12400 6644 12406 6656
rect 12989 6647 13047 6653
rect 12989 6644 13001 6647
rect 12400 6616 13001 6644
rect 12400 6604 12406 6616
rect 12989 6613 13001 6616
rect 13035 6613 13047 6647
rect 12989 6607 13047 6613
rect 13906 6604 13912 6656
rect 13964 6644 13970 6656
rect 14550 6644 14556 6656
rect 13964 6616 14556 6644
rect 13964 6604 13970 6616
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 14660 6644 14688 6684
rect 14728 6681 14740 6715
rect 14774 6712 14786 6715
rect 15286 6712 15292 6724
rect 14774 6684 15292 6712
rect 14774 6681 14786 6684
rect 14728 6675 14786 6681
rect 15286 6672 15292 6684
rect 15344 6672 15350 6724
rect 16393 6715 16451 6721
rect 16393 6681 16405 6715
rect 16439 6712 16451 6715
rect 17494 6712 17500 6724
rect 16439 6684 16896 6712
rect 16439 6681 16451 6684
rect 16393 6675 16451 6681
rect 15562 6644 15568 6656
rect 14660 6616 15568 6644
rect 15562 6604 15568 6616
rect 15620 6604 15626 6656
rect 15838 6644 15844 6656
rect 15799 6616 15844 6644
rect 15838 6604 15844 6616
rect 15896 6604 15902 6656
rect 16298 6644 16304 6656
rect 16259 6616 16304 6644
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 16868 6653 16896 6684
rect 17236 6684 17500 6712
rect 17236 6653 17264 6684
rect 17494 6672 17500 6684
rect 17552 6672 17558 6724
rect 18966 6712 18972 6724
rect 18927 6684 18972 6712
rect 18966 6672 18972 6684
rect 19024 6672 19030 6724
rect 19076 6712 19104 6752
rect 19150 6740 19156 6792
rect 19208 6780 19214 6792
rect 19245 6783 19303 6789
rect 19245 6780 19257 6783
rect 19208 6752 19257 6780
rect 19208 6740 19214 6752
rect 19245 6749 19257 6752
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 19521 6783 19579 6789
rect 19521 6749 19533 6783
rect 19567 6749 19579 6783
rect 19628 6780 19656 6820
rect 21082 6808 21088 6860
rect 21140 6848 21146 6860
rect 21269 6851 21327 6857
rect 21269 6848 21281 6851
rect 21140 6820 21281 6848
rect 21140 6808 21146 6820
rect 21269 6817 21281 6820
rect 21315 6817 21327 6851
rect 21269 6811 21327 6817
rect 21453 6783 21511 6789
rect 19628 6752 20024 6780
rect 19521 6743 19579 6749
rect 19536 6712 19564 6743
rect 19996 6724 20024 6752
rect 21453 6749 21465 6783
rect 21499 6780 21511 6783
rect 21818 6780 21824 6792
rect 21499 6752 21824 6780
rect 21499 6749 21511 6752
rect 21453 6743 21511 6749
rect 21818 6740 21824 6752
rect 21876 6740 21882 6792
rect 19076 6684 19564 6712
rect 19788 6715 19846 6721
rect 19788 6681 19800 6715
rect 19834 6712 19846 6715
rect 19886 6712 19892 6724
rect 19834 6684 19892 6712
rect 19834 6681 19846 6684
rect 19788 6675 19846 6681
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 19978 6672 19984 6724
rect 20036 6672 20042 6724
rect 20714 6672 20720 6724
rect 20772 6712 20778 6724
rect 20993 6715 21051 6721
rect 20993 6712 21005 6715
rect 20772 6684 21005 6712
rect 20772 6672 20778 6684
rect 20993 6681 21005 6684
rect 21039 6681 21051 6715
rect 20993 6675 21051 6681
rect 16853 6647 16911 6653
rect 16853 6613 16865 6647
rect 16899 6613 16911 6647
rect 16853 6607 16911 6613
rect 17221 6647 17279 6653
rect 17221 6613 17233 6647
rect 17267 6613 17279 6647
rect 17221 6607 17279 6613
rect 17402 6604 17408 6656
rect 17460 6644 17466 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17460 6616 17693 6644
rect 17460 6604 17466 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 18049 6647 18107 6653
rect 18049 6613 18061 6647
rect 18095 6644 18107 6647
rect 18138 6644 18144 6656
rect 18095 6616 18144 6644
rect 18095 6613 18107 6616
rect 18049 6607 18107 6613
rect 18138 6604 18144 6616
rect 18196 6604 18202 6656
rect 18506 6604 18512 6656
rect 18564 6644 18570 6656
rect 18877 6647 18935 6653
rect 18877 6644 18889 6647
rect 18564 6616 18889 6644
rect 18564 6604 18570 6616
rect 18877 6613 18889 6616
rect 18923 6613 18935 6647
rect 18877 6607 18935 6613
rect 19429 6647 19487 6653
rect 19429 6613 19441 6647
rect 19475 6644 19487 6647
rect 20438 6644 20444 6656
rect 19475 6616 20444 6644
rect 19475 6613 19487 6616
rect 19429 6607 19487 6613
rect 20438 6604 20444 6616
rect 20496 6604 20502 6656
rect 21450 6604 21456 6656
rect 21508 6644 21514 6656
rect 21818 6644 21824 6656
rect 21508 6616 21824 6644
rect 21508 6604 21514 6616
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 1394 6400 1400 6452
rect 1452 6440 1458 6452
rect 1765 6443 1823 6449
rect 1765 6440 1777 6443
rect 1452 6412 1777 6440
rect 1452 6400 1458 6412
rect 1765 6409 1777 6412
rect 1811 6409 1823 6443
rect 1765 6403 1823 6409
rect 2222 6400 2228 6452
rect 2280 6440 2286 6452
rect 2317 6443 2375 6449
rect 2317 6440 2329 6443
rect 2280 6412 2329 6440
rect 2280 6400 2286 6412
rect 2317 6409 2329 6412
rect 2363 6409 2375 6443
rect 2317 6403 2375 6409
rect 2409 6443 2467 6449
rect 2409 6409 2421 6443
rect 2455 6440 2467 6443
rect 2777 6443 2835 6449
rect 2777 6440 2789 6443
rect 2455 6412 2789 6440
rect 2455 6409 2467 6412
rect 2409 6403 2467 6409
rect 2777 6409 2789 6412
rect 2823 6409 2835 6443
rect 2777 6403 2835 6409
rect 3145 6443 3203 6449
rect 3145 6409 3157 6443
rect 3191 6440 3203 6443
rect 3418 6440 3424 6452
rect 3191 6412 3424 6440
rect 3191 6409 3203 6412
rect 3145 6403 3203 6409
rect 3418 6400 3424 6412
rect 3476 6440 3482 6452
rect 3878 6440 3884 6452
rect 3476 6412 3884 6440
rect 3476 6400 3482 6412
rect 3878 6400 3884 6412
rect 3936 6400 3942 6452
rect 4249 6443 4307 6449
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 5445 6443 5503 6449
rect 5445 6440 5457 6443
rect 4295 6412 5457 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 5445 6409 5457 6412
rect 5491 6409 5503 6443
rect 5445 6403 5503 6409
rect 5718 6400 5724 6452
rect 5776 6400 5782 6452
rect 5810 6400 5816 6452
rect 5868 6400 5874 6452
rect 5994 6400 6000 6452
rect 6052 6440 6058 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 6052 6412 6377 6440
rect 6052 6400 6058 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 6365 6403 6423 6409
rect 6822 6400 6828 6452
rect 6880 6440 6886 6452
rect 6880 6412 6925 6440
rect 6880 6400 6886 6412
rect 7006 6400 7012 6452
rect 7064 6440 7070 6452
rect 7193 6443 7251 6449
rect 7193 6440 7205 6443
rect 7064 6412 7205 6440
rect 7064 6400 7070 6412
rect 7193 6409 7205 6412
rect 7239 6409 7251 6443
rect 7193 6403 7251 6409
rect 8021 6443 8079 6449
rect 8021 6409 8033 6443
rect 8067 6440 8079 6443
rect 8110 6440 8116 6452
rect 8067 6412 8116 6440
rect 8067 6409 8079 6412
rect 8021 6403 8079 6409
rect 8110 6400 8116 6412
rect 8168 6400 8174 6452
rect 8938 6440 8944 6452
rect 8899 6412 8944 6440
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9033 6443 9091 6449
rect 9033 6409 9045 6443
rect 9079 6440 9091 6443
rect 9582 6440 9588 6452
rect 9079 6412 9588 6440
rect 9079 6409 9091 6412
rect 9033 6403 9091 6409
rect 9582 6400 9588 6412
rect 9640 6400 9646 6452
rect 9766 6440 9772 6452
rect 9727 6412 9772 6440
rect 9766 6400 9772 6412
rect 9824 6400 9830 6452
rect 10597 6443 10655 6449
rect 10597 6409 10609 6443
rect 10643 6440 10655 6443
rect 11517 6443 11575 6449
rect 11517 6440 11529 6443
rect 10643 6412 11529 6440
rect 10643 6409 10655 6412
rect 10597 6403 10655 6409
rect 11517 6409 11529 6412
rect 11563 6409 11575 6443
rect 13722 6440 13728 6452
rect 11517 6403 11575 6409
rect 11992 6412 13728 6440
rect 382 6332 388 6384
rect 440 6372 446 6384
rect 934 6372 940 6384
rect 440 6344 940 6372
rect 440 6332 446 6344
rect 934 6332 940 6344
rect 992 6372 998 6384
rect 1489 6375 1547 6381
rect 1489 6372 1501 6375
rect 992 6344 1501 6372
rect 992 6332 998 6344
rect 1489 6341 1501 6344
rect 1535 6341 1547 6375
rect 1489 6335 1547 6341
rect 3050 6332 3056 6384
rect 3108 6372 3114 6384
rect 3237 6375 3295 6381
rect 3237 6372 3249 6375
rect 3108 6344 3249 6372
rect 3108 6332 3114 6344
rect 3237 6341 3249 6344
rect 3283 6341 3295 6375
rect 3237 6335 3295 6341
rect 4522 6332 4528 6384
rect 4580 6372 4586 6384
rect 4580 6344 5304 6372
rect 4580 6332 4586 6344
rect 3694 6304 3700 6316
rect 3655 6276 3700 6304
rect 3694 6264 3700 6276
rect 3752 6264 3758 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4890 6304 4896 6316
rect 4203 6276 4896 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 4985 6307 5043 6313
rect 4985 6273 4997 6307
rect 5031 6304 5043 6307
rect 5166 6304 5172 6316
rect 5031 6276 5172 6304
rect 5031 6273 5043 6276
rect 4985 6267 5043 6273
rect 5166 6264 5172 6276
rect 5224 6264 5230 6316
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6236 1731 6239
rect 2406 6236 2412 6248
rect 1719 6208 2412 6236
rect 1719 6205 1731 6208
rect 1673 6199 1731 6205
rect 2406 6196 2412 6208
rect 2464 6196 2470 6248
rect 2593 6239 2651 6245
rect 2593 6205 2605 6239
rect 2639 6236 2651 6239
rect 2958 6236 2964 6248
rect 2639 6208 2964 6236
rect 2639 6205 2651 6208
rect 2593 6199 2651 6205
rect 2958 6196 2964 6208
rect 3016 6196 3022 6248
rect 3329 6239 3387 6245
rect 3329 6205 3341 6239
rect 3375 6236 3387 6239
rect 4062 6236 4068 6248
rect 3375 6208 4068 6236
rect 3375 6205 3387 6208
rect 3329 6199 3387 6205
rect 3344 6168 3372 6199
rect 4062 6196 4068 6208
rect 4120 6196 4126 6248
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 5276 6245 5304 6344
rect 5350 6332 5356 6384
rect 5408 6372 5414 6384
rect 5736 6372 5764 6400
rect 5408 6344 5764 6372
rect 5828 6372 5856 6400
rect 5905 6375 5963 6381
rect 5905 6372 5917 6375
rect 5828 6344 5917 6372
rect 5408 6332 5414 6344
rect 5905 6341 5917 6344
rect 5951 6341 5963 6375
rect 9306 6372 9312 6384
rect 5905 6335 5963 6341
rect 6380 6344 9312 6372
rect 5813 6307 5871 6313
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6178 6304 6184 6316
rect 5859 6276 6184 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6178 6264 6184 6276
rect 6236 6264 6242 6316
rect 6380 6248 6408 6344
rect 9306 6332 9312 6344
rect 9364 6332 9370 6384
rect 10888 6344 11192 6372
rect 6721 6264 6727 6316
rect 6779 6313 6785 6316
rect 6779 6304 6791 6313
rect 6779 6276 6824 6304
rect 6886 6276 7135 6304
rect 6779 6267 6791 6276
rect 6779 6264 6785 6267
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 4304 6208 4353 6236
rect 4304 6196 4310 6208
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 5077 6239 5135 6245
rect 5077 6205 5089 6239
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5261 6239 5319 6245
rect 5261 6205 5273 6239
rect 5307 6236 5319 6239
rect 5718 6236 5724 6248
rect 5307 6208 5724 6236
rect 5307 6205 5319 6208
rect 5261 6199 5319 6205
rect 3252 6140 3372 6168
rect 3252 6112 3280 6140
rect 3418 6128 3424 6180
rect 3476 6168 3482 6180
rect 3789 6171 3847 6177
rect 3789 6168 3801 6171
rect 3476 6140 3801 6168
rect 3476 6128 3482 6140
rect 3789 6137 3801 6140
rect 3835 6137 3847 6171
rect 5092 6168 5120 6199
rect 5718 6196 5724 6208
rect 5776 6196 5782 6248
rect 6086 6196 6092 6248
rect 6144 6236 6150 6248
rect 6144 6208 6189 6236
rect 6144 6196 6150 6208
rect 6362 6196 6368 6248
rect 6420 6196 6426 6248
rect 6454 6196 6460 6248
rect 6512 6236 6518 6248
rect 6886 6236 6914 6276
rect 6512 6208 6914 6236
rect 7009 6239 7067 6245
rect 6512 6196 6518 6208
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7009 6199 7067 6205
rect 5092 6140 5534 6168
rect 3789 6131 3847 6137
rect 1946 6100 1952 6112
rect 1907 6072 1952 6100
rect 1946 6060 1952 6072
rect 2004 6060 2010 6112
rect 2314 6060 2320 6112
rect 2372 6100 2378 6112
rect 2774 6100 2780 6112
rect 2372 6072 2780 6100
rect 2372 6060 2378 6072
rect 2774 6060 2780 6072
rect 2832 6060 2838 6112
rect 3234 6060 3240 6112
rect 3292 6060 3298 6112
rect 4617 6103 4675 6109
rect 4617 6069 4629 6103
rect 4663 6100 4675 6103
rect 5074 6100 5080 6112
rect 4663 6072 5080 6100
rect 4663 6069 4675 6072
rect 4617 6063 4675 6069
rect 5074 6060 5080 6072
rect 5132 6060 5138 6112
rect 5506 6100 5534 6140
rect 5994 6128 6000 6180
rect 6052 6168 6058 6180
rect 6914 6168 6920 6180
rect 6052 6140 6920 6168
rect 6052 6128 6058 6140
rect 6914 6128 6920 6140
rect 6972 6168 6978 6180
rect 7024 6168 7052 6199
rect 6972 6140 7052 6168
rect 7107 6168 7135 6276
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7377 6307 7435 6313
rect 7377 6304 7389 6307
rect 7248 6276 7389 6304
rect 7248 6264 7254 6276
rect 7377 6273 7389 6276
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 7653 6307 7711 6313
rect 8113 6308 8171 6313
rect 7653 6273 7665 6307
rect 7699 6304 7711 6307
rect 7944 6307 8171 6308
rect 7944 6304 8125 6307
rect 7699 6280 8125 6304
rect 7699 6276 7972 6280
rect 7699 6273 7711 6276
rect 7653 6267 7711 6273
rect 8113 6273 8125 6280
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 9950 6304 9956 6316
rect 8260 6276 9956 6304
rect 8260 6264 8266 6276
rect 9950 6264 9956 6276
rect 10008 6304 10014 6316
rect 10134 6304 10140 6316
rect 10008 6276 10140 6304
rect 10008 6264 10014 6276
rect 10134 6264 10140 6276
rect 10192 6264 10198 6316
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 10778 6304 10784 6316
rect 10735 6276 10784 6304
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 10778 6264 10784 6276
rect 10836 6264 10842 6316
rect 7929 6239 7987 6245
rect 7929 6205 7941 6239
rect 7975 6236 7987 6239
rect 8294 6236 8300 6248
rect 7975 6208 8300 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8294 6196 8300 6208
rect 8352 6236 8358 6248
rect 9217 6239 9275 6245
rect 9217 6236 9229 6239
rect 8352 6208 9229 6236
rect 8352 6196 8358 6208
rect 9217 6205 9229 6208
rect 9263 6236 9275 6239
rect 9493 6239 9551 6245
rect 9263 6208 9343 6236
rect 9263 6205 9275 6208
rect 9217 6199 9275 6205
rect 8018 6168 8024 6180
rect 7107 6140 8024 6168
rect 6972 6128 6978 6140
rect 8018 6128 8024 6140
rect 8076 6128 8082 6180
rect 8202 6128 8208 6180
rect 8260 6168 8266 6180
rect 8260 6140 8616 6168
rect 8260 6128 8266 6140
rect 7926 6100 7932 6112
rect 5506 6072 7932 6100
rect 7926 6060 7932 6072
rect 7984 6060 7990 6112
rect 8110 6060 8116 6112
rect 8168 6100 8174 6112
rect 8588 6109 8616 6140
rect 8481 6103 8539 6109
rect 8481 6100 8493 6103
rect 8168 6072 8493 6100
rect 8168 6060 8174 6072
rect 8481 6069 8493 6072
rect 8527 6069 8539 6103
rect 8481 6063 8539 6069
rect 8573 6103 8631 6109
rect 8573 6069 8585 6103
rect 8619 6069 8631 6103
rect 9315 6100 9343 6208
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9674 6236 9680 6248
rect 9635 6208 9680 6236
rect 9493 6199 9551 6205
rect 9508 6168 9536 6199
rect 9674 6196 9680 6208
rect 9732 6196 9738 6248
rect 10413 6239 10471 6245
rect 10413 6205 10425 6239
rect 10459 6205 10471 6239
rect 10888 6236 10916 6344
rect 11164 6313 11192 6344
rect 11238 6332 11244 6384
rect 11296 6372 11302 6384
rect 11992 6381 12020 6412
rect 13722 6400 13728 6412
rect 13780 6400 13786 6452
rect 13909 6443 13967 6449
rect 13909 6409 13921 6443
rect 13955 6409 13967 6443
rect 13909 6403 13967 6409
rect 15105 6443 15163 6449
rect 15105 6409 15117 6443
rect 15151 6440 15163 6443
rect 16298 6440 16304 6452
rect 15151 6412 16304 6440
rect 15151 6409 15163 6412
rect 15105 6403 15163 6409
rect 11977 6375 12035 6381
rect 11977 6372 11989 6375
rect 11296 6344 11989 6372
rect 11296 6332 11302 6344
rect 11977 6341 11989 6344
rect 12023 6341 12035 6375
rect 11977 6335 12035 6341
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 12774 6375 12832 6381
rect 12774 6372 12786 6375
rect 12400 6344 12786 6372
rect 12400 6332 12406 6344
rect 12774 6341 12786 6344
rect 12820 6341 12832 6375
rect 12774 6335 12832 6341
rect 12986 6332 12992 6384
rect 13044 6372 13050 6384
rect 13630 6372 13636 6384
rect 13044 6344 13636 6372
rect 13044 6332 13050 6344
rect 13630 6332 13636 6344
rect 13688 6332 13694 6384
rect 13924 6372 13952 6403
rect 16298 6400 16304 6412
rect 16356 6400 16362 6452
rect 17221 6443 17279 6449
rect 17221 6409 17233 6443
rect 17267 6440 17279 6443
rect 18138 6440 18144 6452
rect 17267 6412 18144 6440
rect 17267 6409 17279 6412
rect 17221 6403 17279 6409
rect 18138 6400 18144 6412
rect 18196 6400 18202 6452
rect 19058 6440 19064 6452
rect 19019 6412 19064 6440
rect 19058 6400 19064 6412
rect 19116 6400 19122 6452
rect 19610 6400 19616 6452
rect 19668 6440 19674 6452
rect 20165 6443 20223 6449
rect 20165 6440 20177 6443
rect 19668 6412 20177 6440
rect 19668 6400 19674 6412
rect 20165 6409 20177 6412
rect 20211 6409 20223 6443
rect 20622 6440 20628 6452
rect 20583 6412 20628 6440
rect 20165 6403 20223 6409
rect 20622 6400 20628 6412
rect 20680 6400 20686 6452
rect 14185 6375 14243 6381
rect 14185 6372 14197 6375
rect 13924 6344 14197 6372
rect 14185 6341 14197 6344
rect 14231 6372 14243 6375
rect 14642 6372 14648 6384
rect 14231 6344 14648 6372
rect 14231 6341 14243 6344
rect 14185 6335 14243 6341
rect 14642 6332 14648 6344
rect 14700 6332 14706 6384
rect 14737 6375 14795 6381
rect 14737 6341 14749 6375
rect 14783 6372 14795 6375
rect 15470 6372 15476 6384
rect 14783 6344 15476 6372
rect 14783 6341 14795 6344
rect 14737 6335 14795 6341
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 18506 6372 18512 6384
rect 15580 6344 17632 6372
rect 11149 6307 11207 6313
rect 11149 6273 11161 6307
rect 11195 6273 11207 6307
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 11149 6267 11207 6273
rect 11882 6264 11888 6276
rect 11940 6304 11946 6316
rect 12437 6307 12495 6313
rect 12437 6304 12449 6307
rect 11940 6276 12449 6304
rect 11940 6264 11946 6276
rect 12437 6273 12449 6276
rect 12483 6273 12495 6307
rect 12437 6267 12495 6273
rect 12529 6307 12587 6313
rect 12529 6273 12541 6307
rect 12575 6304 12587 6307
rect 14274 6304 14280 6316
rect 12575 6276 14280 6304
rect 12575 6273 12587 6276
rect 12529 6267 12587 6273
rect 14274 6264 14280 6276
rect 14332 6264 14338 6316
rect 15580 6304 15608 6344
rect 15488 6276 15608 6304
rect 10413 6199 10471 6205
rect 10704 6208 10916 6236
rect 9766 6168 9772 6180
rect 9508 6140 9772 6168
rect 9766 6128 9772 6140
rect 9824 6168 9830 6180
rect 10428 6168 10456 6199
rect 10704 6180 10732 6208
rect 11422 6196 11428 6248
rect 11480 6236 11486 6248
rect 11974 6236 11980 6248
rect 11480 6208 11980 6236
rect 11480 6196 11486 6208
rect 11974 6196 11980 6208
rect 12032 6236 12038 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 12032 6208 12081 6236
rect 12032 6196 12038 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12069 6199 12127 6205
rect 14553 6239 14611 6245
rect 14553 6205 14565 6239
rect 14599 6205 14611 6239
rect 14553 6199 14611 6205
rect 14645 6239 14703 6245
rect 14645 6205 14657 6239
rect 14691 6236 14703 6239
rect 15102 6236 15108 6248
rect 14691 6208 15108 6236
rect 14691 6205 14703 6208
rect 14645 6199 14703 6205
rect 10594 6168 10600 6180
rect 9824 6140 10600 6168
rect 9824 6128 9830 6140
rect 10594 6128 10600 6140
rect 10652 6128 10658 6180
rect 10686 6128 10692 6180
rect 10744 6128 10750 6180
rect 11790 6128 11796 6180
rect 11848 6168 11854 6180
rect 12158 6168 12164 6180
rect 11848 6140 12164 6168
rect 11848 6128 11854 6140
rect 12158 6128 12164 6140
rect 12216 6128 12222 6180
rect 13722 6128 13728 6180
rect 13780 6168 13786 6180
rect 14001 6171 14059 6177
rect 14001 6168 14013 6171
rect 13780 6140 14013 6168
rect 13780 6128 13786 6140
rect 14001 6137 14013 6140
rect 14047 6137 14059 6171
rect 14568 6168 14596 6199
rect 15102 6196 15108 6208
rect 15160 6196 15166 6248
rect 15488 6245 15516 6276
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15712 6276 15757 6304
rect 15712 6264 15718 6276
rect 16114 6264 16120 6316
rect 16172 6304 16178 6316
rect 16293 6307 16351 6313
rect 16293 6304 16305 6307
rect 16172 6276 16305 6304
rect 16172 6264 16178 6276
rect 16293 6273 16305 6276
rect 16339 6273 16351 6307
rect 16574 6304 16580 6316
rect 16293 6267 16351 6273
rect 16408 6276 16580 6304
rect 15473 6239 15531 6245
rect 15473 6205 15485 6239
rect 15519 6205 15531 6239
rect 15473 6199 15531 6205
rect 15565 6239 15623 6245
rect 15565 6205 15577 6239
rect 15611 6236 15623 6239
rect 16408 6236 16436 6276
rect 16574 6264 16580 6276
rect 16632 6264 16638 6316
rect 16669 6307 16727 6313
rect 16669 6273 16681 6307
rect 16715 6304 16727 6307
rect 17034 6304 17040 6316
rect 16715 6276 17040 6304
rect 16715 6273 16727 6276
rect 16669 6267 16727 6273
rect 17034 6264 17040 6276
rect 17092 6264 17098 6316
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 17604 6313 17632 6344
rect 17696 6344 18512 6372
rect 17313 6307 17371 6313
rect 17313 6304 17325 6307
rect 17276 6276 17325 6304
rect 17276 6264 17282 6276
rect 17313 6273 17325 6276
rect 17359 6273 17371 6307
rect 17313 6267 17371 6273
rect 17589 6307 17647 6313
rect 17589 6273 17601 6307
rect 17635 6273 17647 6307
rect 17589 6267 17647 6273
rect 15611 6208 16436 6236
rect 15611 6205 15623 6208
rect 15565 6199 15623 6205
rect 15286 6168 15292 6180
rect 14568 6140 15292 6168
rect 14001 6131 14059 6137
rect 15286 6128 15292 6140
rect 15344 6168 15350 6180
rect 15488 6168 15516 6199
rect 16482 6196 16488 6248
rect 16540 6236 16546 6248
rect 17696 6236 17724 6344
rect 18506 6332 18512 6344
rect 18564 6332 18570 6384
rect 19521 6375 19579 6381
rect 19521 6341 19533 6375
rect 19567 6372 19579 6375
rect 22922 6372 22928 6384
rect 19567 6344 22928 6372
rect 19567 6341 19579 6344
rect 19521 6335 19579 6341
rect 22922 6332 22928 6344
rect 22980 6332 22986 6384
rect 18138 6264 18144 6316
rect 18196 6304 18202 6316
rect 18601 6307 18659 6313
rect 18601 6304 18613 6307
rect 18196 6276 18613 6304
rect 18196 6264 18202 6276
rect 18601 6273 18613 6276
rect 18647 6273 18659 6307
rect 19426 6304 19432 6316
rect 19387 6276 19432 6304
rect 18601 6267 18659 6273
rect 19426 6264 19432 6276
rect 19484 6264 19490 6316
rect 19794 6264 19800 6316
rect 19852 6304 19858 6316
rect 20254 6304 20260 6316
rect 19852 6276 20024 6304
rect 20215 6276 20260 6304
rect 19852 6264 19858 6276
rect 18322 6236 18328 6248
rect 16540 6208 17724 6236
rect 18283 6208 18328 6236
rect 16540 6196 16546 6208
rect 18322 6196 18328 6208
rect 18380 6196 18386 6248
rect 18506 6236 18512 6248
rect 18467 6208 18512 6236
rect 18506 6196 18512 6208
rect 18564 6196 18570 6248
rect 19705 6239 19763 6245
rect 18616 6208 19656 6236
rect 18616 6180 18644 6208
rect 15344 6140 15516 6168
rect 16025 6171 16083 6177
rect 15344 6128 15350 6140
rect 16025 6137 16037 6171
rect 16071 6168 16083 6171
rect 17770 6168 17776 6180
rect 16071 6140 17776 6168
rect 16071 6137 16083 6140
rect 16025 6131 16083 6137
rect 17770 6128 17776 6140
rect 17828 6128 17834 6180
rect 18598 6128 18604 6180
rect 18656 6128 18662 6180
rect 18966 6168 18972 6180
rect 18927 6140 18972 6168
rect 18966 6128 18972 6140
rect 19024 6128 19030 6180
rect 19628 6168 19656 6208
rect 19705 6205 19717 6239
rect 19751 6236 19763 6239
rect 19886 6236 19892 6248
rect 19751 6208 19892 6236
rect 19751 6205 19763 6208
rect 19705 6199 19763 6205
rect 19886 6196 19892 6208
rect 19944 6196 19950 6248
rect 19996 6245 20024 6276
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20990 6304 20996 6316
rect 20951 6276 20996 6304
rect 20990 6264 20996 6276
rect 21048 6264 21054 6316
rect 19981 6239 20039 6245
rect 19981 6205 19993 6239
rect 20027 6205 20039 6239
rect 19981 6199 20039 6205
rect 20717 6239 20775 6245
rect 20717 6205 20729 6239
rect 20763 6236 20775 6239
rect 21450 6236 21456 6248
rect 20763 6208 21456 6236
rect 20763 6205 20775 6208
rect 20717 6199 20775 6205
rect 20732 6168 20760 6199
rect 21450 6196 21456 6208
rect 21508 6196 21514 6248
rect 19628 6140 20760 6168
rect 9582 6100 9588 6112
rect 9315 6072 9588 6100
rect 8573 6063 8631 6069
rect 9582 6060 9588 6072
rect 9640 6060 9646 6112
rect 10137 6103 10195 6109
rect 10137 6069 10149 6103
rect 10183 6100 10195 6103
rect 10870 6100 10876 6112
rect 10183 6072 10876 6100
rect 10183 6069 10195 6072
rect 10137 6063 10195 6069
rect 10870 6060 10876 6072
rect 10928 6060 10934 6112
rect 11054 6100 11060 6112
rect 11015 6072 11060 6100
rect 11054 6060 11060 6072
rect 11112 6060 11118 6112
rect 11330 6100 11336 6112
rect 11291 6072 11336 6100
rect 11330 6060 11336 6072
rect 11388 6060 11394 6112
rect 13814 6060 13820 6112
rect 13872 6100 13878 6112
rect 14918 6100 14924 6112
rect 13872 6072 14924 6100
rect 13872 6060 13878 6072
rect 14918 6060 14924 6072
rect 14976 6060 14982 6112
rect 15930 6060 15936 6112
rect 15988 6100 15994 6112
rect 16117 6103 16175 6109
rect 16117 6100 16129 6103
rect 15988 6072 16129 6100
rect 15988 6060 15994 6072
rect 16117 6069 16129 6072
rect 16163 6069 16175 6103
rect 16117 6063 16175 6069
rect 16390 6060 16396 6112
rect 16448 6100 16454 6112
rect 16485 6103 16543 6109
rect 16485 6100 16497 6103
rect 16448 6072 16497 6100
rect 16448 6060 16454 6072
rect 16485 6069 16497 6072
rect 16531 6069 16543 6103
rect 16485 6063 16543 6069
rect 16853 6103 16911 6109
rect 16853 6069 16865 6103
rect 16899 6100 16911 6103
rect 20438 6100 20444 6112
rect 16899 6072 20444 6100
rect 16899 6069 16911 6072
rect 16853 6063 16911 6069
rect 20438 6060 20444 6072
rect 20496 6060 20502 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 2130 5896 2136 5908
rect 2091 5868 2136 5896
rect 2130 5856 2136 5868
rect 2188 5856 2194 5908
rect 4246 5896 4252 5908
rect 4207 5868 4252 5896
rect 4246 5856 4252 5868
rect 4304 5856 4310 5908
rect 4890 5856 4896 5908
rect 4948 5896 4954 5908
rect 6089 5899 6147 5905
rect 6089 5896 6101 5899
rect 4948 5868 6101 5896
rect 4948 5856 4954 5868
rect 6089 5865 6101 5868
rect 6135 5865 6147 5899
rect 6089 5859 6147 5865
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 6917 5899 6975 5905
rect 6917 5896 6929 5899
rect 6604 5868 6929 5896
rect 6604 5856 6610 5868
rect 6917 5865 6929 5868
rect 6963 5865 6975 5899
rect 6917 5859 6975 5865
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7466 5896 7472 5908
rect 7064 5868 7472 5896
rect 7064 5856 7070 5868
rect 7466 5856 7472 5868
rect 7524 5856 7530 5908
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 10594 5896 10600 5908
rect 7984 5868 10272 5896
rect 10555 5868 10600 5896
rect 7984 5856 7990 5868
rect 3602 5788 3608 5840
rect 3660 5828 3666 5840
rect 3973 5831 4031 5837
rect 3973 5828 3985 5831
rect 3660 5800 3985 5828
rect 3660 5788 3666 5800
rect 3973 5797 3985 5800
rect 4019 5828 4031 5831
rect 4062 5828 4068 5840
rect 4019 5800 4068 5828
rect 4019 5797 4031 5800
rect 3973 5791 4031 5797
rect 4062 5788 4068 5800
rect 4120 5788 4126 5840
rect 1578 5760 1584 5772
rect 1539 5732 1584 5760
rect 1578 5720 1584 5732
rect 1636 5720 1642 5772
rect 1673 5763 1731 5769
rect 1673 5729 1685 5763
rect 1719 5760 1731 5763
rect 1946 5760 1952 5772
rect 1719 5732 1952 5760
rect 1719 5729 1731 5732
rect 1673 5723 1731 5729
rect 1946 5720 1952 5732
rect 2004 5720 2010 5772
rect 4264 5760 4292 5856
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 6052 5800 8524 5828
rect 6052 5788 6058 5800
rect 8496 5772 8524 5800
rect 9122 5788 9128 5840
rect 9180 5788 9186 5840
rect 6086 5760 6092 5772
rect 3528 5732 4292 5760
rect 5552 5732 6092 5760
rect 3349 5695 3407 5701
rect 3349 5692 3361 5695
rect 2746 5664 3361 5692
rect 2498 5584 2504 5636
rect 2556 5624 2562 5636
rect 2746 5624 2774 5664
rect 3349 5661 3361 5664
rect 3395 5692 3407 5695
rect 3528 5692 3556 5732
rect 3395 5664 3556 5692
rect 3395 5661 3407 5664
rect 3349 5655 3407 5661
rect 3602 5652 3608 5704
rect 3660 5692 3666 5704
rect 3660 5664 3705 5692
rect 3660 5652 3666 5664
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3844 5664 3889 5692
rect 3844 5652 3850 5664
rect 4338 5652 4344 5704
rect 4396 5692 4402 5704
rect 5373 5695 5431 5701
rect 5373 5692 5385 5695
rect 4396 5664 5385 5692
rect 4396 5652 4402 5664
rect 5373 5661 5385 5664
rect 5419 5692 5431 5695
rect 5552 5692 5580 5732
rect 6086 5720 6092 5732
rect 6144 5760 6150 5772
rect 6733 5763 6791 5769
rect 6733 5760 6745 5763
rect 6144 5732 6745 5760
rect 6144 5720 6150 5732
rect 6733 5729 6745 5732
rect 6779 5760 6791 5763
rect 7098 5760 7104 5772
rect 6779 5732 7104 5760
rect 6779 5729 6791 5732
rect 6733 5723 6791 5729
rect 7098 5720 7104 5732
rect 7156 5720 7162 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 7377 5763 7435 5769
rect 7377 5760 7389 5763
rect 7340 5732 7389 5760
rect 7340 5720 7346 5732
rect 7377 5729 7389 5732
rect 7423 5729 7435 5763
rect 7558 5760 7564 5772
rect 7519 5732 7564 5760
rect 7377 5723 7435 5729
rect 7558 5720 7564 5732
rect 7616 5720 7622 5772
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5760 7987 5763
rect 8294 5760 8300 5772
rect 7975 5732 8300 5760
rect 7975 5729 7987 5732
rect 7929 5723 7987 5729
rect 8294 5720 8300 5732
rect 8352 5720 8358 5772
rect 8478 5720 8484 5772
rect 8536 5720 8542 5772
rect 9140 5760 9168 5788
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 9140 5732 9229 5760
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 5419 5664 5580 5692
rect 5629 5695 5687 5701
rect 5419 5661 5431 5664
rect 5373 5655 5431 5661
rect 5629 5661 5641 5695
rect 5675 5661 5687 5695
rect 5629 5655 5687 5661
rect 2556 5596 2774 5624
rect 2556 5584 2562 5596
rect 3970 5584 3976 5636
rect 4028 5624 4034 5636
rect 5644 5624 5672 5655
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 5902 5692 5908 5704
rect 5863 5664 5908 5692
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 6270 5652 6276 5704
rect 6328 5692 6334 5704
rect 6549 5695 6607 5701
rect 6549 5692 6561 5695
rect 6328 5664 6561 5692
rect 6328 5652 6334 5664
rect 6549 5661 6561 5664
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 6914 5652 6920 5704
rect 6972 5692 6978 5704
rect 7742 5692 7748 5704
rect 6972 5664 7748 5692
rect 6972 5652 6978 5664
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 8021 5695 8079 5701
rect 8021 5692 8033 5695
rect 7852 5664 8033 5692
rect 4028 5596 5672 5624
rect 5736 5624 5764 5652
rect 7285 5627 7343 5633
rect 7285 5624 7297 5627
rect 5736 5596 7297 5624
rect 4028 5584 4034 5596
rect 7285 5593 7297 5596
rect 7331 5593 7343 5627
rect 7285 5587 7343 5593
rect 1762 5556 1768 5568
rect 1723 5528 1768 5556
rect 1762 5516 1768 5528
rect 1820 5516 1826 5568
rect 2225 5559 2283 5565
rect 2225 5525 2237 5559
rect 2271 5556 2283 5559
rect 2314 5556 2320 5568
rect 2271 5528 2320 5556
rect 2271 5525 2283 5528
rect 2225 5519 2283 5525
rect 2314 5516 2320 5528
rect 2372 5516 2378 5568
rect 4890 5516 4896 5568
rect 4948 5556 4954 5568
rect 5442 5556 5448 5568
rect 4948 5528 5448 5556
rect 4948 5516 4954 5528
rect 5442 5516 5448 5528
rect 5500 5516 5506 5568
rect 5718 5556 5724 5568
rect 5679 5528 5724 5556
rect 5718 5516 5724 5528
rect 5776 5516 5782 5568
rect 6457 5559 6515 5565
rect 6457 5525 6469 5559
rect 6503 5556 6515 5559
rect 7098 5556 7104 5568
rect 6503 5528 7104 5556
rect 6503 5525 6515 5528
rect 6457 5519 6515 5525
rect 7098 5516 7104 5528
rect 7156 5516 7162 5568
rect 7300 5556 7328 5587
rect 7466 5584 7472 5636
rect 7524 5624 7530 5636
rect 7852 5624 7880 5664
rect 8021 5661 8033 5664
rect 8067 5661 8079 5695
rect 8021 5655 8079 5661
rect 8110 5652 8116 5704
rect 8168 5692 8174 5704
rect 8496 5692 8524 5720
rect 8757 5695 8815 5701
rect 8757 5692 8769 5695
rect 8168 5664 8213 5692
rect 8496 5664 8769 5692
rect 8168 5652 8174 5664
rect 8757 5661 8769 5664
rect 8803 5661 8815 5695
rect 8757 5655 8815 5661
rect 8846 5652 8852 5704
rect 8904 5692 8910 5704
rect 9125 5695 9183 5701
rect 9125 5692 9137 5695
rect 8904 5664 9137 5692
rect 8904 5652 8910 5664
rect 9125 5661 9137 5664
rect 9171 5661 9183 5695
rect 10244 5692 10272 5868
rect 10594 5856 10600 5868
rect 10652 5856 10658 5908
rect 10778 5896 10784 5908
rect 10739 5868 10784 5896
rect 10778 5856 10784 5868
rect 10836 5856 10842 5908
rect 11330 5896 11336 5908
rect 11164 5868 11336 5896
rect 10318 5788 10324 5840
rect 10376 5828 10382 5840
rect 11164 5828 11192 5868
rect 11330 5856 11336 5868
rect 11388 5856 11394 5908
rect 12618 5856 12624 5908
rect 12676 5856 12682 5908
rect 15013 5899 15071 5905
rect 15013 5865 15025 5899
rect 15059 5896 15071 5899
rect 15470 5896 15476 5908
rect 15059 5868 15476 5896
rect 15059 5865 15071 5868
rect 15013 5859 15071 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 17313 5899 17371 5905
rect 17313 5865 17325 5899
rect 17359 5896 17371 5899
rect 18506 5896 18512 5908
rect 17359 5868 18512 5896
rect 17359 5865 17371 5868
rect 17313 5859 17371 5865
rect 18506 5856 18512 5868
rect 18564 5856 18570 5908
rect 19886 5856 19892 5908
rect 19944 5896 19950 5908
rect 20625 5899 20683 5905
rect 20625 5896 20637 5899
rect 19944 5868 20637 5896
rect 19944 5856 19950 5868
rect 20625 5865 20637 5868
rect 20671 5865 20683 5899
rect 20625 5859 20683 5865
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 20898 5896 20904 5908
rect 20763 5868 20904 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 20898 5856 20904 5868
rect 20956 5856 20962 5908
rect 12636 5828 12664 5856
rect 10376 5800 11192 5828
rect 11256 5800 12664 5828
rect 10376 5788 10382 5800
rect 11256 5769 11284 5800
rect 13538 5788 13544 5840
rect 13596 5828 13602 5840
rect 14093 5831 14151 5837
rect 14093 5828 14105 5831
rect 13596 5800 14105 5828
rect 13596 5788 13602 5800
rect 14093 5797 14105 5800
rect 14139 5797 14151 5831
rect 18417 5831 18475 5837
rect 18417 5828 18429 5831
rect 14093 5791 14151 5797
rect 16408 5800 18429 5828
rect 11241 5763 11299 5769
rect 11241 5729 11253 5763
rect 11287 5729 11299 5763
rect 11422 5760 11428 5772
rect 11383 5732 11428 5760
rect 11241 5723 11299 5729
rect 11422 5720 11428 5732
rect 11480 5720 11486 5772
rect 11793 5763 11851 5769
rect 11793 5729 11805 5763
rect 11839 5760 11851 5763
rect 12526 5760 12532 5772
rect 11839 5732 12532 5760
rect 11839 5729 11851 5732
rect 11793 5723 11851 5729
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 12621 5763 12679 5769
rect 12621 5729 12633 5763
rect 12667 5760 12679 5763
rect 12710 5760 12716 5772
rect 12667 5732 12716 5760
rect 12667 5729 12679 5732
rect 12621 5723 12679 5729
rect 12710 5720 12716 5732
rect 12768 5720 12774 5772
rect 12894 5720 12900 5772
rect 12952 5760 12958 5772
rect 14642 5760 14648 5772
rect 12952 5732 14504 5760
rect 14603 5732 14648 5760
rect 12952 5720 12958 5732
rect 11885 5695 11943 5701
rect 11885 5692 11897 5695
rect 10244 5664 11897 5692
rect 9125 5655 9183 5661
rect 11885 5661 11897 5664
rect 11931 5692 11943 5695
rect 13449 5695 13507 5701
rect 11931 5664 13400 5692
rect 11931 5661 11943 5664
rect 11885 5655 11943 5661
rect 9484 5627 9542 5633
rect 7524 5596 7880 5624
rect 8036 5596 9444 5624
rect 7524 5584 7530 5596
rect 8036 5556 8064 5596
rect 7300 5528 8064 5556
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8481 5559 8539 5565
rect 8481 5556 8493 5559
rect 8352 5528 8493 5556
rect 8352 5516 8358 5528
rect 8481 5525 8493 5528
rect 8527 5525 8539 5559
rect 8481 5519 8539 5525
rect 8573 5559 8631 5565
rect 8573 5525 8585 5559
rect 8619 5556 8631 5559
rect 8662 5556 8668 5568
rect 8619 5528 8668 5556
rect 8619 5525 8631 5528
rect 8573 5519 8631 5525
rect 8662 5516 8668 5528
rect 8720 5516 8726 5568
rect 8941 5559 8999 5565
rect 8941 5525 8953 5559
rect 8987 5556 8999 5559
rect 9306 5556 9312 5568
rect 8987 5528 9312 5556
rect 8987 5525 8999 5528
rect 8941 5519 8999 5525
rect 9306 5516 9312 5528
rect 9364 5516 9370 5568
rect 9416 5556 9444 5596
rect 9484 5593 9496 5627
rect 9530 5624 9542 5627
rect 9950 5624 9956 5636
rect 9530 5596 9956 5624
rect 9530 5593 9542 5596
rect 9484 5587 9542 5593
rect 9950 5584 9956 5596
rect 10008 5624 10014 5636
rect 11422 5624 11428 5636
rect 10008 5596 11428 5624
rect 10008 5584 10014 5596
rect 11422 5584 11428 5596
rect 11480 5584 11486 5636
rect 11974 5624 11980 5636
rect 11935 5596 11980 5624
rect 11974 5584 11980 5596
rect 12032 5584 12038 5636
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12492 5596 13308 5624
rect 12492 5584 12498 5596
rect 9858 5556 9864 5568
rect 9416 5528 9864 5556
rect 9858 5516 9864 5528
rect 9916 5516 9922 5568
rect 10410 5516 10416 5568
rect 10468 5556 10474 5568
rect 10594 5556 10600 5568
rect 10468 5528 10600 5556
rect 10468 5516 10474 5528
rect 10594 5516 10600 5528
rect 10652 5556 10658 5568
rect 11149 5559 11207 5565
rect 11149 5556 11161 5559
rect 10652 5528 11161 5556
rect 10652 5516 10658 5528
rect 11149 5525 11161 5528
rect 11195 5525 11207 5559
rect 11149 5519 11207 5525
rect 11238 5516 11244 5568
rect 11296 5556 11302 5568
rect 11698 5556 11704 5568
rect 11296 5528 11704 5556
rect 11296 5516 11302 5528
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12345 5559 12403 5565
rect 12345 5525 12357 5559
rect 12391 5556 12403 5559
rect 12713 5559 12771 5565
rect 12713 5556 12725 5559
rect 12391 5528 12725 5556
rect 12391 5525 12403 5528
rect 12345 5519 12403 5525
rect 12713 5525 12725 5528
rect 12759 5525 12771 5559
rect 12713 5519 12771 5525
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 13170 5556 13176 5568
rect 12860 5528 12905 5556
rect 13131 5528 13176 5556
rect 12860 5516 12866 5528
rect 13170 5516 13176 5528
rect 13228 5516 13234 5568
rect 13280 5565 13308 5596
rect 13265 5559 13323 5565
rect 13265 5525 13277 5559
rect 13311 5525 13323 5559
rect 13372 5556 13400 5664
rect 13449 5661 13461 5695
rect 13495 5661 13507 5695
rect 13449 5655 13507 5661
rect 13725 5695 13783 5701
rect 13725 5661 13737 5695
rect 13771 5692 13783 5695
rect 13814 5692 13820 5704
rect 13771 5664 13820 5692
rect 13771 5661 13783 5664
rect 13725 5655 13783 5661
rect 13464 5624 13492 5655
rect 13814 5652 13820 5664
rect 13872 5652 13878 5704
rect 14476 5692 14504 5732
rect 14642 5720 14648 5732
rect 14700 5720 14706 5772
rect 14734 5720 14740 5772
rect 14792 5760 14798 5772
rect 15102 5760 15108 5772
rect 14792 5732 15108 5760
rect 14792 5720 14798 5732
rect 15102 5720 15108 5732
rect 15160 5720 15166 5772
rect 14553 5695 14611 5701
rect 14553 5692 14565 5695
rect 14476 5664 14565 5692
rect 14553 5661 14565 5664
rect 14599 5692 14611 5695
rect 15372 5695 15430 5701
rect 14599 5664 15240 5692
rect 14599 5661 14611 5664
rect 14553 5655 14611 5661
rect 14274 5624 14280 5636
rect 13464 5596 14280 5624
rect 14274 5584 14280 5596
rect 14332 5584 14338 5636
rect 15010 5624 15016 5636
rect 14384 5596 15016 5624
rect 13541 5559 13599 5565
rect 13541 5556 13553 5559
rect 13372 5528 13553 5556
rect 13265 5519 13323 5525
rect 13541 5525 13553 5528
rect 13587 5556 13599 5559
rect 13630 5556 13636 5568
rect 13587 5528 13636 5556
rect 13587 5525 13599 5528
rect 13541 5519 13599 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13909 5559 13967 5565
rect 13909 5525 13921 5559
rect 13955 5556 13967 5559
rect 14384 5556 14412 5596
rect 15010 5584 15016 5596
rect 15068 5584 15074 5636
rect 15212 5624 15240 5664
rect 15372 5661 15384 5695
rect 15418 5692 15430 5695
rect 15838 5692 15844 5704
rect 15418 5664 15844 5692
rect 15418 5661 15430 5664
rect 15372 5655 15430 5661
rect 15838 5652 15844 5664
rect 15896 5652 15902 5704
rect 16408 5624 16436 5800
rect 18417 5797 18429 5800
rect 18463 5797 18475 5831
rect 18782 5828 18788 5840
rect 18743 5800 18788 5828
rect 18417 5791 18475 5797
rect 18782 5788 18788 5800
rect 18840 5788 18846 5840
rect 16669 5763 16727 5769
rect 16669 5760 16681 5763
rect 15212 5596 16436 5624
rect 16500 5732 16681 5760
rect 13955 5528 14412 5556
rect 14461 5559 14519 5565
rect 13955 5525 13967 5528
rect 13909 5519 13967 5525
rect 14461 5525 14473 5559
rect 14507 5556 14519 5559
rect 14550 5556 14556 5568
rect 14507 5528 14556 5556
rect 14507 5525 14519 5528
rect 14461 5519 14519 5525
rect 14550 5516 14556 5528
rect 14608 5516 14614 5568
rect 16298 5516 16304 5568
rect 16356 5556 16362 5568
rect 16500 5565 16528 5732
rect 16669 5729 16681 5732
rect 16715 5729 16727 5763
rect 16669 5723 16727 5729
rect 16853 5763 16911 5769
rect 16853 5729 16865 5763
rect 16899 5760 16911 5763
rect 16942 5760 16948 5772
rect 16899 5732 16948 5760
rect 16899 5729 16911 5732
rect 16853 5723 16911 5729
rect 16942 5720 16948 5732
rect 17000 5720 17006 5772
rect 18049 5763 18107 5769
rect 18049 5729 18061 5763
rect 18095 5760 18107 5763
rect 18230 5760 18236 5772
rect 18095 5732 18236 5760
rect 18095 5729 18107 5732
rect 18049 5723 18107 5729
rect 18230 5720 18236 5732
rect 18288 5720 18294 5772
rect 18874 5720 18880 5772
rect 18932 5760 18938 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18932 5732 19257 5760
rect 18932 5720 18938 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5760 21419 5763
rect 21542 5760 21548 5772
rect 21407 5732 21548 5760
rect 21407 5729 21419 5732
rect 21361 5723 21419 5729
rect 21542 5720 21548 5732
rect 21600 5720 21606 5772
rect 17770 5692 17776 5704
rect 17731 5664 17776 5692
rect 17770 5652 17776 5664
rect 17828 5652 17834 5704
rect 18969 5695 19027 5701
rect 17972 5664 18460 5692
rect 16945 5627 17003 5633
rect 16945 5593 16957 5627
rect 16991 5624 17003 5627
rect 16991 5596 17448 5624
rect 16991 5593 17003 5596
rect 16945 5587 17003 5593
rect 17420 5565 17448 5596
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 17972 5624 18000 5664
rect 17736 5596 18000 5624
rect 17736 5584 17742 5596
rect 18046 5584 18052 5636
rect 18104 5624 18110 5636
rect 18233 5627 18291 5633
rect 18233 5624 18245 5627
rect 18104 5596 18245 5624
rect 18104 5584 18110 5596
rect 18233 5593 18245 5596
rect 18279 5593 18291 5627
rect 18233 5587 18291 5593
rect 16485 5559 16543 5565
rect 16485 5556 16497 5559
rect 16356 5528 16497 5556
rect 16356 5516 16362 5528
rect 16485 5525 16497 5528
rect 16531 5525 16543 5559
rect 16485 5519 16543 5525
rect 17405 5559 17463 5565
rect 17405 5525 17417 5559
rect 17451 5525 17463 5559
rect 17405 5519 17463 5525
rect 17862 5516 17868 5568
rect 17920 5556 17926 5568
rect 18432 5556 18460 5664
rect 18969 5661 18981 5695
rect 19015 5692 19027 5695
rect 19334 5692 19340 5704
rect 19015 5664 19340 5692
rect 19015 5661 19027 5664
rect 18969 5655 19027 5661
rect 19334 5652 19340 5664
rect 19392 5652 19398 5704
rect 21082 5692 21088 5704
rect 21043 5664 21088 5692
rect 21082 5652 21088 5664
rect 21140 5652 21146 5704
rect 18598 5624 18604 5636
rect 18559 5596 18604 5624
rect 18598 5584 18604 5596
rect 18656 5584 18662 5636
rect 19512 5627 19570 5633
rect 19512 5593 19524 5627
rect 19558 5624 19570 5627
rect 19886 5624 19892 5636
rect 19558 5596 19892 5624
rect 19558 5593 19570 5596
rect 19512 5587 19570 5593
rect 19886 5584 19892 5596
rect 19944 5584 19950 5636
rect 21177 5559 21235 5565
rect 21177 5556 21189 5559
rect 17920 5528 17965 5556
rect 18432 5528 21189 5556
rect 17920 5516 17926 5528
rect 21177 5525 21189 5528
rect 21223 5525 21235 5559
rect 21177 5519 21235 5525
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 3050 5352 3056 5364
rect 1627 5324 3056 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 3234 5352 3240 5364
rect 3195 5324 3240 5352
rect 3234 5312 3240 5324
rect 3292 5312 3298 5364
rect 3970 5312 3976 5364
rect 4028 5352 4034 5364
rect 5718 5352 5724 5364
rect 4028 5324 5724 5352
rect 4028 5312 4034 5324
rect 5718 5312 5724 5324
rect 5776 5312 5782 5364
rect 6181 5355 6239 5361
rect 6181 5321 6193 5355
rect 6227 5352 6239 5355
rect 6638 5352 6644 5364
rect 6227 5324 6644 5352
rect 6227 5321 6239 5324
rect 6181 5315 6239 5321
rect 1486 5284 1492 5296
rect 1447 5256 1492 5284
rect 1486 5244 1492 5256
rect 1544 5244 1550 5296
rect 3602 5284 3608 5296
rect 2056 5256 3608 5284
rect 2056 5216 2084 5256
rect 3602 5244 3608 5256
rect 3660 5284 3666 5296
rect 4154 5284 4160 5296
rect 3660 5256 4160 5284
rect 3660 5244 3666 5256
rect 4154 5244 4160 5256
rect 4212 5284 4218 5296
rect 4212 5256 5028 5284
rect 4212 5244 4218 5256
rect 2130 5225 2136 5228
rect 1872 5188 2084 5216
rect 1872 5157 1900 5188
rect 2124 5179 2136 5225
rect 2188 5216 2194 5228
rect 2590 5216 2596 5228
rect 2188 5188 2596 5216
rect 2130 5176 2136 5179
rect 2188 5176 2194 5188
rect 2590 5176 2596 5188
rect 2648 5176 2654 5228
rect 3050 5176 3056 5228
rect 3108 5216 3114 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3108 5188 3341 5216
rect 3108 5176 3114 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 5000 5225 5028 5256
rect 5166 5244 5172 5296
rect 5224 5284 5230 5296
rect 6196 5284 6224 5315
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 8110 5312 8116 5364
rect 8168 5352 8174 5364
rect 8297 5355 8355 5361
rect 8297 5352 8309 5355
rect 8168 5324 8309 5352
rect 8168 5312 8174 5324
rect 8297 5321 8309 5324
rect 8343 5321 8355 5355
rect 10413 5355 10471 5361
rect 10413 5352 10425 5355
rect 8297 5315 8355 5321
rect 9232 5324 10425 5352
rect 5224 5256 6224 5284
rect 7500 5287 7558 5293
rect 5224 5244 5230 5256
rect 7500 5253 7512 5287
rect 7546 5284 7558 5287
rect 9232 5284 9260 5324
rect 10413 5321 10425 5324
rect 10459 5321 10471 5355
rect 10413 5315 10471 5321
rect 10781 5355 10839 5361
rect 10781 5321 10793 5355
rect 10827 5352 10839 5355
rect 11054 5352 11060 5364
rect 10827 5324 11060 5352
rect 10827 5321 10839 5324
rect 10781 5315 10839 5321
rect 7546 5256 9260 5284
rect 9300 5287 9358 5293
rect 7546 5253 7558 5256
rect 7500 5247 7558 5253
rect 9300 5253 9312 5287
rect 9346 5284 9358 5287
rect 9766 5284 9772 5296
rect 9346 5256 9772 5284
rect 9346 5253 9358 5256
rect 9300 5247 9358 5253
rect 9766 5244 9772 5256
rect 9824 5244 9830 5296
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3936 5188 4077 5216
rect 3936 5176 3942 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4985 5219 5043 5225
rect 4985 5185 4997 5219
rect 5031 5185 5043 5219
rect 4985 5179 5043 5185
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 5592 5188 5637 5216
rect 5592 5176 5598 5188
rect 5902 5176 5908 5228
rect 5960 5216 5966 5228
rect 5997 5219 6055 5225
rect 5997 5216 6009 5219
rect 5960 5188 6009 5216
rect 5960 5176 5966 5188
rect 5997 5185 6009 5188
rect 6043 5185 6055 5219
rect 5997 5179 6055 5185
rect 7650 5176 7656 5228
rect 7708 5216 7714 5228
rect 7745 5219 7803 5225
rect 7745 5216 7757 5219
rect 7708 5188 7757 5216
rect 7708 5176 7714 5188
rect 7745 5185 7757 5188
rect 7791 5185 7803 5219
rect 7745 5179 7803 5185
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 1857 5151 1915 5157
rect 1857 5117 1869 5151
rect 1903 5117 1915 5151
rect 1857 5111 1915 5117
rect 1872 5012 1900 5111
rect 3234 5108 3240 5160
rect 3292 5148 3298 5160
rect 4157 5151 4215 5157
rect 4157 5148 4169 5151
rect 3292 5120 4169 5148
rect 3292 5108 3298 5120
rect 4157 5117 4169 5120
rect 4203 5117 4215 5151
rect 4338 5148 4344 5160
rect 4299 5120 4344 5148
rect 4157 5111 4215 5117
rect 4338 5108 4344 5120
rect 4396 5108 4402 5160
rect 4522 5148 4528 5160
rect 4483 5120 4528 5148
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 5353 5151 5411 5157
rect 5353 5117 5365 5151
rect 5399 5117 5411 5151
rect 5353 5111 5411 5117
rect 5445 5151 5503 5157
rect 5445 5117 5457 5151
rect 5491 5148 5503 5151
rect 6730 5148 6736 5160
rect 5491 5120 6736 5148
rect 5491 5117 5503 5120
rect 5445 5111 5503 5117
rect 3697 5083 3755 5089
rect 3697 5080 3709 5083
rect 3160 5052 3709 5080
rect 2130 5012 2136 5024
rect 1872 4984 2136 5012
rect 2130 4972 2136 4984
rect 2188 4972 2194 5024
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 3160 5012 3188 5052
rect 3697 5049 3709 5052
rect 3743 5049 3755 5083
rect 4982 5080 4988 5092
rect 3697 5043 3755 5049
rect 4356 5052 4988 5080
rect 2648 4984 3188 5012
rect 3513 5015 3571 5021
rect 2648 4972 2654 4984
rect 3513 4981 3525 5015
rect 3559 5012 3571 5015
rect 4356 5012 4384 5052
rect 4982 5040 4988 5052
rect 5040 5040 5046 5092
rect 5368 5080 5396 5111
rect 6730 5108 6736 5120
rect 6788 5108 6794 5160
rect 7926 5108 7932 5160
rect 7984 5148 7990 5160
rect 8220 5148 8248 5179
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8849 5219 8907 5225
rect 8849 5216 8861 5219
rect 8352 5188 8861 5216
rect 8352 5176 8358 5188
rect 8849 5185 8861 5188
rect 8895 5185 8907 5219
rect 9030 5216 9036 5228
rect 8991 5188 9036 5216
rect 8849 5179 8907 5185
rect 7984 5120 8248 5148
rect 8389 5151 8447 5157
rect 7984 5108 7990 5120
rect 8389 5117 8401 5151
rect 8435 5117 8447 5151
rect 8864 5148 8892 5179
rect 9030 5176 9036 5188
rect 9088 5176 9094 5228
rect 10226 5216 10232 5228
rect 9140 5188 10232 5216
rect 9140 5148 9168 5188
rect 10226 5176 10232 5188
rect 10284 5176 10290 5228
rect 8864 5120 9168 5148
rect 10428 5148 10456 5315
rect 11054 5312 11060 5324
rect 11112 5312 11118 5364
rect 11241 5355 11299 5361
rect 11241 5321 11253 5355
rect 11287 5321 11299 5355
rect 11241 5315 11299 5321
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5352 11575 5355
rect 11882 5352 11888 5364
rect 11563 5324 11888 5352
rect 11563 5321 11575 5324
rect 11517 5315 11575 5321
rect 10870 5284 10876 5296
rect 10831 5256 10876 5284
rect 10870 5244 10876 5256
rect 10928 5244 10934 5296
rect 11256 5284 11284 5315
rect 11882 5312 11888 5324
rect 11940 5312 11946 5364
rect 12161 5355 12219 5361
rect 12161 5321 12173 5355
rect 12207 5352 12219 5355
rect 12250 5352 12256 5364
rect 12207 5324 12256 5352
rect 12207 5321 12219 5324
rect 12161 5315 12219 5321
rect 12250 5312 12256 5324
rect 12308 5312 12314 5364
rect 13630 5312 13636 5364
rect 13688 5352 13694 5364
rect 14461 5355 14519 5361
rect 13688 5324 13952 5352
rect 13688 5312 13694 5324
rect 11330 5284 11336 5296
rect 11256 5256 11336 5284
rect 11330 5244 11336 5256
rect 11388 5244 11394 5296
rect 11422 5244 11428 5296
rect 11480 5284 11486 5296
rect 12526 5284 12532 5296
rect 11480 5256 12532 5284
rect 11480 5244 11486 5256
rect 11701 5219 11759 5225
rect 11882 5220 11888 5228
rect 11701 5185 11713 5219
rect 11747 5216 11759 5219
rect 11808 5216 11888 5220
rect 11747 5192 11888 5216
rect 11747 5188 11836 5192
rect 11880 5188 11888 5192
rect 11747 5185 11759 5188
rect 11701 5179 11759 5185
rect 11882 5176 11888 5188
rect 11940 5176 11946 5228
rect 11992 5157 12020 5256
rect 12526 5244 12532 5256
rect 12584 5284 12590 5296
rect 13722 5284 13728 5296
rect 13780 5293 13786 5296
rect 12584 5256 13728 5284
rect 12584 5244 12590 5256
rect 13722 5244 13728 5256
rect 13780 5247 13792 5293
rect 13924 5284 13952 5324
rect 14461 5321 14473 5355
rect 14507 5352 14519 5355
rect 14918 5352 14924 5364
rect 14507 5324 14924 5352
rect 14507 5321 14519 5324
rect 14461 5315 14519 5321
rect 14918 5312 14924 5324
rect 14976 5312 14982 5364
rect 15286 5352 15292 5364
rect 15247 5324 15292 5352
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15703 5324 16037 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 16485 5355 16543 5361
rect 16485 5321 16497 5355
rect 16531 5352 16543 5355
rect 16945 5355 17003 5361
rect 16945 5352 16957 5355
rect 16531 5324 16957 5352
rect 16531 5321 16543 5324
rect 16485 5315 16543 5321
rect 16945 5321 16957 5324
rect 16991 5321 17003 5355
rect 16945 5315 17003 5321
rect 17037 5355 17095 5361
rect 17037 5321 17049 5355
rect 17083 5352 17095 5355
rect 17402 5352 17408 5364
rect 17083 5324 17408 5352
rect 17083 5321 17095 5324
rect 17037 5315 17095 5321
rect 17402 5312 17408 5324
rect 17460 5312 17466 5364
rect 17497 5355 17555 5361
rect 17497 5321 17509 5355
rect 17543 5352 17555 5355
rect 17862 5352 17868 5364
rect 17543 5324 17868 5352
rect 17543 5321 17555 5324
rect 17497 5315 17555 5321
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 17957 5355 18015 5361
rect 17957 5321 17969 5355
rect 18003 5352 18015 5355
rect 19797 5355 19855 5361
rect 18003 5324 19564 5352
rect 18003 5321 18015 5324
rect 17957 5315 18015 5321
rect 15562 5284 15568 5296
rect 13924 5256 15568 5284
rect 13780 5244 13786 5247
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 15746 5244 15752 5296
rect 15804 5284 15810 5296
rect 16117 5287 16175 5293
rect 16117 5284 16129 5287
rect 15804 5256 16129 5284
rect 15804 5244 15810 5256
rect 16117 5253 16129 5256
rect 16163 5253 16175 5287
rect 18874 5284 18880 5296
rect 16117 5247 16175 5253
rect 18340 5256 18880 5284
rect 12434 5176 12440 5228
rect 12492 5216 12498 5228
rect 14553 5219 14611 5225
rect 12492 5188 14412 5216
rect 12492 5176 12498 5188
rect 10597 5151 10655 5157
rect 10597 5148 10609 5151
rect 10428 5120 10609 5148
rect 8389 5111 8447 5117
rect 10597 5117 10609 5120
rect 10643 5117 10655 5151
rect 10597 5111 10655 5117
rect 11977 5151 12035 5157
rect 11977 5117 11989 5151
rect 12023 5117 12035 5151
rect 11977 5111 12035 5117
rect 12069 5151 12127 5157
rect 12069 5117 12081 5151
rect 12115 5117 12127 5151
rect 12069 5111 12127 5117
rect 14001 5151 14059 5157
rect 14001 5117 14013 5151
rect 14047 5148 14059 5151
rect 14274 5148 14280 5160
rect 14047 5120 14280 5148
rect 14047 5117 14059 5120
rect 14001 5111 14059 5117
rect 5626 5080 5632 5092
rect 5368 5052 5632 5080
rect 5626 5040 5632 5052
rect 5684 5040 5690 5092
rect 5810 5040 5816 5092
rect 5868 5080 5874 5092
rect 5868 5052 6868 5080
rect 5868 5040 5874 5052
rect 6840 5024 6868 5052
rect 8202 5040 8208 5092
rect 8260 5080 8266 5092
rect 8404 5080 8432 5111
rect 8260 5052 8432 5080
rect 8260 5040 8266 5052
rect 3559 4984 4384 5012
rect 3559 4981 3571 4984
rect 3513 4975 3571 4981
rect 4430 4972 4436 5024
rect 4488 5012 4494 5024
rect 4801 5015 4859 5021
rect 4801 5012 4813 5015
rect 4488 4984 4813 5012
rect 4488 4972 4494 4984
rect 4801 4981 4813 4984
rect 4847 4981 4859 5015
rect 5902 5012 5908 5024
rect 5863 4984 5908 5012
rect 4801 4975 4859 4981
rect 5902 4972 5908 4984
rect 5960 4972 5966 5024
rect 6086 4972 6092 5024
rect 6144 5012 6150 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 6144 4984 6377 5012
rect 6144 4972 6150 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6365 4975 6423 4981
rect 6822 4972 6828 5024
rect 6880 5012 6886 5024
rect 7466 5012 7472 5024
rect 6880 4984 7472 5012
rect 6880 4972 6886 4984
rect 7466 4972 7472 4984
rect 7524 4972 7530 5024
rect 7834 5012 7840 5024
rect 7795 4984 7840 5012
rect 7834 4972 7840 4984
rect 7892 4972 7898 5024
rect 8478 4972 8484 5024
rect 8536 5012 8542 5024
rect 8665 5015 8723 5021
rect 8665 5012 8677 5015
rect 8536 4984 8677 5012
rect 8536 4972 8542 4984
rect 8665 4981 8677 4984
rect 8711 5012 8723 5015
rect 9398 5012 9404 5024
rect 8711 4984 9404 5012
rect 8711 4981 8723 4984
rect 8665 4975 8723 4981
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 9766 4972 9772 5024
rect 9824 5012 9830 5024
rect 12084 5012 12112 5111
rect 14274 5108 14280 5120
rect 14332 5108 14338 5160
rect 14384 5080 14412 5188
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 14918 5216 14924 5228
rect 14599 5188 14924 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 14918 5176 14924 5188
rect 14976 5176 14982 5228
rect 15378 5216 15384 5228
rect 15120 5188 15384 5216
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 15120 5157 15148 5188
rect 15378 5176 15384 5188
rect 15436 5176 15442 5228
rect 17678 5176 17684 5228
rect 17736 5216 17742 5228
rect 17865 5219 17923 5225
rect 17865 5216 17877 5219
rect 17736 5188 17877 5216
rect 17736 5176 17742 5188
rect 17865 5185 17877 5188
rect 17911 5185 17923 5219
rect 17865 5179 17923 5185
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 18340 5225 18368 5256
rect 18874 5244 18880 5256
rect 18932 5244 18938 5296
rect 19536 5284 19564 5324
rect 19797 5321 19809 5355
rect 19843 5352 19855 5355
rect 20070 5352 20076 5364
rect 19843 5324 20076 5352
rect 19843 5321 19855 5324
rect 19797 5315 19855 5321
rect 20070 5312 20076 5324
rect 20128 5312 20134 5364
rect 20162 5312 20168 5364
rect 20220 5352 20226 5364
rect 20220 5324 20265 5352
rect 20220 5312 20226 5324
rect 22554 5284 22560 5296
rect 19536 5256 22560 5284
rect 22554 5244 22560 5256
rect 22612 5244 22618 5296
rect 18325 5219 18383 5225
rect 18325 5216 18337 5219
rect 18288 5188 18337 5216
rect 18288 5176 18294 5188
rect 18325 5185 18337 5188
rect 18371 5185 18383 5219
rect 18325 5179 18383 5185
rect 18592 5219 18650 5225
rect 18592 5185 18604 5219
rect 18638 5216 18650 5219
rect 18966 5216 18972 5228
rect 18638 5188 18972 5216
rect 18638 5185 18650 5188
rect 18592 5179 18650 5185
rect 18966 5176 18972 5188
rect 19024 5176 19030 5228
rect 20257 5219 20315 5225
rect 20257 5185 20269 5219
rect 20303 5216 20315 5219
rect 20622 5216 20628 5228
rect 20303 5188 20628 5216
rect 20303 5185 20315 5188
rect 20257 5179 20315 5185
rect 20622 5176 20628 5188
rect 20680 5176 20686 5228
rect 20717 5219 20775 5225
rect 20717 5185 20729 5219
rect 20763 5216 20775 5219
rect 21910 5216 21916 5228
rect 20763 5188 21916 5216
rect 20763 5185 20775 5188
rect 20717 5179 20775 5185
rect 21910 5176 21916 5188
rect 21968 5176 21974 5228
rect 15105 5151 15163 5157
rect 14700 5120 14745 5148
rect 14700 5108 14706 5120
rect 15105 5117 15117 5151
rect 15151 5117 15163 5151
rect 15105 5111 15163 5117
rect 15197 5151 15255 5157
rect 15197 5117 15209 5151
rect 15243 5148 15255 5151
rect 15286 5148 15292 5160
rect 15243 5120 15292 5148
rect 15243 5117 15255 5120
rect 15197 5111 15255 5117
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 15838 5148 15844 5160
rect 15799 5120 15844 5148
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16298 5108 16304 5160
rect 16356 5148 16362 5160
rect 16482 5148 16488 5160
rect 16356 5120 16488 5148
rect 16356 5108 16362 5120
rect 16482 5108 16488 5120
rect 16540 5148 16546 5160
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16540 5120 16773 5148
rect 16540 5108 16546 5120
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 18049 5151 18107 5157
rect 18049 5148 18061 5151
rect 17276 5120 18061 5148
rect 17276 5108 17282 5120
rect 18049 5117 18061 5120
rect 18095 5117 18107 5151
rect 18049 5111 18107 5117
rect 20441 5151 20499 5157
rect 20441 5117 20453 5151
rect 20487 5117 20499 5151
rect 20990 5148 20996 5160
rect 20951 5120 20996 5148
rect 20441 5111 20499 5117
rect 15470 5080 15476 5092
rect 14384 5052 15476 5080
rect 15470 5040 15476 5052
rect 15528 5040 15534 5092
rect 17405 5083 17463 5089
rect 17405 5049 17417 5083
rect 17451 5080 17463 5083
rect 18138 5080 18144 5092
rect 17451 5052 18144 5080
rect 17451 5049 17463 5052
rect 17405 5043 17463 5049
rect 18138 5040 18144 5052
rect 18196 5040 18202 5092
rect 19705 5083 19763 5089
rect 19705 5049 19717 5083
rect 19751 5080 19763 5083
rect 19886 5080 19892 5092
rect 19751 5052 19892 5080
rect 19751 5049 19763 5052
rect 19705 5043 19763 5049
rect 19886 5040 19892 5052
rect 19944 5040 19950 5092
rect 20456 5080 20484 5111
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 21358 5080 21364 5092
rect 20456 5052 21364 5080
rect 21358 5040 21364 5052
rect 21416 5040 21422 5092
rect 12526 5012 12532 5024
rect 9824 4984 12112 5012
rect 12487 4984 12532 5012
rect 9824 4972 9830 4984
rect 12526 4972 12532 4984
rect 12584 4972 12590 5024
rect 12621 5015 12679 5021
rect 12621 4981 12633 5015
rect 12667 5012 12679 5015
rect 12710 5012 12716 5024
rect 12667 4984 12716 5012
rect 12667 4981 12679 4984
rect 12621 4975 12679 4981
rect 12710 4972 12716 4984
rect 12768 4972 12774 5024
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 14093 5015 14151 5021
rect 14093 5012 14105 5015
rect 13688 4984 14105 5012
rect 13688 4972 13694 4984
rect 14093 4981 14105 4984
rect 14139 4981 14151 5015
rect 14093 4975 14151 4981
rect 15378 4972 15384 5024
rect 15436 5012 15442 5024
rect 15654 5012 15660 5024
rect 15436 4984 15660 5012
rect 15436 4972 15442 4984
rect 15654 4972 15660 4984
rect 15712 4972 15718 5024
rect 17494 4972 17500 5024
rect 17552 5012 17558 5024
rect 20898 5012 20904 5024
rect 17552 4984 20904 5012
rect 17552 4972 17558 4984
rect 20898 4972 20904 4984
rect 20956 4972 20962 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 1762 4768 1768 4820
rect 1820 4808 1826 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 1820 4780 2881 4808
rect 1820 4768 1826 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 4614 4808 4620 4820
rect 4575 4780 4620 4808
rect 2869 4771 2927 4777
rect 4614 4768 4620 4780
rect 4672 4768 4678 4820
rect 5902 4768 5908 4820
rect 5960 4808 5966 4820
rect 5960 4780 9628 4808
rect 5960 4768 5966 4780
rect 5997 4743 6055 4749
rect 5997 4709 6009 4743
rect 6043 4740 6055 4743
rect 6043 4712 6500 4740
rect 6043 4709 6055 4712
rect 5997 4703 6055 4709
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 3421 4675 3479 4681
rect 3421 4672 3433 4675
rect 3016 4644 3433 4672
rect 3016 4632 3022 4644
rect 3421 4641 3433 4644
rect 3467 4641 3479 4675
rect 4338 4672 4344 4684
rect 4299 4644 4344 4672
rect 3421 4635 3479 4641
rect 4338 4632 4344 4644
rect 4396 4632 4402 4684
rect 5442 4672 5448 4684
rect 5355 4644 5448 4672
rect 5442 4632 5448 4644
rect 5500 4672 5506 4684
rect 6086 4672 6092 4684
rect 5500 4644 6092 4672
rect 5500 4632 5506 4644
rect 6086 4632 6092 4644
rect 6144 4632 6150 4684
rect 2130 4564 2136 4616
rect 2188 4604 2194 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2188 4576 2789 4604
rect 2188 4564 2194 4576
rect 2777 4573 2789 4576
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3237 4607 3295 4613
rect 3237 4573 3249 4607
rect 3283 4604 3295 4607
rect 3326 4604 3332 4616
rect 3283 4576 3332 4604
rect 3283 4573 3295 4576
rect 3237 4567 3295 4573
rect 3326 4564 3332 4576
rect 3384 4564 3390 4616
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4604 4215 4607
rect 4522 4604 4528 4616
rect 4203 4576 4528 4604
rect 4203 4573 4215 4576
rect 4157 4567 4215 4573
rect 4522 4564 4528 4576
rect 4580 4564 4586 4616
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4604 4859 4607
rect 5258 4604 5264 4616
rect 4847 4576 5264 4604
rect 4847 4573 4859 4576
rect 4801 4567 4859 4573
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5534 4604 5540 4616
rect 5495 4576 5540 4604
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 6362 4604 6368 4616
rect 6323 4576 6368 4604
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 2532 4539 2590 4545
rect 2532 4505 2544 4539
rect 2578 4536 2590 4539
rect 2958 4536 2964 4548
rect 2578 4508 2964 4536
rect 2578 4505 2590 4508
rect 2532 4499 2590 4505
rect 2958 4496 2964 4508
rect 3016 4496 3022 4548
rect 4246 4536 4252 4548
rect 3344 4508 4252 4536
rect 1397 4471 1455 4477
rect 1397 4437 1409 4471
rect 1443 4468 1455 4471
rect 2038 4468 2044 4480
rect 1443 4440 2044 4468
rect 1443 4437 1455 4440
rect 1397 4431 1455 4437
rect 2038 4428 2044 4440
rect 2096 4428 2102 4480
rect 3344 4477 3372 4508
rect 4246 4496 4252 4508
rect 4304 4496 4310 4548
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 4893 4539 4951 4545
rect 4893 4536 4905 4539
rect 4396 4508 4905 4536
rect 4396 4496 4402 4508
rect 4893 4505 4905 4508
rect 4939 4505 4951 4539
rect 4893 4499 4951 4505
rect 5077 4539 5135 4545
rect 5077 4505 5089 4539
rect 5123 4536 5135 4539
rect 5350 4536 5356 4548
rect 5123 4508 5356 4536
rect 5123 4505 5135 4508
rect 5077 4499 5135 4505
rect 5350 4496 5356 4508
rect 5408 4496 5414 4548
rect 6472 4536 6500 4712
rect 6638 4700 6644 4752
rect 6696 4740 6702 4752
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 6696 4712 7205 4740
rect 6696 4700 6702 4712
rect 7193 4709 7205 4712
rect 7239 4709 7251 4743
rect 8478 4740 8484 4752
rect 7193 4703 7251 4709
rect 7668 4712 8484 4740
rect 7006 4672 7012 4684
rect 6967 4644 7012 4672
rect 7006 4632 7012 4644
rect 7064 4632 7070 4684
rect 7668 4681 7696 4712
rect 8478 4700 8484 4712
rect 8536 4700 8542 4752
rect 8941 4743 8999 4749
rect 8941 4709 8953 4743
rect 8987 4740 8999 4743
rect 9306 4740 9312 4752
rect 8987 4712 9312 4740
rect 8987 4709 8999 4712
rect 8941 4703 8999 4709
rect 9306 4700 9312 4712
rect 9364 4700 9370 4752
rect 9600 4740 9628 4780
rect 9674 4768 9680 4820
rect 9732 4808 9738 4820
rect 10045 4811 10103 4817
rect 10045 4808 10057 4811
rect 9732 4780 10057 4808
rect 9732 4768 9738 4780
rect 10045 4777 10057 4780
rect 10091 4777 10103 4811
rect 10045 4771 10103 4777
rect 10870 4768 10876 4820
rect 10928 4808 10934 4820
rect 11054 4808 11060 4820
rect 10928 4780 11060 4808
rect 10928 4768 10934 4780
rect 11054 4768 11060 4780
rect 11112 4768 11118 4820
rect 11422 4768 11428 4820
rect 11480 4768 11486 4820
rect 11882 4768 11888 4820
rect 11940 4808 11946 4820
rect 12342 4808 12348 4820
rect 11940 4780 12348 4808
rect 11940 4768 11946 4780
rect 12342 4768 12348 4780
rect 12400 4768 12406 4820
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 12802 4808 12808 4820
rect 12492 4780 12808 4808
rect 12492 4768 12498 4780
rect 12802 4768 12808 4780
rect 12860 4768 12866 4820
rect 12894 4768 12900 4820
rect 12952 4808 12958 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12952 4780 13093 4808
rect 12952 4768 12958 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13446 4768 13452 4820
rect 13504 4808 13510 4820
rect 17037 4811 17095 4817
rect 13504 4780 15056 4808
rect 13504 4768 13510 4780
rect 11149 4743 11207 4749
rect 9600 4712 10456 4740
rect 7653 4675 7711 4681
rect 7653 4641 7665 4675
rect 7699 4641 7711 4675
rect 7653 4635 7711 4641
rect 7745 4675 7803 4681
rect 7745 4641 7757 4675
rect 7791 4641 7803 4675
rect 7745 4635 7803 4641
rect 6546 4564 6552 4616
rect 6604 4604 6610 4616
rect 7760 4604 7788 4635
rect 8202 4632 8208 4684
rect 8260 4672 8266 4684
rect 8573 4675 8631 4681
rect 8573 4672 8585 4675
rect 8260 4644 8585 4672
rect 8260 4632 8266 4644
rect 8573 4641 8585 4644
rect 8619 4641 8631 4675
rect 8573 4635 8631 4641
rect 9493 4675 9551 4681
rect 9493 4641 9505 4675
rect 9539 4672 9551 4675
rect 9950 4672 9956 4684
rect 9539 4644 9956 4672
rect 9539 4641 9551 4644
rect 9493 4635 9551 4641
rect 9950 4632 9956 4644
rect 10008 4632 10014 4684
rect 10042 4632 10048 4684
rect 10100 4672 10106 4684
rect 10226 4672 10232 4684
rect 10100 4644 10232 4672
rect 10100 4632 10106 4644
rect 10226 4632 10232 4644
rect 10284 4632 10290 4684
rect 10428 4681 10456 4712
rect 11149 4709 11161 4743
rect 11195 4709 11207 4743
rect 11149 4703 11207 4709
rect 10413 4675 10471 4681
rect 10413 4641 10425 4675
rect 10459 4641 10471 4675
rect 10413 4635 10471 4641
rect 7926 4604 7932 4616
rect 6604 4576 7932 4604
rect 6604 4564 6610 4576
rect 7926 4564 7932 4576
rect 7984 4564 7990 4616
rect 10505 4607 10563 4613
rect 10505 4604 10517 4607
rect 8312 4576 10517 4604
rect 8312 4536 8340 4576
rect 10505 4573 10517 4576
rect 10551 4573 10563 4607
rect 10962 4604 10968 4616
rect 10923 4576 10968 4604
rect 10505 4567 10563 4573
rect 10962 4564 10968 4576
rect 11020 4564 11026 4616
rect 11164 4604 11192 4703
rect 11440 4681 11468 4768
rect 12158 4740 12164 4752
rect 12119 4712 12164 4740
rect 12158 4700 12164 4712
rect 12216 4740 12222 4752
rect 14734 4740 14740 4752
rect 12216 4712 14740 4740
rect 12216 4700 12222 4712
rect 14734 4700 14740 4712
rect 14792 4740 14798 4752
rect 14792 4712 14872 4740
rect 14792 4700 14798 4712
rect 11425 4675 11483 4681
rect 11425 4641 11437 4675
rect 11471 4641 11483 4675
rect 11606 4672 11612 4684
rect 11567 4644 11612 4672
rect 11425 4635 11483 4641
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 11698 4632 11704 4684
rect 11756 4672 11762 4684
rect 11974 4672 11980 4684
rect 11756 4644 11980 4672
rect 11756 4632 11762 4644
rect 11974 4632 11980 4644
rect 12032 4632 12038 4684
rect 12437 4675 12495 4681
rect 12437 4641 12449 4675
rect 12483 4641 12495 4675
rect 12437 4635 12495 4641
rect 12342 4604 12348 4616
rect 11164 4576 12348 4604
rect 12342 4564 12348 4576
rect 12400 4564 12406 4616
rect 12452 4604 12480 4635
rect 12526 4632 12532 4684
rect 12584 4672 12590 4684
rect 12621 4675 12679 4681
rect 12621 4672 12633 4675
rect 12584 4644 12633 4672
rect 12584 4632 12590 4644
rect 12621 4641 12633 4644
rect 12667 4641 12679 4675
rect 12802 4672 12808 4684
rect 12621 4635 12679 4641
rect 12728 4644 12808 4672
rect 12728 4604 12756 4644
rect 12802 4632 12808 4644
rect 12860 4632 12866 4684
rect 12894 4632 12900 4684
rect 12952 4672 12958 4684
rect 13170 4672 13176 4684
rect 12952 4644 13176 4672
rect 12952 4632 12958 4644
rect 13170 4632 13176 4644
rect 13228 4632 13234 4684
rect 13630 4672 13636 4684
rect 13591 4644 13636 4672
rect 13630 4632 13636 4644
rect 13688 4632 13694 4684
rect 13817 4675 13875 4681
rect 13817 4641 13829 4675
rect 13863 4672 13875 4675
rect 14182 4672 14188 4684
rect 13863 4644 14188 4672
rect 13863 4641 13875 4644
rect 13817 4635 13875 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 13538 4604 13544 4616
rect 12452 4576 12756 4604
rect 13499 4576 13544 4604
rect 13538 4564 13544 4576
rect 13596 4564 13602 4616
rect 14090 4564 14096 4616
rect 14148 4604 14154 4616
rect 14844 4613 14872 4712
rect 15028 4613 15056 4780
rect 17037 4777 17049 4811
rect 17083 4808 17095 4811
rect 17218 4808 17224 4820
rect 17083 4780 17224 4808
rect 17083 4777 17095 4780
rect 17037 4771 17095 4777
rect 17218 4768 17224 4780
rect 17276 4808 17282 4820
rect 18322 4808 18328 4820
rect 17276 4780 18328 4808
rect 17276 4768 17282 4780
rect 18322 4768 18328 4780
rect 18380 4768 18386 4820
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18472 4780 19012 4808
rect 18472 4768 18478 4780
rect 15197 4743 15255 4749
rect 15197 4709 15209 4743
rect 15243 4740 15255 4743
rect 15654 4740 15660 4752
rect 15243 4712 15660 4740
rect 15243 4709 15255 4712
rect 15197 4703 15255 4709
rect 15654 4700 15660 4712
rect 15712 4700 15718 4752
rect 17129 4743 17187 4749
rect 17129 4709 17141 4743
rect 17175 4740 17187 4743
rect 17402 4740 17408 4752
rect 17175 4712 17408 4740
rect 17175 4709 17187 4712
rect 17129 4703 17187 4709
rect 17402 4700 17408 4712
rect 17460 4700 17466 4752
rect 18984 4740 19012 4780
rect 19058 4768 19064 4820
rect 19116 4808 19122 4820
rect 19245 4811 19303 4817
rect 19245 4808 19257 4811
rect 19116 4780 19257 4808
rect 19116 4768 19122 4780
rect 19245 4777 19257 4780
rect 19291 4777 19303 4811
rect 19245 4771 19303 4777
rect 20254 4768 20260 4820
rect 20312 4808 20318 4820
rect 20441 4811 20499 4817
rect 20441 4808 20453 4811
rect 20312 4780 20453 4808
rect 20312 4768 20318 4780
rect 20441 4777 20453 4780
rect 20487 4777 20499 4811
rect 20441 4771 20499 4777
rect 21361 4811 21419 4817
rect 21361 4777 21373 4811
rect 21407 4808 21419 4811
rect 22738 4808 22744 4820
rect 21407 4780 22744 4808
rect 21407 4777 21419 4780
rect 21361 4771 21419 4777
rect 22738 4768 22744 4780
rect 22796 4768 22802 4820
rect 18984 4712 20208 4740
rect 15102 4632 15108 4684
rect 15160 4672 15166 4684
rect 19886 4672 19892 4684
rect 15160 4644 15700 4672
rect 15160 4632 15166 4644
rect 14369 4607 14427 4613
rect 14369 4604 14381 4607
rect 14148 4576 14381 4604
rect 14148 4564 14154 4576
rect 14369 4573 14381 4576
rect 14415 4573 14427 4607
rect 14369 4567 14427 4573
rect 14829 4607 14887 4613
rect 14829 4573 14841 4607
rect 14875 4573 14887 4607
rect 14829 4567 14887 4573
rect 15013 4607 15071 4613
rect 15013 4573 15025 4607
rect 15059 4573 15071 4607
rect 15013 4567 15071 4573
rect 15289 4607 15347 4613
rect 15289 4573 15301 4607
rect 15335 4604 15347 4607
rect 15378 4604 15384 4616
rect 15335 4576 15384 4604
rect 15335 4573 15347 4576
rect 15289 4567 15347 4573
rect 15378 4564 15384 4576
rect 15436 4564 15442 4616
rect 15672 4613 15700 4644
rect 16684 4644 17816 4672
rect 19847 4644 19892 4672
rect 15657 4607 15715 4613
rect 15657 4573 15669 4607
rect 15703 4573 15715 4607
rect 15657 4567 15715 4573
rect 15924 4607 15982 4613
rect 15924 4573 15936 4607
rect 15970 4604 15982 4607
rect 16482 4604 16488 4616
rect 15970 4576 16488 4604
rect 15970 4573 15982 4576
rect 15924 4567 15982 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 6472 4508 8340 4536
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 8570 4536 8576 4548
rect 8435 4508 8576 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 8570 4496 8576 4508
rect 8628 4496 8634 4548
rect 8754 4496 8760 4548
rect 8812 4536 8818 4548
rect 9125 4539 9183 4545
rect 9125 4536 9137 4539
rect 8812 4508 9137 4536
rect 8812 4496 8818 4508
rect 9125 4505 9137 4508
rect 9171 4536 9183 4539
rect 9490 4536 9496 4548
rect 9171 4508 9496 4536
rect 9171 4505 9183 4508
rect 9125 4499 9183 4505
rect 9490 4496 9496 4508
rect 9548 4496 9554 4548
rect 9677 4539 9735 4545
rect 9677 4505 9689 4539
rect 9723 4536 9735 4539
rect 9858 4536 9864 4548
rect 9723 4508 9864 4536
rect 9723 4505 9735 4508
rect 9677 4499 9735 4505
rect 9858 4496 9864 4508
rect 9916 4496 9922 4548
rect 10226 4496 10232 4548
rect 10284 4536 10290 4548
rect 10284 4508 11008 4536
rect 10284 4496 10290 4508
rect 10980 4480 11008 4508
rect 11606 4496 11612 4548
rect 11664 4536 11670 4548
rect 11974 4536 11980 4548
rect 11664 4508 11980 4536
rect 11664 4496 11670 4508
rect 11974 4496 11980 4508
rect 12032 4496 12038 4548
rect 16684 4536 16712 4644
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4573 17739 4607
rect 17788 4604 17816 4644
rect 19886 4632 19892 4644
rect 19944 4632 19950 4684
rect 20073 4607 20131 4613
rect 20073 4604 20085 4607
rect 17788 4576 20085 4604
rect 17681 4567 17739 4573
rect 20073 4573 20085 4576
rect 20119 4573 20131 4607
rect 20180 4604 20208 4712
rect 20898 4672 20904 4684
rect 20859 4644 20904 4672
rect 20898 4632 20904 4644
rect 20956 4632 20962 4684
rect 21085 4675 21143 4681
rect 21085 4641 21097 4675
rect 21131 4672 21143 4675
rect 21542 4672 21548 4684
rect 21131 4644 21548 4672
rect 21131 4641 21143 4644
rect 21085 4635 21143 4641
rect 21542 4632 21548 4644
rect 21600 4632 21606 4684
rect 20257 4607 20315 4613
rect 20257 4604 20269 4607
rect 20180 4576 20269 4604
rect 20073 4567 20131 4573
rect 20257 4573 20269 4576
rect 20303 4573 20315 4607
rect 20257 4567 20315 4573
rect 21453 4607 21511 4613
rect 21453 4573 21465 4607
rect 21499 4604 21511 4607
rect 22002 4604 22008 4616
rect 21499 4576 22008 4604
rect 21499 4573 21511 4576
rect 21453 4567 21511 4573
rect 17494 4536 17500 4548
rect 12176 4508 16712 4536
rect 17455 4508 17500 4536
rect 12176 4480 12204 4508
rect 17494 4496 17500 4508
rect 17552 4496 17558 4548
rect 17696 4536 17724 4567
rect 22002 4564 22008 4576
rect 22060 4564 22066 4616
rect 17954 4545 17960 4548
rect 17948 4536 17960 4545
rect 17696 4508 17816 4536
rect 17915 4508 17960 4536
rect 3329 4471 3387 4477
rect 3329 4437 3341 4471
rect 3375 4437 3387 4471
rect 3786 4468 3792 4480
rect 3747 4440 3792 4468
rect 3329 4431 3387 4437
rect 3786 4428 3792 4440
rect 3844 4428 3850 4480
rect 5629 4471 5687 4477
rect 5629 4437 5641 4471
rect 5675 4468 5687 4471
rect 5810 4468 5816 4480
rect 5675 4440 5816 4468
rect 5675 4437 5687 4440
rect 5629 4431 5687 4437
rect 5810 4428 5816 4440
rect 5868 4428 5874 4480
rect 7282 4428 7288 4480
rect 7340 4468 7346 4480
rect 7561 4471 7619 4477
rect 7561 4468 7573 4471
rect 7340 4440 7573 4468
rect 7340 4428 7346 4440
rect 7561 4437 7573 4440
rect 7607 4468 7619 4471
rect 7650 4468 7656 4480
rect 7607 4440 7656 4468
rect 7607 4437 7619 4440
rect 7561 4431 7619 4437
rect 7650 4428 7656 4440
rect 7708 4428 7714 4480
rect 8021 4471 8079 4477
rect 8021 4437 8033 4471
rect 8067 4468 8079 4471
rect 8294 4468 8300 4480
rect 8067 4440 8300 4468
rect 8067 4437 8079 4440
rect 8021 4431 8079 4437
rect 8294 4428 8300 4440
rect 8352 4428 8358 4480
rect 8478 4428 8484 4480
rect 8536 4468 8542 4480
rect 8536 4440 8581 4468
rect 8536 4428 8542 4440
rect 9306 4428 9312 4480
rect 9364 4468 9370 4480
rect 9585 4471 9643 4477
rect 9585 4468 9597 4471
rect 9364 4440 9597 4468
rect 9364 4428 9370 4440
rect 9585 4437 9597 4440
rect 9631 4468 9643 4471
rect 9766 4468 9772 4480
rect 9631 4440 9772 4468
rect 9631 4437 9643 4440
rect 9585 4431 9643 4437
rect 9766 4428 9772 4440
rect 9824 4428 9830 4480
rect 10594 4428 10600 4480
rect 10652 4468 10658 4480
rect 10873 4471 10931 4477
rect 10873 4468 10885 4471
rect 10652 4440 10885 4468
rect 10652 4428 10658 4440
rect 10873 4437 10885 4440
rect 10919 4437 10931 4471
rect 10873 4431 10931 4437
rect 10962 4428 10968 4480
rect 11020 4428 11026 4480
rect 11238 4428 11244 4480
rect 11296 4468 11302 4480
rect 11701 4471 11759 4477
rect 11701 4468 11713 4471
rect 11296 4440 11713 4468
rect 11296 4428 11302 4440
rect 11701 4437 11713 4440
rect 11747 4437 11759 4471
rect 12066 4468 12072 4480
rect 12027 4440 12072 4468
rect 11701 4431 11759 4437
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 12158 4428 12164 4480
rect 12216 4428 12222 4480
rect 12526 4428 12532 4480
rect 12584 4468 12590 4480
rect 12713 4471 12771 4477
rect 12713 4468 12725 4471
rect 12584 4440 12725 4468
rect 12584 4428 12590 4440
rect 12713 4437 12725 4440
rect 12759 4437 12771 4471
rect 12713 4431 12771 4437
rect 13170 4428 13176 4480
rect 13228 4468 13234 4480
rect 14274 4468 14280 4480
rect 13228 4440 13273 4468
rect 14235 4440 14280 4468
rect 13228 4428 13234 4440
rect 14274 4428 14280 4440
rect 14332 4428 14338 4480
rect 14550 4468 14556 4480
rect 14511 4440 14556 4468
rect 14550 4428 14556 4440
rect 14608 4428 14614 4480
rect 14645 4471 14703 4477
rect 14645 4437 14657 4471
rect 14691 4468 14703 4471
rect 14734 4468 14740 4480
rect 14691 4440 14740 4468
rect 14691 4437 14703 4440
rect 14645 4431 14703 4437
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 16942 4468 16948 4480
rect 15519 4440 16948 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 17402 4468 17408 4480
rect 17363 4440 17408 4468
rect 17402 4428 17408 4440
rect 17460 4428 17466 4480
rect 17788 4468 17816 4508
rect 17948 4499 17960 4508
rect 17954 4496 17960 4499
rect 18012 4496 18018 4548
rect 18874 4496 18880 4548
rect 18932 4536 18938 4548
rect 19705 4539 19763 4545
rect 19705 4536 19717 4539
rect 18932 4508 19717 4536
rect 18932 4496 18938 4508
rect 19705 4505 19717 4508
rect 19751 4505 19763 4539
rect 19705 4499 19763 4505
rect 20809 4539 20867 4545
rect 20809 4505 20821 4539
rect 20855 4536 20867 4539
rect 20990 4536 20996 4548
rect 20855 4508 20996 4536
rect 20855 4505 20867 4508
rect 20809 4499 20867 4505
rect 20990 4496 20996 4508
rect 21048 4496 21054 4548
rect 21174 4496 21180 4548
rect 21232 4536 21238 4548
rect 21542 4536 21548 4548
rect 21232 4508 21548 4536
rect 21232 4496 21238 4508
rect 21542 4496 21548 4508
rect 21600 4496 21606 4548
rect 18230 4468 18236 4480
rect 17788 4440 18236 4468
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18966 4428 18972 4480
rect 19024 4468 19030 4480
rect 19061 4471 19119 4477
rect 19061 4468 19073 4471
rect 19024 4440 19073 4468
rect 19024 4428 19030 4440
rect 19061 4437 19073 4440
rect 19107 4437 19119 4471
rect 19610 4468 19616 4480
rect 19571 4440 19616 4468
rect 19061 4431 19119 4437
rect 19610 4428 19616 4440
rect 19668 4428 19674 4480
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 3053 4267 3111 4273
rect 3053 4233 3065 4267
rect 3099 4264 3111 4267
rect 3513 4267 3571 4273
rect 3513 4264 3525 4267
rect 3099 4236 3525 4264
rect 3099 4233 3111 4236
rect 3053 4227 3111 4233
rect 3513 4233 3525 4236
rect 3559 4233 3571 4267
rect 3513 4227 3571 4233
rect 4157 4267 4215 4273
rect 4157 4233 4169 4267
rect 4203 4264 4215 4267
rect 5718 4264 5724 4276
rect 4203 4236 5580 4264
rect 5679 4236 5724 4264
rect 4203 4233 4215 4236
rect 4157 4227 4215 4233
rect 2685 4199 2743 4205
rect 2685 4165 2697 4199
rect 2731 4196 2743 4199
rect 3786 4196 3792 4208
rect 2731 4168 3792 4196
rect 2731 4165 2743 4168
rect 2685 4159 2743 4165
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 3878 4156 3884 4208
rect 3936 4196 3942 4208
rect 4246 4196 4252 4208
rect 3936 4168 4252 4196
rect 3936 4156 3942 4168
rect 4246 4156 4252 4168
rect 4304 4196 4310 4208
rect 4341 4199 4399 4205
rect 4341 4196 4353 4199
rect 4304 4168 4353 4196
rect 4304 4156 4310 4168
rect 4341 4165 4353 4168
rect 4387 4165 4399 4199
rect 5552 4196 5580 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 5994 4224 6000 4276
rect 6052 4264 6058 4276
rect 6638 4264 6644 4276
rect 6052 4236 6644 4264
rect 6052 4224 6058 4236
rect 6638 4224 6644 4236
rect 6696 4224 6702 4276
rect 8478 4224 8484 4276
rect 8536 4264 8542 4276
rect 9217 4267 9275 4273
rect 9217 4264 9229 4267
rect 8536 4236 9229 4264
rect 8536 4224 8542 4236
rect 9217 4233 9229 4236
rect 9263 4233 9275 4267
rect 9217 4227 9275 4233
rect 9490 4224 9496 4276
rect 9548 4264 9554 4276
rect 9585 4267 9643 4273
rect 9585 4264 9597 4267
rect 9548 4236 9597 4264
rect 9548 4224 9554 4236
rect 9585 4233 9597 4236
rect 9631 4233 9643 4267
rect 9585 4227 9643 4233
rect 9950 4224 9956 4276
rect 10008 4264 10014 4276
rect 10008 4236 10732 4264
rect 10008 4224 10014 4236
rect 6730 4196 6736 4208
rect 5552 4168 6736 4196
rect 4341 4159 4399 4165
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 7190 4196 7196 4208
rect 7024 4168 7196 4196
rect 198 4088 204 4140
rect 256 4128 262 4140
rect 934 4128 940 4140
rect 256 4100 940 4128
rect 256 4088 262 4100
rect 934 4088 940 4100
rect 992 4088 998 4140
rect 1946 4128 1952 4140
rect 1907 4100 1952 4128
rect 1946 4088 1952 4100
rect 2004 4088 2010 4140
rect 2222 4128 2228 4140
rect 2183 4100 2228 4128
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2590 4128 2596 4140
rect 2551 4100 2596 4128
rect 2590 4088 2596 4100
rect 2648 4088 2654 4140
rect 3418 4128 3424 4140
rect 3379 4100 3424 4128
rect 3418 4088 3424 4100
rect 3476 4088 3482 4140
rect 4525 4131 4583 4137
rect 4525 4097 4537 4131
rect 4571 4128 4583 4131
rect 4798 4128 4804 4140
rect 4571 4100 4804 4128
rect 4571 4097 4583 4100
rect 4525 4091 4583 4097
rect 4798 4088 4804 4100
rect 4856 4088 4862 4140
rect 4985 4131 5043 4137
rect 4985 4128 4997 4131
rect 4908 4100 4997 4128
rect 2498 4060 2504 4072
rect 2459 4032 2504 4060
rect 2498 4020 2504 4032
rect 2556 4020 2562 4072
rect 3237 4063 3295 4069
rect 3237 4060 3249 4063
rect 2746 4032 3249 4060
rect 1762 3952 1768 4004
rect 1820 3992 1826 4004
rect 2314 3992 2320 4004
rect 1820 3964 2320 3992
rect 1820 3952 1826 3964
rect 2314 3952 2320 3964
rect 2372 3992 2378 4004
rect 2746 3992 2774 4032
rect 3237 4029 3249 4032
rect 3283 4029 3295 4063
rect 4614 4060 4620 4072
rect 3237 4023 3295 4029
rect 3712 4032 4620 4060
rect 2372 3964 2774 3992
rect 2372 3952 2378 3964
rect 3050 3952 3056 4004
rect 3108 3992 3114 4004
rect 3712 3992 3740 4032
rect 4614 4020 4620 4032
rect 4672 4060 4678 4072
rect 4908 4060 4936 4100
rect 4985 4097 4997 4100
rect 5031 4097 5043 4131
rect 4985 4091 5043 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 6457 4131 6515 4137
rect 6457 4128 6469 4131
rect 5813 4091 5871 4097
rect 6012 4100 6469 4128
rect 5074 4060 5080 4072
rect 4672 4032 4936 4060
rect 5035 4032 5080 4060
rect 4672 4020 4678 4032
rect 5074 4020 5080 4032
rect 5132 4020 5138 4072
rect 5258 4060 5264 4072
rect 5219 4032 5264 4060
rect 5258 4020 5264 4032
rect 5316 4020 5322 4072
rect 5537 4063 5595 4069
rect 5537 4029 5549 4063
rect 5583 4029 5595 4063
rect 5537 4023 5595 4029
rect 3878 3992 3884 4004
rect 3108 3964 3740 3992
rect 3839 3964 3884 3992
rect 3108 3952 3114 3964
rect 3878 3952 3884 3964
rect 3936 3952 3942 4004
rect 4448 3964 4752 3992
rect 1210 3884 1216 3936
rect 1268 3924 1274 3936
rect 4448 3924 4476 3964
rect 4614 3924 4620 3936
rect 1268 3896 4476 3924
rect 4575 3896 4620 3924
rect 1268 3884 1274 3896
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 4724 3924 4752 3964
rect 4798 3952 4804 4004
rect 4856 3992 4862 4004
rect 5276 3992 5304 4020
rect 4856 3964 5304 3992
rect 4856 3952 4862 3964
rect 5350 3924 5356 3936
rect 4724 3896 5356 3924
rect 5350 3884 5356 3896
rect 5408 3884 5414 3936
rect 5552 3924 5580 4023
rect 5718 4020 5724 4072
rect 5776 4060 5782 4072
rect 5828 4060 5856 4091
rect 5776 4032 5856 4060
rect 5776 4020 5782 4032
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 6012 3992 6040 4100
rect 6457 4097 6469 4100
rect 6503 4097 6515 4131
rect 6457 4091 6515 4097
rect 6641 4131 6699 4137
rect 6641 4097 6653 4131
rect 6687 4128 6699 4131
rect 7024 4128 7052 4168
rect 7190 4156 7196 4168
rect 7248 4196 7254 4208
rect 7374 4196 7380 4208
rect 7248 4168 7380 4196
rect 7248 4156 7254 4168
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 10594 4156 10600 4208
rect 10652 4156 10658 4208
rect 7098 4137 7104 4140
rect 6687 4100 7052 4128
rect 6687 4097 6699 4100
rect 6641 4091 6699 4097
rect 7092 4091 7104 4137
rect 7156 4128 7162 4140
rect 7156 4100 7192 4128
rect 7098 4088 7104 4091
rect 7156 4088 7162 4100
rect 8478 4088 8484 4140
rect 8536 4128 8542 4140
rect 8665 4131 8723 4137
rect 8665 4128 8677 4131
rect 8536 4100 8677 4128
rect 8536 4088 8542 4100
rect 8665 4097 8677 4100
rect 8711 4097 8723 4131
rect 8665 4091 8723 4097
rect 8846 4088 8852 4140
rect 8904 4128 8910 4140
rect 10226 4128 10232 4140
rect 8904 4100 10232 4128
rect 8904 4088 8910 4100
rect 10226 4088 10232 4100
rect 10284 4088 10290 4140
rect 10410 4128 10416 4140
rect 10371 4100 10416 4128
rect 10410 4088 10416 4100
rect 10468 4088 10474 4140
rect 6822 4060 6828 4072
rect 6783 4032 6828 4060
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 8386 4060 8392 4072
rect 8220 4032 8392 4060
rect 5684 3964 6040 3992
rect 6181 3995 6239 4001
rect 5684 3952 5690 3964
rect 6181 3961 6193 3995
rect 6227 3992 6239 3995
rect 6730 3992 6736 4004
rect 6227 3964 6736 3992
rect 6227 3961 6239 3964
rect 6181 3955 6239 3961
rect 6730 3952 6736 3964
rect 6788 3952 6794 4004
rect 8220 4001 8248 4032
rect 8386 4020 8392 4032
rect 8444 4020 8450 4072
rect 8570 4060 8576 4072
rect 8531 4032 8576 4060
rect 8570 4020 8576 4032
rect 8628 4020 8634 4072
rect 9677 4063 9735 4069
rect 9677 4029 9689 4063
rect 9723 4029 9735 4063
rect 9677 4023 9735 4029
rect 8205 3995 8263 4001
rect 8205 3961 8217 3995
rect 8251 3961 8263 3995
rect 9692 3992 9720 4023
rect 9766 4020 9772 4072
rect 9824 4060 9830 4072
rect 10505 4063 10563 4069
rect 9824 4032 9869 4060
rect 9824 4020 9830 4032
rect 10505 4029 10517 4063
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 10045 3995 10103 4001
rect 10045 3992 10057 3995
rect 9692 3964 10057 3992
rect 8205 3955 8263 3961
rect 10045 3961 10057 3964
rect 10091 3961 10103 3995
rect 10045 3955 10103 3961
rect 10410 3952 10416 4004
rect 10468 3992 10474 4004
rect 10520 3992 10548 4023
rect 10468 3964 10548 3992
rect 10612 3992 10640 4156
rect 10704 4069 10732 4236
rect 10870 4224 10876 4276
rect 10928 4264 10934 4276
rect 11885 4267 11943 4273
rect 10928 4236 11192 4264
rect 10928 4224 10934 4236
rect 10873 4131 10931 4137
rect 10873 4097 10885 4131
rect 10919 4097 10931 4131
rect 10873 4091 10931 4097
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4029 10747 4063
rect 10689 4023 10747 4029
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10897 4060 10925 4091
rect 11054 4088 11060 4140
rect 11112 4088 11118 4140
rect 11164 4137 11192 4236
rect 11885 4233 11897 4267
rect 11931 4233 11943 4267
rect 11885 4227 11943 4233
rect 11900 4196 11928 4227
rect 12066 4224 12072 4276
rect 12124 4264 12130 4276
rect 12434 4264 12440 4276
rect 12124 4236 12440 4264
rect 12124 4224 12130 4236
rect 12434 4224 12440 4236
rect 12492 4224 12498 4276
rect 12805 4267 12863 4273
rect 12805 4233 12817 4267
rect 12851 4264 12863 4267
rect 13170 4264 13176 4276
rect 12851 4236 13176 4264
rect 12851 4233 12863 4236
rect 12805 4227 12863 4233
rect 13170 4224 13176 4236
rect 13228 4224 13234 4276
rect 13265 4267 13323 4273
rect 13265 4233 13277 4267
rect 13311 4264 13323 4267
rect 13538 4264 13544 4276
rect 13311 4236 13544 4264
rect 13311 4233 13323 4236
rect 13265 4227 13323 4233
rect 13538 4224 13544 4236
rect 13596 4224 13602 4276
rect 13725 4267 13783 4273
rect 13725 4233 13737 4267
rect 13771 4264 13783 4267
rect 14185 4267 14243 4273
rect 14185 4264 14197 4267
rect 13771 4236 14197 4264
rect 13771 4233 13783 4236
rect 13725 4227 13783 4233
rect 14185 4233 14197 4236
rect 14231 4233 14243 4267
rect 14185 4227 14243 4233
rect 14274 4224 14280 4276
rect 14332 4264 14338 4276
rect 14553 4267 14611 4273
rect 14553 4264 14565 4267
rect 14332 4236 14565 4264
rect 14332 4224 14338 4236
rect 14553 4233 14565 4236
rect 14599 4233 14611 4267
rect 15470 4264 15476 4276
rect 15431 4236 15476 4264
rect 14553 4227 14611 4233
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 18874 4264 18880 4276
rect 18835 4236 18880 4264
rect 18874 4224 18880 4236
rect 18932 4224 18938 4276
rect 19610 4224 19616 4276
rect 19668 4264 19674 4276
rect 19705 4267 19763 4273
rect 19705 4264 19717 4267
rect 19668 4236 19717 4264
rect 19668 4224 19674 4236
rect 19705 4233 19717 4236
rect 19751 4233 19763 4267
rect 19705 4227 19763 4233
rect 19797 4267 19855 4273
rect 19797 4233 19809 4267
rect 19843 4233 19855 4267
rect 19797 4227 19855 4233
rect 20165 4267 20223 4273
rect 20165 4233 20177 4267
rect 20211 4264 20223 4267
rect 20714 4264 20720 4276
rect 20211 4236 20720 4264
rect 20211 4233 20223 4236
rect 20165 4227 20223 4233
rect 12894 4196 12900 4208
rect 11256 4168 11928 4196
rect 12855 4168 12900 4196
rect 11149 4131 11207 4137
rect 11149 4097 11161 4131
rect 11195 4097 11207 4131
rect 11149 4091 11207 4097
rect 10836 4032 10925 4060
rect 11072 4060 11100 4088
rect 11256 4060 11284 4168
rect 12894 4156 12900 4168
rect 12952 4156 12958 4208
rect 13633 4199 13691 4205
rect 13633 4165 13645 4199
rect 13679 4196 13691 4199
rect 13998 4196 14004 4208
rect 13679 4168 14004 4196
rect 13679 4165 13691 4168
rect 13633 4159 13691 4165
rect 13998 4156 14004 4168
rect 14056 4156 14062 4208
rect 15562 4156 15568 4208
rect 15620 4196 15626 4208
rect 17494 4196 17500 4208
rect 15620 4168 16252 4196
rect 15620 4156 15626 4168
rect 11422 4088 11428 4140
rect 11480 4128 11486 4140
rect 12158 4128 12164 4140
rect 11480 4100 12164 4128
rect 11480 4088 11486 4100
rect 12158 4088 12164 4100
rect 12216 4088 12222 4140
rect 12434 4088 12440 4140
rect 12492 4128 12498 4140
rect 12802 4128 12808 4140
rect 12492 4100 12808 4128
rect 12492 4088 12498 4100
rect 12802 4088 12808 4100
rect 12860 4128 12866 4140
rect 12860 4100 13584 4128
rect 12860 4088 12866 4100
rect 11072 4032 11284 4060
rect 10836 4020 10842 4032
rect 11514 4020 11520 4072
rect 11572 4060 11578 4072
rect 11977 4063 12035 4069
rect 11977 4060 11989 4063
rect 11572 4032 11989 4060
rect 11572 4020 11578 4032
rect 11977 4029 11989 4032
rect 12023 4029 12035 4063
rect 11977 4023 12035 4029
rect 12069 4063 12127 4069
rect 12069 4029 12081 4063
rect 12115 4060 12127 4063
rect 12250 4060 12256 4072
rect 12115 4032 12256 4060
rect 12115 4029 12127 4032
rect 12069 4023 12127 4029
rect 12250 4020 12256 4032
rect 12308 4060 12314 4072
rect 12526 4060 12532 4072
rect 12308 4032 12532 4060
rect 12308 4020 12314 4032
rect 12526 4020 12532 4032
rect 12584 4020 12590 4072
rect 12713 4063 12771 4069
rect 12713 4029 12725 4063
rect 12759 4060 12771 4063
rect 13354 4060 13360 4072
rect 12759 4032 13360 4060
rect 12759 4029 12771 4032
rect 12713 4023 12771 4029
rect 13354 4020 13360 4032
rect 13412 4060 13418 4072
rect 13449 4063 13507 4069
rect 13449 4060 13461 4063
rect 13412 4032 13461 4060
rect 13412 4020 13418 4032
rect 13449 4029 13461 4032
rect 13495 4029 13507 4063
rect 13556 4060 13584 4100
rect 13906 4088 13912 4140
rect 13964 4128 13970 4140
rect 15381 4131 15439 4137
rect 15381 4128 15393 4131
rect 13964 4100 15393 4128
rect 13964 4088 13970 4100
rect 15381 4097 15393 4100
rect 15427 4097 15439 4131
rect 15381 4091 15439 4097
rect 15470 4088 15476 4140
rect 15528 4128 15534 4140
rect 16224 4137 16252 4168
rect 16592 4168 17500 4196
rect 15933 4131 15991 4137
rect 15933 4128 15945 4131
rect 15528 4100 15945 4128
rect 15528 4088 15534 4100
rect 15933 4097 15945 4100
rect 15979 4097 15991 4131
rect 15933 4091 15991 4097
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 13556 4032 14228 4060
rect 13449 4023 13507 4029
rect 14200 4004 14228 4032
rect 14366 4020 14372 4072
rect 14424 4060 14430 4072
rect 14642 4060 14648 4072
rect 14424 4032 14648 4060
rect 14424 4020 14430 4032
rect 14642 4020 14648 4032
rect 14700 4020 14706 4072
rect 14737 4063 14795 4069
rect 14737 4029 14749 4063
rect 14783 4029 14795 4063
rect 15286 4060 15292 4072
rect 15247 4032 15292 4060
rect 14737 4023 14795 4029
rect 11057 3995 11115 4001
rect 10612 3964 11008 3992
rect 10468 3952 10474 3964
rect 6454 3924 6460 3936
rect 5552 3896 6460 3924
rect 6454 3884 6460 3896
rect 6512 3884 6518 3936
rect 9033 3927 9091 3933
rect 9033 3893 9045 3927
rect 9079 3924 9091 3927
rect 10778 3924 10784 3936
rect 9079 3896 10784 3924
rect 9079 3893 9091 3896
rect 9033 3887 9091 3893
rect 10778 3884 10784 3896
rect 10836 3884 10842 3936
rect 10980 3924 11008 3964
rect 11057 3961 11069 3995
rect 11103 3992 11115 3995
rect 13722 3992 13728 4004
rect 11103 3964 13728 3992
rect 11103 3961 11115 3964
rect 11057 3955 11115 3961
rect 13722 3952 13728 3964
rect 13780 3952 13786 4004
rect 14182 3952 14188 4004
rect 14240 3992 14246 4004
rect 14752 3992 14780 4023
rect 15286 4020 15292 4032
rect 15344 4060 15350 4072
rect 16592 4060 16620 4168
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 18046 4156 18052 4208
rect 18104 4196 18110 4208
rect 19337 4199 19395 4205
rect 18104 4168 18635 4196
rect 18104 4156 18110 4168
rect 16936 4131 16994 4137
rect 16936 4097 16948 4131
rect 16982 4128 16994 4131
rect 17218 4128 17224 4140
rect 16982 4100 17224 4128
rect 16982 4097 16994 4100
rect 16936 4091 16994 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17512 4128 17540 4156
rect 18506 4128 18512 4140
rect 17512 4100 17724 4128
rect 18467 4100 18512 4128
rect 15344 4032 16620 4060
rect 16669 4063 16727 4069
rect 15344 4020 15350 4032
rect 16669 4029 16681 4063
rect 16715 4029 16727 4063
rect 16669 4023 16727 4029
rect 14240 3964 14780 3992
rect 14240 3952 14246 3964
rect 15102 3952 15108 4004
rect 15160 3992 15166 4004
rect 16114 3992 16120 4004
rect 15160 3964 15976 3992
rect 16075 3964 16120 3992
rect 15160 3952 15166 3964
rect 11146 3924 11152 3936
rect 10980 3896 11152 3924
rect 11146 3884 11152 3896
rect 11204 3884 11210 3936
rect 11238 3884 11244 3936
rect 11296 3924 11302 3936
rect 11333 3927 11391 3933
rect 11333 3924 11345 3927
rect 11296 3896 11345 3924
rect 11296 3884 11302 3896
rect 11333 3893 11345 3896
rect 11379 3893 11391 3927
rect 11333 3887 11391 3893
rect 11517 3927 11575 3933
rect 11517 3893 11529 3927
rect 11563 3924 11575 3927
rect 11698 3924 11704 3936
rect 11563 3896 11704 3924
rect 11563 3893 11575 3896
rect 11517 3887 11575 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 12437 3927 12495 3933
rect 12437 3893 12449 3927
rect 12483 3924 12495 3927
rect 13814 3924 13820 3936
rect 12483 3896 13820 3924
rect 12483 3893 12495 3896
rect 12437 3887 12495 3893
rect 13814 3884 13820 3896
rect 13872 3884 13878 3936
rect 14093 3927 14151 3933
rect 14093 3893 14105 3927
rect 14139 3924 14151 3927
rect 14458 3924 14464 3936
rect 14139 3896 14464 3924
rect 14139 3893 14151 3896
rect 14093 3887 14151 3893
rect 14458 3884 14464 3896
rect 14516 3884 14522 3936
rect 15838 3924 15844 3936
rect 15799 3896 15844 3924
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 15948 3924 15976 3964
rect 16114 3952 16120 3964
rect 16172 3952 16178 4004
rect 16574 3992 16580 4004
rect 16316 3964 16580 3992
rect 16316 3924 16344 3964
rect 16574 3952 16580 3964
rect 16632 3992 16638 4004
rect 16684 3992 16712 4023
rect 16632 3964 16712 3992
rect 17696 3992 17724 4100
rect 18506 4088 18512 4100
rect 18564 4088 18570 4140
rect 18607 4128 18635 4168
rect 19337 4165 19349 4199
rect 19383 4196 19395 4199
rect 19812 4196 19840 4227
rect 20714 4224 20720 4236
rect 20772 4224 20778 4276
rect 19383 4168 19840 4196
rect 19383 4165 19395 4168
rect 19337 4159 19395 4165
rect 20162 4128 20168 4140
rect 18607 4100 20168 4128
rect 20162 4088 20168 4100
rect 20220 4088 20226 4140
rect 20717 4131 20775 4137
rect 20717 4097 20729 4131
rect 20763 4128 20775 4131
rect 21634 4128 21640 4140
rect 20763 4100 21640 4128
rect 20763 4097 20775 4100
rect 20717 4091 20775 4097
rect 21634 4088 21640 4100
rect 21692 4088 21698 4140
rect 18325 4063 18383 4069
rect 18325 4029 18337 4063
rect 18371 4029 18383 4063
rect 18325 4023 18383 4029
rect 18417 4063 18475 4069
rect 18417 4029 18429 4063
rect 18463 4060 18475 4063
rect 18782 4060 18788 4072
rect 18463 4032 18788 4060
rect 18463 4029 18475 4032
rect 18417 4023 18475 4029
rect 18049 3995 18107 4001
rect 18049 3992 18061 3995
rect 17696 3964 18061 3992
rect 16632 3952 16638 3964
rect 18049 3961 18061 3964
rect 18095 3961 18107 3995
rect 18340 3992 18368 4023
rect 18782 4020 18788 4032
rect 18840 4020 18846 4072
rect 18966 4020 18972 4072
rect 19024 4060 19030 4072
rect 19061 4063 19119 4069
rect 19061 4060 19073 4063
rect 19024 4032 19073 4060
rect 19024 4020 19030 4032
rect 19061 4029 19073 4032
rect 19107 4029 19119 4063
rect 19061 4023 19119 4029
rect 19245 4063 19303 4069
rect 19245 4029 19257 4063
rect 19291 4029 19303 4063
rect 19245 4023 19303 4029
rect 18984 3992 19012 4020
rect 18340 3964 19012 3992
rect 18049 3955 18107 3961
rect 15948 3896 16344 3924
rect 16393 3927 16451 3933
rect 16393 3893 16405 3927
rect 16439 3924 16451 3927
rect 17034 3924 17040 3936
rect 16439 3896 17040 3924
rect 16439 3893 16451 3896
rect 16393 3887 16451 3893
rect 17034 3884 17040 3896
rect 17092 3884 17098 3936
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 18966 3924 18972 3936
rect 18288 3896 18972 3924
rect 18288 3884 18294 3896
rect 18966 3884 18972 3896
rect 19024 3884 19030 3936
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 19260 3924 19288 4023
rect 19334 4020 19340 4072
rect 19392 4060 19398 4072
rect 19610 4060 19616 4072
rect 19392 4032 19616 4060
rect 19392 4020 19398 4032
rect 19610 4020 19616 4032
rect 19668 4020 19674 4072
rect 20254 4060 20260 4072
rect 20215 4032 20260 4060
rect 20254 4020 20260 4032
rect 20312 4020 20318 4072
rect 20346 4020 20352 4072
rect 20404 4060 20410 4072
rect 20993 4063 21051 4069
rect 20404 4032 20449 4060
rect 20404 4020 20410 4032
rect 20993 4029 21005 4063
rect 21039 4060 21051 4063
rect 21818 4060 21824 4072
rect 21039 4032 21824 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 21818 4020 21824 4032
rect 21876 4020 21882 4072
rect 19116 3896 19288 3924
rect 19116 3884 19122 3896
rect 20714 3884 20720 3936
rect 20772 3924 20778 3936
rect 21726 3924 21732 3936
rect 20772 3896 21732 3924
rect 20772 3884 20778 3896
rect 21726 3884 21732 3896
rect 21784 3884 21790 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 5166 3720 5172 3732
rect 3016 3692 5172 3720
rect 3016 3680 3022 3692
rect 5166 3680 5172 3692
rect 5224 3680 5230 3732
rect 5629 3723 5687 3729
rect 5629 3689 5641 3723
rect 5675 3720 5687 3723
rect 5718 3720 5724 3732
rect 5675 3692 5724 3720
rect 5675 3689 5687 3692
rect 5629 3683 5687 3689
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6822 3720 6828 3732
rect 6472 3692 6828 3720
rect 2774 3612 2780 3664
rect 2832 3652 2838 3664
rect 5994 3652 6000 3664
rect 2832 3624 6000 3652
rect 2832 3612 2838 3624
rect 5994 3612 6000 3624
rect 6052 3612 6058 3664
rect 1949 3587 2007 3593
rect 1949 3553 1961 3587
rect 1995 3584 2007 3587
rect 2682 3584 2688 3596
rect 1995 3556 2688 3584
rect 1995 3553 2007 3556
rect 1949 3547 2007 3553
rect 2682 3544 2688 3556
rect 2740 3544 2746 3596
rect 4154 3584 4160 3596
rect 4115 3556 4160 3584
rect 4154 3544 4160 3556
rect 4212 3544 4218 3596
rect 4249 3587 4307 3593
rect 4249 3553 4261 3587
rect 4295 3584 4307 3587
rect 4614 3584 4620 3596
rect 4295 3556 4620 3584
rect 4295 3553 4307 3556
rect 4249 3547 4307 3553
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5442 3584 5448 3596
rect 5403 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3544 5506 3596
rect 5718 3544 5724 3596
rect 5776 3584 5782 3596
rect 6086 3584 6092 3596
rect 5776 3556 6092 3584
rect 5776 3544 5782 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 6270 3584 6276 3596
rect 6231 3556 6276 3584
rect 6270 3544 6276 3556
rect 6328 3544 6334 3596
rect 6472 3593 6500 3692
rect 6822 3680 6828 3692
rect 6880 3680 6886 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 7156 3692 7849 3720
rect 7156 3680 7162 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 6457 3587 6515 3593
rect 6457 3553 6469 3587
rect 6503 3553 6515 3587
rect 7852 3584 7880 3683
rect 8570 3680 8576 3732
rect 8628 3720 8634 3732
rect 8757 3723 8815 3729
rect 8757 3720 8769 3723
rect 8628 3692 8769 3720
rect 8628 3680 8634 3692
rect 8757 3689 8769 3692
rect 8803 3689 8815 3723
rect 8757 3683 8815 3689
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 10502 3720 10508 3732
rect 9916 3692 10508 3720
rect 9916 3680 9922 3692
rect 10502 3680 10508 3692
rect 10560 3680 10566 3732
rect 10778 3680 10784 3732
rect 10836 3720 10842 3732
rect 11701 3723 11759 3729
rect 11701 3720 11713 3723
rect 10836 3692 11713 3720
rect 10836 3680 10842 3692
rect 11701 3689 11713 3692
rect 11747 3689 11759 3723
rect 11701 3683 11759 3689
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 13354 3720 13360 3732
rect 12308 3692 13216 3720
rect 13315 3692 13360 3720
rect 12308 3680 12314 3692
rect 7926 3612 7932 3664
rect 7984 3652 7990 3664
rect 10134 3652 10140 3664
rect 7984 3624 10140 3652
rect 7984 3612 7990 3624
rect 10134 3612 10140 3624
rect 10192 3612 10198 3664
rect 11425 3655 11483 3661
rect 11425 3621 11437 3655
rect 11471 3652 11483 3655
rect 11790 3652 11796 3664
rect 11471 3624 11796 3652
rect 11471 3621 11483 3624
rect 11425 3615 11483 3621
rect 11790 3612 11796 3624
rect 11848 3612 11854 3664
rect 13188 3652 13216 3692
rect 13354 3680 13360 3692
rect 13412 3680 13418 3732
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 15470 3720 15476 3732
rect 13504 3692 15476 3720
rect 13504 3680 13510 3692
rect 15470 3680 15476 3692
rect 15528 3680 15534 3732
rect 15657 3723 15715 3729
rect 15657 3689 15669 3723
rect 15703 3720 15715 3723
rect 18782 3720 18788 3732
rect 15703 3692 18276 3720
rect 18743 3692 18788 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 14826 3652 14832 3664
rect 13188 3624 14832 3652
rect 14826 3612 14832 3624
rect 14884 3612 14890 3664
rect 17954 3652 17960 3664
rect 17867 3624 17960 3652
rect 17954 3612 17960 3624
rect 18012 3612 18018 3664
rect 8113 3587 8171 3593
rect 8113 3584 8125 3587
rect 7852 3556 8125 3584
rect 6457 3547 6515 3553
rect 8113 3553 8125 3556
rect 8159 3553 8171 3587
rect 8294 3584 8300 3596
rect 8255 3556 8300 3584
rect 8113 3547 8171 3553
rect 8294 3544 8300 3556
rect 8352 3544 8358 3596
rect 9306 3584 9312 3596
rect 8404 3556 9312 3584
rect 934 3476 940 3528
rect 992 3516 998 3528
rect 2225 3519 2283 3525
rect 2225 3516 2237 3519
rect 992 3488 2237 3516
rect 992 3476 998 3488
rect 2225 3485 2237 3488
rect 2271 3485 2283 3519
rect 2866 3516 2872 3528
rect 2827 3488 2872 3516
rect 2225 3479 2283 3485
rect 2866 3476 2872 3488
rect 2924 3476 2930 3528
rect 3145 3519 3203 3525
rect 3145 3485 3157 3519
rect 3191 3485 3203 3519
rect 3145 3479 3203 3485
rect 3605 3519 3663 3525
rect 3605 3485 3617 3519
rect 3651 3516 3663 3519
rect 4522 3516 4528 3528
rect 3651 3488 4528 3516
rect 3651 3485 3663 3488
rect 3605 3479 3663 3485
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 3160 3448 3188 3479
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 4706 3476 4712 3528
rect 4764 3516 4770 3528
rect 5997 3519 6055 3525
rect 5997 3516 6009 3519
rect 4764 3488 6009 3516
rect 4764 3476 4770 3488
rect 5997 3485 6009 3488
rect 6043 3516 6055 3519
rect 8404 3516 8432 3556
rect 9306 3544 9312 3556
rect 9364 3544 9370 3596
rect 9493 3587 9551 3593
rect 9493 3553 9505 3587
rect 9539 3553 9551 3587
rect 9493 3547 9551 3553
rect 11149 3587 11207 3593
rect 11149 3553 11161 3587
rect 11195 3584 11207 3587
rect 11606 3584 11612 3596
rect 11195 3556 11612 3584
rect 11195 3553 11207 3556
rect 11149 3547 11207 3553
rect 6043 3488 8432 3516
rect 6043 3485 6055 3488
rect 5997 3479 6055 3485
rect 8938 3476 8944 3528
rect 8996 3516 9002 3528
rect 9508 3516 9536 3547
rect 11164 3516 11192 3547
rect 11606 3544 11612 3556
rect 11664 3544 11670 3596
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 11977 3587 12035 3593
rect 11977 3584 11989 3587
rect 11940 3556 11989 3584
rect 11940 3544 11946 3556
rect 11977 3553 11989 3556
rect 12023 3584 12035 3587
rect 12023 3556 12112 3584
rect 12023 3553 12035 3556
rect 11977 3547 12035 3553
rect 8996 3488 9536 3516
rect 9600 3488 11192 3516
rect 11241 3519 11299 3525
rect 8996 3476 9002 3488
rect 1084 3420 3188 3448
rect 3421 3451 3479 3457
rect 1084 3408 1090 3420
rect 3421 3417 3433 3451
rect 3467 3448 3479 3451
rect 4246 3448 4252 3460
rect 3467 3420 4252 3448
rect 3467 3417 3479 3420
rect 3421 3411 3479 3417
rect 4246 3408 4252 3420
rect 4304 3408 4310 3460
rect 4341 3451 4399 3457
rect 4341 3417 4353 3451
rect 4387 3448 4399 3451
rect 4387 3420 4844 3448
rect 4387 3417 4399 3420
rect 4341 3411 4399 3417
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 3970 3380 3976 3392
rect 3927 3352 3976 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 3970 3340 3976 3352
rect 4028 3340 4034 3392
rect 4706 3380 4712 3392
rect 4667 3352 4712 3380
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 4816 3389 4844 3420
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 6724 3451 6782 3457
rect 6724 3448 6736 3451
rect 6512 3420 6736 3448
rect 6512 3408 6518 3420
rect 6724 3417 6736 3420
rect 6770 3448 6782 3451
rect 7742 3448 7748 3460
rect 6770 3420 7748 3448
rect 6770 3417 6782 3420
rect 6724 3411 6782 3417
rect 7742 3408 7748 3420
rect 7800 3448 7806 3460
rect 8202 3448 8208 3460
rect 7800 3420 8208 3448
rect 7800 3408 7806 3420
rect 8202 3408 8208 3420
rect 8260 3408 8266 3460
rect 9122 3448 9128 3460
rect 8312 3420 9128 3448
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3349 4859 3383
rect 5166 3380 5172 3392
rect 5127 3352 5172 3380
rect 4801 3343 4859 3349
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5261 3383 5319 3389
rect 5261 3349 5273 3383
rect 5307 3380 5319 3383
rect 5442 3380 5448 3392
rect 5307 3352 5448 3380
rect 5307 3349 5319 3352
rect 5261 3343 5319 3349
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5810 3340 5816 3392
rect 5868 3380 5874 3392
rect 6638 3380 6644 3392
rect 5868 3352 6644 3380
rect 5868 3340 5874 3352
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6822 3340 6828 3392
rect 6880 3380 6886 3392
rect 8312 3380 8340 3420
rect 9122 3408 9128 3420
rect 9180 3448 9186 3460
rect 9600 3448 9628 3488
rect 11241 3485 11253 3519
rect 11287 3485 11299 3519
rect 12084 3516 12112 3556
rect 13538 3544 13544 3596
rect 13596 3584 13602 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 13596 3556 14565 3584
rect 13596 3544 13602 3556
rect 14553 3553 14565 3556
rect 14599 3553 14611 3587
rect 14553 3547 14611 3553
rect 14642 3544 14648 3596
rect 14700 3584 14706 3596
rect 15105 3587 15163 3593
rect 14700 3556 14745 3584
rect 14700 3544 14706 3556
rect 15105 3553 15117 3587
rect 15151 3584 15163 3587
rect 15286 3584 15292 3596
rect 15151 3556 15292 3584
rect 15151 3553 15163 3556
rect 15105 3547 15163 3553
rect 15286 3544 15292 3556
rect 15344 3544 15350 3596
rect 16574 3584 16580 3596
rect 16535 3556 16580 3584
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 17972 3584 18000 3612
rect 18141 3587 18199 3593
rect 18141 3584 18153 3587
rect 17972 3556 18153 3584
rect 18141 3553 18153 3556
rect 18187 3553 18199 3587
rect 18248 3584 18276 3692
rect 18782 3680 18788 3692
rect 18840 3680 18846 3732
rect 19058 3680 19064 3732
rect 19116 3720 19122 3732
rect 19245 3723 19303 3729
rect 19245 3720 19257 3723
rect 19116 3692 19257 3720
rect 19116 3680 19122 3692
rect 19245 3689 19257 3692
rect 19291 3689 19303 3723
rect 19245 3683 19303 3689
rect 19610 3680 19616 3732
rect 19668 3720 19674 3732
rect 22830 3720 22836 3732
rect 19668 3692 22836 3720
rect 19668 3680 19674 3692
rect 22830 3680 22836 3692
rect 22888 3680 22894 3732
rect 19518 3612 19524 3664
rect 19576 3652 19582 3664
rect 20070 3652 20076 3664
rect 19576 3624 20076 3652
rect 19576 3612 19582 3624
rect 20070 3612 20076 3624
rect 20128 3612 20134 3664
rect 20254 3612 20260 3664
rect 20312 3652 20318 3664
rect 20993 3655 21051 3661
rect 20993 3652 21005 3655
rect 20312 3624 21005 3652
rect 20312 3612 20318 3624
rect 20993 3621 21005 3624
rect 21039 3621 21051 3655
rect 20993 3615 21051 3621
rect 18325 3587 18383 3593
rect 18325 3584 18337 3587
rect 18248 3556 18337 3584
rect 18141 3547 18199 3553
rect 18325 3553 18337 3556
rect 18371 3553 18383 3587
rect 19702 3584 19708 3596
rect 18325 3547 18383 3553
rect 18432 3556 19196 3584
rect 19663 3556 19708 3584
rect 12710 3516 12716 3528
rect 12084 3488 12716 3516
rect 11241 3479 11299 3485
rect 9180 3420 9628 3448
rect 9180 3408 9186 3420
rect 9674 3408 9680 3460
rect 9732 3448 9738 3460
rect 9732 3420 9904 3448
rect 9732 3408 9738 3420
rect 6880 3352 8340 3380
rect 8389 3383 8447 3389
rect 6880 3340 6886 3352
rect 8389 3349 8401 3383
rect 8435 3380 8447 3383
rect 8941 3383 8999 3389
rect 8941 3380 8953 3383
rect 8435 3352 8953 3380
rect 8435 3349 8447 3352
rect 8389 3343 8447 3349
rect 8941 3349 8953 3352
rect 8987 3349 8999 3383
rect 9306 3380 9312 3392
rect 9267 3352 9312 3380
rect 8941 3343 8999 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9398 3340 9404 3392
rect 9456 3380 9462 3392
rect 9766 3380 9772 3392
rect 9456 3352 9501 3380
rect 9727 3352 9772 3380
rect 9456 3340 9462 3352
rect 9766 3340 9772 3352
rect 9824 3340 9830 3392
rect 9876 3380 9904 3420
rect 9950 3408 9956 3460
rect 10008 3448 10014 3460
rect 10882 3451 10940 3457
rect 10882 3448 10894 3451
rect 10008 3420 10894 3448
rect 10008 3408 10014 3420
rect 10882 3417 10894 3420
rect 10928 3417 10940 3451
rect 10882 3411 10940 3417
rect 11054 3408 11060 3460
rect 11112 3448 11118 3460
rect 11256 3448 11284 3479
rect 12710 3476 12716 3488
rect 12768 3476 12774 3528
rect 13449 3519 13507 3525
rect 13449 3485 13461 3519
rect 13495 3485 13507 3519
rect 13722 3516 13728 3528
rect 13683 3488 13728 3516
rect 13449 3479 13507 3485
rect 11112 3420 11284 3448
rect 11793 3451 11851 3457
rect 11112 3408 11118 3420
rect 11793 3417 11805 3451
rect 11839 3417 11851 3451
rect 11793 3411 11851 3417
rect 12244 3451 12302 3457
rect 12244 3417 12256 3451
rect 12290 3448 12302 3451
rect 12434 3448 12440 3460
rect 12290 3420 12440 3448
rect 12290 3417 12302 3420
rect 12244 3411 12302 3417
rect 11808 3380 11836 3411
rect 12434 3408 12440 3420
rect 12492 3408 12498 3460
rect 13464 3448 13492 3479
rect 13722 3476 13728 3488
rect 13780 3476 13786 3528
rect 14458 3516 14464 3528
rect 14419 3488 14464 3516
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 15197 3519 15255 3525
rect 15197 3485 15209 3519
rect 15243 3516 15255 3519
rect 15470 3516 15476 3528
rect 15243 3488 15476 3516
rect 15243 3485 15255 3488
rect 15197 3479 15255 3485
rect 15470 3476 15476 3488
rect 15528 3476 15534 3528
rect 15749 3519 15807 3525
rect 15749 3485 15761 3519
rect 15795 3516 15807 3519
rect 15930 3516 15936 3528
rect 15795 3488 15936 3516
rect 15795 3485 15807 3488
rect 15749 3479 15807 3485
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 16485 3519 16543 3525
rect 16485 3485 16497 3519
rect 16531 3485 16543 3519
rect 16485 3479 16543 3485
rect 16844 3519 16902 3525
rect 16844 3485 16856 3519
rect 16890 3516 16902 3519
rect 17402 3516 17408 3528
rect 16890 3488 17408 3516
rect 16890 3485 16902 3488
rect 16844 3479 16902 3485
rect 13464 3420 14136 3448
rect 9876 3352 11836 3380
rect 13633 3383 13691 3389
rect 13633 3349 13645 3383
rect 13679 3380 13691 3383
rect 13722 3380 13728 3392
rect 13679 3352 13728 3380
rect 13679 3349 13691 3352
rect 13633 3343 13691 3349
rect 13722 3340 13728 3352
rect 13780 3340 13786 3392
rect 13814 3340 13820 3392
rect 13872 3380 13878 3392
rect 14108 3389 14136 3420
rect 14918 3408 14924 3460
rect 14976 3448 14982 3460
rect 15289 3451 15347 3457
rect 15289 3448 15301 3451
rect 14976 3420 15301 3448
rect 14976 3408 14982 3420
rect 15289 3417 15301 3420
rect 15335 3448 15347 3451
rect 16022 3448 16028 3460
rect 15335 3420 16028 3448
rect 15335 3417 15347 3420
rect 15289 3411 15347 3417
rect 16022 3408 16028 3420
rect 16080 3408 16086 3460
rect 16500 3448 16528 3479
rect 17402 3476 17408 3488
rect 17460 3516 17466 3528
rect 17770 3516 17776 3528
rect 17460 3488 17776 3516
rect 17460 3476 17466 3488
rect 17770 3476 17776 3488
rect 17828 3476 17834 3528
rect 18156 3516 18184 3547
rect 18432 3516 18460 3556
rect 19168 3528 19196 3556
rect 19702 3544 19708 3556
rect 19760 3544 19766 3596
rect 19889 3587 19947 3593
rect 19889 3553 19901 3587
rect 19935 3584 19947 3587
rect 20346 3584 20352 3596
rect 19935 3556 20352 3584
rect 19935 3553 19947 3556
rect 19889 3547 19947 3553
rect 18156 3488 18460 3516
rect 18598 3476 18604 3528
rect 18656 3516 18662 3528
rect 19061 3519 19119 3525
rect 19061 3516 19073 3519
rect 18656 3488 19073 3516
rect 18656 3476 18662 3488
rect 19061 3485 19073 3488
rect 19107 3485 19119 3519
rect 19061 3479 19119 3485
rect 19150 3476 19156 3528
rect 19208 3516 19214 3528
rect 19904 3516 19932 3547
rect 20346 3544 20352 3556
rect 20404 3544 20410 3596
rect 20070 3516 20076 3528
rect 19208 3488 19932 3516
rect 20031 3488 20076 3516
rect 19208 3476 19214 3488
rect 20070 3476 20076 3488
rect 20128 3476 20134 3528
rect 20438 3516 20444 3528
rect 20399 3488 20444 3516
rect 20438 3476 20444 3488
rect 20496 3476 20502 3528
rect 20806 3516 20812 3528
rect 20767 3488 20812 3516
rect 20806 3476 20812 3488
rect 20864 3476 20870 3528
rect 21453 3519 21511 3525
rect 21453 3485 21465 3519
rect 21499 3516 21511 3519
rect 22002 3516 22008 3528
rect 21499 3488 22008 3516
rect 21499 3485 21511 3488
rect 21453 3479 21511 3485
rect 22002 3476 22008 3488
rect 22060 3476 22066 3528
rect 17954 3448 17960 3460
rect 16500 3420 17960 3448
rect 17954 3408 17960 3420
rect 18012 3408 18018 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 19576 3420 20668 3448
rect 19576 3408 19582 3420
rect 13909 3383 13967 3389
rect 13909 3380 13921 3383
rect 13872 3352 13921 3380
rect 13872 3340 13878 3352
rect 13909 3349 13921 3352
rect 13955 3349 13967 3383
rect 13909 3343 13967 3349
rect 14093 3383 14151 3389
rect 14093 3349 14105 3383
rect 14139 3349 14151 3383
rect 15930 3380 15936 3392
rect 15891 3352 15936 3380
rect 14093 3343 14151 3349
rect 15930 3340 15936 3352
rect 15988 3340 15994 3392
rect 16298 3380 16304 3392
rect 16259 3352 16304 3380
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 18414 3340 18420 3392
rect 18472 3380 18478 3392
rect 18472 3352 18517 3380
rect 18472 3340 18478 3352
rect 18782 3340 18788 3392
rect 18840 3380 18846 3392
rect 18877 3383 18935 3389
rect 18877 3380 18889 3383
rect 18840 3352 18889 3380
rect 18840 3340 18846 3352
rect 18877 3349 18889 3352
rect 18923 3349 18935 3383
rect 19610 3380 19616 3392
rect 19571 3352 19616 3380
rect 18877 3343 18935 3349
rect 19610 3340 19616 3352
rect 19668 3340 19674 3392
rect 19794 3340 19800 3392
rect 19852 3380 19858 3392
rect 20640 3389 20668 3420
rect 20257 3383 20315 3389
rect 20257 3380 20269 3383
rect 19852 3352 20269 3380
rect 19852 3340 19858 3352
rect 20257 3349 20269 3352
rect 20303 3349 20315 3383
rect 20257 3343 20315 3349
rect 20625 3383 20683 3389
rect 20625 3349 20637 3383
rect 20671 3349 20683 3383
rect 21358 3380 21364 3392
rect 21319 3352 21364 3380
rect 20625 3343 20683 3349
rect 21358 3340 21364 3352
rect 21416 3340 21422 3392
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 5810 3136 5816 3188
rect 5868 3176 5874 3188
rect 6181 3179 6239 3185
rect 6181 3176 6193 3179
rect 5868 3148 6193 3176
rect 5868 3136 5874 3148
rect 6181 3145 6193 3148
rect 6227 3176 6239 3179
rect 6546 3176 6552 3188
rect 6227 3148 6552 3176
rect 6227 3145 6239 3148
rect 6181 3139 6239 3145
rect 6546 3136 6552 3148
rect 6604 3136 6610 3188
rect 6730 3136 6736 3188
rect 6788 3176 6794 3188
rect 7193 3179 7251 3185
rect 7193 3176 7205 3179
rect 6788 3148 7205 3176
rect 6788 3136 6794 3148
rect 7193 3145 7205 3148
rect 7239 3145 7251 3179
rect 7193 3139 7251 3145
rect 7285 3179 7343 3185
rect 7285 3145 7297 3179
rect 7331 3176 7343 3179
rect 7834 3176 7840 3188
rect 7331 3148 7840 3176
rect 7331 3145 7343 3148
rect 7285 3139 7343 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8202 3136 8208 3188
rect 8260 3176 8266 3188
rect 8938 3176 8944 3188
rect 8260 3148 8944 3176
rect 8260 3136 8266 3148
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9030 3136 9036 3188
rect 9088 3176 9094 3188
rect 9490 3176 9496 3188
rect 9088 3148 9496 3176
rect 9088 3136 9094 3148
rect 9490 3136 9496 3148
rect 9548 3136 9554 3188
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9950 3176 9956 3188
rect 9911 3148 9956 3176
rect 9950 3136 9956 3148
rect 10008 3136 10014 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 10778 3176 10784 3188
rect 10192 3148 10784 3176
rect 10192 3136 10198 3148
rect 10778 3136 10784 3148
rect 10836 3136 10842 3188
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 14918 3176 14924 3188
rect 11296 3148 14412 3176
rect 14831 3148 14924 3176
rect 11296 3136 11302 3148
rect 2590 3108 2596 3120
rect 2551 3080 2596 3108
rect 2590 3068 2596 3080
rect 2648 3068 2654 3120
rect 2777 3111 2835 3117
rect 2777 3077 2789 3111
rect 2823 3108 2835 3111
rect 3050 3108 3056 3120
rect 2823 3080 3056 3108
rect 2823 3077 2835 3080
rect 2777 3071 2835 3077
rect 3050 3068 3056 3080
rect 3108 3068 3114 3120
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 8294 3108 8300 3120
rect 4387 3080 8300 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 9766 3108 9772 3120
rect 9727 3080 9772 3108
rect 9766 3068 9772 3080
rect 9824 3068 9830 3120
rect 11330 3068 11336 3120
rect 11388 3108 11394 3120
rect 11790 3108 11796 3120
rect 11388 3080 11796 3108
rect 11388 3068 11394 3080
rect 11790 3068 11796 3080
rect 11848 3068 11854 3120
rect 11885 3111 11943 3117
rect 11885 3077 11897 3111
rect 11931 3108 11943 3111
rect 12342 3108 12348 3120
rect 11931 3080 12348 3108
rect 11931 3077 11943 3080
rect 11885 3071 11943 3077
rect 12342 3068 12348 3080
rect 12400 3068 12406 3120
rect 12437 3111 12495 3117
rect 12437 3077 12449 3111
rect 12483 3108 12495 3111
rect 12980 3111 13038 3117
rect 12483 3080 12572 3108
rect 12483 3077 12495 3080
rect 12437 3071 12495 3077
rect 566 3000 572 3052
rect 624 3040 630 3052
rect 2225 3043 2283 3049
rect 2225 3040 2237 3043
rect 624 3012 2237 3040
rect 624 3000 630 3012
rect 2225 3009 2237 3012
rect 2271 3040 2283 3043
rect 2406 3040 2412 3052
rect 2271 3012 2412 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2406 3000 2412 3012
rect 2464 3000 2470 3052
rect 3993 3043 4051 3049
rect 3993 3009 4005 3043
rect 4039 3040 4051 3043
rect 4154 3040 4160 3052
rect 4039 3012 4160 3040
rect 4039 3009 4051 3012
rect 3993 3003 4051 3009
rect 4154 3000 4160 3012
rect 4212 3000 4218 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3040 4307 3043
rect 4430 3040 4436 3052
rect 4295 3012 4436 3040
rect 4295 3009 4307 3012
rect 4249 3003 4307 3009
rect 4430 3000 4436 3012
rect 4488 3040 4494 3052
rect 4798 3049 4804 3052
rect 4525 3043 4583 3049
rect 4525 3040 4537 3043
rect 4488 3012 4537 3040
rect 4488 3000 4494 3012
rect 4525 3009 4537 3012
rect 4571 3009 4583 3043
rect 4792 3040 4804 3049
rect 4759 3012 4804 3040
rect 4525 3003 4583 3009
rect 4792 3003 4804 3012
rect 4798 3000 4804 3003
rect 4856 3000 4862 3052
rect 5350 3000 5356 3052
rect 5408 3040 5414 3052
rect 5997 3043 6055 3049
rect 5408 3012 5580 3040
rect 5408 3000 5414 3012
rect 1946 2972 1952 2984
rect 1907 2944 1952 2972
rect 1946 2932 1952 2944
rect 2004 2932 2010 2984
rect 4172 2972 4200 3000
rect 4172 2944 4283 2972
rect 2869 2907 2927 2913
rect 2869 2873 2881 2907
rect 2915 2904 2927 2907
rect 2958 2904 2964 2916
rect 2915 2876 2964 2904
rect 2915 2873 2927 2876
rect 2869 2867 2927 2873
rect 2958 2864 2964 2876
rect 3016 2864 3022 2916
rect 2409 2839 2467 2845
rect 2409 2805 2421 2839
rect 2455 2836 2467 2839
rect 4062 2836 4068 2848
rect 2455 2808 4068 2836
rect 2455 2805 2467 2808
rect 2409 2799 2467 2805
rect 4062 2796 4068 2808
rect 4120 2796 4126 2848
rect 4255 2836 4283 2944
rect 5552 2904 5580 3012
rect 5997 3009 6009 3043
rect 6043 3040 6055 3043
rect 6086 3040 6092 3052
rect 6043 3012 6092 3040
rect 6043 3009 6055 3012
rect 5997 3003 6055 3009
rect 6086 3000 6092 3012
rect 6144 3000 6150 3052
rect 6641 3043 6699 3049
rect 6641 3009 6653 3043
rect 6687 3040 6699 3043
rect 7650 3040 7656 3052
rect 6687 3012 7656 3040
rect 6687 3009 6699 3012
rect 6641 3003 6699 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7926 3000 7932 3052
rect 7984 3040 7990 3052
rect 8858 3043 8916 3049
rect 8858 3040 8870 3043
rect 7984 3012 8870 3040
rect 7984 3000 7990 3012
rect 8858 3009 8870 3012
rect 8904 3009 8916 3043
rect 9122 3040 9128 3052
rect 9083 3012 9128 3040
rect 8858 3003 8916 3009
rect 9122 3000 9128 3012
rect 9180 3000 9186 3052
rect 9401 3043 9459 3049
rect 9401 3009 9413 3043
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 11077 3043 11135 3049
rect 11077 3009 11089 3043
rect 11123 3040 11135 3043
rect 11123 3012 11468 3040
rect 11123 3009 11135 3012
rect 11077 3003 11135 3009
rect 5626 2932 5632 2984
rect 5684 2972 5690 2984
rect 6822 2972 6828 2984
rect 5684 2944 6828 2972
rect 5684 2932 5690 2944
rect 6822 2932 6828 2944
rect 6880 2932 6886 2984
rect 7098 2932 7104 2984
rect 7156 2972 7162 2984
rect 7668 2972 7696 3000
rect 8018 2972 8024 2984
rect 7156 2944 7201 2972
rect 7668 2944 8024 2972
rect 7156 2932 7162 2944
rect 8018 2932 8024 2944
rect 8076 2932 8082 2984
rect 6546 2904 6552 2916
rect 5552 2876 6552 2904
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 7653 2907 7711 2913
rect 7653 2873 7665 2907
rect 7699 2904 7711 2907
rect 9416 2904 9444 3003
rect 11330 2972 11336 2984
rect 11291 2944 11336 2972
rect 11330 2932 11336 2944
rect 11388 2932 11394 2984
rect 9858 2904 9864 2916
rect 7699 2876 8156 2904
rect 9416 2876 9864 2904
rect 7699 2873 7711 2876
rect 7653 2867 7711 2873
rect 5902 2836 5908 2848
rect 4255 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 5994 2796 6000 2848
rect 6052 2836 6058 2848
rect 6365 2839 6423 2845
rect 6365 2836 6377 2839
rect 6052 2808 6377 2836
rect 6052 2796 6058 2808
rect 6365 2805 6377 2808
rect 6411 2805 6423 2839
rect 6365 2799 6423 2805
rect 6733 2839 6791 2845
rect 6733 2805 6745 2839
rect 6779 2836 6791 2839
rect 7006 2836 7012 2848
rect 6779 2808 7012 2836
rect 6779 2805 6791 2808
rect 6733 2799 6791 2805
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 7742 2836 7748 2848
rect 7703 2808 7748 2836
rect 7742 2796 7748 2808
rect 7800 2796 7806 2848
rect 8128 2836 8156 2876
rect 9858 2864 9864 2876
rect 9916 2864 9922 2916
rect 11440 2904 11468 3012
rect 11514 3000 11520 3052
rect 11572 3040 11578 3052
rect 11572 3012 12112 3040
rect 11572 3000 11578 3012
rect 11790 2932 11796 2984
rect 11848 2972 11854 2984
rect 12084 2981 12112 3012
rect 11977 2975 12035 2981
rect 11977 2972 11989 2975
rect 11848 2944 11989 2972
rect 11848 2932 11854 2944
rect 11977 2941 11989 2944
rect 12023 2941 12035 2975
rect 11977 2935 12035 2941
rect 12069 2975 12127 2981
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12544 2972 12572 3080
rect 12980 3077 12992 3111
rect 13026 3108 13038 3111
rect 13354 3108 13360 3120
rect 13026 3080 13360 3108
rect 13026 3077 13038 3080
rect 12980 3071 13038 3077
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 12710 3040 12716 3052
rect 12671 3012 12716 3040
rect 12710 3000 12716 3012
rect 12768 3000 12774 3052
rect 14384 3049 14412 3148
rect 14918 3136 14924 3148
rect 14976 3176 14982 3188
rect 15194 3176 15200 3188
rect 14976 3148 15200 3176
rect 14976 3136 14982 3148
rect 15194 3136 15200 3148
rect 15252 3136 15258 3188
rect 16025 3179 16083 3185
rect 16025 3145 16037 3179
rect 16071 3145 16083 3179
rect 16025 3139 16083 3145
rect 16393 3179 16451 3185
rect 16393 3145 16405 3179
rect 16439 3176 16451 3179
rect 18506 3176 18512 3188
rect 16439 3148 18368 3176
rect 18467 3148 18512 3176
rect 16439 3145 16451 3148
rect 16393 3139 16451 3145
rect 15010 3068 15016 3120
rect 15068 3108 15074 3120
rect 16040 3108 16068 3139
rect 15068 3080 15884 3108
rect 16040 3080 18000 3108
rect 15068 3068 15074 3080
rect 14369 3043 14427 3049
rect 14369 3009 14381 3043
rect 14415 3009 14427 3043
rect 14369 3003 14427 3009
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 14737 3043 14795 3049
rect 14737 3009 14749 3043
rect 14783 3040 14795 3043
rect 14826 3040 14832 3052
rect 14783 3012 14832 3040
rect 14783 3009 14795 3012
rect 14737 3003 14795 3009
rect 12618 2972 12624 2984
rect 12544 2944 12624 2972
rect 12069 2935 12127 2941
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 13722 2932 13728 2984
rect 13780 2972 13786 2984
rect 14660 2972 14688 3003
rect 14826 3000 14832 3012
rect 14884 3000 14890 3052
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15746 3040 15752 3052
rect 15707 3012 15752 3040
rect 15746 3000 15752 3012
rect 15804 3000 15810 3052
rect 15856 3049 15884 3080
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3009 15899 3043
rect 16206 3040 16212 3052
rect 16167 3012 16212 3040
rect 15841 3003 15899 3009
rect 16206 3000 16212 3012
rect 16264 3000 16270 3052
rect 16853 3043 16911 3049
rect 16853 3009 16865 3043
rect 16899 3009 16911 3043
rect 16853 3003 16911 3009
rect 13780 2944 14688 2972
rect 13780 2932 13786 2944
rect 16022 2932 16028 2984
rect 16080 2972 16086 2984
rect 16868 2972 16896 3003
rect 16942 3000 16948 3052
rect 17000 3040 17006 3052
rect 17310 3040 17316 3052
rect 17000 3012 17045 3040
rect 17271 3012 17316 3040
rect 17000 3000 17006 3012
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 17586 3000 17592 3052
rect 17644 3040 17650 3052
rect 17972 3040 18000 3080
rect 18046 3068 18052 3120
rect 18104 3108 18110 3120
rect 18104 3080 18149 3108
rect 18104 3068 18110 3080
rect 18230 3040 18236 3052
rect 17644 3012 17908 3040
rect 17972 3012 18236 3040
rect 17644 3000 17650 3012
rect 17770 2972 17776 2984
rect 16080 2944 16896 2972
rect 17731 2944 17776 2972
rect 16080 2932 16086 2944
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 17880 2972 17908 3012
rect 18230 3000 18236 3012
rect 18288 3000 18294 3052
rect 17957 2975 18015 2981
rect 17957 2972 17969 2975
rect 17880 2944 17969 2972
rect 17957 2941 17969 2944
rect 18003 2941 18015 2975
rect 17957 2935 18015 2941
rect 14642 2904 14648 2916
rect 11440 2876 12756 2904
rect 8478 2836 8484 2848
rect 8128 2808 8484 2836
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 9309 2839 9367 2845
rect 9309 2805 9321 2839
rect 9355 2836 9367 2839
rect 10042 2836 10048 2848
rect 9355 2808 10048 2836
rect 9355 2805 9367 2808
rect 9309 2799 9367 2805
rect 10042 2796 10048 2808
rect 10100 2796 10106 2848
rect 10134 2796 10140 2848
rect 10192 2836 10198 2848
rect 11422 2836 11428 2848
rect 10192 2808 11428 2836
rect 10192 2796 10198 2808
rect 11422 2796 11428 2808
rect 11480 2796 11486 2848
rect 11517 2839 11575 2845
rect 11517 2805 11529 2839
rect 11563 2836 11575 2839
rect 11698 2836 11704 2848
rect 11563 2808 11704 2836
rect 11563 2805 11575 2808
rect 11517 2799 11575 2805
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 12434 2796 12440 2848
rect 12492 2836 12498 2848
rect 12529 2839 12587 2845
rect 12529 2836 12541 2839
rect 12492 2808 12541 2836
rect 12492 2796 12498 2808
rect 12529 2805 12541 2808
rect 12575 2805 12587 2839
rect 12728 2836 12756 2876
rect 14108 2876 14648 2904
rect 14108 2845 14136 2876
rect 14642 2864 14648 2876
rect 14700 2864 14706 2916
rect 15194 2904 15200 2916
rect 15155 2876 15200 2904
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 15562 2904 15568 2916
rect 15523 2876 15568 2904
rect 15562 2864 15568 2876
rect 15620 2864 15626 2916
rect 14093 2839 14151 2845
rect 14093 2836 14105 2839
rect 12728 2808 14105 2836
rect 12529 2799 12587 2805
rect 14093 2805 14105 2808
rect 14139 2805 14151 2839
rect 14093 2799 14151 2805
rect 14185 2839 14243 2845
rect 14185 2805 14197 2839
rect 14231 2836 14243 2839
rect 14274 2836 14280 2848
rect 14231 2808 14280 2836
rect 14231 2805 14243 2808
rect 14185 2799 14243 2805
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 14458 2836 14464 2848
rect 14419 2808 14464 2836
rect 14458 2796 14464 2808
rect 14516 2796 14522 2848
rect 16666 2836 16672 2848
rect 16627 2808 16672 2836
rect 16666 2796 16672 2808
rect 16724 2796 16730 2848
rect 17129 2839 17187 2845
rect 17129 2805 17141 2839
rect 17175 2836 17187 2839
rect 17218 2836 17224 2848
rect 17175 2808 17224 2836
rect 17175 2805 17187 2808
rect 17129 2799 17187 2805
rect 17218 2796 17224 2808
rect 17276 2796 17282 2848
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 17497 2839 17555 2845
rect 17497 2836 17509 2839
rect 17368 2808 17509 2836
rect 17368 2796 17374 2808
rect 17497 2805 17509 2808
rect 17543 2805 17555 2839
rect 18340 2836 18368 3148
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 18874 3136 18880 3188
rect 18932 3136 18938 3188
rect 18969 3179 19027 3185
rect 18969 3145 18981 3179
rect 19015 3176 19027 3179
rect 19337 3179 19395 3185
rect 19337 3176 19349 3179
rect 19015 3148 19349 3176
rect 19015 3145 19027 3148
rect 18969 3139 19027 3145
rect 19337 3145 19349 3148
rect 19383 3145 19395 3179
rect 19337 3139 19395 3145
rect 19705 3179 19763 3185
rect 19705 3145 19717 3179
rect 19751 3176 19763 3179
rect 21082 3176 21088 3188
rect 19751 3148 21088 3176
rect 19751 3145 19763 3148
rect 19705 3139 19763 3145
rect 21082 3136 21088 3148
rect 21140 3136 21146 3188
rect 18892 3108 18920 3136
rect 19794 3108 19800 3120
rect 18892 3080 19800 3108
rect 19794 3068 19800 3080
rect 19852 3068 19858 3120
rect 20622 3108 20628 3120
rect 20583 3080 20628 3108
rect 20622 3068 20628 3080
rect 20680 3068 20686 3120
rect 18877 3043 18935 3049
rect 18877 3040 18889 3043
rect 18524 3012 18889 3040
rect 18417 2907 18475 2913
rect 18417 2873 18429 2907
rect 18463 2904 18475 2907
rect 18524 2904 18552 3012
rect 18877 3009 18889 3012
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 18966 3000 18972 3052
rect 19024 3040 19030 3052
rect 19024 3012 19932 3040
rect 19024 3000 19030 3012
rect 19150 2972 19156 2984
rect 19111 2944 19156 2972
rect 19150 2932 19156 2944
rect 19208 2932 19214 2984
rect 19702 2932 19708 2984
rect 19760 2972 19766 2984
rect 19904 2981 19932 3012
rect 19978 3000 19984 3052
rect 20036 3040 20042 3052
rect 20165 3043 20223 3049
rect 20165 3040 20177 3043
rect 20036 3012 20177 3040
rect 20036 3000 20042 3012
rect 20165 3009 20177 3012
rect 20211 3009 20223 3043
rect 20714 3040 20720 3052
rect 20675 3012 20720 3040
rect 20165 3003 20223 3009
rect 20714 3000 20720 3012
rect 20772 3000 20778 3052
rect 19797 2975 19855 2981
rect 19797 2972 19809 2975
rect 19760 2944 19809 2972
rect 19760 2932 19766 2944
rect 19797 2941 19809 2944
rect 19843 2941 19855 2975
rect 19797 2935 19855 2941
rect 19889 2975 19947 2981
rect 19889 2941 19901 2975
rect 19935 2941 19947 2975
rect 19889 2935 19947 2941
rect 20530 2932 20536 2984
rect 20588 2972 20594 2984
rect 20993 2975 21051 2981
rect 20993 2972 21005 2975
rect 20588 2944 21005 2972
rect 20588 2932 20594 2944
rect 20993 2941 21005 2944
rect 21039 2941 21051 2975
rect 20993 2935 21051 2941
rect 18463 2876 18552 2904
rect 18463 2873 18475 2876
rect 18417 2867 18475 2873
rect 19058 2864 19064 2916
rect 19116 2904 19122 2916
rect 20622 2904 20628 2916
rect 19116 2876 20628 2904
rect 19116 2864 19122 2876
rect 20622 2864 20628 2876
rect 20680 2864 20686 2916
rect 18506 2836 18512 2848
rect 18340 2808 18512 2836
rect 17497 2799 17555 2805
rect 18506 2796 18512 2808
rect 18564 2796 18570 2848
rect 18598 2796 18604 2848
rect 18656 2836 18662 2848
rect 20349 2839 20407 2845
rect 20349 2836 20361 2839
rect 18656 2808 20361 2836
rect 18656 2796 18662 2808
rect 20349 2805 20361 2808
rect 20395 2805 20407 2839
rect 20349 2799 20407 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3375 2635 3433 2641
rect 3375 2601 3387 2635
rect 3421 2632 3433 2635
rect 5718 2632 5724 2644
rect 3421 2604 5724 2632
rect 3421 2601 3433 2604
rect 3375 2595 3433 2601
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 6086 2592 6092 2644
rect 6144 2632 6150 2644
rect 6914 2632 6920 2644
rect 6144 2604 6920 2632
rect 6144 2592 6150 2604
rect 6914 2592 6920 2604
rect 6972 2592 6978 2644
rect 9122 2632 9128 2644
rect 9083 2604 9128 2632
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 12345 2635 12403 2641
rect 12345 2632 12357 2635
rect 9232 2604 12357 2632
rect 5169 2567 5227 2573
rect 5169 2533 5181 2567
rect 5215 2564 5227 2567
rect 7558 2564 7564 2576
rect 5215 2536 7564 2564
rect 5215 2533 5227 2536
rect 5169 2527 5227 2533
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 7650 2524 7656 2576
rect 7708 2564 7714 2576
rect 9232 2564 9260 2604
rect 12345 2601 12357 2604
rect 12391 2601 12403 2635
rect 12345 2595 12403 2601
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 13265 2635 13323 2641
rect 13265 2632 13277 2635
rect 12768 2604 13277 2632
rect 12768 2592 12774 2604
rect 13265 2601 13277 2604
rect 13311 2601 13323 2635
rect 14274 2632 14280 2644
rect 13265 2595 13323 2601
rect 13740 2604 14280 2632
rect 7708 2536 9260 2564
rect 7708 2524 7714 2536
rect 9306 2524 9312 2576
rect 9364 2564 9370 2576
rect 10229 2567 10287 2573
rect 10229 2564 10241 2567
rect 9364 2536 10241 2564
rect 9364 2524 9370 2536
rect 10229 2533 10241 2536
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 12066 2564 12072 2576
rect 10744 2536 12072 2564
rect 10744 2524 10750 2536
rect 12066 2524 12072 2536
rect 12124 2524 12130 2576
rect 12253 2567 12311 2573
rect 12253 2533 12265 2567
rect 12299 2564 12311 2567
rect 12299 2536 12434 2564
rect 12299 2533 12311 2536
rect 12253 2527 12311 2533
rect 2222 2456 2228 2508
rect 2280 2496 2286 2508
rect 2682 2496 2688 2508
rect 2280 2468 2688 2496
rect 2280 2456 2286 2468
rect 2682 2456 2688 2468
rect 2740 2456 2746 2508
rect 2774 2456 2780 2508
rect 2832 2496 2838 2508
rect 3605 2499 3663 2505
rect 3605 2496 3617 2499
rect 2832 2468 3617 2496
rect 2832 2456 2838 2468
rect 3605 2465 3617 2468
rect 3651 2465 3663 2499
rect 5810 2496 5816 2508
rect 5771 2468 5816 2496
rect 3605 2459 3663 2465
rect 5810 2456 5816 2468
rect 5868 2456 5874 2508
rect 6917 2499 6975 2505
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 7006 2496 7012 2508
rect 6963 2468 7012 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8168 2468 9720 2496
rect 8168 2456 8174 2468
rect 1762 2428 1768 2440
rect 1723 2400 1768 2428
rect 1762 2388 1768 2400
rect 1820 2388 1826 2440
rect 2406 2428 2412 2440
rect 2367 2400 2412 2428
rect 2406 2388 2412 2400
rect 2464 2388 2470 2440
rect 3789 2431 3847 2437
rect 3789 2397 3801 2431
rect 3835 2397 3847 2431
rect 3789 2391 3847 2397
rect 3804 2360 3832 2391
rect 3878 2388 3884 2440
rect 3936 2428 3942 2440
rect 4045 2431 4103 2437
rect 4045 2428 4057 2431
rect 3936 2400 4057 2428
rect 3936 2388 3942 2400
rect 4045 2397 4057 2400
rect 4091 2397 4103 2431
rect 4045 2391 4103 2397
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 6089 2431 6147 2437
rect 6089 2428 6101 2431
rect 4856 2400 6101 2428
rect 4856 2388 4862 2400
rect 6089 2397 6101 2400
rect 6135 2397 6147 2431
rect 7190 2428 7196 2440
rect 7151 2400 7196 2428
rect 6089 2391 6147 2397
rect 7190 2388 7196 2400
rect 7248 2388 7254 2440
rect 7926 2428 7932 2440
rect 7887 2400 7932 2428
rect 7926 2388 7932 2400
rect 7984 2388 7990 2440
rect 8205 2431 8263 2437
rect 8205 2397 8217 2431
rect 8251 2397 8263 2431
rect 8205 2391 8263 2397
rect 8665 2431 8723 2437
rect 8665 2397 8677 2431
rect 8711 2428 8723 2431
rect 8754 2428 8760 2440
rect 8711 2400 8760 2428
rect 8711 2397 8723 2400
rect 8665 2391 8723 2397
rect 4430 2360 4436 2372
rect 3804 2332 4436 2360
rect 4430 2320 4436 2332
rect 4488 2320 4494 2372
rect 7282 2320 7288 2372
rect 7340 2360 7346 2372
rect 8220 2360 8248 2391
rect 8754 2388 8760 2400
rect 8812 2388 8818 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9490 2428 9496 2440
rect 9355 2400 9496 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9490 2388 9496 2400
rect 9548 2388 9554 2440
rect 9692 2428 9720 2468
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 9953 2499 10011 2505
rect 9953 2496 9965 2499
rect 9824 2468 9965 2496
rect 9824 2456 9830 2468
rect 9953 2465 9965 2468
rect 9999 2465 10011 2499
rect 10778 2496 10784 2508
rect 10739 2468 10784 2496
rect 9953 2459 10011 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 11609 2499 11667 2505
rect 11609 2496 11621 2499
rect 10928 2468 11621 2496
rect 10928 2456 10934 2468
rect 11609 2465 11621 2468
rect 11655 2465 11667 2499
rect 11609 2459 11667 2465
rect 11698 2456 11704 2508
rect 11756 2496 11762 2508
rect 11793 2499 11851 2505
rect 11793 2496 11805 2499
rect 11756 2468 11805 2496
rect 11756 2456 11762 2468
rect 11793 2465 11805 2468
rect 11839 2465 11851 2499
rect 12406 2496 12434 2536
rect 13078 2524 13084 2576
rect 13136 2564 13142 2576
rect 13633 2567 13691 2573
rect 13633 2564 13645 2567
rect 13136 2536 13645 2564
rect 13136 2524 13142 2536
rect 13633 2533 13645 2536
rect 13679 2533 13691 2567
rect 13633 2527 13691 2533
rect 12406 2468 12480 2496
rect 11793 2459 11851 2465
rect 9692 2400 9996 2428
rect 7340 2332 8248 2360
rect 7340 2320 7346 2332
rect 9582 2320 9588 2372
rect 9640 2360 9646 2372
rect 9861 2363 9919 2369
rect 9861 2360 9873 2363
rect 9640 2332 9873 2360
rect 9640 2320 9646 2332
rect 9861 2329 9873 2332
rect 9907 2329 9919 2363
rect 9968 2360 9996 2400
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 10597 2431 10655 2437
rect 10597 2428 10609 2431
rect 10560 2400 10609 2428
rect 10560 2388 10566 2400
rect 10597 2397 10609 2400
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10686 2388 10692 2440
rect 10744 2428 10750 2440
rect 10744 2400 10789 2428
rect 10744 2388 10750 2400
rect 11146 2388 11152 2440
rect 11204 2428 11210 2440
rect 11241 2431 11299 2437
rect 11241 2428 11253 2431
rect 11204 2400 11253 2428
rect 11204 2388 11210 2400
rect 11241 2397 11253 2400
rect 11287 2397 11299 2431
rect 11882 2428 11888 2440
rect 11843 2400 11888 2428
rect 11241 2391 11299 2397
rect 11882 2388 11888 2400
rect 11940 2388 11946 2440
rect 11057 2363 11115 2369
rect 11057 2360 11069 2363
rect 9968 2332 11069 2360
rect 9861 2323 9919 2329
rect 11057 2329 11069 2332
rect 11103 2329 11115 2363
rect 12452 2360 12480 2468
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12584 2468 12909 2496
rect 12584 2456 12590 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 13449 2431 13507 2437
rect 13449 2397 13461 2431
rect 13495 2428 13507 2431
rect 13740 2428 13768 2604
rect 14274 2592 14280 2604
rect 14332 2592 14338 2644
rect 15930 2592 15936 2644
rect 15988 2632 15994 2644
rect 15988 2604 18000 2632
rect 15988 2592 15994 2604
rect 13814 2524 13820 2576
rect 13872 2524 13878 2576
rect 13998 2524 14004 2576
rect 14056 2564 14062 2576
rect 14553 2567 14611 2573
rect 14553 2564 14565 2567
rect 14056 2536 14565 2564
rect 14056 2524 14062 2536
rect 14553 2533 14565 2536
rect 14599 2533 14611 2567
rect 14553 2527 14611 2533
rect 14826 2524 14832 2576
rect 14884 2564 14890 2576
rect 15289 2567 15347 2573
rect 15289 2564 15301 2567
rect 14884 2536 15301 2564
rect 14884 2524 14890 2536
rect 15289 2533 15301 2536
rect 15335 2533 15347 2567
rect 15289 2527 15347 2533
rect 16022 2524 16028 2576
rect 16080 2564 16086 2576
rect 16761 2567 16819 2573
rect 16761 2564 16773 2567
rect 16080 2536 16773 2564
rect 16080 2524 16086 2536
rect 16761 2533 16773 2536
rect 16807 2533 16819 2567
rect 16761 2527 16819 2533
rect 16942 2524 16948 2576
rect 17000 2564 17006 2576
rect 17497 2567 17555 2573
rect 17497 2564 17509 2567
rect 17000 2536 17509 2564
rect 17000 2524 17006 2536
rect 17497 2533 17509 2536
rect 17543 2533 17555 2567
rect 17497 2527 17555 2533
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2533 17831 2567
rect 17773 2527 17831 2533
rect 13832 2496 13860 2524
rect 16666 2496 16672 2508
rect 13832 2468 14136 2496
rect 14108 2437 14136 2468
rect 15488 2468 16672 2496
rect 13495 2400 13768 2428
rect 13817 2431 13875 2437
rect 13495 2397 13507 2400
rect 13449 2391 13507 2397
rect 13817 2397 13829 2431
rect 13863 2397 13875 2431
rect 13817 2391 13875 2397
rect 14093 2431 14151 2437
rect 14093 2397 14105 2431
rect 14139 2397 14151 2431
rect 14734 2428 14740 2440
rect 14695 2400 14740 2428
rect 14093 2391 14151 2397
rect 12805 2363 12863 2369
rect 12805 2360 12817 2363
rect 12452 2332 12817 2360
rect 11057 2323 11115 2329
rect 12805 2329 12817 2332
rect 12851 2329 12863 2363
rect 13832 2360 13860 2391
rect 14734 2388 14740 2400
rect 14792 2388 14798 2440
rect 15488 2437 15516 2468
rect 16666 2456 16672 2468
rect 16724 2456 16730 2508
rect 17788 2496 17816 2527
rect 16960 2468 17816 2496
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2397 14887 2431
rect 14829 2391 14887 2397
rect 15473 2431 15531 2437
rect 15473 2397 15485 2431
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 15841 2431 15899 2437
rect 15841 2397 15853 2431
rect 15887 2397 15899 2431
rect 15841 2391 15899 2397
rect 14458 2360 14464 2372
rect 13832 2332 14464 2360
rect 12805 2323 12863 2329
rect 14458 2320 14464 2332
rect 14516 2320 14522 2372
rect 14550 2320 14556 2372
rect 14608 2360 14614 2372
rect 14844 2360 14872 2391
rect 14608 2332 14872 2360
rect 15856 2360 15884 2391
rect 15930 2388 15936 2440
rect 15988 2428 15994 2440
rect 15988 2400 16033 2428
rect 15988 2388 15994 2400
rect 16206 2388 16212 2440
rect 16264 2428 16270 2440
rect 16960 2437 16988 2468
rect 17972 2437 18000 2604
rect 18414 2592 18420 2644
rect 18472 2632 18478 2644
rect 18785 2635 18843 2641
rect 18785 2632 18797 2635
rect 18472 2604 18797 2632
rect 18472 2592 18478 2604
rect 18785 2601 18797 2604
rect 18831 2601 18843 2635
rect 18785 2595 18843 2601
rect 19705 2635 19763 2641
rect 19705 2601 19717 2635
rect 19751 2632 19763 2635
rect 19886 2632 19892 2644
rect 19751 2604 19892 2632
rect 19751 2601 19763 2604
rect 19705 2595 19763 2601
rect 19886 2592 19892 2604
rect 19944 2592 19950 2644
rect 20990 2564 20996 2576
rect 20640 2536 20996 2564
rect 18230 2505 18236 2508
rect 18187 2499 18236 2505
rect 18187 2465 18199 2499
rect 18233 2465 18236 2499
rect 18187 2459 18236 2465
rect 18230 2456 18236 2459
rect 18288 2456 18294 2508
rect 18322 2456 18328 2508
rect 18380 2496 18386 2508
rect 20640 2496 20668 2536
rect 20990 2524 20996 2536
rect 21048 2524 21054 2576
rect 21726 2524 21732 2576
rect 21784 2564 21790 2576
rect 22646 2564 22652 2576
rect 21784 2536 22652 2564
rect 21784 2524 21790 2536
rect 22646 2524 22652 2536
rect 22704 2524 22710 2576
rect 22186 2496 22192 2508
rect 18380 2468 18425 2496
rect 18892 2468 20668 2496
rect 20732 2468 22192 2496
rect 18380 2456 18386 2468
rect 16485 2431 16543 2437
rect 16485 2428 16497 2431
rect 16264 2400 16497 2428
rect 16264 2388 16270 2400
rect 16485 2397 16497 2400
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 16945 2431 17003 2437
rect 16945 2397 16957 2431
rect 16991 2397 17003 2431
rect 16945 2391 17003 2397
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2397 17371 2431
rect 17313 2391 17371 2397
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2397 17739 2431
rect 17681 2391 17739 2397
rect 17957 2431 18015 2437
rect 17957 2397 17969 2431
rect 18003 2397 18015 2431
rect 18414 2428 18420 2440
rect 18375 2400 18420 2428
rect 17957 2391 18015 2397
rect 15856 2332 16344 2360
rect 14608 2320 14614 2332
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 3878 2292 3884 2304
rect 1627 2264 3884 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 7466 2292 7472 2304
rect 4120 2264 7472 2292
rect 4120 2252 4126 2264
rect 7466 2252 7472 2264
rect 7524 2252 7530 2304
rect 8202 2252 8208 2304
rect 8260 2292 8266 2304
rect 8297 2295 8355 2301
rect 8297 2292 8309 2295
rect 8260 2264 8309 2292
rect 8260 2252 8266 2264
rect 8297 2261 8309 2264
rect 8343 2261 8355 2295
rect 8570 2292 8576 2304
rect 8531 2264 8576 2292
rect 8297 2255 8355 2261
rect 8570 2252 8576 2264
rect 8628 2252 8634 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9401 2295 9459 2301
rect 9401 2292 9413 2295
rect 9364 2264 9413 2292
rect 9364 2252 9370 2264
rect 9401 2261 9413 2264
rect 9447 2261 9459 2295
rect 9766 2292 9772 2304
rect 9727 2264 9772 2292
rect 9401 2255 9459 2261
rect 9766 2252 9772 2264
rect 9824 2292 9830 2304
rect 12158 2292 12164 2304
rect 9824 2264 12164 2292
rect 9824 2252 9830 2264
rect 12158 2252 12164 2264
rect 12216 2252 12222 2304
rect 12434 2252 12440 2304
rect 12492 2292 12498 2304
rect 12713 2295 12771 2301
rect 12713 2292 12725 2295
rect 12492 2264 12725 2292
rect 12492 2252 12498 2264
rect 12713 2261 12725 2264
rect 12759 2261 12771 2295
rect 12713 2255 12771 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13596 2264 14289 2292
rect 13596 2252 13602 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 14366 2252 14372 2304
rect 14424 2292 14430 2304
rect 15013 2295 15071 2301
rect 15013 2292 15025 2295
rect 14424 2264 15025 2292
rect 14424 2252 14430 2264
rect 15013 2261 15025 2264
rect 15059 2261 15071 2295
rect 15013 2255 15071 2261
rect 15194 2252 15200 2304
rect 15252 2292 15258 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15252 2264 15669 2292
rect 15252 2252 15258 2264
rect 15657 2261 15669 2264
rect 15703 2261 15715 2295
rect 15657 2255 15715 2261
rect 15746 2252 15752 2304
rect 15804 2292 15810 2304
rect 16316 2301 16344 2332
rect 16390 2320 16396 2372
rect 16448 2360 16454 2372
rect 16448 2332 17172 2360
rect 16448 2320 16454 2332
rect 17144 2301 17172 2332
rect 16117 2295 16175 2301
rect 16117 2292 16129 2295
rect 15804 2264 16129 2292
rect 15804 2252 15810 2264
rect 16117 2261 16129 2264
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 16301 2295 16359 2301
rect 16301 2261 16313 2295
rect 16347 2261 16359 2295
rect 16301 2255 16359 2261
rect 17129 2295 17187 2301
rect 17129 2261 17141 2295
rect 17175 2261 17187 2295
rect 17328 2292 17356 2391
rect 17696 2360 17724 2391
rect 18414 2388 18420 2400
rect 18472 2428 18478 2440
rect 18892 2428 18920 2468
rect 20732 2440 20760 2468
rect 22186 2456 22192 2468
rect 22244 2456 22250 2508
rect 19058 2428 19064 2440
rect 18472 2400 18920 2428
rect 19019 2400 19064 2428
rect 18472 2388 18478 2400
rect 19058 2388 19064 2400
rect 19116 2388 19122 2440
rect 19242 2428 19248 2440
rect 19203 2400 19248 2428
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 20346 2428 20352 2440
rect 20307 2400 20352 2428
rect 20346 2388 20352 2400
rect 20404 2388 20410 2440
rect 20625 2431 20683 2437
rect 20625 2397 20637 2431
rect 20671 2397 20683 2431
rect 20625 2391 20683 2397
rect 20640 2360 20668 2391
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20993 2431 21051 2437
rect 20772 2400 20817 2428
rect 20772 2388 20778 2400
rect 20993 2397 21005 2431
rect 21039 2428 21051 2431
rect 22554 2428 22560 2440
rect 21039 2400 22560 2428
rect 21039 2397 21051 2400
rect 20993 2391 21051 2397
rect 22554 2388 22560 2400
rect 22612 2388 22618 2440
rect 21818 2360 21824 2372
rect 17696 2332 18920 2360
rect 20640 2332 21824 2360
rect 18690 2292 18696 2304
rect 17328 2264 18696 2292
rect 17129 2255 17187 2261
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 18892 2301 18920 2332
rect 21818 2320 21824 2332
rect 21876 2320 21882 2372
rect 18877 2295 18935 2301
rect 18877 2261 18889 2295
rect 18923 2261 18935 2295
rect 18877 2255 18935 2261
rect 18966 2252 18972 2304
rect 19024 2292 19030 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19024 2264 19441 2292
rect 19024 2252 19030 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
rect 5994 2048 6000 2100
rect 6052 2088 6058 2100
rect 11698 2088 11704 2100
rect 6052 2060 11704 2088
rect 6052 2048 6058 2060
rect 11698 2048 11704 2060
rect 11756 2048 11762 2100
rect 12434 2088 12440 2100
rect 12406 2048 12440 2088
rect 12492 2048 12498 2100
rect 16298 2048 16304 2100
rect 16356 2088 16362 2100
rect 19242 2088 19248 2100
rect 16356 2060 19248 2088
rect 16356 2048 16362 2060
rect 19242 2048 19248 2060
rect 19300 2048 19306 2100
rect 2406 1980 2412 2032
rect 2464 2020 2470 2032
rect 7098 2020 7104 2032
rect 2464 1992 7104 2020
rect 2464 1980 2470 1992
rect 7098 1980 7104 1992
rect 7156 2020 7162 2032
rect 8202 2020 8208 2032
rect 7156 1992 8208 2020
rect 7156 1980 7162 1992
rect 8202 1980 8208 1992
rect 8260 1980 8266 2032
rect 9214 1980 9220 2032
rect 9272 2020 9278 2032
rect 12406 2020 12434 2048
rect 9272 1992 12434 2020
rect 9272 1980 9278 1992
rect 17770 1980 17776 2032
rect 17828 2020 17834 2032
rect 20346 2020 20352 2032
rect 17828 1992 20352 2020
rect 17828 1980 17834 1992
rect 20346 1980 20352 1992
rect 20404 1980 20410 2032
rect 842 1912 848 1964
rect 900 1952 906 1964
rect 4798 1952 4804 1964
rect 900 1924 4804 1952
rect 900 1912 906 1924
rect 4798 1912 4804 1924
rect 4856 1912 4862 1964
rect 8294 1912 8300 1964
rect 8352 1952 8358 1964
rect 11882 1952 11888 1964
rect 8352 1924 11888 1952
rect 8352 1912 8358 1924
rect 11882 1912 11888 1924
rect 11940 1952 11946 1964
rect 12618 1952 12624 1964
rect 11940 1924 12624 1952
rect 11940 1912 11946 1924
rect 12618 1912 12624 1924
rect 12676 1912 12682 1964
rect 1946 1844 1952 1896
rect 2004 1884 2010 1896
rect 2004 1856 2774 1884
rect 2004 1844 2010 1856
rect 2746 1680 2774 1856
rect 5902 1844 5908 1896
rect 5960 1884 5966 1896
rect 10870 1884 10876 1896
rect 5960 1856 10876 1884
rect 5960 1844 5966 1856
rect 10870 1844 10876 1856
rect 10928 1844 10934 1896
rect 16114 1844 16120 1896
rect 16172 1884 16178 1896
rect 19242 1884 19248 1896
rect 16172 1856 19248 1884
rect 16172 1844 16178 1856
rect 19242 1844 19248 1856
rect 19300 1844 19306 1896
rect 21818 1844 21824 1896
rect 21876 1884 21882 1896
rect 22370 1884 22376 1896
rect 21876 1856 22376 1884
rect 21876 1844 21882 1856
rect 22370 1844 22376 1856
rect 22428 1844 22434 1896
rect 2866 1776 2872 1828
rect 2924 1816 2930 1828
rect 10686 1816 10692 1828
rect 2924 1788 10692 1816
rect 2924 1776 2930 1788
rect 10686 1776 10692 1788
rect 10744 1776 10750 1828
rect 15010 1776 15016 1828
rect 15068 1816 15074 1828
rect 19058 1816 19064 1828
rect 15068 1788 19064 1816
rect 15068 1776 15074 1788
rect 19058 1776 19064 1788
rect 19116 1776 19122 1828
rect 3970 1708 3976 1760
rect 4028 1748 4034 1760
rect 11054 1748 11060 1760
rect 4028 1720 11060 1748
rect 4028 1708 4034 1720
rect 11054 1708 11060 1720
rect 11112 1708 11118 1760
rect 9766 1680 9772 1692
rect 2746 1652 9772 1680
rect 9766 1640 9772 1652
rect 9824 1640 9830 1692
rect 10502 1640 10508 1692
rect 10560 1680 10566 1692
rect 11974 1680 11980 1692
rect 10560 1652 11980 1680
rect 10560 1640 10566 1652
rect 11974 1640 11980 1652
rect 12032 1640 12038 1692
rect 17218 1436 17224 1488
rect 17276 1476 17282 1488
rect 18138 1476 18144 1488
rect 17276 1448 18144 1476
rect 17276 1436 17282 1448
rect 18138 1436 18144 1448
rect 18196 1436 18202 1488
rect 17678 1368 17684 1420
rect 17736 1408 17742 1420
rect 18966 1408 18972 1420
rect 17736 1380 18972 1408
rect 17736 1368 17742 1380
rect 18966 1368 18972 1380
rect 19024 1368 19030 1420
rect 22002 1368 22008 1420
rect 22060 1408 22066 1420
rect 22738 1408 22744 1420
rect 22060 1380 22744 1408
rect 22060 1368 22066 1380
rect 22738 1368 22744 1380
rect 22796 1368 22802 1420
rect 3234 1300 3240 1352
rect 3292 1340 3298 1352
rect 10318 1340 10324 1352
rect 3292 1312 10324 1340
rect 3292 1300 3298 1312
rect 10318 1300 10324 1312
rect 10376 1300 10382 1352
rect 17126 1300 17132 1352
rect 17184 1340 17190 1352
rect 18690 1340 18696 1352
rect 17184 1312 18696 1340
rect 17184 1300 17190 1312
rect 18690 1300 18696 1312
rect 18748 1300 18754 1352
rect 3510 1232 3516 1284
rect 3568 1272 3574 1284
rect 5718 1272 5724 1284
rect 3568 1244 5724 1272
rect 3568 1232 3574 1244
rect 5718 1232 5724 1244
rect 5776 1272 5782 1284
rect 13170 1272 13176 1284
rect 5776 1244 13176 1272
rect 5776 1232 5782 1244
rect 13170 1232 13176 1244
rect 13228 1232 13234 1284
rect 18506 1232 18512 1284
rect 18564 1272 18570 1284
rect 20254 1272 20260 1284
rect 18564 1244 20260 1272
rect 18564 1232 18570 1244
rect 20254 1232 20260 1244
rect 20312 1232 20318 1284
rect 3234 1164 3240 1216
rect 3292 1204 3298 1216
rect 4522 1204 4528 1216
rect 3292 1176 4528 1204
rect 3292 1164 3298 1176
rect 4522 1164 4528 1176
rect 4580 1164 4586 1216
rect 1026 1028 1032 1080
rect 1084 1068 1090 1080
rect 12802 1068 12808 1080
rect 1084 1040 12808 1068
rect 1084 1028 1090 1040
rect 12802 1028 12808 1040
rect 12860 1028 12866 1080
rect 7834 960 7840 1012
rect 7892 1000 7898 1012
rect 17954 1000 17960 1012
rect 7892 972 17960 1000
rect 7892 960 7898 972
rect 17954 960 17960 972
rect 18012 960 18018 1012
rect 6638 892 6644 944
rect 6696 932 6702 944
rect 14642 932 14648 944
rect 6696 904 14648 932
rect 6696 892 6702 904
rect 14642 892 14648 904
rect 14700 932 14706 944
rect 21358 932 21364 944
rect 14700 904 21364 932
rect 14700 892 14706 904
rect 21358 892 21364 904
rect 21416 892 21422 944
<< via1 >>
rect 848 22040 900 22092
rect 1032 22040 1084 22092
rect 20 21632 72 21684
rect 14280 21632 14332 21684
rect 7564 21564 7616 21616
rect 16212 21564 16264 21616
rect 1400 21496 1452 21548
rect 2504 21496 2556 21548
rect 4712 21496 4764 21548
rect 15660 21496 15712 21548
rect 2596 21428 2648 21480
rect 16120 21428 16172 21480
rect 4804 21360 4856 21412
rect 5080 21360 5132 21412
rect 12900 21360 12952 21412
rect 2780 21292 2832 21344
rect 17868 21292 17920 21344
rect 4068 21224 4120 21276
rect 12164 21224 12216 21276
rect 3608 21156 3660 21208
rect 13268 21156 13320 21208
rect 4436 21088 4488 21140
rect 16028 21088 16080 21140
rect 2688 21020 2740 21072
rect 7564 21020 7616 21072
rect 3332 20952 3384 21004
rect 13084 21020 13136 21072
rect 3148 20884 3200 20936
rect 11980 20884 12032 20936
rect 12164 20884 12216 20936
rect 14924 20884 14976 20936
rect 8208 20816 8260 20868
rect 12992 20816 13044 20868
rect 940 20748 992 20800
rect 3056 20748 3108 20800
rect 4252 20748 4304 20800
rect 10692 20748 10744 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 5172 20544 5224 20596
rect 6920 20544 6972 20596
rect 7380 20544 7432 20596
rect 8208 20544 8260 20596
rect 8668 20544 8720 20596
rect 9312 20544 9364 20596
rect 6000 20476 6052 20528
rect 1308 20408 1360 20460
rect 3332 20451 3384 20460
rect 3332 20417 3341 20451
rect 3341 20417 3375 20451
rect 3375 20417 3384 20451
rect 3332 20408 3384 20417
rect 3608 20451 3660 20460
rect 3608 20417 3617 20451
rect 3617 20417 3651 20451
rect 3651 20417 3660 20451
rect 3608 20408 3660 20417
rect 1952 20383 2004 20392
rect 1952 20349 1961 20383
rect 1961 20349 1995 20383
rect 1995 20349 2004 20383
rect 1952 20340 2004 20349
rect 4620 20340 4672 20392
rect 4988 20383 5040 20392
rect 4988 20349 4997 20383
rect 4997 20349 5031 20383
rect 5031 20349 5040 20383
rect 4988 20340 5040 20349
rect 4344 20272 4396 20324
rect 5632 20408 5684 20460
rect 5540 20383 5592 20392
rect 5540 20349 5549 20383
rect 5549 20349 5583 20383
rect 5583 20349 5592 20383
rect 5540 20340 5592 20349
rect 3884 20204 3936 20256
rect 4896 20204 4948 20256
rect 5816 20272 5868 20324
rect 9496 20476 9548 20528
rect 6828 20408 6880 20460
rect 7472 20408 7524 20460
rect 6920 20340 6972 20392
rect 7840 20408 7892 20460
rect 8208 20451 8260 20460
rect 8208 20417 8217 20451
rect 8217 20417 8251 20451
rect 8251 20417 8260 20451
rect 8208 20408 8260 20417
rect 8484 20408 8536 20460
rect 8944 20408 8996 20460
rect 9680 20408 9732 20460
rect 10876 20544 10928 20596
rect 6736 20272 6788 20324
rect 8024 20340 8076 20392
rect 9128 20340 9180 20392
rect 10508 20451 10560 20460
rect 10508 20417 10517 20451
rect 10517 20417 10551 20451
rect 10551 20417 10560 20451
rect 10508 20408 10560 20417
rect 10692 20408 10744 20460
rect 11796 20544 11848 20596
rect 12072 20544 12124 20596
rect 12440 20544 12492 20596
rect 12808 20544 12860 20596
rect 13176 20544 13228 20596
rect 13544 20544 13596 20596
rect 14004 20544 14056 20596
rect 14372 20544 14424 20596
rect 14740 20544 14792 20596
rect 15200 20544 15252 20596
rect 15476 20544 15528 20596
rect 15844 20544 15896 20596
rect 17960 20544 18012 20596
rect 18144 20544 18196 20596
rect 19524 20544 19576 20596
rect 19800 20544 19852 20596
rect 19984 20544 20036 20596
rect 20536 20587 20588 20596
rect 11888 20408 11940 20460
rect 10784 20383 10836 20392
rect 10784 20349 10793 20383
rect 10793 20349 10827 20383
rect 10827 20349 10836 20383
rect 10784 20340 10836 20349
rect 10876 20340 10928 20392
rect 12808 20408 12860 20460
rect 13176 20408 13228 20460
rect 13728 20408 13780 20460
rect 14464 20451 14516 20460
rect 13452 20340 13504 20392
rect 14464 20417 14473 20451
rect 14473 20417 14507 20451
rect 14507 20417 14516 20451
rect 14464 20408 14516 20417
rect 14648 20408 14700 20460
rect 15016 20408 15068 20460
rect 15568 20451 15620 20460
rect 15568 20417 15577 20451
rect 15577 20417 15611 20451
rect 15611 20417 15620 20451
rect 15568 20408 15620 20417
rect 15936 20451 15988 20460
rect 15936 20417 15945 20451
rect 15945 20417 15979 20451
rect 15979 20417 15988 20451
rect 15936 20408 15988 20417
rect 16672 20451 16724 20460
rect 16672 20417 16681 20451
rect 16681 20417 16715 20451
rect 16715 20417 16724 20451
rect 16672 20408 16724 20417
rect 17500 20476 17552 20528
rect 18972 20476 19024 20528
rect 17132 20408 17184 20460
rect 19524 20408 19576 20460
rect 20536 20553 20545 20587
rect 20545 20553 20579 20587
rect 20579 20553 20588 20587
rect 20536 20544 20588 20553
rect 20904 20544 20956 20596
rect 21640 20476 21692 20528
rect 19432 20340 19484 20392
rect 5356 20204 5408 20256
rect 6460 20204 6512 20256
rect 6828 20204 6880 20256
rect 7012 20204 7064 20256
rect 7380 20204 7432 20256
rect 12624 20272 12676 20324
rect 16580 20272 16632 20324
rect 18604 20272 18656 20324
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 9404 20204 9456 20256
rect 10508 20204 10560 20256
rect 10692 20204 10744 20256
rect 12256 20204 12308 20256
rect 16028 20204 16080 20256
rect 16396 20204 16448 20256
rect 17224 20247 17276 20256
rect 17224 20213 17233 20247
rect 17233 20213 17267 20247
rect 17267 20213 17276 20247
rect 17224 20204 17276 20213
rect 19616 20204 19668 20256
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 20168 20272 20220 20324
rect 21364 20408 21416 20460
rect 20996 20272 21048 20324
rect 21088 20204 21140 20256
rect 21456 20247 21508 20256
rect 21456 20213 21465 20247
rect 21465 20213 21499 20247
rect 21499 20213 21508 20247
rect 21456 20204 21508 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 1584 20000 1636 20052
rect 2688 19975 2740 19984
rect 2688 19941 2697 19975
rect 2697 19941 2731 19975
rect 2731 19941 2740 19975
rect 2688 19932 2740 19941
rect 3608 19932 3660 19984
rect 3792 19932 3844 19984
rect 3976 19932 4028 19984
rect 1492 19796 1544 19848
rect 2044 19839 2096 19848
rect 2044 19805 2053 19839
rect 2053 19805 2087 19839
rect 2087 19805 2096 19839
rect 2044 19796 2096 19805
rect 4068 19864 4120 19916
rect 3240 19796 3292 19848
rect 3700 19796 3752 19848
rect 5540 19864 5592 19916
rect 6828 19907 6880 19916
rect 5448 19796 5500 19848
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 1676 19660 1728 19712
rect 5540 19728 5592 19780
rect 3332 19660 3384 19712
rect 3792 19660 3844 19712
rect 4896 19660 4948 19712
rect 6828 19873 6837 19907
rect 6837 19873 6871 19907
rect 6871 19873 6880 19907
rect 6828 19864 6880 19873
rect 6736 19796 6788 19848
rect 7564 20000 7616 20052
rect 7104 19932 7156 19984
rect 8300 19907 8352 19916
rect 7104 19796 7156 19848
rect 6828 19728 6880 19780
rect 8300 19873 8309 19907
rect 8309 19873 8343 19907
rect 8343 19873 8352 19907
rect 8300 19864 8352 19873
rect 7748 19796 7800 19848
rect 7932 19728 7984 19780
rect 10692 20000 10744 20052
rect 10876 20043 10928 20052
rect 10876 20009 10885 20043
rect 10885 20009 10919 20043
rect 10919 20009 10928 20043
rect 10876 20000 10928 20009
rect 11888 20000 11940 20052
rect 12440 20043 12492 20052
rect 12440 20009 12449 20043
rect 12449 20009 12483 20043
rect 12483 20009 12492 20043
rect 12808 20043 12860 20052
rect 12440 20000 12492 20009
rect 12808 20009 12817 20043
rect 12817 20009 12851 20043
rect 12851 20009 12860 20043
rect 12808 20000 12860 20009
rect 13176 20043 13228 20052
rect 13176 20009 13185 20043
rect 13185 20009 13219 20043
rect 13219 20009 13228 20043
rect 13176 20000 13228 20009
rect 13452 20043 13504 20052
rect 13452 20009 13461 20043
rect 13461 20009 13495 20043
rect 13495 20009 13504 20043
rect 13452 20000 13504 20009
rect 13728 20043 13780 20052
rect 13728 20009 13737 20043
rect 13737 20009 13771 20043
rect 13771 20009 13780 20043
rect 13728 20000 13780 20009
rect 14648 20043 14700 20052
rect 14648 20009 14657 20043
rect 14657 20009 14691 20043
rect 14691 20009 14700 20043
rect 14648 20000 14700 20009
rect 15016 20043 15068 20052
rect 15016 20009 15025 20043
rect 15025 20009 15059 20043
rect 15059 20009 15068 20043
rect 15016 20000 15068 20009
rect 15936 20000 15988 20052
rect 16120 20043 16172 20052
rect 16120 20009 16129 20043
rect 16129 20009 16163 20043
rect 16163 20009 16172 20043
rect 16120 20000 16172 20009
rect 17040 20000 17092 20052
rect 17776 20000 17828 20052
rect 11244 19932 11296 19984
rect 12348 19932 12400 19984
rect 15844 19932 15896 19984
rect 16948 19932 17000 19984
rect 17408 19932 17460 19984
rect 8760 19796 8812 19848
rect 9588 19796 9640 19848
rect 9128 19771 9180 19780
rect 6920 19703 6972 19712
rect 6920 19669 6929 19703
rect 6929 19669 6963 19703
rect 6963 19669 6972 19703
rect 6920 19660 6972 19669
rect 7288 19703 7340 19712
rect 7288 19669 7297 19703
rect 7297 19669 7331 19703
rect 7331 19669 7340 19703
rect 7288 19660 7340 19669
rect 8116 19703 8168 19712
rect 8116 19669 8125 19703
rect 8125 19669 8159 19703
rect 8159 19669 8168 19703
rect 8116 19660 8168 19669
rect 9128 19737 9137 19771
rect 9137 19737 9171 19771
rect 9171 19737 9180 19771
rect 9128 19728 9180 19737
rect 9404 19728 9456 19780
rect 9772 19728 9824 19780
rect 10140 19728 10192 19780
rect 11704 19864 11756 19916
rect 10968 19839 11020 19848
rect 10968 19805 10977 19839
rect 10977 19805 11011 19839
rect 11011 19805 11020 19839
rect 10968 19796 11020 19805
rect 11060 19796 11112 19848
rect 9220 19660 9272 19712
rect 9956 19703 10008 19712
rect 9956 19669 9965 19703
rect 9965 19669 9999 19703
rect 9999 19669 10008 19703
rect 9956 19660 10008 19669
rect 10324 19703 10376 19712
rect 10324 19669 10333 19703
rect 10333 19669 10367 19703
rect 10367 19669 10376 19703
rect 10324 19660 10376 19669
rect 11244 19728 11296 19780
rect 12440 19796 12492 19848
rect 13360 19864 13412 19916
rect 18696 20000 18748 20052
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 13176 19796 13228 19848
rect 14832 19839 14884 19848
rect 11888 19728 11940 19780
rect 12164 19660 12216 19712
rect 12348 19728 12400 19780
rect 14832 19805 14841 19839
rect 14841 19805 14875 19839
rect 14875 19805 14884 19839
rect 14832 19796 14884 19805
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 15936 19796 15988 19848
rect 16396 19796 16448 19848
rect 14556 19728 14608 19780
rect 16672 19796 16724 19848
rect 16948 19796 17000 19848
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 17592 19796 17644 19848
rect 18788 19932 18840 19984
rect 20352 20000 20404 20052
rect 20536 20043 20588 20052
rect 20536 20009 20545 20043
rect 20545 20009 20579 20043
rect 20579 20009 20588 20043
rect 20536 20000 20588 20009
rect 19064 19932 19116 19984
rect 19616 19864 19668 19916
rect 20536 19864 20588 19916
rect 20812 19864 20864 19916
rect 18880 19796 18932 19848
rect 20352 19839 20404 19848
rect 20352 19805 20383 19839
rect 20383 19805 20404 19839
rect 18604 19728 18656 19780
rect 19432 19771 19484 19780
rect 19432 19737 19441 19771
rect 19441 19737 19475 19771
rect 19475 19737 19484 19771
rect 19432 19728 19484 19737
rect 20352 19796 20404 19805
rect 20720 19839 20772 19848
rect 20720 19805 20729 19839
rect 20729 19805 20763 19839
rect 20763 19805 20772 19839
rect 20720 19796 20772 19805
rect 21272 19839 21324 19848
rect 21272 19805 21281 19839
rect 21281 19805 21315 19839
rect 21315 19805 21324 19839
rect 21272 19796 21324 19805
rect 17132 19660 17184 19712
rect 18512 19660 18564 19712
rect 19616 19660 19668 19712
rect 22008 19728 22060 19780
rect 21548 19660 21600 19712
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 2596 19456 2648 19508
rect 2872 19388 2924 19440
rect 1952 19320 2004 19372
rect 2044 19363 2096 19372
rect 2044 19329 2053 19363
rect 2053 19329 2087 19363
rect 2087 19329 2096 19363
rect 2044 19320 2096 19329
rect 2320 19320 2372 19372
rect 2504 19320 2556 19372
rect 1860 19227 1912 19236
rect 1860 19193 1869 19227
rect 1869 19193 1903 19227
rect 1903 19193 1912 19227
rect 1860 19184 1912 19193
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3240 19320 3292 19372
rect 2872 19252 2924 19304
rect 3516 19252 3568 19304
rect 3976 19388 4028 19440
rect 4896 19388 4948 19440
rect 5632 19456 5684 19508
rect 5908 19388 5960 19440
rect 3700 19320 3752 19372
rect 2964 19184 3016 19236
rect 4068 19252 4120 19304
rect 5448 19320 5500 19372
rect 7012 19388 7064 19440
rect 7288 19456 7340 19508
rect 9312 19499 9364 19508
rect 9312 19465 9321 19499
rect 9321 19465 9355 19499
rect 9355 19465 9364 19499
rect 9312 19456 9364 19465
rect 9588 19499 9640 19508
rect 9588 19465 9597 19499
rect 9597 19465 9631 19499
rect 9631 19465 9640 19499
rect 9588 19456 9640 19465
rect 9864 19456 9916 19508
rect 11060 19456 11112 19508
rect 11244 19499 11296 19508
rect 11244 19465 11253 19499
rect 11253 19465 11287 19499
rect 11287 19465 11296 19499
rect 11244 19456 11296 19465
rect 11704 19456 11756 19508
rect 12440 19456 12492 19508
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 6460 19320 6512 19372
rect 6644 19363 6696 19372
rect 6644 19329 6653 19363
rect 6653 19329 6687 19363
rect 6687 19329 6696 19363
rect 6644 19320 6696 19329
rect 8300 19320 8352 19372
rect 8576 19320 8628 19372
rect 9128 19363 9180 19372
rect 9128 19329 9137 19363
rect 9137 19329 9171 19363
rect 9171 19329 9180 19363
rect 9128 19320 9180 19329
rect 10140 19388 10192 19440
rect 10784 19431 10836 19440
rect 10784 19397 10793 19431
rect 10793 19397 10827 19431
rect 10827 19397 10836 19431
rect 10784 19388 10836 19397
rect 11152 19388 11204 19440
rect 11888 19388 11940 19440
rect 12256 19388 12308 19440
rect 17316 19456 17368 19508
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 17868 19456 17920 19508
rect 18512 19499 18564 19508
rect 5908 19295 5960 19304
rect 4160 19184 4212 19236
rect 5908 19261 5917 19295
rect 5917 19261 5951 19295
rect 5951 19261 5960 19295
rect 5908 19252 5960 19261
rect 6092 19295 6144 19304
rect 6092 19261 6101 19295
rect 6101 19261 6135 19295
rect 6135 19261 6144 19295
rect 6092 19252 6144 19261
rect 6736 19252 6788 19304
rect 7012 19252 7064 19304
rect 10232 19320 10284 19372
rect 10876 19363 10928 19372
rect 10876 19329 10885 19363
rect 10885 19329 10919 19363
rect 10919 19329 10928 19363
rect 10876 19320 10928 19329
rect 6368 19184 6420 19236
rect 8300 19184 8352 19236
rect 9496 19252 9548 19304
rect 12164 19320 12216 19372
rect 13636 19320 13688 19372
rect 18144 19388 18196 19440
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 18788 19499 18840 19508
rect 18788 19465 18797 19499
rect 18797 19465 18831 19499
rect 18831 19465 18840 19499
rect 18788 19456 18840 19465
rect 19156 19499 19208 19508
rect 19156 19465 19165 19499
rect 19165 19465 19199 19499
rect 19199 19465 19208 19499
rect 19156 19456 19208 19465
rect 19248 19456 19300 19508
rect 11520 19295 11572 19304
rect 10324 19184 10376 19236
rect 11520 19261 11529 19295
rect 11529 19261 11563 19295
rect 11563 19261 11572 19295
rect 11520 19252 11572 19261
rect 12532 19252 12584 19304
rect 17960 19363 18012 19372
rect 14740 19295 14792 19304
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 15292 19295 15344 19304
rect 15292 19261 15301 19295
rect 15301 19261 15335 19295
rect 15335 19261 15344 19295
rect 15292 19252 15344 19261
rect 16304 19252 16356 19304
rect 13544 19184 13596 19236
rect 13728 19184 13780 19236
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 3976 19159 4028 19168
rect 3976 19125 3985 19159
rect 3985 19125 4019 19159
rect 4019 19125 4028 19159
rect 3976 19116 4028 19125
rect 6552 19159 6604 19168
rect 6552 19125 6561 19159
rect 6561 19125 6595 19159
rect 6595 19125 6604 19159
rect 6828 19159 6880 19168
rect 6552 19116 6604 19125
rect 6828 19125 6837 19159
rect 6837 19125 6871 19159
rect 6871 19125 6880 19159
rect 6828 19116 6880 19125
rect 6920 19116 6972 19168
rect 7932 19116 7984 19168
rect 8024 19116 8076 19168
rect 8208 19116 8260 19168
rect 8484 19116 8536 19168
rect 12256 19116 12308 19168
rect 12440 19116 12492 19168
rect 12624 19116 12676 19168
rect 13360 19159 13412 19168
rect 13360 19125 13369 19159
rect 13369 19125 13403 19159
rect 13403 19125 13412 19159
rect 13360 19116 13412 19125
rect 13452 19159 13504 19168
rect 13452 19125 13461 19159
rect 13461 19125 13495 19159
rect 13495 19125 13504 19159
rect 13820 19159 13872 19168
rect 13452 19116 13504 19125
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 14372 19159 14424 19168
rect 14372 19125 14381 19159
rect 14381 19125 14415 19159
rect 14415 19125 14424 19159
rect 14372 19116 14424 19125
rect 15016 19159 15068 19168
rect 15016 19125 15025 19159
rect 15025 19125 15059 19159
rect 15059 19125 15068 19159
rect 15016 19116 15068 19125
rect 15292 19116 15344 19168
rect 15936 19184 15988 19236
rect 17960 19329 17969 19363
rect 17969 19329 18003 19363
rect 18003 19329 18012 19363
rect 17960 19320 18012 19329
rect 18236 19320 18288 19372
rect 17592 19252 17644 19304
rect 18420 19320 18472 19372
rect 18972 19320 19024 19372
rect 20904 19388 20956 19440
rect 19524 19320 19576 19372
rect 19616 19320 19668 19372
rect 19800 19295 19852 19304
rect 17316 19184 17368 19236
rect 19340 19184 19392 19236
rect 19800 19261 19809 19295
rect 19809 19261 19843 19295
rect 19843 19261 19852 19295
rect 19800 19252 19852 19261
rect 20352 19184 20404 19236
rect 15752 19159 15804 19168
rect 15752 19125 15761 19159
rect 15761 19125 15795 19159
rect 15795 19125 15804 19159
rect 15752 19116 15804 19125
rect 16396 19159 16448 19168
rect 16396 19125 16405 19159
rect 16405 19125 16439 19159
rect 16439 19125 16448 19159
rect 16396 19116 16448 19125
rect 17040 19116 17092 19168
rect 18788 19116 18840 19168
rect 21180 19116 21232 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1768 18912 1820 18964
rect 2228 18955 2280 18964
rect 2228 18921 2237 18955
rect 2237 18921 2271 18955
rect 2271 18921 2280 18955
rect 2228 18912 2280 18921
rect 2412 18912 2464 18964
rect 848 18844 900 18896
rect 1124 18844 1176 18896
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 2320 18708 2372 18760
rect 2688 18708 2740 18760
rect 3424 18912 3476 18964
rect 4252 18912 4304 18964
rect 6092 18912 6144 18964
rect 3700 18844 3752 18896
rect 5356 18844 5408 18896
rect 6736 18912 6788 18964
rect 7288 18912 7340 18964
rect 7472 18955 7524 18964
rect 7472 18921 7481 18955
rect 7481 18921 7515 18955
rect 7515 18921 7524 18955
rect 7472 18912 7524 18921
rect 4528 18776 4580 18828
rect 4896 18819 4948 18828
rect 4896 18785 4905 18819
rect 4905 18785 4939 18819
rect 4939 18785 4948 18819
rect 4896 18776 4948 18785
rect 8116 18912 8168 18964
rect 8484 18955 8536 18964
rect 8484 18921 8493 18955
rect 8493 18921 8527 18955
rect 8527 18921 8536 18955
rect 8484 18912 8536 18921
rect 8668 18912 8720 18964
rect 9864 18912 9916 18964
rect 10232 18912 10284 18964
rect 10508 18912 10560 18964
rect 13820 18912 13872 18964
rect 14464 18912 14516 18964
rect 15568 18912 15620 18964
rect 17408 18912 17460 18964
rect 17500 18955 17552 18964
rect 17500 18921 17509 18955
rect 17509 18921 17543 18955
rect 17543 18921 17552 18955
rect 17500 18912 17552 18921
rect 18052 18912 18104 18964
rect 18236 18955 18288 18964
rect 18236 18921 18245 18955
rect 18245 18921 18279 18955
rect 18279 18921 18288 18955
rect 18236 18912 18288 18921
rect 19064 18955 19116 18964
rect 19064 18921 19073 18955
rect 19073 18921 19107 18955
rect 19107 18921 19116 18955
rect 19064 18912 19116 18921
rect 19984 18912 20036 18964
rect 20444 18912 20496 18964
rect 3700 18708 3752 18760
rect 3884 18708 3936 18760
rect 3976 18708 4028 18760
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 3608 18615 3660 18624
rect 3608 18581 3617 18615
rect 3617 18581 3651 18615
rect 3651 18581 3660 18615
rect 3608 18572 3660 18581
rect 4160 18615 4212 18624
rect 4160 18581 4169 18615
rect 4169 18581 4203 18615
rect 4203 18581 4212 18615
rect 4160 18572 4212 18581
rect 6460 18708 6512 18760
rect 7380 18708 7432 18760
rect 8024 18708 8076 18760
rect 5448 18683 5500 18692
rect 5448 18649 5457 18683
rect 5457 18649 5491 18683
rect 5491 18649 5500 18683
rect 5448 18640 5500 18649
rect 5724 18640 5776 18692
rect 6184 18640 6236 18692
rect 6736 18640 6788 18692
rect 6828 18683 6880 18692
rect 6828 18649 6846 18683
rect 6846 18649 6880 18683
rect 8392 18844 8444 18896
rect 8392 18708 8444 18760
rect 9128 18887 9180 18896
rect 9128 18853 9137 18887
rect 9137 18853 9171 18887
rect 9171 18853 9180 18887
rect 9128 18844 9180 18853
rect 12992 18844 13044 18896
rect 13728 18844 13780 18896
rect 15292 18844 15344 18896
rect 17316 18844 17368 18896
rect 17960 18887 18012 18896
rect 17960 18853 17969 18887
rect 17969 18853 18003 18887
rect 18003 18853 18012 18887
rect 17960 18844 18012 18853
rect 18880 18844 18932 18896
rect 19708 18887 19760 18896
rect 19708 18853 19717 18887
rect 19717 18853 19751 18887
rect 19751 18853 19760 18887
rect 19708 18844 19760 18853
rect 19892 18844 19944 18896
rect 22744 18844 22796 18896
rect 12808 18776 12860 18828
rect 13176 18776 13228 18828
rect 9496 18708 9548 18760
rect 9772 18708 9824 18760
rect 10324 18708 10376 18760
rect 11612 18708 11664 18760
rect 12532 18708 12584 18760
rect 6828 18640 6880 18649
rect 10968 18640 11020 18692
rect 14556 18751 14608 18760
rect 4804 18572 4856 18624
rect 5816 18572 5868 18624
rect 7840 18615 7892 18624
rect 7840 18581 7849 18615
rect 7849 18581 7883 18615
rect 7883 18581 7892 18615
rect 7840 18572 7892 18581
rect 8024 18572 8076 18624
rect 8116 18572 8168 18624
rect 10140 18572 10192 18624
rect 10692 18572 10744 18624
rect 11244 18615 11296 18624
rect 11244 18581 11253 18615
rect 11253 18581 11287 18615
rect 11287 18581 11296 18615
rect 11244 18572 11296 18581
rect 12440 18572 12492 18624
rect 13820 18683 13872 18692
rect 13820 18649 13829 18683
rect 13829 18649 13863 18683
rect 13863 18649 13872 18683
rect 13820 18640 13872 18649
rect 14556 18717 14565 18751
rect 14565 18717 14599 18751
rect 14599 18717 14608 18751
rect 14556 18708 14608 18717
rect 15936 18708 15988 18760
rect 17224 18708 17276 18760
rect 20444 18776 20496 18828
rect 18236 18708 18288 18760
rect 18788 18751 18840 18760
rect 18788 18717 18797 18751
rect 18797 18717 18831 18751
rect 18831 18717 18840 18751
rect 18788 18708 18840 18717
rect 18880 18751 18932 18760
rect 18880 18717 18889 18751
rect 18889 18717 18923 18751
rect 18923 18717 18932 18751
rect 18880 18708 18932 18717
rect 19064 18708 19116 18760
rect 19892 18751 19944 18760
rect 19892 18717 19901 18751
rect 19901 18717 19935 18751
rect 19935 18717 19944 18751
rect 19892 18708 19944 18717
rect 20352 18751 20404 18760
rect 20352 18717 20361 18751
rect 20361 18717 20395 18751
rect 20395 18717 20404 18751
rect 20720 18751 20772 18760
rect 20352 18708 20404 18717
rect 20720 18717 20729 18751
rect 20729 18717 20763 18751
rect 20763 18717 20772 18751
rect 20720 18708 20772 18717
rect 20812 18640 20864 18692
rect 20996 18683 21048 18692
rect 20996 18649 21005 18683
rect 21005 18649 21039 18683
rect 21039 18649 21048 18683
rect 20996 18640 21048 18649
rect 13176 18615 13228 18624
rect 13176 18581 13185 18615
rect 13185 18581 13219 18615
rect 13219 18581 13228 18615
rect 13176 18572 13228 18581
rect 17408 18615 17460 18624
rect 17408 18581 17417 18615
rect 17417 18581 17451 18615
rect 17451 18581 17460 18615
rect 17408 18572 17460 18581
rect 18328 18572 18380 18624
rect 18696 18572 18748 18624
rect 21456 18615 21508 18624
rect 21456 18581 21465 18615
rect 21465 18581 21499 18615
rect 21499 18581 21508 18615
rect 21456 18572 21508 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 2596 18368 2648 18420
rect 3608 18411 3660 18420
rect 3608 18377 3617 18411
rect 3617 18377 3651 18411
rect 3651 18377 3660 18411
rect 3608 18368 3660 18377
rect 2872 18300 2924 18352
rect 4068 18368 4120 18420
rect 5816 18411 5868 18420
rect 4436 18343 4488 18352
rect 4436 18309 4445 18343
rect 4445 18309 4479 18343
rect 4479 18309 4488 18343
rect 4436 18300 4488 18309
rect 4712 18300 4764 18352
rect 5080 18343 5132 18352
rect 5080 18309 5089 18343
rect 5089 18309 5123 18343
rect 5123 18309 5132 18343
rect 5080 18300 5132 18309
rect 5816 18377 5825 18411
rect 5825 18377 5859 18411
rect 5859 18377 5868 18411
rect 5816 18368 5868 18377
rect 5908 18368 5960 18420
rect 7196 18411 7248 18420
rect 6920 18300 6972 18352
rect 7196 18377 7205 18411
rect 7205 18377 7239 18411
rect 7239 18377 7248 18411
rect 7196 18368 7248 18377
rect 7288 18368 7340 18420
rect 7656 18368 7708 18420
rect 7932 18368 7984 18420
rect 1676 18275 1728 18284
rect 1676 18241 1685 18275
rect 1685 18241 1719 18275
rect 1719 18241 1728 18275
rect 1676 18232 1728 18241
rect 4068 18232 4120 18284
rect 2504 18164 2556 18216
rect 572 18096 624 18148
rect 5448 18232 5500 18284
rect 4804 18164 4856 18216
rect 4896 18164 4948 18216
rect 5172 18164 5224 18216
rect 5264 18164 5316 18216
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 1860 18071 1912 18080
rect 1860 18037 1869 18071
rect 1869 18037 1903 18071
rect 1903 18037 1912 18071
rect 1860 18028 1912 18037
rect 2136 18071 2188 18080
rect 2136 18037 2145 18071
rect 2145 18037 2179 18071
rect 2179 18037 2188 18071
rect 2136 18028 2188 18037
rect 2320 18071 2372 18080
rect 2320 18037 2329 18071
rect 2329 18037 2363 18071
rect 2363 18037 2372 18071
rect 2320 18028 2372 18037
rect 2780 18028 2832 18080
rect 4712 18096 4764 18148
rect 5724 18207 5776 18216
rect 5724 18173 5733 18207
rect 5733 18173 5767 18207
rect 5767 18173 5776 18207
rect 6736 18275 6788 18284
rect 6736 18241 6745 18275
rect 6745 18241 6779 18275
rect 6779 18241 6788 18275
rect 6736 18232 6788 18241
rect 7012 18232 7064 18284
rect 7472 18232 7524 18284
rect 5724 18164 5776 18173
rect 6000 18096 6052 18148
rect 6828 18164 6880 18216
rect 7656 18207 7708 18216
rect 7656 18173 7665 18207
rect 7665 18173 7699 18207
rect 7699 18173 7708 18207
rect 7656 18164 7708 18173
rect 7748 18164 7800 18216
rect 8300 18300 8352 18352
rect 8116 18232 8168 18284
rect 8760 18300 8812 18352
rect 9036 18300 9088 18352
rect 9956 18368 10008 18420
rect 10508 18368 10560 18420
rect 10876 18368 10928 18420
rect 10968 18411 11020 18420
rect 10968 18377 10977 18411
rect 10977 18377 11011 18411
rect 11011 18377 11020 18411
rect 10968 18368 11020 18377
rect 12440 18368 12492 18420
rect 12716 18411 12768 18420
rect 12716 18377 12725 18411
rect 12725 18377 12759 18411
rect 12759 18377 12768 18411
rect 12716 18368 12768 18377
rect 12900 18411 12952 18420
rect 12900 18377 12909 18411
rect 12909 18377 12943 18411
rect 12943 18377 12952 18411
rect 12900 18368 12952 18377
rect 13268 18411 13320 18420
rect 13268 18377 13277 18411
rect 13277 18377 13311 18411
rect 13311 18377 13320 18411
rect 13268 18368 13320 18377
rect 13544 18368 13596 18420
rect 14556 18368 14608 18420
rect 14648 18411 14700 18420
rect 14648 18377 14657 18411
rect 14657 18377 14691 18411
rect 14691 18377 14700 18411
rect 14924 18411 14976 18420
rect 14648 18368 14700 18377
rect 14924 18377 14933 18411
rect 14933 18377 14967 18411
rect 14967 18377 14976 18411
rect 14924 18368 14976 18377
rect 15200 18411 15252 18420
rect 15200 18377 15209 18411
rect 15209 18377 15243 18411
rect 15243 18377 15252 18411
rect 15200 18368 15252 18377
rect 15292 18411 15344 18420
rect 15292 18377 15301 18411
rect 15301 18377 15335 18411
rect 15335 18377 15344 18411
rect 15936 18411 15988 18420
rect 15292 18368 15344 18377
rect 15936 18377 15945 18411
rect 15945 18377 15979 18411
rect 15979 18377 15988 18411
rect 15936 18368 15988 18377
rect 16396 18368 16448 18420
rect 17592 18368 17644 18420
rect 18236 18411 18288 18420
rect 18236 18377 18245 18411
rect 18245 18377 18279 18411
rect 18279 18377 18288 18411
rect 18236 18368 18288 18377
rect 18512 18411 18564 18420
rect 18512 18377 18521 18411
rect 18521 18377 18555 18411
rect 18555 18377 18564 18411
rect 18512 18368 18564 18377
rect 19524 18368 19576 18420
rect 20720 18368 20772 18420
rect 11428 18300 11480 18352
rect 12532 18343 12584 18352
rect 12532 18309 12541 18343
rect 12541 18309 12575 18343
rect 12575 18309 12584 18343
rect 12532 18300 12584 18309
rect 8300 18207 8352 18216
rect 8300 18173 8309 18207
rect 8309 18173 8343 18207
rect 8343 18173 8352 18207
rect 8668 18232 8720 18284
rect 8300 18164 8352 18173
rect 8760 18164 8812 18216
rect 8116 18096 8168 18148
rect 9312 18164 9364 18216
rect 9588 18232 9640 18284
rect 10324 18207 10376 18216
rect 10324 18173 10333 18207
rect 10333 18173 10367 18207
rect 10367 18173 10376 18207
rect 10324 18164 10376 18173
rect 10508 18164 10560 18216
rect 11060 18207 11112 18216
rect 11060 18173 11069 18207
rect 11069 18173 11103 18207
rect 11103 18173 11112 18207
rect 11060 18164 11112 18173
rect 11980 18207 12032 18216
rect 11980 18173 11989 18207
rect 11989 18173 12023 18207
rect 12023 18173 12032 18207
rect 11980 18164 12032 18173
rect 11244 18096 11296 18148
rect 12348 18096 12400 18148
rect 14280 18300 14332 18352
rect 14372 18343 14424 18352
rect 14372 18309 14381 18343
rect 14381 18309 14415 18343
rect 14415 18309 14424 18343
rect 14740 18343 14792 18352
rect 14372 18300 14424 18309
rect 14740 18309 14749 18343
rect 14749 18309 14783 18343
rect 14783 18309 14792 18343
rect 14740 18300 14792 18309
rect 15384 18300 15436 18352
rect 19800 18343 19852 18352
rect 13544 18275 13596 18284
rect 13544 18241 13553 18275
rect 13553 18241 13587 18275
rect 13587 18241 13596 18275
rect 13544 18232 13596 18241
rect 16948 18232 17000 18284
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 18696 18275 18748 18284
rect 18696 18241 18705 18275
rect 18705 18241 18739 18275
rect 18739 18241 18748 18275
rect 18696 18232 18748 18241
rect 19064 18232 19116 18284
rect 19800 18309 19809 18343
rect 19809 18309 19843 18343
rect 19843 18309 19852 18343
rect 19800 18300 19852 18309
rect 14556 18164 14608 18216
rect 18788 18164 18840 18216
rect 20260 18232 20312 18284
rect 13452 18096 13504 18148
rect 16396 18096 16448 18148
rect 21364 18096 21416 18148
rect 4896 18028 4948 18080
rect 5448 18028 5500 18080
rect 9864 18028 9916 18080
rect 10968 18028 11020 18080
rect 11060 18028 11112 18080
rect 11980 18028 12032 18080
rect 14280 18028 14332 18080
rect 15016 18028 15068 18080
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 19524 18071 19576 18080
rect 19524 18037 19533 18071
rect 19533 18037 19567 18071
rect 19567 18037 19576 18071
rect 19524 18028 19576 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1676 17824 1728 17876
rect 2044 17824 2096 17876
rect 3332 17824 3384 17876
rect 3884 17824 3936 17876
rect 4068 17824 4120 17876
rect 1768 17688 1820 17740
rect 2688 17688 2740 17740
rect 2872 17799 2924 17808
rect 2872 17765 2881 17799
rect 2881 17765 2915 17799
rect 2915 17765 2924 17799
rect 5356 17824 5408 17876
rect 2872 17756 2924 17765
rect 6276 17824 6328 17876
rect 6920 17867 6972 17876
rect 6920 17833 6929 17867
rect 6929 17833 6963 17867
rect 6963 17833 6972 17867
rect 6920 17824 6972 17833
rect 7840 17824 7892 17876
rect 8300 17824 8352 17876
rect 8484 17824 8536 17876
rect 2320 17620 2372 17672
rect 3332 17620 3384 17672
rect 3976 17688 4028 17740
rect 4436 17731 4488 17740
rect 4436 17697 4445 17731
rect 4445 17697 4479 17731
rect 4479 17697 4488 17731
rect 4436 17688 4488 17697
rect 4620 17663 4672 17672
rect 4620 17629 4629 17663
rect 4629 17629 4663 17663
rect 4663 17629 4672 17663
rect 4620 17620 4672 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 2044 17552 2096 17604
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2780 17552 2832 17604
rect 5356 17731 5408 17740
rect 5356 17697 5365 17731
rect 5365 17697 5399 17731
rect 5399 17697 5408 17731
rect 5356 17688 5408 17697
rect 5448 17663 5500 17672
rect 5448 17629 5457 17663
rect 5457 17629 5491 17663
rect 5491 17629 5500 17663
rect 5448 17620 5500 17629
rect 5632 17620 5684 17672
rect 6828 17688 6880 17740
rect 8576 17756 8628 17808
rect 7748 17731 7800 17740
rect 7748 17697 7757 17731
rect 7757 17697 7791 17731
rect 7791 17697 7800 17731
rect 7748 17688 7800 17697
rect 7932 17688 7984 17740
rect 8484 17731 8536 17740
rect 8484 17697 8493 17731
rect 8493 17697 8527 17731
rect 8527 17697 8536 17731
rect 8484 17688 8536 17697
rect 7012 17620 7064 17672
rect 7288 17663 7340 17672
rect 7288 17629 7297 17663
rect 7297 17629 7331 17663
rect 7331 17629 7340 17663
rect 7288 17620 7340 17629
rect 9864 17824 9916 17876
rect 10048 17824 10100 17876
rect 10692 17824 10744 17876
rect 11888 17824 11940 17876
rect 13360 17824 13412 17876
rect 13544 17824 13596 17876
rect 10140 17756 10192 17808
rect 9956 17688 10008 17740
rect 10876 17688 10928 17740
rect 11060 17731 11112 17740
rect 11060 17697 11069 17731
rect 11069 17697 11103 17731
rect 11103 17697 11112 17731
rect 11060 17688 11112 17697
rect 11704 17756 11756 17808
rect 12992 17756 13044 17808
rect 13820 17799 13872 17808
rect 13820 17765 13829 17799
rect 13829 17765 13863 17799
rect 13863 17765 13872 17799
rect 13820 17756 13872 17765
rect 17408 17824 17460 17876
rect 19064 17824 19116 17876
rect 19616 17824 19668 17876
rect 18052 17756 18104 17808
rect 2596 17484 2648 17536
rect 6276 17552 6328 17604
rect 9496 17620 9548 17672
rect 10324 17620 10376 17672
rect 11244 17620 11296 17672
rect 11428 17620 11480 17672
rect 3976 17484 4028 17536
rect 4160 17527 4212 17536
rect 4160 17493 4169 17527
rect 4169 17493 4203 17527
rect 4203 17493 4212 17527
rect 4160 17484 4212 17493
rect 5080 17484 5132 17536
rect 5724 17484 5776 17536
rect 5908 17527 5960 17536
rect 5908 17493 5917 17527
rect 5917 17493 5951 17527
rect 5951 17493 5960 17527
rect 5908 17484 5960 17493
rect 6000 17527 6052 17536
rect 6000 17493 6009 17527
rect 6009 17493 6043 17527
rect 6043 17493 6052 17527
rect 7656 17552 7708 17604
rect 10876 17552 10928 17604
rect 6000 17484 6052 17493
rect 7288 17484 7340 17536
rect 7748 17484 7800 17536
rect 10324 17527 10376 17536
rect 10324 17493 10333 17527
rect 10333 17493 10367 17527
rect 10367 17493 10376 17527
rect 10324 17484 10376 17493
rect 10508 17527 10560 17536
rect 10508 17493 10517 17527
rect 10517 17493 10551 17527
rect 10551 17493 10560 17527
rect 10508 17484 10560 17493
rect 10692 17484 10744 17536
rect 12164 17527 12216 17536
rect 12164 17493 12173 17527
rect 12173 17493 12207 17527
rect 12207 17493 12216 17527
rect 12164 17484 12216 17493
rect 12348 17552 12400 17604
rect 13728 17620 13780 17672
rect 16028 17688 16080 17740
rect 16856 17731 16908 17740
rect 16856 17697 16865 17731
rect 16865 17697 16899 17731
rect 16899 17697 16908 17731
rect 16856 17688 16908 17697
rect 17040 17620 17092 17672
rect 18696 17620 18748 17672
rect 19064 17663 19116 17672
rect 19064 17629 19073 17663
rect 19073 17629 19107 17663
rect 19107 17629 19116 17663
rect 19064 17620 19116 17629
rect 19616 17688 19668 17740
rect 20076 17824 20128 17876
rect 20444 17824 20496 17876
rect 21272 17756 21324 17808
rect 19708 17663 19760 17672
rect 19708 17629 19717 17663
rect 19717 17629 19751 17663
rect 19751 17629 19760 17663
rect 19708 17620 19760 17629
rect 19800 17663 19852 17672
rect 19800 17629 19809 17663
rect 19809 17629 19843 17663
rect 19843 17629 19852 17663
rect 20076 17663 20128 17672
rect 19800 17620 19852 17629
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 20352 17663 20404 17672
rect 20352 17629 20361 17663
rect 20361 17629 20395 17663
rect 20395 17629 20404 17663
rect 20352 17620 20404 17629
rect 20720 17663 20772 17672
rect 20720 17629 20729 17663
rect 20729 17629 20763 17663
rect 20763 17629 20772 17663
rect 20720 17620 20772 17629
rect 21088 17620 21140 17672
rect 13820 17552 13872 17604
rect 16212 17552 16264 17604
rect 12532 17484 12584 17536
rect 13084 17527 13136 17536
rect 13084 17493 13093 17527
rect 13093 17493 13127 17527
rect 13127 17493 13136 17527
rect 13084 17484 13136 17493
rect 13268 17484 13320 17536
rect 15108 17484 15160 17536
rect 15568 17484 15620 17536
rect 15936 17527 15988 17536
rect 15936 17493 15945 17527
rect 15945 17493 15979 17527
rect 15979 17493 15988 17527
rect 16304 17527 16356 17536
rect 15936 17484 15988 17493
rect 16304 17493 16313 17527
rect 16313 17493 16347 17527
rect 16347 17493 16356 17527
rect 16304 17484 16356 17493
rect 18144 17484 18196 17536
rect 20536 17527 20588 17536
rect 20536 17493 20545 17527
rect 20545 17493 20579 17527
rect 20579 17493 20588 17527
rect 20536 17484 20588 17493
rect 20904 17552 20956 17604
rect 22652 17552 22704 17604
rect 21456 17527 21508 17536
rect 21456 17493 21465 17527
rect 21465 17493 21499 17527
rect 21499 17493 21508 17527
rect 21456 17484 21508 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 1768 17280 1820 17332
rect 4436 17255 4488 17264
rect 4436 17221 4470 17255
rect 4470 17221 4488 17255
rect 4436 17212 4488 17221
rect 5080 17212 5132 17264
rect 5724 17280 5776 17332
rect 6552 17280 6604 17332
rect 7104 17280 7156 17332
rect 8392 17280 8444 17332
rect 8668 17280 8720 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 9956 17280 10008 17332
rect 10508 17323 10560 17332
rect 10508 17289 10517 17323
rect 10517 17289 10551 17323
rect 10551 17289 10560 17323
rect 10508 17280 10560 17289
rect 10784 17280 10836 17332
rect 12348 17323 12400 17332
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 1860 17144 1912 17196
rect 2412 17187 2464 17196
rect 2412 17153 2421 17187
rect 2421 17153 2455 17187
rect 2455 17153 2464 17187
rect 2412 17144 2464 17153
rect 3240 17144 3292 17196
rect 5724 17144 5776 17196
rect 6184 17212 6236 17264
rect 6368 17144 6420 17196
rect 1952 17008 2004 17060
rect 1492 16983 1544 16992
rect 1492 16949 1501 16983
rect 1501 16949 1535 16983
rect 1535 16949 1544 16983
rect 1492 16940 1544 16949
rect 2136 16983 2188 16992
rect 2136 16949 2145 16983
rect 2145 16949 2179 16983
rect 2179 16949 2188 16983
rect 2136 16940 2188 16949
rect 2228 16983 2280 16992
rect 2228 16949 2237 16983
rect 2237 16949 2271 16983
rect 2271 16949 2280 16983
rect 2228 16940 2280 16949
rect 5540 17076 5592 17128
rect 6460 17076 6512 17128
rect 8208 17212 8260 17264
rect 8300 17212 8352 17264
rect 9128 17212 9180 17264
rect 12348 17289 12357 17323
rect 12357 17289 12391 17323
rect 12391 17289 12400 17323
rect 12348 17280 12400 17289
rect 12440 17280 12492 17332
rect 15568 17280 15620 17332
rect 16212 17323 16264 17332
rect 7380 17144 7432 17196
rect 7840 17144 7892 17196
rect 6736 17119 6788 17128
rect 6736 17085 6745 17119
rect 6745 17085 6779 17119
rect 6779 17085 6788 17119
rect 6736 17076 6788 17085
rect 8668 17144 8720 17196
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 9772 17187 9824 17196
rect 9772 17153 9781 17187
rect 9781 17153 9815 17187
rect 9815 17153 9824 17187
rect 9772 17144 9824 17153
rect 10692 17144 10744 17196
rect 10968 17144 11020 17196
rect 12072 17212 12124 17264
rect 12992 17212 13044 17264
rect 13360 17212 13412 17264
rect 14648 17212 14700 17264
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 16304 17280 16356 17332
rect 19616 17323 19668 17332
rect 19616 17289 19625 17323
rect 19625 17289 19659 17323
rect 19659 17289 19668 17323
rect 19616 17280 19668 17289
rect 19892 17323 19944 17332
rect 19892 17289 19901 17323
rect 19901 17289 19935 17323
rect 19935 17289 19944 17323
rect 19892 17280 19944 17289
rect 20812 17280 20864 17332
rect 22376 17280 22428 17332
rect 4436 16940 4488 16992
rect 7104 16940 7156 16992
rect 8484 17008 8536 17060
rect 9128 17076 9180 17128
rect 10048 17119 10100 17128
rect 10048 17085 10057 17119
rect 10057 17085 10091 17119
rect 10091 17085 10100 17119
rect 10048 17076 10100 17085
rect 10324 17119 10376 17128
rect 10324 17085 10333 17119
rect 10333 17085 10367 17119
rect 10367 17085 10376 17119
rect 10324 17076 10376 17085
rect 8852 17008 8904 17060
rect 11244 17051 11296 17060
rect 11244 17017 11253 17051
rect 11253 17017 11287 17051
rect 11287 17017 11296 17051
rect 12716 17144 12768 17196
rect 13176 17144 13228 17196
rect 13452 17187 13504 17196
rect 13452 17153 13470 17187
rect 13470 17153 13504 17187
rect 13728 17187 13780 17196
rect 13452 17144 13504 17153
rect 13728 17153 13737 17187
rect 13737 17153 13771 17187
rect 13771 17153 13780 17187
rect 13728 17144 13780 17153
rect 15200 17144 15252 17196
rect 15384 17187 15436 17196
rect 15384 17153 15393 17187
rect 15393 17153 15427 17187
rect 15427 17153 15436 17187
rect 15384 17144 15436 17153
rect 18880 17212 18932 17264
rect 16396 17187 16448 17196
rect 15016 17076 15068 17128
rect 15292 17119 15344 17128
rect 11244 17008 11296 17017
rect 14280 17008 14332 17060
rect 15292 17085 15301 17119
rect 15301 17085 15335 17119
rect 15335 17085 15344 17119
rect 15292 17076 15344 17085
rect 16396 17153 16405 17187
rect 16405 17153 16439 17187
rect 16439 17153 16448 17187
rect 16396 17144 16448 17153
rect 19432 17144 19484 17196
rect 19524 17144 19576 17196
rect 15660 17008 15712 17060
rect 8576 16940 8628 16992
rect 10140 16940 10192 16992
rect 10692 16940 10744 16992
rect 12072 16940 12124 16992
rect 12256 16983 12308 16992
rect 12256 16949 12265 16983
rect 12265 16949 12299 16983
rect 12299 16949 12308 16983
rect 12256 16940 12308 16949
rect 12348 16940 12400 16992
rect 14648 16940 14700 16992
rect 14924 16940 14976 16992
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 19064 17076 19116 17128
rect 16948 17008 17000 17060
rect 18512 17008 18564 17060
rect 20996 17187 21048 17196
rect 20996 17153 21005 17187
rect 21005 17153 21039 17187
rect 21039 17153 21048 17187
rect 21272 17187 21324 17196
rect 20996 17144 21048 17153
rect 21272 17153 21281 17187
rect 21281 17153 21315 17187
rect 21315 17153 21324 17187
rect 21272 17144 21324 17153
rect 16396 16940 16448 16992
rect 17132 16940 17184 16992
rect 19616 16940 19668 16992
rect 19800 16983 19852 16992
rect 19800 16949 19809 16983
rect 19809 16949 19843 16983
rect 19843 16949 19852 16983
rect 19800 16940 19852 16949
rect 20076 16940 20128 16992
rect 20168 16983 20220 16992
rect 20168 16949 20177 16983
rect 20177 16949 20211 16983
rect 20211 16949 20220 16983
rect 20168 16940 20220 16949
rect 20628 16940 20680 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1676 16736 1728 16788
rect 5356 16736 5408 16788
rect 6460 16779 6512 16788
rect 1768 16668 1820 16720
rect 3240 16643 3292 16652
rect 3240 16609 3249 16643
rect 3249 16609 3283 16643
rect 3283 16609 3292 16643
rect 3240 16600 3292 16609
rect 2228 16532 2280 16584
rect 2044 16464 2096 16516
rect 2964 16507 3016 16516
rect 2964 16473 2982 16507
rect 2982 16473 3016 16507
rect 2964 16464 3016 16473
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 5632 16668 5684 16720
rect 6000 16668 6052 16720
rect 6184 16711 6236 16720
rect 6184 16677 6193 16711
rect 6193 16677 6227 16711
rect 6227 16677 6236 16711
rect 6184 16668 6236 16677
rect 6460 16745 6469 16779
rect 6469 16745 6503 16779
rect 6503 16745 6512 16779
rect 6460 16736 6512 16745
rect 9404 16736 9456 16788
rect 10876 16779 10928 16788
rect 6828 16668 6880 16720
rect 7932 16668 7984 16720
rect 8852 16668 8904 16720
rect 10876 16745 10885 16779
rect 10885 16745 10919 16779
rect 10919 16745 10928 16779
rect 10876 16736 10928 16745
rect 12348 16736 12400 16788
rect 12440 16736 12492 16788
rect 13544 16779 13596 16788
rect 13544 16745 13553 16779
rect 13553 16745 13587 16779
rect 13587 16745 13596 16779
rect 13544 16736 13596 16745
rect 15660 16711 15712 16720
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4712 16575 4764 16584
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 1676 16396 1728 16448
rect 4252 16396 4304 16448
rect 4712 16541 4721 16575
rect 4721 16541 4755 16575
rect 4755 16541 4764 16575
rect 4712 16532 4764 16541
rect 7840 16643 7892 16652
rect 7840 16609 7849 16643
rect 7849 16609 7883 16643
rect 7883 16609 7892 16643
rect 7840 16600 7892 16609
rect 8576 16643 8628 16652
rect 8576 16609 8585 16643
rect 8585 16609 8619 16643
rect 8619 16609 8628 16643
rect 8576 16600 8628 16609
rect 5908 16532 5960 16584
rect 6000 16575 6052 16584
rect 6000 16541 6009 16575
rect 6009 16541 6043 16575
rect 6043 16541 6052 16575
rect 6276 16575 6328 16584
rect 6000 16532 6052 16541
rect 6276 16541 6285 16575
rect 6285 16541 6319 16575
rect 6319 16541 6328 16575
rect 6276 16532 6328 16541
rect 6368 16532 6420 16584
rect 7012 16532 7064 16584
rect 7288 16532 7340 16584
rect 8484 16575 8536 16584
rect 8484 16541 8493 16575
rect 8493 16541 8527 16575
rect 8527 16541 8536 16575
rect 9496 16643 9548 16652
rect 9496 16609 9505 16643
rect 9505 16609 9539 16643
rect 9539 16609 9548 16643
rect 9496 16600 9548 16609
rect 11152 16600 11204 16652
rect 11520 16643 11572 16652
rect 11520 16609 11529 16643
rect 11529 16609 11563 16643
rect 11563 16609 11572 16643
rect 11520 16600 11572 16609
rect 11704 16643 11756 16652
rect 11704 16609 11713 16643
rect 11713 16609 11747 16643
rect 11747 16609 11756 16643
rect 11704 16600 11756 16609
rect 15660 16677 15669 16711
rect 15669 16677 15703 16711
rect 15703 16677 15712 16711
rect 15660 16668 15712 16677
rect 17224 16736 17276 16788
rect 17316 16779 17368 16788
rect 17316 16745 17325 16779
rect 17325 16745 17359 16779
rect 17359 16745 17368 16779
rect 17316 16736 17368 16745
rect 18696 16736 18748 16788
rect 20168 16736 20220 16788
rect 17500 16668 17552 16720
rect 17776 16711 17828 16720
rect 17776 16677 17785 16711
rect 17785 16677 17819 16711
rect 17819 16677 17828 16711
rect 17776 16668 17828 16677
rect 17960 16711 18012 16720
rect 17960 16677 17969 16711
rect 17969 16677 18003 16711
rect 18003 16677 18012 16711
rect 17960 16668 18012 16677
rect 18604 16668 18656 16720
rect 20260 16668 20312 16720
rect 13544 16600 13596 16652
rect 14280 16643 14332 16652
rect 14280 16609 14289 16643
rect 14289 16609 14323 16643
rect 14323 16609 14332 16643
rect 14280 16600 14332 16609
rect 8484 16532 8536 16541
rect 10508 16532 10560 16584
rect 11244 16575 11296 16584
rect 11244 16541 11253 16575
rect 11253 16541 11287 16575
rect 11287 16541 11296 16575
rect 11244 16532 11296 16541
rect 12992 16532 13044 16584
rect 13636 16532 13688 16584
rect 17316 16600 17368 16652
rect 17868 16600 17920 16652
rect 19984 16643 20036 16652
rect 19984 16609 19993 16643
rect 19993 16609 20027 16643
rect 20027 16609 20036 16643
rect 19984 16600 20036 16609
rect 21272 16736 21324 16788
rect 21088 16668 21140 16720
rect 21732 16600 21784 16652
rect 16028 16575 16080 16584
rect 16028 16541 16051 16575
rect 16051 16541 16080 16575
rect 5448 16464 5500 16516
rect 8116 16464 8168 16516
rect 8208 16464 8260 16516
rect 4528 16396 4580 16448
rect 5080 16439 5132 16448
rect 5080 16405 5089 16439
rect 5089 16405 5123 16439
rect 5123 16405 5132 16439
rect 5080 16396 5132 16405
rect 5540 16396 5592 16448
rect 5908 16439 5960 16448
rect 5908 16405 5917 16439
rect 5917 16405 5951 16439
rect 5951 16405 5960 16439
rect 5908 16396 5960 16405
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 8392 16439 8444 16448
rect 8392 16405 8401 16439
rect 8401 16405 8435 16439
rect 8435 16405 8444 16439
rect 8392 16396 8444 16405
rect 10048 16464 10100 16516
rect 10324 16464 10376 16516
rect 10784 16464 10836 16516
rect 12440 16464 12492 16516
rect 12624 16464 12676 16516
rect 15108 16464 15160 16516
rect 15200 16464 15252 16516
rect 16028 16532 16080 16541
rect 16948 16464 17000 16516
rect 10692 16396 10744 16448
rect 11888 16396 11940 16448
rect 12808 16396 12860 16448
rect 13728 16396 13780 16448
rect 13912 16439 13964 16448
rect 13912 16405 13921 16439
rect 13921 16405 13955 16439
rect 13955 16405 13964 16439
rect 13912 16396 13964 16405
rect 14372 16396 14424 16448
rect 14740 16396 14792 16448
rect 19892 16532 19944 16584
rect 18052 16464 18104 16516
rect 20168 16464 20220 16516
rect 17500 16396 17552 16448
rect 18420 16396 18472 16448
rect 18880 16396 18932 16448
rect 20812 16575 20864 16584
rect 20812 16541 20821 16575
rect 20821 16541 20855 16575
rect 20855 16541 20864 16575
rect 20812 16532 20864 16541
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 21456 16439 21508 16448
rect 21456 16405 21465 16439
rect 21465 16405 21499 16439
rect 21499 16405 21508 16439
rect 21456 16396 21508 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 2964 16192 3016 16244
rect 4896 16192 4948 16244
rect 5264 16235 5316 16244
rect 5264 16201 5273 16235
rect 5273 16201 5307 16235
rect 5307 16201 5316 16235
rect 5264 16192 5316 16201
rect 5908 16192 5960 16244
rect 6736 16192 6788 16244
rect 7196 16235 7248 16244
rect 7196 16201 7205 16235
rect 7205 16201 7239 16235
rect 7239 16201 7248 16235
rect 7196 16192 7248 16201
rect 8208 16192 8260 16244
rect 10324 16235 10376 16244
rect 2228 16124 2280 16176
rect 2412 16124 2464 16176
rect 1676 16099 1728 16108
rect 1676 16065 1685 16099
rect 1685 16065 1719 16099
rect 1719 16065 1728 16099
rect 1676 16056 1728 16065
rect 2964 16099 3016 16108
rect 2964 16065 2973 16099
rect 2973 16065 3007 16099
rect 3007 16065 3016 16099
rect 2964 16056 3016 16065
rect 6092 16124 6144 16176
rect 1768 15988 1820 16040
rect 3056 16031 3108 16040
rect 3056 15997 3065 16031
rect 3065 15997 3099 16031
rect 3099 15997 3108 16031
rect 3056 15988 3108 15997
rect 4068 16031 4120 16040
rect 4068 15997 4077 16031
rect 4077 15997 4111 16031
rect 4111 15997 4120 16031
rect 4068 15988 4120 15997
rect 4344 16056 4396 16108
rect 4896 16031 4948 16040
rect 4896 15997 4905 16031
rect 4905 15997 4939 16031
rect 4939 15997 4948 16031
rect 4896 15988 4948 15997
rect 5264 16056 5316 16108
rect 3976 15920 4028 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 2504 15895 2556 15904
rect 2504 15861 2513 15895
rect 2513 15861 2547 15895
rect 2547 15861 2556 15895
rect 2504 15852 2556 15861
rect 4344 15852 4396 15904
rect 4804 15920 4856 15972
rect 5356 15988 5408 16040
rect 5540 16031 5592 16040
rect 5540 15997 5549 16031
rect 5549 15997 5583 16031
rect 5583 15997 5592 16031
rect 5540 15988 5592 15997
rect 5908 16056 5960 16108
rect 8116 16056 8168 16108
rect 9496 16124 9548 16176
rect 10324 16201 10333 16235
rect 10333 16201 10367 16235
rect 10367 16201 10376 16235
rect 10324 16192 10376 16201
rect 10600 16235 10652 16244
rect 10600 16201 10609 16235
rect 10609 16201 10643 16235
rect 10643 16201 10652 16235
rect 10600 16192 10652 16201
rect 11244 16192 11296 16244
rect 12624 16235 12676 16244
rect 12624 16201 12633 16235
rect 12633 16201 12667 16235
rect 12667 16201 12676 16235
rect 12624 16192 12676 16201
rect 13084 16192 13136 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 13912 16192 13964 16244
rect 15292 16192 15344 16244
rect 15660 16192 15712 16244
rect 12164 16124 12216 16176
rect 12348 16124 12400 16176
rect 14372 16124 14424 16176
rect 14832 16124 14884 16176
rect 15936 16192 15988 16244
rect 17224 16192 17276 16244
rect 18052 16192 18104 16244
rect 18236 16192 18288 16244
rect 19156 16235 19208 16244
rect 19156 16201 19165 16235
rect 19165 16201 19199 16235
rect 19199 16201 19208 16235
rect 19156 16192 19208 16201
rect 19892 16235 19944 16244
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 20352 16192 20404 16244
rect 18328 16167 18380 16176
rect 18328 16133 18337 16167
rect 18337 16133 18371 16167
rect 18371 16133 18380 16167
rect 18328 16124 18380 16133
rect 21088 16167 21140 16176
rect 6184 15988 6236 16040
rect 6552 15988 6604 16040
rect 8208 16031 8260 16040
rect 8208 15997 8217 16031
rect 8217 15997 8251 16031
rect 8251 15997 8260 16031
rect 8208 15988 8260 15997
rect 8392 15988 8444 16040
rect 9588 16056 9640 16108
rect 10968 16099 11020 16108
rect 10968 16065 10977 16099
rect 10977 16065 11011 16099
rect 11011 16065 11020 16099
rect 10968 16056 11020 16065
rect 11336 16056 11388 16108
rect 12808 16056 12860 16108
rect 13176 16056 13228 16108
rect 13636 16056 13688 16108
rect 16764 16056 16816 16108
rect 10876 15988 10928 16040
rect 12716 16031 12768 16040
rect 12716 15997 12725 16031
rect 12725 15997 12759 16031
rect 12759 15997 12768 16031
rect 12716 15988 12768 15997
rect 13452 16031 13504 16040
rect 13452 15997 13461 16031
rect 13461 15997 13495 16031
rect 13495 15997 13504 16031
rect 13452 15988 13504 15997
rect 13544 16031 13596 16040
rect 13544 15997 13553 16031
rect 13553 15997 13587 16031
rect 13587 15997 13596 16031
rect 13544 15988 13596 15997
rect 5908 15920 5960 15972
rect 6460 15920 6512 15972
rect 6736 15920 6788 15972
rect 6920 15920 6972 15972
rect 7380 15920 7432 15972
rect 8852 15920 8904 15972
rect 6092 15852 6144 15904
rect 6644 15852 6696 15904
rect 8576 15895 8628 15904
rect 8576 15861 8585 15895
rect 8585 15861 8619 15895
rect 8619 15861 8628 15895
rect 8576 15852 8628 15861
rect 13084 15920 13136 15972
rect 15108 15988 15160 16040
rect 16028 15988 16080 16040
rect 10232 15852 10284 15904
rect 10784 15852 10836 15904
rect 11336 15852 11388 15904
rect 11704 15895 11756 15904
rect 11704 15861 11713 15895
rect 11713 15861 11747 15895
rect 11747 15861 11756 15895
rect 11704 15852 11756 15861
rect 11888 15895 11940 15904
rect 11888 15861 11897 15895
rect 11897 15861 11931 15895
rect 11931 15861 11940 15895
rect 11888 15852 11940 15861
rect 12164 15895 12216 15904
rect 12164 15861 12173 15895
rect 12173 15861 12207 15895
rect 12207 15861 12216 15895
rect 12164 15852 12216 15861
rect 14648 15852 14700 15904
rect 19800 15988 19852 16040
rect 18328 15920 18380 15972
rect 19616 15920 19668 15972
rect 20168 16056 20220 16108
rect 21088 16133 21097 16167
rect 21097 16133 21131 16167
rect 21131 16133 21140 16167
rect 21088 16124 21140 16133
rect 20996 16056 21048 16108
rect 20352 15963 20404 15972
rect 17960 15852 18012 15904
rect 18512 15895 18564 15904
rect 18512 15861 18521 15895
rect 18521 15861 18555 15895
rect 18555 15861 18564 15895
rect 18512 15852 18564 15861
rect 19524 15895 19576 15904
rect 19524 15861 19533 15895
rect 19533 15861 19567 15895
rect 19567 15861 19576 15895
rect 19524 15852 19576 15861
rect 20352 15929 20361 15963
rect 20361 15929 20395 15963
rect 20395 15929 20404 15963
rect 20352 15920 20404 15929
rect 20536 15852 20588 15904
rect 21916 15920 21968 15972
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 2228 15691 2280 15700
rect 2228 15657 2237 15691
rect 2237 15657 2271 15691
rect 2271 15657 2280 15691
rect 2228 15648 2280 15657
rect 3240 15648 3292 15700
rect 5540 15648 5592 15700
rect 5632 15648 5684 15700
rect 6184 15648 6236 15700
rect 9128 15648 9180 15700
rect 4804 15580 4856 15632
rect 8668 15580 8720 15632
rect 1676 15487 1728 15496
rect 1676 15453 1685 15487
rect 1685 15453 1719 15487
rect 1719 15453 1728 15487
rect 1676 15444 1728 15453
rect 2044 15487 2096 15496
rect 2044 15453 2053 15487
rect 2053 15453 2087 15487
rect 2087 15453 2096 15487
rect 2044 15444 2096 15453
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 4620 15444 4672 15496
rect 5816 15444 5868 15496
rect 6276 15444 6328 15496
rect 6552 15487 6604 15496
rect 6552 15453 6570 15487
rect 6570 15453 6604 15487
rect 6552 15444 6604 15453
rect 7840 15512 7892 15564
rect 8392 15512 8444 15564
rect 9496 15648 9548 15700
rect 9588 15648 9640 15700
rect 9772 15648 9824 15700
rect 12348 15648 12400 15700
rect 13176 15691 13228 15700
rect 13176 15657 13185 15691
rect 13185 15657 13219 15691
rect 13219 15657 13228 15691
rect 13176 15648 13228 15657
rect 14648 15648 14700 15700
rect 15384 15648 15436 15700
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 9588 15512 9640 15564
rect 12440 15580 12492 15632
rect 12256 15512 12308 15564
rect 13636 15580 13688 15632
rect 15108 15512 15160 15564
rect 15292 15512 15344 15564
rect 9864 15444 9916 15496
rect 10508 15444 10560 15496
rect 6460 15376 6512 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 1860 15351 1912 15360
rect 1860 15317 1869 15351
rect 1869 15317 1903 15351
rect 1903 15317 1912 15351
rect 1860 15308 1912 15317
rect 2688 15308 2740 15360
rect 4712 15308 4764 15360
rect 5080 15308 5132 15360
rect 5540 15308 5592 15360
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 7380 15351 7432 15360
rect 7380 15317 7389 15351
rect 7389 15317 7423 15351
rect 7423 15317 7432 15351
rect 7748 15351 7800 15360
rect 7380 15308 7432 15317
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 8300 15351 8352 15360
rect 8300 15317 8309 15351
rect 8309 15317 8343 15351
rect 8343 15317 8352 15351
rect 8300 15308 8352 15317
rect 9772 15308 9824 15360
rect 12164 15444 12216 15496
rect 14372 15444 14424 15496
rect 14924 15487 14976 15496
rect 14924 15453 14933 15487
rect 14933 15453 14967 15487
rect 14967 15453 14976 15487
rect 14924 15444 14976 15453
rect 15660 15444 15712 15496
rect 16396 15444 16448 15496
rect 16764 15648 16816 15700
rect 17408 15648 17460 15700
rect 17500 15648 17552 15700
rect 18972 15648 19024 15700
rect 19064 15691 19116 15700
rect 19064 15657 19073 15691
rect 19073 15657 19107 15691
rect 19107 15657 19116 15691
rect 19064 15648 19116 15657
rect 19984 15648 20036 15700
rect 20168 15691 20220 15700
rect 20168 15657 20177 15691
rect 20177 15657 20211 15691
rect 20211 15657 20220 15691
rect 20168 15648 20220 15657
rect 20260 15648 20312 15700
rect 21272 15648 21324 15700
rect 17408 15512 17460 15564
rect 19892 15580 19944 15632
rect 22376 15580 22428 15632
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 17868 15512 17920 15564
rect 18420 15512 18472 15564
rect 19616 15512 19668 15564
rect 19800 15512 19852 15564
rect 22008 15512 22060 15564
rect 14280 15376 14332 15428
rect 18236 15444 18288 15496
rect 19340 15444 19392 15496
rect 20536 15487 20588 15496
rect 20536 15453 20545 15487
rect 20545 15453 20579 15487
rect 20579 15453 20588 15487
rect 20536 15444 20588 15453
rect 20720 15444 20772 15496
rect 21272 15487 21324 15496
rect 21272 15453 21281 15487
rect 21281 15453 21315 15487
rect 21315 15453 21324 15487
rect 21272 15444 21324 15453
rect 20996 15376 21048 15428
rect 22192 15376 22244 15428
rect 10048 15351 10100 15360
rect 10048 15317 10057 15351
rect 10057 15317 10091 15351
rect 10091 15317 10100 15351
rect 10048 15308 10100 15317
rect 10324 15308 10376 15360
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 12624 15351 12676 15360
rect 10876 15308 10928 15317
rect 12624 15317 12633 15351
rect 12633 15317 12667 15351
rect 12667 15317 12676 15351
rect 12624 15308 12676 15317
rect 13360 15308 13412 15360
rect 14648 15308 14700 15360
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 15200 15308 15252 15360
rect 15660 15351 15712 15360
rect 15660 15317 15669 15351
rect 15669 15317 15703 15351
rect 15703 15317 15712 15351
rect 15660 15308 15712 15317
rect 16120 15351 16172 15360
rect 16120 15317 16129 15351
rect 16129 15317 16163 15351
rect 16163 15317 16172 15351
rect 16120 15308 16172 15317
rect 16304 15308 16356 15360
rect 17776 15351 17828 15360
rect 17776 15317 17785 15351
rect 17785 15317 17819 15351
rect 17819 15317 17828 15351
rect 17776 15308 17828 15317
rect 17868 15308 17920 15360
rect 18696 15308 18748 15360
rect 20812 15308 20864 15360
rect 21088 15351 21140 15360
rect 21088 15317 21097 15351
rect 21097 15317 21131 15351
rect 21131 15317 21140 15351
rect 21088 15308 21140 15317
rect 21456 15351 21508 15360
rect 21456 15317 21465 15351
rect 21465 15317 21499 15351
rect 21499 15317 21508 15351
rect 21456 15308 21508 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 2044 15104 2096 15156
rect 2596 15104 2648 15156
rect 2964 15104 3016 15156
rect 4068 15104 4120 15156
rect 5172 15104 5224 15156
rect 6552 15104 6604 15156
rect 4252 15036 4304 15088
rect 7932 15104 7984 15156
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 8760 15104 8812 15156
rect 9588 15079 9640 15088
rect 2320 15011 2372 15020
rect 1584 14900 1636 14952
rect 2320 14977 2329 15011
rect 2329 14977 2363 15011
rect 2363 14977 2372 15011
rect 2320 14968 2372 14977
rect 2596 15011 2648 15020
rect 2596 14977 2605 15011
rect 2605 14977 2639 15011
rect 2639 14977 2648 15011
rect 2596 14968 2648 14977
rect 3240 14943 3292 14952
rect 3240 14909 3249 14943
rect 3249 14909 3283 14943
rect 3283 14909 3292 14943
rect 3240 14900 3292 14909
rect 4620 14943 4672 14952
rect 1400 14832 1452 14884
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1676 14832 1728 14884
rect 4620 14909 4629 14943
rect 4629 14909 4663 14943
rect 4663 14909 4672 14943
rect 4620 14900 4672 14909
rect 4160 14832 4212 14884
rect 6736 14968 6788 15020
rect 7104 14968 7156 15020
rect 9588 15045 9606 15079
rect 9606 15045 9640 15079
rect 10048 15104 10100 15156
rect 10416 15104 10468 15156
rect 10600 15104 10652 15156
rect 9588 15036 9640 15045
rect 8668 14968 8720 15020
rect 11060 15036 11112 15088
rect 8024 14900 8076 14952
rect 9864 14943 9916 14952
rect 9864 14909 9873 14943
rect 9873 14909 9907 14943
rect 9907 14909 9916 14943
rect 9864 14900 9916 14909
rect 10048 14900 10100 14952
rect 10968 14968 11020 15020
rect 12624 15104 12676 15156
rect 13360 15104 13412 15156
rect 12716 15036 12768 15088
rect 16120 15104 16172 15156
rect 17592 15104 17644 15156
rect 18880 15104 18932 15156
rect 20720 15104 20772 15156
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 15200 15036 15252 15088
rect 11520 14943 11572 14952
rect 4804 14832 4856 14884
rect 6092 14832 6144 14884
rect 7012 14832 7064 14884
rect 6000 14764 6052 14816
rect 6644 14807 6696 14816
rect 6644 14773 6653 14807
rect 6653 14773 6687 14807
rect 6687 14773 6696 14807
rect 6644 14764 6696 14773
rect 7196 14764 7248 14816
rect 10600 14764 10652 14816
rect 10784 14764 10836 14816
rect 11520 14909 11529 14943
rect 11529 14909 11563 14943
rect 11563 14909 11572 14943
rect 11520 14900 11572 14909
rect 13268 14900 13320 14952
rect 10968 14764 11020 14816
rect 11428 14764 11480 14816
rect 12440 14764 12492 14816
rect 13360 14764 13412 14816
rect 13728 14764 13780 14816
rect 14464 14900 14516 14952
rect 14740 14943 14792 14952
rect 14740 14909 14749 14943
rect 14749 14909 14783 14943
rect 14783 14909 14792 14943
rect 14740 14900 14792 14909
rect 15200 14900 15252 14952
rect 19340 15036 19392 15088
rect 15752 15011 15804 15020
rect 15752 14977 15761 15011
rect 15761 14977 15795 15011
rect 15795 14977 15804 15011
rect 15752 14968 15804 14977
rect 18236 14968 18288 15020
rect 18420 15011 18472 15020
rect 18420 14977 18454 15011
rect 18454 14977 18472 15011
rect 18420 14968 18472 14977
rect 18972 14968 19024 15020
rect 19984 15011 20036 15020
rect 19984 14977 19993 15011
rect 19993 14977 20027 15011
rect 20027 14977 20036 15011
rect 19984 14968 20036 14977
rect 15936 14943 15988 14952
rect 15936 14909 15945 14943
rect 15945 14909 15979 14943
rect 15979 14909 15988 14943
rect 15936 14900 15988 14909
rect 16396 14943 16448 14952
rect 16396 14909 16405 14943
rect 16405 14909 16439 14943
rect 16439 14909 16448 14943
rect 16396 14900 16448 14909
rect 19800 14943 19852 14952
rect 14464 14807 14516 14816
rect 14464 14773 14473 14807
rect 14473 14773 14507 14807
rect 14507 14773 14516 14807
rect 14464 14764 14516 14773
rect 14832 14764 14884 14816
rect 16948 14764 17000 14816
rect 17408 14764 17460 14816
rect 19800 14909 19809 14943
rect 19809 14909 19843 14943
rect 19843 14909 19852 14943
rect 19800 14900 19852 14909
rect 20444 14968 20496 15020
rect 20812 15011 20864 15020
rect 20812 14977 20821 15011
rect 20821 14977 20855 15011
rect 20855 14977 20864 15011
rect 20812 14968 20864 14977
rect 21180 14968 21232 15020
rect 22744 14900 22796 14952
rect 21272 14832 21324 14884
rect 19892 14764 19944 14816
rect 20996 14807 21048 14816
rect 20996 14773 21005 14807
rect 21005 14773 21039 14807
rect 21039 14773 21048 14807
rect 20996 14764 21048 14773
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 3056 14560 3108 14612
rect 4528 14560 4580 14612
rect 4804 14560 4856 14612
rect 5264 14560 5316 14612
rect 5724 14560 5776 14612
rect 6644 14560 6696 14612
rect 2964 14492 3016 14544
rect 6828 14492 6880 14544
rect 8208 14492 8260 14544
rect 112 14424 164 14476
rect 2228 14356 2280 14408
rect 2688 14356 2740 14408
rect 4160 14424 4212 14476
rect 5908 14424 5960 14476
rect 6552 14467 6604 14476
rect 6552 14433 6561 14467
rect 6561 14433 6595 14467
rect 6595 14433 6604 14467
rect 6552 14424 6604 14433
rect 6736 14424 6788 14476
rect 8024 14424 8076 14476
rect 10876 14560 10928 14612
rect 8484 14492 8536 14544
rect 11796 14560 11848 14612
rect 12164 14560 12216 14612
rect 12348 14560 12400 14612
rect 12624 14560 12676 14612
rect 13452 14560 13504 14612
rect 11520 14492 11572 14544
rect 8760 14424 8812 14476
rect 9220 14424 9272 14476
rect 9588 14424 9640 14476
rect 10600 14467 10652 14476
rect 10600 14433 10609 14467
rect 10609 14433 10643 14467
rect 10643 14433 10652 14467
rect 10600 14424 10652 14433
rect 12440 14467 12492 14476
rect 3884 14356 3936 14408
rect 5172 14356 5224 14408
rect 5264 14356 5316 14408
rect 6092 14356 6144 14408
rect 8116 14356 8168 14408
rect 8392 14356 8444 14408
rect 9128 14356 9180 14408
rect 9312 14356 9364 14408
rect 11152 14356 11204 14408
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 12624 14467 12676 14476
rect 12624 14433 12633 14467
rect 12633 14433 12667 14467
rect 12667 14433 12676 14467
rect 13360 14492 13412 14544
rect 14004 14492 14056 14544
rect 15936 14560 15988 14612
rect 18236 14560 18288 14612
rect 19984 14603 20036 14612
rect 12624 14424 12676 14433
rect 11428 14356 11480 14408
rect 13452 14399 13504 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2044 14263 2096 14272
rect 2044 14229 2053 14263
rect 2053 14229 2087 14263
rect 2087 14229 2096 14263
rect 2044 14220 2096 14229
rect 2412 14263 2464 14272
rect 2412 14229 2421 14263
rect 2421 14229 2455 14263
rect 2455 14229 2464 14263
rect 2412 14220 2464 14229
rect 3148 14263 3200 14272
rect 3148 14229 3157 14263
rect 3157 14229 3191 14263
rect 3191 14229 3200 14263
rect 3148 14220 3200 14229
rect 3516 14220 3568 14272
rect 4068 14263 4120 14272
rect 4068 14229 4077 14263
rect 4077 14229 4111 14263
rect 4111 14229 4120 14263
rect 4068 14220 4120 14229
rect 4436 14263 4488 14272
rect 4436 14229 4445 14263
rect 4445 14229 4479 14263
rect 4479 14229 4488 14263
rect 4436 14220 4488 14229
rect 4528 14263 4580 14272
rect 4528 14229 4537 14263
rect 4537 14229 4571 14263
rect 4571 14229 4580 14263
rect 4896 14288 4948 14340
rect 6736 14331 6788 14340
rect 6736 14297 6745 14331
rect 6745 14297 6779 14331
rect 6779 14297 6788 14331
rect 6736 14288 6788 14297
rect 7840 14288 7892 14340
rect 9404 14288 9456 14340
rect 12900 14288 12952 14340
rect 13452 14365 13461 14399
rect 13461 14365 13495 14399
rect 13495 14365 13504 14399
rect 13452 14356 13504 14365
rect 14280 14424 14332 14476
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 19984 14569 19993 14603
rect 19993 14569 20027 14603
rect 20027 14569 20036 14603
rect 19984 14560 20036 14569
rect 21088 14560 21140 14612
rect 18972 14492 19024 14544
rect 19156 14492 19208 14544
rect 19708 14424 19760 14476
rect 20536 14424 20588 14476
rect 20996 14424 21048 14476
rect 15476 14399 15528 14408
rect 15476 14365 15485 14399
rect 15485 14365 15519 14399
rect 15519 14365 15528 14399
rect 15476 14356 15528 14365
rect 16304 14356 16356 14408
rect 18788 14356 18840 14408
rect 19432 14356 19484 14408
rect 19800 14356 19852 14408
rect 4528 14220 4580 14229
rect 5264 14220 5316 14272
rect 5540 14263 5592 14272
rect 5540 14229 5549 14263
rect 5549 14229 5583 14263
rect 5583 14229 5592 14263
rect 5540 14220 5592 14229
rect 6552 14220 6604 14272
rect 7196 14263 7248 14272
rect 7196 14229 7205 14263
rect 7205 14229 7239 14263
rect 7239 14229 7248 14263
rect 7196 14220 7248 14229
rect 7288 14220 7340 14272
rect 7932 14220 7984 14272
rect 9220 14220 9272 14272
rect 9496 14263 9548 14272
rect 9496 14229 9505 14263
rect 9505 14229 9539 14263
rect 9539 14229 9548 14263
rect 9496 14220 9548 14229
rect 10048 14263 10100 14272
rect 10048 14229 10057 14263
rect 10057 14229 10091 14263
rect 10091 14229 10100 14263
rect 10048 14220 10100 14229
rect 10876 14220 10928 14272
rect 11244 14220 11296 14272
rect 11704 14220 11756 14272
rect 11888 14220 11940 14272
rect 13360 14220 13412 14272
rect 13544 14263 13596 14272
rect 13544 14229 13553 14263
rect 13553 14229 13587 14263
rect 13587 14229 13596 14263
rect 13544 14220 13596 14229
rect 14832 14220 14884 14272
rect 15292 14288 15344 14340
rect 15384 14220 15436 14272
rect 17868 14288 17920 14340
rect 19340 14288 19392 14340
rect 20168 14288 20220 14340
rect 16120 14220 16172 14272
rect 16948 14220 17000 14272
rect 17224 14220 17276 14272
rect 17408 14263 17460 14272
rect 17408 14229 17417 14263
rect 17417 14229 17451 14263
rect 17451 14229 17460 14263
rect 17408 14220 17460 14229
rect 18604 14220 18656 14272
rect 19524 14263 19576 14272
rect 19524 14229 19533 14263
rect 19533 14229 19567 14263
rect 19567 14229 19576 14263
rect 19524 14220 19576 14229
rect 19708 14220 19760 14272
rect 20536 14263 20588 14272
rect 20536 14229 20545 14263
rect 20545 14229 20579 14263
rect 20579 14229 20588 14263
rect 20536 14220 20588 14229
rect 21456 14263 21508 14272
rect 21456 14229 21465 14263
rect 21465 14229 21499 14263
rect 21499 14229 21508 14263
rect 21456 14220 21508 14229
rect 21824 14220 21876 14272
rect 22468 14220 22520 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 2596 14016 2648 14068
rect 2412 13948 2464 14000
rect 5264 14016 5316 14068
rect 5908 14059 5960 14068
rect 5908 14025 5917 14059
rect 5917 14025 5951 14059
rect 5951 14025 5960 14059
rect 5908 14016 5960 14025
rect 7104 14016 7156 14068
rect 8300 14016 8352 14068
rect 10048 14016 10100 14068
rect 10324 14059 10376 14068
rect 10324 14025 10333 14059
rect 10333 14025 10367 14059
rect 10367 14025 10376 14059
rect 10324 14016 10376 14025
rect 10876 14059 10928 14068
rect 10876 14025 10885 14059
rect 10885 14025 10919 14059
rect 10919 14025 10928 14059
rect 10876 14016 10928 14025
rect 11060 14016 11112 14068
rect 2044 13923 2096 13932
rect 2044 13889 2053 13923
rect 2053 13889 2087 13923
rect 2087 13889 2096 13923
rect 2044 13880 2096 13889
rect 2688 13880 2740 13932
rect 4620 13948 4672 14000
rect 6000 13948 6052 14000
rect 6644 13948 6696 14000
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 8484 13991 8536 14000
rect 6828 13948 6880 13957
rect 8484 13957 8493 13991
rect 8493 13957 8527 13991
rect 8527 13957 8536 13991
rect 8484 13948 8536 13957
rect 8576 13948 8628 14000
rect 10784 13948 10836 14000
rect 3332 13923 3384 13932
rect 2228 13812 2280 13864
rect 3332 13889 3366 13923
rect 3366 13889 3384 13923
rect 3332 13880 3384 13889
rect 1860 13787 1912 13796
rect 1860 13753 1869 13787
rect 1869 13753 1903 13787
rect 1903 13753 1912 13787
rect 1860 13744 1912 13753
rect 4068 13812 4120 13864
rect 1492 13719 1544 13728
rect 1492 13685 1501 13719
rect 1501 13685 1535 13719
rect 1535 13685 1544 13719
rect 1492 13676 1544 13685
rect 2688 13676 2740 13728
rect 4344 13676 4396 13728
rect 7012 13880 7064 13932
rect 5908 13812 5960 13864
rect 6460 13812 6512 13864
rect 9312 13880 9364 13932
rect 9496 13880 9548 13932
rect 6368 13744 6420 13796
rect 4712 13676 4764 13728
rect 6552 13676 6604 13728
rect 6828 13744 6880 13796
rect 8576 13812 8628 13864
rect 8760 13812 8812 13864
rect 9588 13812 9640 13864
rect 10416 13855 10468 13864
rect 10416 13821 10425 13855
rect 10425 13821 10459 13855
rect 10459 13821 10468 13855
rect 10416 13812 10468 13821
rect 10692 13855 10744 13864
rect 10692 13821 10701 13855
rect 10701 13821 10735 13855
rect 10735 13821 10744 13855
rect 10692 13812 10744 13821
rect 11152 13855 11204 13864
rect 11152 13821 11161 13855
rect 11161 13821 11195 13855
rect 11195 13821 11204 13855
rect 11152 13812 11204 13821
rect 11704 14016 11756 14068
rect 11796 14016 11848 14068
rect 11980 14016 12032 14068
rect 12992 14016 13044 14068
rect 15200 14059 15252 14068
rect 15200 14025 15209 14059
rect 15209 14025 15243 14059
rect 15243 14025 15252 14059
rect 15200 14016 15252 14025
rect 15476 14016 15528 14068
rect 17132 14016 17184 14068
rect 19340 14059 19392 14068
rect 19340 14025 19349 14059
rect 19349 14025 19383 14059
rect 19383 14025 19392 14059
rect 19340 14016 19392 14025
rect 19708 14059 19760 14068
rect 19708 14025 19717 14059
rect 19717 14025 19751 14059
rect 19751 14025 19760 14059
rect 19708 14016 19760 14025
rect 21088 14059 21140 14068
rect 12072 13948 12124 14000
rect 12532 13948 12584 14000
rect 13452 13948 13504 14000
rect 11336 13880 11388 13932
rect 11796 13880 11848 13932
rect 15660 13948 15712 14000
rect 18420 13948 18472 14000
rect 14004 13923 14056 13932
rect 14004 13889 14038 13923
rect 14038 13889 14056 13923
rect 14004 13880 14056 13889
rect 15108 13880 15160 13932
rect 16304 13880 16356 13932
rect 17224 13923 17276 13932
rect 17224 13889 17233 13923
rect 17233 13889 17267 13923
rect 17267 13889 17276 13923
rect 17224 13880 17276 13889
rect 18052 13923 18104 13932
rect 18052 13889 18061 13923
rect 18061 13889 18095 13923
rect 18095 13889 18104 13923
rect 18052 13880 18104 13889
rect 11612 13812 11664 13864
rect 12992 13855 13044 13864
rect 7932 13744 7984 13796
rect 8300 13787 8352 13796
rect 8300 13753 8309 13787
rect 8309 13753 8343 13787
rect 8343 13753 8352 13787
rect 8300 13744 8352 13753
rect 10140 13744 10192 13796
rect 6920 13676 6972 13728
rect 7656 13676 7708 13728
rect 8484 13676 8536 13728
rect 11520 13676 11572 13728
rect 11796 13744 11848 13796
rect 12992 13821 13001 13855
rect 13001 13821 13035 13855
rect 13035 13821 13044 13855
rect 12992 13812 13044 13821
rect 13176 13855 13228 13864
rect 13176 13821 13185 13855
rect 13185 13821 13219 13855
rect 13219 13821 13228 13855
rect 13176 13812 13228 13821
rect 14740 13812 14792 13864
rect 15660 13855 15712 13864
rect 15660 13821 15669 13855
rect 15669 13821 15703 13855
rect 15703 13821 15712 13855
rect 15660 13812 15712 13821
rect 15936 13812 15988 13864
rect 16580 13812 16632 13864
rect 17132 13855 17184 13864
rect 17132 13821 17141 13855
rect 17141 13821 17175 13855
rect 17175 13821 17184 13855
rect 17132 13812 17184 13821
rect 17592 13812 17644 13864
rect 17868 13855 17920 13864
rect 17868 13821 17877 13855
rect 17877 13821 17911 13855
rect 17911 13821 17920 13855
rect 19524 13948 19576 14000
rect 19616 13948 19668 14000
rect 21088 14025 21097 14059
rect 21097 14025 21131 14059
rect 21131 14025 21140 14059
rect 21088 14016 21140 14025
rect 21180 13948 21232 14000
rect 18880 13923 18932 13932
rect 18880 13889 18889 13923
rect 18889 13889 18923 13923
rect 18923 13889 18932 13923
rect 18880 13880 18932 13889
rect 20444 13923 20496 13932
rect 20444 13889 20453 13923
rect 20453 13889 20487 13923
rect 20487 13889 20496 13923
rect 20444 13880 20496 13889
rect 20720 13880 20772 13932
rect 21272 13923 21324 13932
rect 21272 13889 21281 13923
rect 21281 13889 21315 13923
rect 21315 13889 21324 13923
rect 21272 13880 21324 13889
rect 18972 13855 19024 13864
rect 17868 13812 17920 13821
rect 12624 13719 12676 13728
rect 12624 13685 12633 13719
rect 12633 13685 12667 13719
rect 12667 13685 12676 13719
rect 12624 13676 12676 13685
rect 12716 13676 12768 13728
rect 17224 13744 17276 13796
rect 14832 13676 14884 13728
rect 16212 13676 16264 13728
rect 16672 13676 16724 13728
rect 18972 13821 18981 13855
rect 18981 13821 19015 13855
rect 19015 13821 19024 13855
rect 18972 13812 19024 13821
rect 19156 13855 19208 13864
rect 19156 13821 19165 13855
rect 19165 13821 19199 13855
rect 19199 13821 19208 13855
rect 19156 13812 19208 13821
rect 19892 13855 19944 13864
rect 19892 13821 19901 13855
rect 19901 13821 19935 13855
rect 19935 13821 19944 13855
rect 19892 13812 19944 13821
rect 20076 13812 20128 13864
rect 20536 13812 20588 13864
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 3332 13472 3384 13524
rect 3424 13472 3476 13524
rect 3884 13515 3936 13524
rect 3884 13481 3893 13515
rect 3893 13481 3927 13515
rect 3927 13481 3936 13515
rect 3884 13472 3936 13481
rect 4528 13472 4580 13524
rect 4988 13472 5040 13524
rect 6736 13472 6788 13524
rect 7012 13515 7064 13524
rect 7012 13481 7021 13515
rect 7021 13481 7055 13515
rect 7055 13481 7064 13515
rect 7012 13472 7064 13481
rect 1676 13311 1728 13320
rect 1676 13277 1685 13311
rect 1685 13277 1719 13311
rect 1719 13277 1728 13311
rect 1676 13268 1728 13277
rect 4068 13336 4120 13388
rect 4344 13336 4396 13388
rect 5724 13336 5776 13388
rect 6368 13379 6420 13388
rect 6368 13345 6377 13379
rect 6377 13345 6411 13379
rect 6411 13345 6420 13379
rect 6368 13336 6420 13345
rect 4712 13268 4764 13320
rect 6920 13404 6972 13456
rect 7748 13472 7800 13524
rect 8024 13472 8076 13524
rect 9128 13404 9180 13456
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 6552 13268 6604 13320
rect 7196 13268 7248 13320
rect 11336 13472 11388 13524
rect 11520 13472 11572 13524
rect 15108 13515 15160 13524
rect 13084 13404 13136 13456
rect 13360 13404 13412 13456
rect 13820 13404 13872 13456
rect 14372 13404 14424 13456
rect 15108 13481 15117 13515
rect 15117 13481 15151 13515
rect 15151 13481 15160 13515
rect 15108 13472 15160 13481
rect 15752 13472 15804 13524
rect 18052 13515 18104 13524
rect 18052 13481 18061 13515
rect 18061 13481 18095 13515
rect 18095 13481 18104 13515
rect 18052 13472 18104 13481
rect 18420 13472 18472 13524
rect 20720 13515 20772 13524
rect 20720 13481 20729 13515
rect 20729 13481 20763 13515
rect 20763 13481 20772 13515
rect 20720 13472 20772 13481
rect 21272 13472 21324 13524
rect 9680 13379 9732 13388
rect 9680 13345 9689 13379
rect 9689 13345 9723 13379
rect 9723 13345 9732 13379
rect 11612 13379 11664 13388
rect 9680 13336 9732 13345
rect 11612 13345 11621 13379
rect 11621 13345 11655 13379
rect 11655 13345 11664 13379
rect 11612 13336 11664 13345
rect 15292 13336 15344 13388
rect 2320 13200 2372 13252
rect 3332 13243 3384 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 1860 13175 1912 13184
rect 1860 13141 1869 13175
rect 1869 13141 1903 13175
rect 1903 13141 1912 13175
rect 1860 13132 1912 13141
rect 3332 13209 3350 13243
rect 3350 13209 3384 13243
rect 3332 13200 3384 13209
rect 3148 13132 3200 13184
rect 3516 13132 3568 13184
rect 8208 13200 8260 13252
rect 9496 13243 9548 13252
rect 9496 13209 9505 13243
rect 9505 13209 9539 13243
rect 9539 13209 9548 13243
rect 9496 13200 9548 13209
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 4988 13175 5040 13184
rect 4988 13141 4997 13175
rect 4997 13141 5031 13175
rect 5031 13141 5040 13175
rect 4988 13132 5040 13141
rect 5448 13175 5500 13184
rect 5448 13141 5457 13175
rect 5457 13141 5491 13175
rect 5491 13141 5500 13175
rect 5448 13132 5500 13141
rect 6000 13132 6052 13184
rect 7564 13132 7616 13184
rect 7932 13132 7984 13184
rect 8668 13175 8720 13184
rect 8668 13141 8677 13175
rect 8677 13141 8711 13175
rect 8711 13141 8720 13175
rect 8668 13132 8720 13141
rect 8760 13132 8812 13184
rect 9956 13268 10008 13320
rect 10876 13200 10928 13252
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 10324 13132 10376 13184
rect 11060 13132 11112 13184
rect 15200 13268 15252 13320
rect 15476 13268 15528 13320
rect 16120 13336 16172 13388
rect 16212 13268 16264 13320
rect 16396 13311 16448 13320
rect 16396 13277 16405 13311
rect 16405 13277 16439 13311
rect 16439 13277 16448 13311
rect 16396 13268 16448 13277
rect 18972 13404 19024 13456
rect 19524 13404 19576 13456
rect 19616 13447 19668 13456
rect 19616 13413 19625 13447
rect 19625 13413 19659 13447
rect 19659 13413 19668 13447
rect 19616 13404 19668 13413
rect 22928 13404 22980 13456
rect 18144 13336 18196 13388
rect 19064 13336 19116 13388
rect 11980 13200 12032 13252
rect 12532 13200 12584 13252
rect 12256 13132 12308 13184
rect 12992 13175 13044 13184
rect 12992 13141 13001 13175
rect 13001 13141 13035 13175
rect 13035 13141 13044 13175
rect 12992 13132 13044 13141
rect 13084 13175 13136 13184
rect 13084 13141 13093 13175
rect 13093 13141 13127 13175
rect 13127 13141 13136 13175
rect 13360 13243 13412 13252
rect 13360 13209 13369 13243
rect 13369 13209 13403 13243
rect 13403 13209 13412 13243
rect 13820 13243 13872 13252
rect 13360 13200 13412 13209
rect 13820 13209 13829 13243
rect 13829 13209 13863 13243
rect 13863 13209 13872 13243
rect 13820 13200 13872 13209
rect 13084 13132 13136 13141
rect 13728 13132 13780 13184
rect 14648 13132 14700 13184
rect 15108 13200 15160 13252
rect 15936 13200 15988 13252
rect 19524 13200 19576 13252
rect 20536 13311 20588 13320
rect 20536 13277 20545 13311
rect 20545 13277 20579 13311
rect 20579 13277 20588 13311
rect 20536 13268 20588 13277
rect 21272 13311 21324 13320
rect 21272 13277 21281 13311
rect 21281 13277 21315 13311
rect 21315 13277 21324 13311
rect 21272 13268 21324 13277
rect 21824 13200 21876 13252
rect 15292 13132 15344 13184
rect 15568 13175 15620 13184
rect 15568 13141 15577 13175
rect 15577 13141 15611 13175
rect 15611 13141 15620 13175
rect 15568 13132 15620 13141
rect 16212 13132 16264 13184
rect 16396 13132 16448 13184
rect 17592 13175 17644 13184
rect 17592 13141 17601 13175
rect 17601 13141 17635 13175
rect 17635 13141 17644 13175
rect 17592 13132 17644 13141
rect 18420 13175 18472 13184
rect 18420 13141 18429 13175
rect 18429 13141 18463 13175
rect 18463 13141 18472 13175
rect 18420 13132 18472 13141
rect 18512 13175 18564 13184
rect 18512 13141 18521 13175
rect 18521 13141 18555 13175
rect 18555 13141 18564 13175
rect 19892 13175 19944 13184
rect 18512 13132 18564 13141
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 20076 13175 20128 13184
rect 20076 13141 20085 13175
rect 20085 13141 20119 13175
rect 20119 13141 20128 13175
rect 20076 13132 20128 13141
rect 21456 13175 21508 13184
rect 21456 13141 21465 13175
rect 21465 13141 21499 13175
rect 21499 13141 21508 13175
rect 21456 13132 21508 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 1676 12928 1728 12980
rect 4436 12971 4488 12980
rect 4436 12937 4445 12971
rect 4445 12937 4479 12971
rect 4479 12937 4488 12971
rect 4436 12928 4488 12937
rect 4896 12928 4948 12980
rect 2044 12860 2096 12912
rect 2780 12860 2832 12912
rect 3516 12860 3568 12912
rect 1676 12835 1728 12844
rect 1676 12801 1685 12835
rect 1685 12801 1719 12835
rect 1719 12801 1728 12835
rect 1676 12792 1728 12801
rect 1768 12792 1820 12844
rect 3240 12792 3292 12844
rect 4068 12835 4120 12844
rect 4068 12801 4077 12835
rect 4077 12801 4111 12835
rect 4111 12801 4120 12835
rect 4068 12792 4120 12801
rect 4344 12792 4396 12844
rect 5080 12792 5132 12844
rect 5448 12928 5500 12980
rect 6000 12928 6052 12980
rect 7380 12928 7432 12980
rect 8024 12971 8076 12980
rect 8024 12937 8033 12971
rect 8033 12937 8067 12971
rect 8067 12937 8076 12971
rect 8024 12928 8076 12937
rect 8668 12928 8720 12980
rect 6460 12860 6512 12912
rect 6736 12860 6788 12912
rect 7196 12835 7248 12844
rect 3884 12767 3936 12776
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 3884 12733 3893 12767
rect 3893 12733 3927 12767
rect 3927 12733 3936 12767
rect 3884 12724 3936 12733
rect 3332 12699 3384 12708
rect 3332 12665 3341 12699
rect 3341 12665 3375 12699
rect 3375 12665 3384 12699
rect 3332 12656 3384 12665
rect 2228 12588 2280 12640
rect 2688 12588 2740 12640
rect 3976 12588 4028 12640
rect 6828 12724 6880 12776
rect 4988 12656 5040 12708
rect 6460 12656 6512 12708
rect 6920 12656 6972 12708
rect 7196 12801 7205 12835
rect 7205 12801 7239 12835
rect 7239 12801 7248 12835
rect 7196 12792 7248 12801
rect 7748 12860 7800 12912
rect 8760 12860 8812 12912
rect 9772 12928 9824 12980
rect 10048 12928 10100 12980
rect 10968 12928 11020 12980
rect 9036 12860 9088 12912
rect 10140 12860 10192 12912
rect 11244 12928 11296 12980
rect 12348 12928 12400 12980
rect 13268 12928 13320 12980
rect 14924 12928 14976 12980
rect 15292 12971 15344 12980
rect 15292 12937 15301 12971
rect 15301 12937 15335 12971
rect 15335 12937 15344 12971
rect 15292 12928 15344 12937
rect 15660 12928 15712 12980
rect 15936 12928 15988 12980
rect 12992 12903 13044 12912
rect 7288 12767 7340 12776
rect 7288 12733 7297 12767
rect 7297 12733 7331 12767
rect 7331 12733 7340 12767
rect 7288 12724 7340 12733
rect 7380 12767 7432 12776
rect 7380 12733 7389 12767
rect 7389 12733 7423 12767
rect 7423 12733 7432 12767
rect 7380 12724 7432 12733
rect 7564 12724 7616 12776
rect 8208 12767 8260 12776
rect 8208 12733 8217 12767
rect 8217 12733 8251 12767
rect 8251 12733 8260 12767
rect 8208 12724 8260 12733
rect 8484 12724 8536 12776
rect 8852 12656 8904 12708
rect 5540 12588 5592 12640
rect 5816 12588 5868 12640
rect 6552 12588 6604 12640
rect 6828 12631 6880 12640
rect 6828 12597 6837 12631
rect 6837 12597 6871 12631
rect 6871 12597 6880 12631
rect 6828 12588 6880 12597
rect 8484 12588 8536 12640
rect 9128 12767 9180 12776
rect 9128 12733 9137 12767
rect 9137 12733 9171 12767
rect 9171 12733 9180 12767
rect 9128 12724 9180 12733
rect 9220 12656 9272 12708
rect 9772 12767 9824 12776
rect 9772 12733 9781 12767
rect 9781 12733 9815 12767
rect 9815 12733 9824 12767
rect 9772 12724 9824 12733
rect 10876 12724 10928 12776
rect 11704 12724 11756 12776
rect 12992 12869 13026 12903
rect 13026 12869 13044 12903
rect 12992 12860 13044 12869
rect 17592 12928 17644 12980
rect 12532 12792 12584 12844
rect 13544 12792 13596 12844
rect 13728 12792 13780 12844
rect 15476 12792 15528 12844
rect 15936 12835 15988 12844
rect 15936 12801 15945 12835
rect 15945 12801 15979 12835
rect 15979 12801 15988 12835
rect 15936 12792 15988 12801
rect 16396 12792 16448 12844
rect 16948 12792 17000 12844
rect 17592 12835 17644 12844
rect 12164 12767 12216 12776
rect 12164 12733 12173 12767
rect 12173 12733 12207 12767
rect 12207 12733 12216 12767
rect 12164 12724 12216 12733
rect 11244 12656 11296 12708
rect 16120 12724 16172 12776
rect 16212 12724 16264 12776
rect 17040 12724 17092 12776
rect 17592 12801 17601 12835
rect 17601 12801 17635 12835
rect 17635 12801 17644 12835
rect 17592 12792 17644 12801
rect 14280 12656 14332 12708
rect 15568 12656 15620 12708
rect 18144 12903 18196 12912
rect 18144 12869 18178 12903
rect 18178 12869 18196 12903
rect 18144 12860 18196 12869
rect 18696 12860 18748 12912
rect 17776 12792 17828 12844
rect 21548 12928 21600 12980
rect 21640 12860 21692 12912
rect 21180 12792 21232 12844
rect 10048 12631 10100 12640
rect 10048 12597 10057 12631
rect 10057 12597 10091 12631
rect 10091 12597 10100 12631
rect 10048 12588 10100 12597
rect 10508 12588 10560 12640
rect 11796 12631 11848 12640
rect 11796 12597 11805 12631
rect 11805 12597 11839 12631
rect 11839 12597 11848 12631
rect 11796 12588 11848 12597
rect 12624 12588 12676 12640
rect 14464 12631 14516 12640
rect 14464 12597 14473 12631
rect 14473 12597 14507 12631
rect 14507 12597 14516 12631
rect 14464 12588 14516 12597
rect 14648 12588 14700 12640
rect 15016 12588 15068 12640
rect 16120 12588 16172 12640
rect 17776 12631 17828 12640
rect 17776 12597 17785 12631
rect 17785 12597 17819 12631
rect 17819 12597 17828 12631
rect 17776 12588 17828 12597
rect 20720 12724 20772 12776
rect 18972 12656 19024 12708
rect 21088 12656 21140 12708
rect 21364 12656 21416 12708
rect 19064 12588 19116 12640
rect 19708 12631 19760 12640
rect 19708 12597 19717 12631
rect 19717 12597 19751 12631
rect 19751 12597 19760 12631
rect 19708 12588 19760 12597
rect 20260 12631 20312 12640
rect 20260 12597 20269 12631
rect 20269 12597 20303 12631
rect 20303 12597 20312 12631
rect 20260 12588 20312 12597
rect 20996 12631 21048 12640
rect 20996 12597 21005 12631
rect 21005 12597 21039 12631
rect 21039 12597 21048 12631
rect 20996 12588 21048 12597
rect 21456 12631 21508 12640
rect 21456 12597 21465 12631
rect 21465 12597 21499 12631
rect 21499 12597 21508 12631
rect 21456 12588 21508 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1768 12384 1820 12436
rect 2688 12384 2740 12436
rect 3240 12427 3292 12436
rect 3240 12393 3249 12427
rect 3249 12393 3283 12427
rect 3283 12393 3292 12427
rect 3240 12384 3292 12393
rect 4068 12384 4120 12436
rect 5080 12384 5132 12436
rect 5356 12427 5408 12436
rect 5356 12393 5365 12427
rect 5365 12393 5399 12427
rect 5399 12393 5408 12427
rect 5356 12384 5408 12393
rect 3056 12316 3108 12368
rect 3976 12248 4028 12300
rect 4620 12316 4672 12368
rect 7012 12384 7064 12436
rect 7196 12427 7248 12436
rect 7196 12393 7205 12427
rect 7205 12393 7239 12427
rect 7239 12393 7248 12427
rect 7196 12384 7248 12393
rect 7288 12384 7340 12436
rect 8116 12384 8168 12436
rect 9220 12384 9272 12436
rect 10324 12384 10376 12436
rect 11704 12384 11756 12436
rect 1308 12180 1360 12232
rect 2412 12112 2464 12164
rect 2504 12112 2556 12164
rect 2872 12180 2924 12232
rect 3884 12180 3936 12232
rect 4252 12180 4304 12232
rect 4528 12112 4580 12164
rect 4988 12112 5040 12164
rect 5724 12248 5776 12300
rect 6000 12248 6052 12300
rect 7196 12248 7248 12300
rect 8484 12291 8536 12300
rect 8484 12257 8493 12291
rect 8493 12257 8527 12291
rect 8527 12257 8536 12291
rect 8484 12248 8536 12257
rect 12164 12384 12216 12436
rect 14372 12384 14424 12436
rect 12072 12316 12124 12368
rect 12256 12316 12308 12368
rect 10416 12291 10468 12300
rect 10416 12257 10425 12291
rect 10425 12257 10459 12291
rect 10459 12257 10468 12291
rect 10416 12248 10468 12257
rect 11796 12248 11848 12300
rect 12164 12248 12216 12300
rect 5908 12180 5960 12232
rect 6736 12223 6788 12232
rect 6736 12189 6754 12223
rect 6754 12189 6788 12223
rect 6736 12180 6788 12189
rect 7104 12180 7156 12232
rect 9772 12180 9824 12232
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 1676 12044 1728 12096
rect 4620 12044 4672 12096
rect 4896 12087 4948 12096
rect 4896 12053 4905 12087
rect 4905 12053 4939 12087
rect 4939 12053 4948 12087
rect 4896 12044 4948 12053
rect 5356 12044 5408 12096
rect 6000 12044 6052 12096
rect 6828 12112 6880 12164
rect 7380 12044 7432 12096
rect 7656 12087 7708 12096
rect 7656 12053 7665 12087
rect 7665 12053 7699 12087
rect 7699 12053 7708 12087
rect 7656 12044 7708 12053
rect 8852 12044 8904 12096
rect 9128 12112 9180 12164
rect 10508 12180 10560 12232
rect 10968 12180 11020 12232
rect 11888 12180 11940 12232
rect 12532 12180 12584 12232
rect 11152 12112 11204 12164
rect 11612 12112 11664 12164
rect 12992 12316 13044 12368
rect 13636 12316 13688 12368
rect 15752 12384 15804 12436
rect 15844 12384 15896 12436
rect 16396 12384 16448 12436
rect 17224 12384 17276 12436
rect 18880 12384 18932 12436
rect 20536 12384 20588 12436
rect 20628 12384 20680 12436
rect 21272 12384 21324 12436
rect 16120 12316 16172 12368
rect 17316 12316 17368 12368
rect 13728 12248 13780 12300
rect 16580 12291 16632 12300
rect 16580 12257 16589 12291
rect 16589 12257 16623 12291
rect 16623 12257 16632 12291
rect 16580 12248 16632 12257
rect 17040 12248 17092 12300
rect 17408 12248 17460 12300
rect 17684 12291 17736 12300
rect 17684 12257 17693 12291
rect 17693 12257 17727 12291
rect 17727 12257 17736 12291
rect 17684 12248 17736 12257
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 14372 12180 14424 12232
rect 15384 12180 15436 12232
rect 16304 12180 16356 12232
rect 16396 12180 16448 12232
rect 9956 12044 10008 12096
rect 10508 12044 10560 12096
rect 11244 12044 11296 12096
rect 12348 12087 12400 12096
rect 12348 12053 12357 12087
rect 12357 12053 12391 12087
rect 12391 12053 12400 12087
rect 12348 12044 12400 12053
rect 13544 12044 13596 12096
rect 14096 12087 14148 12096
rect 14096 12053 14105 12087
rect 14105 12053 14139 12087
rect 14139 12053 14148 12087
rect 14096 12044 14148 12053
rect 14464 12044 14516 12096
rect 14740 12112 14792 12164
rect 16672 12112 16724 12164
rect 16764 12112 16816 12164
rect 16948 12155 17000 12164
rect 16948 12121 16957 12155
rect 16957 12121 16991 12155
rect 16991 12121 17000 12155
rect 16948 12112 17000 12121
rect 17684 12112 17736 12164
rect 18236 12112 18288 12164
rect 15292 12044 15344 12096
rect 15660 12044 15712 12096
rect 16212 12087 16264 12096
rect 16212 12053 16221 12087
rect 16221 12053 16255 12087
rect 16255 12053 16264 12087
rect 16212 12044 16264 12053
rect 17224 12087 17276 12096
rect 17224 12053 17233 12087
rect 17233 12053 17267 12087
rect 17267 12053 17276 12087
rect 17224 12044 17276 12053
rect 17500 12087 17552 12096
rect 17500 12053 17509 12087
rect 17509 12053 17543 12087
rect 17543 12053 17552 12087
rect 17500 12044 17552 12053
rect 18144 12044 18196 12096
rect 19248 12248 19300 12300
rect 19616 12155 19668 12164
rect 19616 12121 19625 12155
rect 19625 12121 19659 12155
rect 19659 12121 19668 12155
rect 19616 12112 19668 12121
rect 19708 12155 19760 12164
rect 19708 12121 19717 12155
rect 19717 12121 19751 12155
rect 19751 12121 19760 12155
rect 20812 12316 20864 12368
rect 19984 12248 20036 12300
rect 21088 12248 21140 12300
rect 21548 12248 21600 12300
rect 22192 12248 22244 12300
rect 19708 12112 19760 12121
rect 19156 12044 19208 12096
rect 20260 12112 20312 12164
rect 20352 12112 20404 12164
rect 21456 12180 21508 12232
rect 21548 12112 21600 12164
rect 20536 12087 20588 12096
rect 20536 12053 20545 12087
rect 20545 12053 20579 12087
rect 20579 12053 20588 12087
rect 20536 12044 20588 12053
rect 21088 12044 21140 12096
rect 21456 12087 21508 12096
rect 21456 12053 21465 12087
rect 21465 12053 21499 12087
rect 21499 12053 21508 12087
rect 21456 12044 21508 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 1676 11840 1728 11892
rect 3056 11840 3108 11892
rect 4160 11840 4212 11892
rect 5264 11840 5316 11892
rect 1860 11704 1912 11756
rect 2136 11704 2188 11756
rect 2412 11500 2464 11552
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 4252 11704 4304 11756
rect 4620 11747 4672 11756
rect 4620 11713 4629 11747
rect 4629 11713 4663 11747
rect 4663 11713 4672 11747
rect 4620 11704 4672 11713
rect 5264 11704 5316 11756
rect 5908 11815 5960 11824
rect 5908 11781 5917 11815
rect 5917 11781 5951 11815
rect 5951 11781 5960 11815
rect 5908 11772 5960 11781
rect 5816 11747 5868 11756
rect 4068 11679 4120 11688
rect 4068 11645 4077 11679
rect 4077 11645 4111 11679
rect 4111 11645 4120 11679
rect 4068 11636 4120 11645
rect 4160 11679 4212 11688
rect 4160 11645 4169 11679
rect 4169 11645 4203 11679
rect 4203 11645 4212 11679
rect 4160 11636 4212 11645
rect 4988 11636 5040 11688
rect 5816 11713 5825 11747
rect 5825 11713 5859 11747
rect 5859 11713 5868 11747
rect 5816 11704 5868 11713
rect 6000 11704 6052 11756
rect 6368 11772 6420 11824
rect 6736 11772 6788 11824
rect 7288 11840 7340 11892
rect 7656 11840 7708 11892
rect 8852 11883 8904 11892
rect 8852 11849 8861 11883
rect 8861 11849 8895 11883
rect 8895 11849 8904 11883
rect 8852 11840 8904 11849
rect 10324 11883 10376 11892
rect 7104 11772 7156 11824
rect 5540 11636 5592 11688
rect 5908 11636 5960 11688
rect 6644 11704 6696 11756
rect 7196 11704 7248 11756
rect 8668 11772 8720 11824
rect 8760 11772 8812 11824
rect 10048 11772 10100 11824
rect 10324 11849 10333 11883
rect 10333 11849 10367 11883
rect 10367 11849 10376 11883
rect 10324 11840 10376 11849
rect 12348 11840 12400 11892
rect 8392 11747 8444 11756
rect 8392 11713 8401 11747
rect 8401 11713 8435 11747
rect 8435 11713 8444 11747
rect 8392 11704 8444 11713
rect 9036 11704 9088 11756
rect 9128 11636 9180 11688
rect 10416 11704 10468 11756
rect 10232 11636 10284 11688
rect 4528 11500 4580 11552
rect 4712 11543 4764 11552
rect 4712 11509 4721 11543
rect 4721 11509 4755 11543
rect 4755 11509 4764 11543
rect 4712 11500 4764 11509
rect 5080 11500 5132 11552
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 10140 11543 10192 11552
rect 10140 11509 10149 11543
rect 10149 11509 10183 11543
rect 10183 11509 10192 11543
rect 10140 11500 10192 11509
rect 11152 11568 11204 11620
rect 11888 11704 11940 11756
rect 12072 11704 12124 11756
rect 11704 11636 11756 11688
rect 12348 11704 12400 11756
rect 12808 11840 12860 11892
rect 15200 11840 15252 11892
rect 15752 11840 15804 11892
rect 15936 11772 15988 11824
rect 16304 11772 16356 11824
rect 17592 11772 17644 11824
rect 18236 11840 18288 11892
rect 18512 11840 18564 11892
rect 19340 11883 19392 11892
rect 19340 11849 19349 11883
rect 19349 11849 19383 11883
rect 19383 11849 19392 11883
rect 19340 11840 19392 11849
rect 19524 11840 19576 11892
rect 20352 11883 20404 11892
rect 20352 11849 20361 11883
rect 20361 11849 20395 11883
rect 20395 11849 20404 11883
rect 20352 11840 20404 11849
rect 20628 11883 20680 11892
rect 20628 11849 20637 11883
rect 20637 11849 20671 11883
rect 20671 11849 20680 11883
rect 20628 11840 20680 11849
rect 21456 11772 21508 11824
rect 12808 11704 12860 11756
rect 13544 11704 13596 11756
rect 14924 11747 14976 11756
rect 14924 11713 14953 11747
rect 14953 11713 14976 11747
rect 14924 11704 14976 11713
rect 15108 11704 15160 11756
rect 15384 11704 15436 11756
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 16488 11704 16540 11756
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 17960 11704 18012 11756
rect 18512 11747 18564 11756
rect 18512 11713 18521 11747
rect 18521 11713 18555 11747
rect 18555 11713 18564 11747
rect 18512 11704 18564 11713
rect 19800 11704 19852 11756
rect 20352 11704 20404 11756
rect 20444 11747 20496 11756
rect 20444 11713 20453 11747
rect 20453 11713 20487 11747
rect 20487 11713 20496 11747
rect 20444 11704 20496 11713
rect 12348 11568 12400 11620
rect 13452 11636 13504 11688
rect 15844 11679 15896 11688
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 13636 11568 13688 11620
rect 13544 11500 13596 11552
rect 13728 11543 13780 11552
rect 13728 11509 13737 11543
rect 13737 11509 13771 11543
rect 13771 11509 13780 11543
rect 13728 11500 13780 11509
rect 15844 11645 15853 11679
rect 15853 11645 15887 11679
rect 15887 11645 15896 11679
rect 15844 11636 15896 11645
rect 18236 11679 18288 11688
rect 18236 11645 18245 11679
rect 18245 11645 18279 11679
rect 18279 11645 18288 11679
rect 18236 11636 18288 11645
rect 18420 11679 18472 11688
rect 18420 11645 18429 11679
rect 18429 11645 18463 11679
rect 18463 11645 18472 11679
rect 18420 11636 18472 11645
rect 19156 11636 19208 11688
rect 19248 11636 19300 11688
rect 21548 11679 21600 11688
rect 21548 11645 21557 11679
rect 21557 11645 21591 11679
rect 21591 11645 21600 11679
rect 21548 11636 21600 11645
rect 17408 11500 17460 11552
rect 20628 11568 20680 11620
rect 20812 11568 20864 11620
rect 22744 11568 22796 11620
rect 19892 11500 19944 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2872 11296 2924 11348
rect 3976 11296 4028 11348
rect 4068 11296 4120 11348
rect 1768 11228 1820 11280
rect 5816 11271 5868 11280
rect 5816 11237 5825 11271
rect 5825 11237 5859 11271
rect 5859 11237 5868 11271
rect 5816 11228 5868 11237
rect 1676 11203 1728 11212
rect 1676 11169 1685 11203
rect 1685 11169 1719 11203
rect 1719 11169 1728 11203
rect 1676 11160 1728 11169
rect 2228 11203 2280 11212
rect 2228 11169 2237 11203
rect 2237 11169 2271 11203
rect 2271 11169 2280 11203
rect 2228 11160 2280 11169
rect 4068 11160 4120 11212
rect 4712 11160 4764 11212
rect 4896 11160 4948 11212
rect 3792 11135 3844 11144
rect 3792 11101 3801 11135
rect 3801 11101 3835 11135
rect 3835 11101 3844 11135
rect 3792 11092 3844 11101
rect 4988 11092 5040 11144
rect 5264 11160 5316 11212
rect 8668 11296 8720 11348
rect 9864 11339 9916 11348
rect 9864 11305 9873 11339
rect 9873 11305 9907 11339
rect 9907 11305 9916 11339
rect 9864 11296 9916 11305
rect 11244 11296 11296 11348
rect 11704 11339 11756 11348
rect 11704 11305 11713 11339
rect 11713 11305 11747 11339
rect 11747 11305 11756 11339
rect 11704 11296 11756 11305
rect 12348 11296 12400 11348
rect 12808 11296 12860 11348
rect 13176 11296 13228 11348
rect 13544 11296 13596 11348
rect 15016 11339 15068 11348
rect 15016 11305 15025 11339
rect 15025 11305 15059 11339
rect 15059 11305 15068 11339
rect 15016 11296 15068 11305
rect 15200 11296 15252 11348
rect 16120 11296 16172 11348
rect 9956 11271 10008 11280
rect 9956 11237 9965 11271
rect 9965 11237 9999 11271
rect 9999 11237 10008 11271
rect 9956 11228 10008 11237
rect 10600 11228 10652 11280
rect 10784 11228 10836 11280
rect 6000 11160 6052 11212
rect 6368 11203 6420 11212
rect 6368 11169 6377 11203
rect 6377 11169 6411 11203
rect 6411 11169 6420 11203
rect 6368 11160 6420 11169
rect 7748 11160 7800 11212
rect 10048 11160 10100 11212
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 11888 11203 11940 11212
rect 11888 11169 11897 11203
rect 11897 11169 11931 11203
rect 11931 11169 11940 11203
rect 11888 11160 11940 11169
rect 12256 11228 12308 11280
rect 13360 11228 13412 11280
rect 14372 11228 14424 11280
rect 14740 11228 14792 11280
rect 15292 11228 15344 11280
rect 15844 11228 15896 11280
rect 16672 11296 16724 11348
rect 18420 11296 18472 11348
rect 5816 11092 5868 11144
rect 3424 11024 3476 11076
rect 4160 11024 4212 11076
rect 5080 11024 5132 11076
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6736 11135 6788 11144
rect 6276 11092 6328 11101
rect 6736 11101 6745 11135
rect 6745 11101 6779 11135
rect 6779 11101 6788 11135
rect 6736 11092 6788 11101
rect 9220 11092 9272 11144
rect 10968 11092 11020 11144
rect 1768 10999 1820 11008
rect 1768 10965 1777 10999
rect 1777 10965 1811 10999
rect 1811 10965 1820 10999
rect 1768 10956 1820 10965
rect 2964 10956 3016 11008
rect 5264 10999 5316 11008
rect 5264 10965 5273 10999
rect 5273 10965 5307 10999
rect 5307 10965 5316 10999
rect 5264 10956 5316 10965
rect 5632 10956 5684 11008
rect 7380 11024 7432 11076
rect 9128 11024 9180 11076
rect 8116 10999 8168 11008
rect 8116 10965 8125 10999
rect 8125 10965 8159 10999
rect 8159 10965 8168 10999
rect 8116 10956 8168 10965
rect 8484 10956 8536 11008
rect 9312 10956 9364 11008
rect 9956 11024 10008 11076
rect 12992 11092 13044 11144
rect 10600 10956 10652 11008
rect 11244 10999 11296 11008
rect 11244 10965 11253 10999
rect 11253 10965 11287 10999
rect 11287 10965 11296 10999
rect 11796 11024 11848 11076
rect 11888 11024 11940 11076
rect 12624 11024 12676 11076
rect 13544 11203 13596 11212
rect 13544 11169 13553 11203
rect 13553 11169 13587 11203
rect 13587 11169 13596 11203
rect 13820 11203 13872 11212
rect 13544 11160 13596 11169
rect 13820 11169 13829 11203
rect 13829 11169 13863 11203
rect 13863 11169 13872 11203
rect 13820 11160 13872 11169
rect 13912 11160 13964 11212
rect 14924 11160 14976 11212
rect 15752 11160 15804 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 20168 11296 20220 11348
rect 20352 11339 20404 11348
rect 20352 11305 20361 11339
rect 20361 11305 20395 11339
rect 20395 11305 20404 11339
rect 20352 11296 20404 11305
rect 20628 11296 20680 11348
rect 21456 11296 21508 11348
rect 19708 11228 19760 11280
rect 20260 11271 20312 11280
rect 20260 11237 20269 11271
rect 20269 11237 20303 11271
rect 20303 11237 20312 11271
rect 20260 11228 20312 11237
rect 20812 11271 20864 11280
rect 20812 11237 20821 11271
rect 20821 11237 20855 11271
rect 20855 11237 20864 11271
rect 20812 11228 20864 11237
rect 19524 11160 19576 11212
rect 20168 11160 20220 11212
rect 13728 11092 13780 11144
rect 15200 11135 15252 11144
rect 15200 11101 15209 11135
rect 15209 11101 15243 11135
rect 15243 11101 15252 11135
rect 16120 11135 16172 11144
rect 15200 11092 15252 11101
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 17500 11092 17552 11144
rect 17776 11092 17828 11144
rect 19340 11092 19392 11144
rect 11244 10956 11296 10965
rect 13912 10956 13964 11008
rect 15016 11024 15068 11076
rect 16396 11024 16448 11076
rect 16948 11024 17000 11076
rect 17316 11024 17368 11076
rect 20352 11024 20404 11076
rect 20904 11092 20956 11144
rect 21456 11135 21508 11144
rect 21456 11101 21465 11135
rect 21465 11101 21499 11135
rect 21499 11101 21508 11135
rect 21456 11092 21508 11101
rect 21088 11067 21140 11076
rect 21088 11033 21097 11067
rect 21097 11033 21131 11067
rect 21131 11033 21140 11067
rect 21088 11024 21140 11033
rect 15292 10956 15344 11008
rect 15660 10956 15712 11008
rect 15752 10999 15804 11008
rect 15752 10965 15761 10999
rect 15761 10965 15795 10999
rect 15795 10965 15804 10999
rect 15752 10956 15804 10965
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 18052 10999 18104 11008
rect 15936 10956 15988 10965
rect 18052 10965 18061 10999
rect 18061 10965 18095 10999
rect 18095 10965 18104 10999
rect 18052 10956 18104 10965
rect 18788 10999 18840 11008
rect 18788 10965 18797 10999
rect 18797 10965 18831 10999
rect 18831 10965 18840 10999
rect 18788 10956 18840 10965
rect 19616 10956 19668 11008
rect 20628 10956 20680 11008
rect 20812 10956 20864 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 388 10752 440 10804
rect 3148 10752 3200 10804
rect 4068 10752 4120 10804
rect 5632 10752 5684 10804
rect 1492 10727 1544 10736
rect 1492 10693 1501 10727
rect 1501 10693 1535 10727
rect 1535 10693 1544 10727
rect 1492 10684 1544 10693
rect 2228 10684 2280 10736
rect 2688 10684 2740 10736
rect 3976 10684 4028 10736
rect 1860 10616 1912 10668
rect 4344 10616 4396 10668
rect 4988 10684 5040 10736
rect 5816 10684 5868 10736
rect 7288 10752 7340 10804
rect 7748 10752 7800 10804
rect 8024 10752 8076 10804
rect 4712 10591 4764 10600
rect 1952 10412 2004 10464
rect 2504 10412 2556 10464
rect 3332 10412 3384 10464
rect 4712 10557 4721 10591
rect 4721 10557 4755 10591
rect 4755 10557 4764 10591
rect 4712 10548 4764 10557
rect 4896 10591 4948 10600
rect 4896 10557 4905 10591
rect 4905 10557 4939 10591
rect 4939 10557 4948 10591
rect 4896 10548 4948 10557
rect 5172 10548 5224 10600
rect 7196 10684 7248 10736
rect 10232 10752 10284 10804
rect 8576 10684 8628 10736
rect 10324 10684 10376 10736
rect 11152 10752 11204 10804
rect 11888 10752 11940 10804
rect 12072 10752 12124 10804
rect 12992 10684 13044 10736
rect 15936 10752 15988 10804
rect 16120 10752 16172 10804
rect 18052 10752 18104 10804
rect 18512 10752 18564 10804
rect 19524 10795 19576 10804
rect 19524 10761 19533 10795
rect 19533 10761 19567 10795
rect 19567 10761 19576 10795
rect 19524 10752 19576 10761
rect 20352 10795 20404 10804
rect 13544 10684 13596 10736
rect 13728 10684 13780 10736
rect 15292 10684 15344 10736
rect 15568 10684 15620 10736
rect 15752 10684 15804 10736
rect 20352 10761 20361 10795
rect 20361 10761 20395 10795
rect 20395 10761 20404 10795
rect 20352 10752 20404 10761
rect 20628 10752 20680 10804
rect 4252 10523 4304 10532
rect 4252 10489 4261 10523
rect 4261 10489 4295 10523
rect 4295 10489 4304 10523
rect 4252 10480 4304 10489
rect 4528 10480 4580 10532
rect 6000 10480 6052 10532
rect 7196 10548 7248 10600
rect 7840 10548 7892 10600
rect 8116 10548 8168 10600
rect 7472 10480 7524 10532
rect 8024 10480 8076 10532
rect 9220 10548 9272 10600
rect 10508 10616 10560 10668
rect 10600 10616 10652 10668
rect 12532 10616 12584 10668
rect 9680 10548 9732 10600
rect 10968 10548 11020 10600
rect 12808 10548 12860 10600
rect 9864 10480 9916 10532
rect 11888 10480 11940 10532
rect 13268 10616 13320 10668
rect 14372 10659 14424 10668
rect 14372 10625 14381 10659
rect 14381 10625 14415 10659
rect 14415 10625 14424 10659
rect 17868 10659 17920 10668
rect 14372 10616 14424 10625
rect 17868 10625 17877 10659
rect 17877 10625 17911 10659
rect 17911 10625 17920 10659
rect 17868 10616 17920 10625
rect 13912 10591 13964 10600
rect 13912 10557 13921 10591
rect 13921 10557 13955 10591
rect 13955 10557 13964 10591
rect 13912 10548 13964 10557
rect 14004 10548 14056 10600
rect 14924 10548 14976 10600
rect 15384 10591 15436 10600
rect 15384 10557 15393 10591
rect 15393 10557 15427 10591
rect 15427 10557 15436 10591
rect 15384 10548 15436 10557
rect 16028 10480 16080 10532
rect 4896 10412 4948 10464
rect 5264 10412 5316 10464
rect 5632 10412 5684 10464
rect 7840 10455 7892 10464
rect 7840 10421 7849 10455
rect 7849 10421 7883 10455
rect 7883 10421 7892 10455
rect 7840 10412 7892 10421
rect 9128 10412 9180 10464
rect 10324 10412 10376 10464
rect 12072 10455 12124 10464
rect 12072 10421 12081 10455
rect 12081 10421 12115 10455
rect 12115 10421 12124 10455
rect 12072 10412 12124 10421
rect 12164 10455 12216 10464
rect 12164 10421 12173 10455
rect 12173 10421 12207 10455
rect 12207 10421 12216 10455
rect 12164 10412 12216 10421
rect 13268 10412 13320 10464
rect 15108 10412 15160 10464
rect 16948 10548 17000 10600
rect 17960 10548 18012 10600
rect 18972 10548 19024 10600
rect 19708 10591 19760 10600
rect 19708 10557 19717 10591
rect 19717 10557 19751 10591
rect 19751 10557 19760 10591
rect 20904 10616 20956 10668
rect 22192 10616 22244 10668
rect 22560 10616 22612 10668
rect 19708 10548 19760 10557
rect 21548 10548 21600 10600
rect 18236 10480 18288 10532
rect 19616 10412 19668 10464
rect 20720 10412 20772 10464
rect 21272 10412 21324 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1768 10208 1820 10260
rect 3976 10251 4028 10260
rect 3976 10217 3985 10251
rect 3985 10217 4019 10251
rect 4019 10217 4028 10251
rect 3976 10208 4028 10217
rect 4988 10208 5040 10260
rect 5172 10251 5224 10260
rect 5172 10217 5181 10251
rect 5181 10217 5215 10251
rect 5215 10217 5224 10251
rect 5172 10208 5224 10217
rect 5264 10208 5316 10260
rect 2504 10115 2556 10124
rect 2504 10081 2513 10115
rect 2513 10081 2547 10115
rect 2547 10081 2556 10115
rect 2504 10072 2556 10081
rect 4712 10140 4764 10192
rect 5448 10140 5500 10192
rect 6920 10208 6972 10260
rect 7380 10140 7432 10192
rect 3424 10072 3476 10124
rect 2780 10004 2832 10056
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 2228 9911 2280 9920
rect 2228 9877 2237 9911
rect 2237 9877 2271 9911
rect 2271 9877 2280 9911
rect 2228 9868 2280 9877
rect 2320 9911 2372 9920
rect 2320 9877 2329 9911
rect 2329 9877 2363 9911
rect 2363 9877 2372 9911
rect 2688 9911 2740 9920
rect 2320 9868 2372 9877
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 2780 9868 2832 9920
rect 2964 9868 3016 9920
rect 3332 9868 3384 9920
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 4252 10047 4304 10056
rect 4252 10013 4261 10047
rect 4261 10013 4295 10047
rect 4295 10013 4304 10047
rect 4252 10004 4304 10013
rect 4896 10072 4948 10124
rect 6000 10072 6052 10124
rect 7104 10072 7156 10124
rect 9128 10208 9180 10260
rect 10508 10251 10560 10260
rect 10508 10217 10517 10251
rect 10517 10217 10551 10251
rect 10551 10217 10560 10251
rect 10508 10208 10560 10217
rect 10784 10208 10836 10260
rect 11980 10208 12032 10260
rect 8852 10140 8904 10192
rect 10600 10183 10652 10192
rect 10600 10149 10609 10183
rect 10609 10149 10643 10183
rect 10643 10149 10652 10183
rect 10600 10140 10652 10149
rect 11796 10183 11848 10192
rect 11796 10149 11805 10183
rect 11805 10149 11839 10183
rect 11839 10149 11848 10183
rect 13636 10208 13688 10260
rect 14372 10208 14424 10260
rect 14924 10251 14976 10260
rect 14924 10217 14933 10251
rect 14933 10217 14967 10251
rect 14967 10217 14976 10251
rect 14924 10208 14976 10217
rect 15752 10208 15804 10260
rect 15936 10208 15988 10260
rect 16120 10208 16172 10260
rect 17316 10251 17368 10260
rect 17316 10217 17325 10251
rect 17325 10217 17359 10251
rect 17359 10217 17368 10251
rect 17316 10208 17368 10217
rect 11796 10140 11848 10149
rect 13820 10140 13872 10192
rect 14188 10140 14240 10192
rect 14556 10140 14608 10192
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 6920 10047 6972 10056
rect 6920 10013 6929 10047
rect 6929 10013 6963 10047
rect 6963 10013 6972 10047
rect 6920 10004 6972 10013
rect 8116 10047 8168 10056
rect 8116 10013 8134 10047
rect 8134 10013 8168 10047
rect 8116 10004 8168 10013
rect 8300 10004 8352 10056
rect 10140 10072 10192 10124
rect 12256 10115 12308 10124
rect 12256 10081 12265 10115
rect 12265 10081 12299 10115
rect 12299 10081 12308 10115
rect 12256 10072 12308 10081
rect 13360 10072 13412 10124
rect 13636 10072 13688 10124
rect 13728 10072 13780 10124
rect 15384 10140 15436 10192
rect 15108 10072 15160 10124
rect 15936 10115 15988 10124
rect 15936 10081 15945 10115
rect 15945 10081 15979 10115
rect 15979 10081 15988 10115
rect 15936 10072 15988 10081
rect 16212 10072 16264 10124
rect 16948 10140 17000 10192
rect 19708 10208 19760 10260
rect 20536 10208 20588 10260
rect 18972 10183 19024 10192
rect 18972 10149 18981 10183
rect 18981 10149 19015 10183
rect 19015 10149 19024 10183
rect 18972 10140 19024 10149
rect 19800 10140 19852 10192
rect 20996 10183 21048 10192
rect 20996 10149 21005 10183
rect 21005 10149 21039 10183
rect 21039 10149 21048 10183
rect 20996 10140 21048 10149
rect 17500 10115 17552 10124
rect 17500 10081 17509 10115
rect 17509 10081 17543 10115
rect 17543 10081 17552 10115
rect 17500 10072 17552 10081
rect 18788 10072 18840 10124
rect 19708 10072 19760 10124
rect 21088 10072 21140 10124
rect 3608 9936 3660 9988
rect 4068 9868 4120 9920
rect 4528 9868 4580 9920
rect 4712 9911 4764 9920
rect 4712 9877 4721 9911
rect 4721 9877 4755 9911
rect 4755 9877 4764 9911
rect 4712 9868 4764 9877
rect 5172 9868 5224 9920
rect 5356 9936 5408 9988
rect 7380 9936 7432 9988
rect 8392 9936 8444 9988
rect 5540 9911 5592 9920
rect 5540 9877 5549 9911
rect 5549 9877 5583 9911
rect 5583 9877 5592 9911
rect 5540 9868 5592 9877
rect 5908 9911 5960 9920
rect 5908 9877 5917 9911
rect 5917 9877 5951 9911
rect 5951 9877 5960 9911
rect 5908 9868 5960 9877
rect 6644 9868 6696 9920
rect 7104 9868 7156 9920
rect 7932 9868 7984 9920
rect 8576 9911 8628 9920
rect 8576 9877 8585 9911
rect 8585 9877 8619 9911
rect 8619 9877 8628 9911
rect 8576 9868 8628 9877
rect 8944 9868 8996 9920
rect 9680 10004 9732 10056
rect 9864 10004 9916 10056
rect 9128 9936 9180 9988
rect 10876 9936 10928 9988
rect 13544 10004 13596 10056
rect 14004 10004 14056 10056
rect 15384 10004 15436 10056
rect 16396 10004 16448 10056
rect 16948 10004 17000 10056
rect 18052 10004 18104 10056
rect 19432 10047 19484 10056
rect 19432 10013 19441 10047
rect 19441 10013 19475 10047
rect 19475 10013 19484 10047
rect 19432 10004 19484 10013
rect 21180 10047 21232 10056
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 21456 10047 21508 10056
rect 21456 10013 21465 10047
rect 21465 10013 21499 10047
rect 21499 10013 21508 10047
rect 21456 10004 21508 10013
rect 15752 9936 15804 9988
rect 16212 9936 16264 9988
rect 16304 9936 16356 9988
rect 9588 9868 9640 9920
rect 9680 9868 9732 9920
rect 10048 9868 10100 9920
rect 10784 9868 10836 9920
rect 11060 9911 11112 9920
rect 11060 9877 11069 9911
rect 11069 9877 11103 9911
rect 11103 9877 11112 9911
rect 11060 9868 11112 9877
rect 11796 9868 11848 9920
rect 13176 9868 13228 9920
rect 14188 9868 14240 9920
rect 14556 9911 14608 9920
rect 14556 9877 14565 9911
rect 14565 9877 14599 9911
rect 14599 9877 14608 9911
rect 14556 9868 14608 9877
rect 14924 9868 14976 9920
rect 15292 9911 15344 9920
rect 15292 9877 15301 9911
rect 15301 9877 15335 9911
rect 15335 9877 15344 9911
rect 15292 9868 15344 9877
rect 15568 9868 15620 9920
rect 15660 9868 15712 9920
rect 16396 9868 16448 9920
rect 20536 9936 20588 9988
rect 20812 9936 20864 9988
rect 18236 9868 18288 9920
rect 20352 9868 20404 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 2320 9664 2372 9716
rect 2688 9664 2740 9716
rect 2964 9664 3016 9716
rect 3792 9664 3844 9716
rect 4344 9664 4396 9716
rect 4712 9664 4764 9716
rect 4896 9707 4948 9716
rect 4896 9673 4905 9707
rect 4905 9673 4939 9707
rect 4939 9673 4948 9707
rect 4896 9664 4948 9673
rect 4988 9664 5040 9716
rect 5356 9664 5408 9716
rect 5816 9707 5868 9716
rect 5816 9673 5825 9707
rect 5825 9673 5859 9707
rect 5859 9673 5868 9707
rect 5816 9664 5868 9673
rect 5908 9664 5960 9716
rect 7840 9664 7892 9716
rect 1308 9596 1360 9648
rect 1676 9596 1728 9648
rect 3700 9596 3752 9648
rect 848 9460 900 9512
rect 1032 9460 1084 9512
rect 2872 9528 2924 9580
rect 9496 9664 9548 9716
rect 1860 9460 1912 9512
rect 2688 9503 2740 9512
rect 2688 9469 2697 9503
rect 2697 9469 2731 9503
rect 2731 9469 2740 9503
rect 2688 9460 2740 9469
rect 1952 9435 2004 9444
rect 1952 9401 1961 9435
rect 1961 9401 1995 9435
rect 1995 9401 2004 9435
rect 1952 9392 2004 9401
rect 2320 9392 2372 9444
rect 2412 9392 2464 9444
rect 4252 9528 4304 9580
rect 4436 9528 4488 9580
rect 1400 9324 1452 9376
rect 2136 9324 2188 9376
rect 3240 9324 3292 9376
rect 4712 9460 4764 9512
rect 5080 9503 5132 9512
rect 5080 9469 5089 9503
rect 5089 9469 5123 9503
rect 5123 9469 5132 9503
rect 5448 9528 5500 9580
rect 5080 9460 5132 9469
rect 6460 9528 6512 9580
rect 8392 9596 8444 9648
rect 10416 9664 10468 9716
rect 10600 9664 10652 9716
rect 11980 9664 12032 9716
rect 12716 9664 12768 9716
rect 14556 9707 14608 9716
rect 9956 9596 10008 9648
rect 14556 9673 14565 9707
rect 14565 9673 14599 9707
rect 14599 9673 14608 9707
rect 14556 9664 14608 9673
rect 15016 9707 15068 9716
rect 15016 9673 15025 9707
rect 15025 9673 15059 9707
rect 15059 9673 15068 9707
rect 15016 9664 15068 9673
rect 15384 9707 15436 9716
rect 15384 9673 15393 9707
rect 15393 9673 15427 9707
rect 15427 9673 15436 9707
rect 15384 9664 15436 9673
rect 15660 9707 15712 9716
rect 15660 9673 15669 9707
rect 15669 9673 15703 9707
rect 15703 9673 15712 9707
rect 15660 9664 15712 9673
rect 16212 9664 16264 9716
rect 16948 9664 17000 9716
rect 17868 9664 17920 9716
rect 19524 9664 19576 9716
rect 20536 9664 20588 9716
rect 8852 9571 8904 9580
rect 3700 9392 3752 9444
rect 4436 9392 4488 9444
rect 4252 9324 4304 9376
rect 4896 9324 4948 9376
rect 5172 9392 5224 9444
rect 5724 9392 5776 9444
rect 6920 9460 6972 9512
rect 7472 9503 7524 9512
rect 7472 9469 7481 9503
rect 7481 9469 7515 9503
rect 7515 9469 7524 9503
rect 7472 9460 7524 9469
rect 7932 9460 7984 9512
rect 8116 9460 8168 9512
rect 6000 9392 6052 9444
rect 8300 9392 8352 9444
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 10140 9528 10192 9580
rect 12256 9528 12308 9580
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 13544 9528 13596 9580
rect 13636 9528 13688 9580
rect 10416 9503 10468 9512
rect 10416 9469 10425 9503
rect 10425 9469 10459 9503
rect 10459 9469 10468 9503
rect 10416 9460 10468 9469
rect 10600 9503 10652 9512
rect 10600 9469 10609 9503
rect 10609 9469 10643 9503
rect 10643 9469 10652 9503
rect 10600 9460 10652 9469
rect 13176 9503 13228 9512
rect 9864 9392 9916 9444
rect 7012 9367 7064 9376
rect 7012 9333 7021 9367
rect 7021 9333 7055 9367
rect 7055 9333 7064 9367
rect 7840 9367 7892 9376
rect 7012 9324 7064 9333
rect 7840 9333 7849 9367
rect 7849 9333 7883 9367
rect 7883 9333 7892 9367
rect 7840 9324 7892 9333
rect 8668 9367 8720 9376
rect 8668 9333 8677 9367
rect 8677 9333 8711 9367
rect 8711 9333 8720 9367
rect 8668 9324 8720 9333
rect 9128 9324 9180 9376
rect 10416 9324 10468 9376
rect 10784 9324 10836 9376
rect 11152 9367 11204 9376
rect 11152 9333 11161 9367
rect 11161 9333 11195 9367
rect 11195 9333 11204 9367
rect 11152 9324 11204 9333
rect 12256 9324 12308 9376
rect 13176 9469 13185 9503
rect 13185 9469 13219 9503
rect 13219 9469 13228 9503
rect 13176 9460 13228 9469
rect 14004 9503 14056 9512
rect 14004 9469 14013 9503
rect 14013 9469 14047 9503
rect 14047 9469 14056 9503
rect 14004 9460 14056 9469
rect 12992 9392 13044 9444
rect 15016 9460 15068 9512
rect 14556 9392 14608 9444
rect 14832 9392 14884 9444
rect 15476 9596 15528 9648
rect 16304 9596 16356 9648
rect 16488 9596 16540 9648
rect 16212 9571 16264 9580
rect 16212 9537 16221 9571
rect 16221 9537 16255 9571
rect 16255 9537 16264 9571
rect 16212 9528 16264 9537
rect 17316 9596 17368 9648
rect 15660 9460 15712 9512
rect 17224 9503 17276 9512
rect 17224 9469 17233 9503
rect 17233 9469 17267 9503
rect 17267 9469 17276 9503
rect 17224 9460 17276 9469
rect 17684 9528 17736 9580
rect 20352 9596 20404 9648
rect 18696 9528 18748 9580
rect 19064 9571 19116 9580
rect 19064 9537 19073 9571
rect 19073 9537 19107 9571
rect 19107 9537 19116 9571
rect 19064 9528 19116 9537
rect 19524 9571 19576 9580
rect 19524 9537 19558 9571
rect 19558 9537 19576 9571
rect 19524 9528 19576 9537
rect 19984 9528 20036 9580
rect 18236 9503 18288 9512
rect 17316 9392 17368 9444
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18788 9460 18840 9512
rect 20720 9460 20772 9512
rect 19156 9392 19208 9444
rect 13360 9324 13412 9376
rect 14648 9367 14700 9376
rect 14648 9333 14657 9367
rect 14657 9333 14691 9367
rect 14691 9333 14700 9367
rect 14648 9324 14700 9333
rect 14924 9367 14976 9376
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 15752 9367 15804 9376
rect 15752 9333 15761 9367
rect 15761 9333 15795 9367
rect 15795 9333 15804 9367
rect 15752 9324 15804 9333
rect 17224 9324 17276 9376
rect 17684 9324 17736 9376
rect 20168 9324 20220 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 2228 9120 2280 9172
rect 2412 9120 2464 9172
rect 2872 9163 2924 9172
rect 2504 9052 2556 9104
rect 2872 9129 2881 9163
rect 2881 9129 2915 9163
rect 2915 9129 2924 9163
rect 2872 9120 2924 9129
rect 3884 9120 3936 9172
rect 4068 9120 4120 9172
rect 4712 9120 4764 9172
rect 2688 9027 2740 9036
rect 2688 8993 2697 9027
rect 2697 8993 2731 9027
rect 2731 8993 2740 9027
rect 2688 8984 2740 8993
rect 3424 8984 3476 9036
rect 3516 9027 3568 9036
rect 3516 8993 3525 9027
rect 3525 8993 3559 9027
rect 3559 8993 3568 9027
rect 4344 9052 4396 9104
rect 6920 9052 6972 9104
rect 7472 9120 7524 9172
rect 7748 9120 7800 9172
rect 9312 9120 9364 9172
rect 10600 9120 10652 9172
rect 10876 9120 10928 9172
rect 11796 9120 11848 9172
rect 11980 9163 12032 9172
rect 11980 9129 11989 9163
rect 11989 9129 12023 9163
rect 12023 9129 12032 9163
rect 11980 9120 12032 9129
rect 12900 9120 12952 9172
rect 13544 9120 13596 9172
rect 14372 9120 14424 9172
rect 15108 9120 15160 9172
rect 8484 9052 8536 9104
rect 8668 9052 8720 9104
rect 3516 8984 3568 8993
rect 1492 8916 1544 8968
rect 1584 8916 1636 8968
rect 2780 8916 2832 8968
rect 4068 8959 4120 8968
rect 4068 8925 4077 8959
rect 4077 8925 4111 8959
rect 4111 8925 4120 8959
rect 4344 8959 4396 8968
rect 4068 8916 4120 8925
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 4436 8916 4488 8968
rect 2872 8848 2924 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2412 8823 2464 8832
rect 2412 8789 2421 8823
rect 2421 8789 2455 8823
rect 2455 8789 2464 8823
rect 2412 8780 2464 8789
rect 2504 8823 2556 8832
rect 2504 8789 2513 8823
rect 2513 8789 2547 8823
rect 2547 8789 2556 8823
rect 3240 8823 3292 8832
rect 2504 8780 2556 8789
rect 3240 8789 3249 8823
rect 3249 8789 3283 8823
rect 3283 8789 3292 8823
rect 3240 8780 3292 8789
rect 4068 8780 4120 8832
rect 4344 8780 4396 8832
rect 6644 8916 6696 8968
rect 7748 8916 7800 8968
rect 5632 8848 5684 8900
rect 5724 8823 5776 8832
rect 5724 8789 5733 8823
rect 5733 8789 5767 8823
rect 5767 8789 5776 8823
rect 5724 8780 5776 8789
rect 5908 8848 5960 8900
rect 7932 8916 7984 8968
rect 8116 9027 8168 9036
rect 8116 8993 8125 9027
rect 8125 8993 8159 9027
rect 8159 8993 8168 9027
rect 8392 9027 8444 9036
rect 8116 8984 8168 8993
rect 8392 8993 8401 9027
rect 8401 8993 8435 9027
rect 8435 8993 8444 9027
rect 8392 8984 8444 8993
rect 9036 8916 9088 8968
rect 10140 8984 10192 9036
rect 10508 9027 10560 9036
rect 10508 8993 10517 9027
rect 10517 8993 10551 9027
rect 10551 8993 10560 9027
rect 10508 8984 10560 8993
rect 10784 8959 10836 8968
rect 10784 8925 10793 8959
rect 10793 8925 10827 8959
rect 10827 8925 10836 8959
rect 10784 8916 10836 8925
rect 11152 8984 11204 9036
rect 11612 9052 11664 9104
rect 12992 9052 13044 9104
rect 12808 8984 12860 9036
rect 11520 8916 11572 8968
rect 12440 8959 12492 8968
rect 7288 8780 7340 8832
rect 9588 8848 9640 8900
rect 10324 8848 10376 8900
rect 12440 8925 12449 8959
rect 12449 8925 12483 8959
rect 12483 8925 12492 8959
rect 12440 8916 12492 8925
rect 13176 8916 13228 8968
rect 14188 8984 14240 9036
rect 14832 8916 14884 8968
rect 15568 8984 15620 9036
rect 11796 8848 11848 8900
rect 13636 8891 13688 8900
rect 13636 8857 13645 8891
rect 13645 8857 13679 8891
rect 13679 8857 13688 8891
rect 13636 8848 13688 8857
rect 8116 8780 8168 8832
rect 8392 8780 8444 8832
rect 8668 8780 8720 8832
rect 9312 8780 9364 8832
rect 10416 8780 10468 8832
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 10968 8780 11020 8832
rect 11244 8780 11296 8832
rect 11704 8780 11756 8832
rect 12532 8823 12584 8832
rect 12532 8789 12541 8823
rect 12541 8789 12575 8823
rect 12575 8789 12584 8823
rect 12532 8780 12584 8789
rect 13084 8823 13136 8832
rect 13084 8789 13093 8823
rect 13093 8789 13127 8823
rect 13127 8789 13136 8823
rect 13084 8780 13136 8789
rect 13452 8780 13504 8832
rect 14372 8780 14424 8832
rect 14464 8780 14516 8832
rect 15016 8780 15068 8832
rect 15844 8916 15896 8968
rect 17132 9120 17184 9172
rect 17316 9120 17368 9172
rect 19524 9120 19576 9172
rect 20720 9163 20772 9172
rect 17040 9052 17092 9104
rect 17776 9052 17828 9104
rect 16212 8984 16264 9036
rect 16488 8984 16540 9036
rect 17224 9027 17276 9036
rect 17224 8993 17233 9027
rect 17233 8993 17267 9027
rect 17267 8993 17276 9027
rect 17224 8984 17276 8993
rect 18696 9052 18748 9104
rect 18972 9052 19024 9104
rect 20720 9129 20729 9163
rect 20729 9129 20763 9163
rect 20763 9129 20772 9163
rect 20720 9120 20772 9129
rect 18052 8916 18104 8968
rect 18788 8984 18840 9036
rect 19892 8916 19944 8968
rect 20628 8916 20680 8968
rect 16120 8823 16172 8832
rect 16120 8789 16129 8823
rect 16129 8789 16163 8823
rect 16163 8789 16172 8823
rect 16120 8780 16172 8789
rect 17592 8848 17644 8900
rect 19800 8848 19852 8900
rect 17040 8823 17092 8832
rect 17040 8789 17049 8823
rect 17049 8789 17083 8823
rect 17083 8789 17092 8823
rect 17040 8780 17092 8789
rect 17500 8780 17552 8832
rect 18420 8780 18472 8832
rect 18972 8780 19024 8832
rect 19708 8780 19760 8832
rect 21088 8823 21140 8832
rect 21088 8789 21097 8823
rect 21097 8789 21131 8823
rect 21131 8789 21140 8823
rect 21088 8780 21140 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 2504 8576 2556 8628
rect 4988 8576 5040 8628
rect 5172 8619 5224 8628
rect 5172 8585 5181 8619
rect 5181 8585 5215 8619
rect 5215 8585 5224 8619
rect 5172 8576 5224 8585
rect 5264 8576 5316 8628
rect 5816 8576 5868 8628
rect 7840 8619 7892 8628
rect 7840 8585 7849 8619
rect 7849 8585 7883 8619
rect 7883 8585 7892 8619
rect 7840 8576 7892 8585
rect 9956 8619 10008 8628
rect 1952 8440 2004 8492
rect 1676 8415 1728 8424
rect 1676 8381 1685 8415
rect 1685 8381 1719 8415
rect 1719 8381 1728 8415
rect 1676 8372 1728 8381
rect 2228 8372 2280 8424
rect 4344 8440 4396 8492
rect 5264 8483 5316 8492
rect 5264 8449 5273 8483
rect 5273 8449 5307 8483
rect 5307 8449 5316 8483
rect 5264 8440 5316 8449
rect 5908 8508 5960 8560
rect 8300 8508 8352 8560
rect 9496 8508 9548 8560
rect 6092 8440 6144 8492
rect 6368 8440 6420 8492
rect 3976 8236 4028 8288
rect 6460 8372 6512 8424
rect 6736 8372 6788 8424
rect 6552 8304 6604 8356
rect 7840 8440 7892 8492
rect 8024 8440 8076 8492
rect 9404 8440 9456 8492
rect 9956 8585 9965 8619
rect 9965 8585 9999 8619
rect 9999 8585 10008 8619
rect 9956 8576 10008 8585
rect 10692 8576 10744 8628
rect 10876 8619 10928 8628
rect 10876 8585 10885 8619
rect 10885 8585 10919 8619
rect 10919 8585 10928 8619
rect 10876 8576 10928 8585
rect 11244 8576 11296 8628
rect 10600 8508 10652 8560
rect 11152 8508 11204 8560
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 12808 8576 12860 8628
rect 14188 8619 14240 8628
rect 14188 8585 14197 8619
rect 14197 8585 14231 8619
rect 14231 8585 14240 8619
rect 14188 8576 14240 8585
rect 12256 8508 12308 8560
rect 13728 8508 13780 8560
rect 14832 8576 14884 8628
rect 15476 8576 15528 8628
rect 16120 8576 16172 8628
rect 17040 8576 17092 8628
rect 17960 8576 18012 8628
rect 19248 8576 19300 8628
rect 19984 8619 20036 8628
rect 7932 8415 7984 8424
rect 7932 8381 7941 8415
rect 7941 8381 7975 8415
rect 7975 8381 7984 8415
rect 7932 8372 7984 8381
rect 7380 8304 7432 8356
rect 8024 8304 8076 8356
rect 8300 8304 8352 8356
rect 8484 8415 8536 8424
rect 8484 8381 8493 8415
rect 8493 8381 8527 8415
rect 8527 8381 8536 8415
rect 9128 8415 9180 8424
rect 8484 8372 8536 8381
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 9312 8415 9364 8424
rect 9312 8381 9321 8415
rect 9321 8381 9355 8415
rect 9355 8381 9364 8415
rect 9312 8372 9364 8381
rect 10048 8415 10100 8424
rect 10048 8381 10057 8415
rect 10057 8381 10091 8415
rect 10091 8381 10100 8415
rect 10048 8372 10100 8381
rect 15936 8508 15988 8560
rect 16764 8508 16816 8560
rect 18512 8508 18564 8560
rect 13544 8415 13596 8424
rect 13544 8381 13553 8415
rect 13553 8381 13587 8415
rect 13587 8381 13596 8415
rect 13544 8372 13596 8381
rect 14372 8415 14424 8424
rect 14372 8381 14381 8415
rect 14381 8381 14415 8415
rect 14415 8381 14424 8415
rect 14372 8372 14424 8381
rect 17040 8483 17092 8492
rect 14556 8372 14608 8424
rect 15016 8415 15068 8424
rect 10140 8304 10192 8356
rect 10324 8347 10376 8356
rect 10324 8313 10333 8347
rect 10333 8313 10367 8347
rect 10367 8313 10376 8347
rect 10324 8304 10376 8313
rect 5724 8236 5776 8288
rect 7196 8236 7248 8288
rect 7472 8236 7524 8288
rect 10692 8236 10744 8288
rect 10876 8304 10928 8356
rect 11060 8304 11112 8356
rect 11152 8304 11204 8356
rect 13268 8304 13320 8356
rect 13452 8304 13504 8356
rect 15016 8381 15025 8415
rect 15025 8381 15059 8415
rect 15059 8381 15068 8415
rect 15016 8372 15068 8381
rect 14832 8304 14884 8356
rect 17040 8449 17049 8483
rect 17049 8449 17083 8483
rect 17083 8449 17092 8483
rect 17040 8440 17092 8449
rect 17316 8440 17368 8492
rect 18236 8440 18288 8492
rect 16856 8372 16908 8424
rect 17224 8415 17276 8424
rect 17224 8381 17233 8415
rect 17233 8381 17267 8415
rect 17267 8381 17276 8415
rect 17224 8372 17276 8381
rect 18512 8415 18564 8424
rect 18512 8381 18521 8415
rect 18521 8381 18555 8415
rect 18555 8381 18564 8415
rect 18512 8372 18564 8381
rect 19524 8508 19576 8560
rect 19984 8585 19993 8619
rect 19993 8585 20027 8619
rect 20027 8585 20036 8619
rect 19984 8576 20036 8585
rect 20720 8508 20772 8560
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 20352 8440 20404 8492
rect 21272 8440 21324 8492
rect 19524 8415 19576 8424
rect 19524 8381 19533 8415
rect 19533 8381 19567 8415
rect 19567 8381 19576 8415
rect 19524 8372 19576 8381
rect 20168 8372 20220 8424
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 11336 8236 11388 8288
rect 11796 8236 11848 8288
rect 12532 8236 12584 8288
rect 12624 8236 12676 8288
rect 13176 8236 13228 8288
rect 15384 8236 15436 8288
rect 15936 8236 15988 8288
rect 20076 8304 20128 8356
rect 18972 8236 19024 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1952 8032 2004 8084
rect 2412 8032 2464 8084
rect 5448 8075 5500 8084
rect 5448 8041 5457 8075
rect 5457 8041 5491 8075
rect 5491 8041 5500 8075
rect 5448 8032 5500 8041
rect 3240 7964 3292 8016
rect 4896 7964 4948 8016
rect 5632 7964 5684 8016
rect 3976 7896 4028 7948
rect 4252 7896 4304 7948
rect 5172 7939 5224 7948
rect 5172 7905 5181 7939
rect 5181 7905 5215 7939
rect 5215 7905 5224 7939
rect 5172 7896 5224 7905
rect 5724 7896 5776 7948
rect 6368 7964 6420 8016
rect 7656 8032 7708 8084
rect 7380 7964 7432 8016
rect 8668 8032 8720 8084
rect 9312 8032 9364 8084
rect 10140 8032 10192 8084
rect 10784 8032 10836 8084
rect 10876 8032 10928 8084
rect 8576 7964 8628 8016
rect 8300 7896 8352 7948
rect 11612 8032 11664 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 12440 8032 12492 8041
rect 12716 8032 12768 8084
rect 12808 8032 12860 8084
rect 20 7828 72 7880
rect 1032 7828 1084 7880
rect 1584 7828 1636 7880
rect 1676 7803 1728 7812
rect 1676 7769 1685 7803
rect 1685 7769 1719 7803
rect 1719 7769 1728 7803
rect 1676 7760 1728 7769
rect 3516 7828 3568 7880
rect 4160 7871 4212 7880
rect 4160 7837 4169 7871
rect 4169 7837 4203 7871
rect 4203 7837 4212 7871
rect 4160 7828 4212 7837
rect 5264 7828 5316 7880
rect 3700 7760 3752 7812
rect 6000 7760 6052 7812
rect 4068 7692 4120 7744
rect 4344 7692 4396 7744
rect 5080 7735 5132 7744
rect 5080 7701 5089 7735
rect 5089 7701 5123 7735
rect 5123 7701 5132 7735
rect 5080 7692 5132 7701
rect 5724 7692 5776 7744
rect 6644 7828 6696 7880
rect 7656 7828 7708 7880
rect 6828 7760 6880 7812
rect 7380 7692 7432 7744
rect 7472 7692 7524 7744
rect 9036 7828 9088 7880
rect 11244 7871 11296 7880
rect 11244 7837 11278 7871
rect 11278 7837 11296 7871
rect 12532 7896 12584 7948
rect 13544 7896 13596 7948
rect 12808 7871 12860 7880
rect 11244 7828 11296 7837
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 13728 8032 13780 8084
rect 14556 8032 14608 8084
rect 15016 8032 15068 8084
rect 15568 8075 15620 8084
rect 15568 8041 15577 8075
rect 15577 8041 15611 8075
rect 15611 8041 15620 8075
rect 15568 8032 15620 8041
rect 15844 8032 15896 8084
rect 14464 7964 14516 8016
rect 14832 7964 14884 8016
rect 13912 7896 13964 7948
rect 14372 7896 14424 7948
rect 15844 7896 15896 7948
rect 17316 7896 17368 7948
rect 9588 7760 9640 7812
rect 9864 7760 9916 7812
rect 10140 7760 10192 7812
rect 10692 7760 10744 7812
rect 12256 7760 12308 7812
rect 12624 7760 12676 7812
rect 13084 7760 13136 7812
rect 13176 7803 13228 7812
rect 13176 7769 13185 7803
rect 13185 7769 13219 7803
rect 13219 7769 13228 7803
rect 13176 7760 13228 7769
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8576 7692 8628 7744
rect 9312 7692 9364 7744
rect 9496 7692 9548 7744
rect 10416 7692 10468 7744
rect 10876 7735 10928 7744
rect 10876 7701 10885 7735
rect 10885 7701 10919 7735
rect 10919 7701 10928 7735
rect 10876 7692 10928 7701
rect 11888 7692 11940 7744
rect 12348 7735 12400 7744
rect 12348 7701 12357 7735
rect 12357 7701 12391 7735
rect 12391 7701 12400 7735
rect 12348 7692 12400 7701
rect 13544 7692 13596 7744
rect 14832 7692 14884 7744
rect 15384 7828 15436 7880
rect 16212 7828 16264 7880
rect 16856 7828 16908 7880
rect 17408 7871 17460 7880
rect 17408 7837 17417 7871
rect 17417 7837 17451 7871
rect 17451 7837 17460 7871
rect 17408 7828 17460 7837
rect 18052 8032 18104 8084
rect 19524 8032 19576 8084
rect 21364 8075 21416 8084
rect 21364 8041 21373 8075
rect 21373 8041 21407 8075
rect 21407 8041 21416 8075
rect 21364 8032 21416 8041
rect 19800 7964 19852 8016
rect 19708 7896 19760 7948
rect 19892 7896 19944 7948
rect 21364 7896 21416 7948
rect 19984 7828 20036 7880
rect 15752 7760 15804 7812
rect 16948 7760 17000 7812
rect 18512 7760 18564 7812
rect 18972 7760 19024 7812
rect 20536 7828 20588 7880
rect 20720 7760 20772 7812
rect 15476 7692 15528 7744
rect 16212 7692 16264 7744
rect 18236 7692 18288 7744
rect 19156 7692 19208 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 756 7488 808 7540
rect 2964 7488 3016 7540
rect 1492 7463 1544 7472
rect 1492 7429 1501 7463
rect 1501 7429 1535 7463
rect 1535 7429 1544 7463
rect 1492 7420 1544 7429
rect 2964 7395 3016 7404
rect 2964 7361 2982 7395
rect 2982 7361 3016 7395
rect 5172 7488 5224 7540
rect 7288 7488 7340 7540
rect 7656 7531 7708 7540
rect 7656 7497 7665 7531
rect 7665 7497 7699 7531
rect 7699 7497 7708 7531
rect 7656 7488 7708 7497
rect 8392 7488 8444 7540
rect 8484 7488 8536 7540
rect 10232 7488 10284 7540
rect 11980 7531 12032 7540
rect 11980 7497 11989 7531
rect 11989 7497 12023 7531
rect 12023 7497 12032 7531
rect 11980 7488 12032 7497
rect 12256 7488 12308 7540
rect 12716 7531 12768 7540
rect 12716 7497 12725 7531
rect 12725 7497 12759 7531
rect 12759 7497 12768 7531
rect 12716 7488 12768 7497
rect 13084 7488 13136 7540
rect 13176 7488 13228 7540
rect 13636 7531 13688 7540
rect 13636 7497 13645 7531
rect 13645 7497 13679 7531
rect 13679 7497 13688 7531
rect 13636 7488 13688 7497
rect 6184 7420 6236 7472
rect 6460 7420 6512 7472
rect 6644 7420 6696 7472
rect 6828 7463 6880 7472
rect 6828 7429 6837 7463
rect 6837 7429 6871 7463
rect 6871 7429 6880 7463
rect 6828 7420 6880 7429
rect 2964 7352 3016 7361
rect 3700 7352 3752 7404
rect 4068 7352 4120 7404
rect 4252 7395 4304 7404
rect 4252 7361 4286 7395
rect 4286 7361 4304 7395
rect 4252 7352 4304 7361
rect 4988 7352 5040 7404
rect 5172 7352 5224 7404
rect 3332 7327 3384 7336
rect 3332 7293 3341 7327
rect 3341 7293 3375 7327
rect 3375 7293 3384 7327
rect 3332 7284 3384 7293
rect 3608 7284 3660 7336
rect 1584 7148 1636 7200
rect 4988 7216 5040 7268
rect 7472 7352 7524 7404
rect 8392 7352 8444 7404
rect 9312 7420 9364 7472
rect 10600 7420 10652 7472
rect 9128 7352 9180 7404
rect 6644 7284 6696 7336
rect 9588 7284 9640 7336
rect 10232 7327 10284 7336
rect 10232 7293 10241 7327
rect 10241 7293 10275 7327
rect 10275 7293 10284 7327
rect 10232 7284 10284 7293
rect 11796 7284 11848 7336
rect 12348 7284 12400 7336
rect 12532 7327 12584 7336
rect 12532 7293 12541 7327
rect 12541 7293 12575 7327
rect 12575 7293 12584 7327
rect 12532 7284 12584 7293
rect 3976 7148 4028 7200
rect 4344 7148 4396 7200
rect 6920 7148 6972 7200
rect 7656 7148 7708 7200
rect 10876 7216 10928 7268
rect 9312 7148 9364 7200
rect 10140 7148 10192 7200
rect 10600 7148 10652 7200
rect 11152 7148 11204 7200
rect 12532 7148 12584 7200
rect 12900 7352 12952 7404
rect 13084 7352 13136 7404
rect 13636 7352 13688 7404
rect 13820 7488 13872 7540
rect 15108 7488 15160 7540
rect 16028 7531 16080 7540
rect 16028 7497 16037 7531
rect 16037 7497 16071 7531
rect 16071 7497 16080 7531
rect 16028 7488 16080 7497
rect 16304 7488 16356 7540
rect 13360 7284 13412 7336
rect 13912 7327 13964 7336
rect 13912 7293 13921 7327
rect 13921 7293 13955 7327
rect 13955 7293 13964 7327
rect 13912 7284 13964 7293
rect 12716 7216 12768 7268
rect 13728 7216 13780 7268
rect 14464 7395 14516 7404
rect 14464 7361 14473 7395
rect 14473 7361 14507 7395
rect 14507 7361 14516 7395
rect 14464 7352 14516 7361
rect 14280 7259 14332 7268
rect 14280 7225 14289 7259
rect 14289 7225 14323 7259
rect 14323 7225 14332 7259
rect 14832 7352 14884 7404
rect 15200 7395 15252 7404
rect 15200 7361 15209 7395
rect 15209 7361 15243 7395
rect 15243 7361 15252 7395
rect 15200 7352 15252 7361
rect 14280 7216 14332 7225
rect 12992 7148 13044 7200
rect 13176 7191 13228 7200
rect 13176 7157 13185 7191
rect 13185 7157 13219 7191
rect 13219 7157 13228 7191
rect 13176 7148 13228 7157
rect 13360 7148 13412 7200
rect 14740 7191 14792 7200
rect 14740 7157 14749 7191
rect 14749 7157 14783 7191
rect 14783 7157 14792 7191
rect 14740 7148 14792 7157
rect 15384 7420 15436 7472
rect 15752 7395 15804 7404
rect 15752 7361 15761 7395
rect 15761 7361 15795 7395
rect 15795 7361 15804 7395
rect 15752 7352 15804 7361
rect 16212 7395 16264 7404
rect 16212 7361 16221 7395
rect 16221 7361 16255 7395
rect 16255 7361 16264 7395
rect 17040 7488 17092 7540
rect 17960 7488 18012 7540
rect 19156 7488 19208 7540
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 19616 7488 19668 7540
rect 20076 7488 20128 7540
rect 20812 7531 20864 7540
rect 20812 7497 20821 7531
rect 20821 7497 20855 7531
rect 20855 7497 20864 7531
rect 20812 7488 20864 7497
rect 20904 7488 20956 7540
rect 21088 7488 21140 7540
rect 21364 7531 21416 7540
rect 21364 7497 21373 7531
rect 21373 7497 21407 7531
rect 21407 7497 21416 7531
rect 21364 7488 21416 7497
rect 16580 7420 16632 7472
rect 17776 7420 17828 7472
rect 19064 7420 19116 7472
rect 20536 7420 20588 7472
rect 16212 7352 16264 7361
rect 16672 7395 16724 7404
rect 16672 7361 16681 7395
rect 16681 7361 16715 7395
rect 16715 7361 16724 7395
rect 16672 7352 16724 7361
rect 17224 7352 17276 7404
rect 17592 7395 17644 7404
rect 17592 7361 17601 7395
rect 17601 7361 17635 7395
rect 17635 7361 17644 7395
rect 17592 7352 17644 7361
rect 15936 7284 15988 7336
rect 16212 7216 16264 7268
rect 17316 7216 17368 7268
rect 17408 7216 17460 7268
rect 18512 7352 18564 7404
rect 20076 7395 20128 7404
rect 20076 7361 20085 7395
rect 20085 7361 20119 7395
rect 20119 7361 20128 7395
rect 20076 7352 20128 7361
rect 18972 7327 19024 7336
rect 18972 7293 18981 7327
rect 18981 7293 19015 7327
rect 19015 7293 19024 7327
rect 18972 7284 19024 7293
rect 19064 7284 19116 7336
rect 19800 7284 19852 7336
rect 19708 7216 19760 7268
rect 20904 7395 20956 7404
rect 20904 7361 20913 7395
rect 20913 7361 20947 7395
rect 20947 7361 20956 7395
rect 20904 7352 20956 7361
rect 21548 7395 21600 7404
rect 21548 7361 21557 7395
rect 21557 7361 21591 7395
rect 21591 7361 21600 7395
rect 21548 7352 21600 7361
rect 15108 7148 15160 7200
rect 15936 7191 15988 7200
rect 15936 7157 15945 7191
rect 15945 7157 15979 7191
rect 15979 7157 15988 7191
rect 15936 7148 15988 7157
rect 16488 7148 16540 7200
rect 16580 7148 16632 7200
rect 17868 7148 17920 7200
rect 19616 7191 19668 7200
rect 19616 7157 19625 7191
rect 19625 7157 19659 7191
rect 19659 7157 19668 7191
rect 19616 7148 19668 7157
rect 19984 7148 20036 7200
rect 20812 7148 20864 7200
rect 21732 7148 21784 7200
rect 22008 7148 22060 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 22008 7012 22060 7064
rect 22376 7012 22428 7064
rect 4068 6944 4120 6996
rect 1032 6808 1084 6860
rect 1308 6740 1360 6792
rect 1952 6808 2004 6860
rect 2596 6808 2648 6860
rect 4896 6876 4948 6928
rect 3516 6851 3568 6860
rect 3516 6817 3525 6851
rect 3525 6817 3559 6851
rect 3559 6817 3568 6851
rect 3516 6808 3568 6817
rect 7104 6919 7156 6928
rect 7104 6885 7113 6919
rect 7113 6885 7147 6919
rect 7147 6885 7156 6919
rect 7104 6876 7156 6885
rect 7288 6944 7340 6996
rect 8208 6944 8260 6996
rect 8300 6944 8352 6996
rect 9404 6944 9456 6996
rect 7656 6876 7708 6928
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 3976 6783 4028 6792
rect 3976 6749 3985 6783
rect 3985 6749 4019 6783
rect 4019 6749 4028 6783
rect 3976 6740 4028 6749
rect 4068 6740 4120 6792
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 4528 6783 4580 6792
rect 4528 6749 4537 6783
rect 4537 6749 4571 6783
rect 4571 6749 4580 6783
rect 4528 6740 4580 6749
rect 4896 6740 4948 6792
rect 5172 6783 5224 6792
rect 5172 6749 5181 6783
rect 5181 6749 5215 6783
rect 5215 6749 5224 6783
rect 5172 6740 5224 6749
rect 5448 6783 5500 6792
rect 5448 6749 5457 6783
rect 5457 6749 5491 6783
rect 5491 6749 5500 6783
rect 5448 6740 5500 6749
rect 2044 6672 2096 6724
rect 4988 6672 5040 6724
rect 6736 6808 6788 6860
rect 8300 6851 8352 6860
rect 8300 6817 8309 6851
rect 8309 6817 8343 6851
rect 8343 6817 8352 6851
rect 8300 6808 8352 6817
rect 8668 6808 8720 6860
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 10600 6876 10652 6928
rect 11980 6944 12032 6996
rect 12992 6944 13044 6996
rect 15660 6944 15712 6996
rect 15752 6944 15804 6996
rect 18052 6944 18104 6996
rect 18236 6944 18288 6996
rect 21548 6944 21600 6996
rect 5816 6740 5868 6792
rect 8116 6740 8168 6792
rect 8484 6740 8536 6792
rect 9220 6740 9272 6792
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 10048 6740 10100 6792
rect 10232 6740 10284 6792
rect 15936 6876 15988 6928
rect 16488 6876 16540 6928
rect 11060 6808 11112 6860
rect 11244 6808 11296 6860
rect 13544 6851 13596 6860
rect 13544 6817 13553 6851
rect 13553 6817 13587 6851
rect 13587 6817 13596 6851
rect 13544 6808 13596 6817
rect 14464 6851 14516 6860
rect 6552 6672 6604 6724
rect 11244 6672 11296 6724
rect 1860 6604 1912 6656
rect 2136 6604 2188 6656
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 4160 6647 4212 6656
rect 2780 6604 2832 6613
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4712 6604 4764 6656
rect 5632 6647 5684 6656
rect 5632 6613 5641 6647
rect 5641 6613 5675 6647
rect 5675 6613 5684 6647
rect 5632 6604 5684 6613
rect 5908 6604 5960 6656
rect 7472 6604 7524 6656
rect 7932 6604 7984 6656
rect 9220 6604 9272 6656
rect 9312 6604 9364 6656
rect 9772 6647 9824 6656
rect 9772 6613 9781 6647
rect 9781 6613 9815 6647
rect 9815 6613 9824 6647
rect 9772 6604 9824 6613
rect 10140 6604 10192 6656
rect 10876 6604 10928 6656
rect 12440 6740 12492 6792
rect 13176 6740 13228 6792
rect 12072 6672 12124 6724
rect 14464 6817 14473 6851
rect 14473 6817 14507 6851
rect 14507 6817 14516 6851
rect 14464 6808 14516 6817
rect 17224 6876 17276 6928
rect 15936 6740 15988 6792
rect 16120 6740 16172 6792
rect 16948 6808 17000 6860
rect 17132 6808 17184 6860
rect 18144 6876 18196 6928
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 18420 6808 18472 6860
rect 19248 6876 19300 6928
rect 17960 6740 18012 6792
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18880 6740 18932 6792
rect 13728 6672 13780 6724
rect 11704 6604 11756 6656
rect 11796 6604 11848 6656
rect 12348 6604 12400 6656
rect 13912 6604 13964 6656
rect 14556 6604 14608 6656
rect 15292 6672 15344 6724
rect 15568 6604 15620 6656
rect 15844 6647 15896 6656
rect 15844 6613 15853 6647
rect 15853 6613 15887 6647
rect 15887 6613 15896 6647
rect 15844 6604 15896 6613
rect 16304 6647 16356 6656
rect 16304 6613 16313 6647
rect 16313 6613 16347 6647
rect 16347 6613 16356 6647
rect 16304 6604 16356 6613
rect 17500 6672 17552 6724
rect 18972 6715 19024 6724
rect 18972 6681 18981 6715
rect 18981 6681 19015 6715
rect 19015 6681 19024 6715
rect 18972 6672 19024 6681
rect 19156 6740 19208 6792
rect 21088 6808 21140 6860
rect 21824 6740 21876 6792
rect 19892 6672 19944 6724
rect 19984 6672 20036 6724
rect 20720 6672 20772 6724
rect 17408 6604 17460 6656
rect 18144 6604 18196 6656
rect 18512 6604 18564 6656
rect 20444 6604 20496 6656
rect 21456 6604 21508 6656
rect 21824 6604 21876 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 1400 6400 1452 6452
rect 2228 6400 2280 6452
rect 3424 6400 3476 6452
rect 3884 6400 3936 6452
rect 5724 6400 5776 6452
rect 5816 6400 5868 6452
rect 6000 6400 6052 6452
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 7012 6400 7064 6452
rect 8116 6400 8168 6452
rect 8944 6443 8996 6452
rect 8944 6409 8953 6443
rect 8953 6409 8987 6443
rect 8987 6409 8996 6443
rect 8944 6400 8996 6409
rect 9588 6400 9640 6452
rect 9772 6443 9824 6452
rect 9772 6409 9781 6443
rect 9781 6409 9815 6443
rect 9815 6409 9824 6443
rect 9772 6400 9824 6409
rect 388 6332 440 6384
rect 940 6332 992 6384
rect 3056 6332 3108 6384
rect 4528 6332 4580 6384
rect 3700 6307 3752 6316
rect 3700 6273 3709 6307
rect 3709 6273 3743 6307
rect 3743 6273 3752 6307
rect 3700 6264 3752 6273
rect 4896 6264 4948 6316
rect 5172 6264 5224 6316
rect 2412 6196 2464 6248
rect 2964 6196 3016 6248
rect 4068 6196 4120 6248
rect 4252 6196 4304 6248
rect 5356 6332 5408 6384
rect 6184 6264 6236 6316
rect 9312 6332 9364 6384
rect 6727 6307 6779 6316
rect 6727 6273 6745 6307
rect 6745 6273 6779 6307
rect 6727 6264 6779 6273
rect 3424 6128 3476 6180
rect 5724 6196 5776 6248
rect 6092 6239 6144 6248
rect 6092 6205 6101 6239
rect 6101 6205 6135 6239
rect 6135 6205 6144 6239
rect 6092 6196 6144 6205
rect 6368 6196 6420 6248
rect 6460 6196 6512 6248
rect 1952 6103 2004 6112
rect 1952 6069 1961 6103
rect 1961 6069 1995 6103
rect 1995 6069 2004 6103
rect 1952 6060 2004 6069
rect 2320 6060 2372 6112
rect 2780 6060 2832 6112
rect 3240 6060 3292 6112
rect 5080 6060 5132 6112
rect 6000 6128 6052 6180
rect 6920 6128 6972 6180
rect 7196 6264 7248 6316
rect 8208 6264 8260 6316
rect 9956 6264 10008 6316
rect 10140 6264 10192 6316
rect 10784 6264 10836 6316
rect 8300 6196 8352 6248
rect 8024 6128 8076 6180
rect 8208 6128 8260 6180
rect 7932 6060 7984 6112
rect 8116 6060 8168 6112
rect 9680 6239 9732 6248
rect 9680 6205 9689 6239
rect 9689 6205 9723 6239
rect 9723 6205 9732 6239
rect 9680 6196 9732 6205
rect 11244 6332 11296 6384
rect 13728 6400 13780 6452
rect 12348 6332 12400 6384
rect 12992 6332 13044 6384
rect 13636 6332 13688 6384
rect 16304 6400 16356 6452
rect 18144 6400 18196 6452
rect 19064 6443 19116 6452
rect 19064 6409 19073 6443
rect 19073 6409 19107 6443
rect 19107 6409 19116 6443
rect 19064 6400 19116 6409
rect 19616 6400 19668 6452
rect 20628 6443 20680 6452
rect 20628 6409 20637 6443
rect 20637 6409 20671 6443
rect 20671 6409 20680 6443
rect 20628 6400 20680 6409
rect 14648 6332 14700 6384
rect 15476 6332 15528 6384
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 14280 6264 14332 6316
rect 9772 6128 9824 6180
rect 11428 6196 11480 6248
rect 11980 6196 12032 6248
rect 10600 6128 10652 6180
rect 10692 6128 10744 6180
rect 11796 6128 11848 6180
rect 12164 6128 12216 6180
rect 13728 6128 13780 6180
rect 15108 6196 15160 6248
rect 15660 6307 15712 6316
rect 15660 6273 15669 6307
rect 15669 6273 15703 6307
rect 15703 6273 15712 6307
rect 15660 6264 15712 6273
rect 16120 6264 16172 6316
rect 16580 6264 16632 6316
rect 17040 6264 17092 6316
rect 17224 6264 17276 6316
rect 15292 6128 15344 6180
rect 16488 6196 16540 6248
rect 18512 6332 18564 6384
rect 22928 6332 22980 6384
rect 18144 6264 18196 6316
rect 19432 6307 19484 6316
rect 19432 6273 19441 6307
rect 19441 6273 19475 6307
rect 19475 6273 19484 6307
rect 19432 6264 19484 6273
rect 19800 6264 19852 6316
rect 20260 6307 20312 6316
rect 18328 6239 18380 6248
rect 18328 6205 18337 6239
rect 18337 6205 18371 6239
rect 18371 6205 18380 6239
rect 18328 6196 18380 6205
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 17776 6128 17828 6180
rect 18604 6128 18656 6180
rect 18972 6171 19024 6180
rect 18972 6137 18981 6171
rect 18981 6137 19015 6171
rect 19015 6137 19024 6171
rect 18972 6128 19024 6137
rect 19892 6196 19944 6248
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20996 6307 21048 6316
rect 20996 6273 21005 6307
rect 21005 6273 21039 6307
rect 21039 6273 21048 6307
rect 20996 6264 21048 6273
rect 21456 6196 21508 6248
rect 9588 6060 9640 6112
rect 10876 6060 10928 6112
rect 11060 6103 11112 6112
rect 11060 6069 11069 6103
rect 11069 6069 11103 6103
rect 11103 6069 11112 6103
rect 11060 6060 11112 6069
rect 11336 6103 11388 6112
rect 11336 6069 11345 6103
rect 11345 6069 11379 6103
rect 11379 6069 11388 6103
rect 11336 6060 11388 6069
rect 13820 6060 13872 6112
rect 14924 6060 14976 6112
rect 15936 6060 15988 6112
rect 16396 6060 16448 6112
rect 20444 6060 20496 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 2136 5899 2188 5908
rect 2136 5865 2145 5899
rect 2145 5865 2179 5899
rect 2179 5865 2188 5899
rect 2136 5856 2188 5865
rect 4252 5899 4304 5908
rect 4252 5865 4261 5899
rect 4261 5865 4295 5899
rect 4295 5865 4304 5899
rect 4252 5856 4304 5865
rect 4896 5856 4948 5908
rect 6552 5856 6604 5908
rect 7012 5856 7064 5908
rect 7472 5856 7524 5908
rect 7932 5856 7984 5908
rect 10600 5899 10652 5908
rect 3608 5788 3660 5840
rect 4068 5788 4120 5840
rect 1584 5763 1636 5772
rect 1584 5729 1593 5763
rect 1593 5729 1627 5763
rect 1627 5729 1636 5763
rect 1584 5720 1636 5729
rect 1952 5720 2004 5772
rect 6000 5788 6052 5840
rect 9128 5788 9180 5840
rect 2504 5584 2556 5636
rect 3608 5695 3660 5704
rect 3608 5661 3617 5695
rect 3617 5661 3651 5695
rect 3651 5661 3660 5695
rect 3608 5652 3660 5661
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 4344 5652 4396 5704
rect 6092 5720 6144 5772
rect 7104 5720 7156 5772
rect 7288 5720 7340 5772
rect 7564 5763 7616 5772
rect 7564 5729 7573 5763
rect 7573 5729 7607 5763
rect 7607 5729 7616 5763
rect 7564 5720 7616 5729
rect 8300 5720 8352 5772
rect 8484 5720 8536 5772
rect 3976 5584 4028 5636
rect 5724 5652 5776 5704
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 6276 5652 6328 5704
rect 6920 5652 6972 5704
rect 7748 5652 7800 5704
rect 1768 5559 1820 5568
rect 1768 5525 1777 5559
rect 1777 5525 1811 5559
rect 1811 5525 1820 5559
rect 1768 5516 1820 5525
rect 2320 5516 2372 5568
rect 4896 5516 4948 5568
rect 5448 5516 5500 5568
rect 5724 5559 5776 5568
rect 5724 5525 5733 5559
rect 5733 5525 5767 5559
rect 5767 5525 5776 5559
rect 5724 5516 5776 5525
rect 7104 5516 7156 5568
rect 7472 5584 7524 5636
rect 8116 5695 8168 5704
rect 8116 5661 8125 5695
rect 8125 5661 8159 5695
rect 8159 5661 8168 5695
rect 8116 5652 8168 5661
rect 8852 5652 8904 5704
rect 10600 5865 10609 5899
rect 10609 5865 10643 5899
rect 10643 5865 10652 5899
rect 10600 5856 10652 5865
rect 10784 5899 10836 5908
rect 10784 5865 10793 5899
rect 10793 5865 10827 5899
rect 10827 5865 10836 5899
rect 10784 5856 10836 5865
rect 10324 5788 10376 5840
rect 11336 5856 11388 5908
rect 12624 5856 12676 5908
rect 15476 5856 15528 5908
rect 18512 5856 18564 5908
rect 19892 5856 19944 5908
rect 20904 5856 20956 5908
rect 13544 5788 13596 5840
rect 11428 5763 11480 5772
rect 11428 5729 11437 5763
rect 11437 5729 11471 5763
rect 11471 5729 11480 5763
rect 11428 5720 11480 5729
rect 12532 5720 12584 5772
rect 12716 5720 12768 5772
rect 12900 5720 12952 5772
rect 14648 5763 14700 5772
rect 8300 5516 8352 5568
rect 8668 5516 8720 5568
rect 9312 5516 9364 5568
rect 9956 5584 10008 5636
rect 11428 5584 11480 5636
rect 11980 5627 12032 5636
rect 11980 5593 11989 5627
rect 11989 5593 12023 5627
rect 12023 5593 12032 5627
rect 11980 5584 12032 5593
rect 12440 5584 12492 5636
rect 9864 5516 9916 5568
rect 10416 5516 10468 5568
rect 10600 5516 10652 5568
rect 11244 5516 11296 5568
rect 11704 5516 11756 5568
rect 12808 5559 12860 5568
rect 12808 5525 12817 5559
rect 12817 5525 12851 5559
rect 12851 5525 12860 5559
rect 13176 5559 13228 5568
rect 12808 5516 12860 5525
rect 13176 5525 13185 5559
rect 13185 5525 13219 5559
rect 13219 5525 13228 5559
rect 13176 5516 13228 5525
rect 13820 5652 13872 5704
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 14740 5720 14792 5772
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 14280 5584 14332 5636
rect 13636 5516 13688 5568
rect 15016 5584 15068 5636
rect 15844 5652 15896 5704
rect 18788 5831 18840 5840
rect 18788 5797 18797 5831
rect 18797 5797 18831 5831
rect 18831 5797 18840 5831
rect 18788 5788 18840 5797
rect 14556 5516 14608 5568
rect 16304 5516 16356 5568
rect 16948 5720 17000 5772
rect 18236 5720 18288 5772
rect 18880 5720 18932 5772
rect 21548 5720 21600 5772
rect 17776 5695 17828 5704
rect 17776 5661 17785 5695
rect 17785 5661 17819 5695
rect 17819 5661 17828 5695
rect 17776 5652 17828 5661
rect 17684 5584 17736 5636
rect 18052 5584 18104 5636
rect 17868 5559 17920 5568
rect 17868 5525 17877 5559
rect 17877 5525 17911 5559
rect 17911 5525 17920 5559
rect 19340 5652 19392 5704
rect 21088 5695 21140 5704
rect 21088 5661 21097 5695
rect 21097 5661 21131 5695
rect 21131 5661 21140 5695
rect 21088 5652 21140 5661
rect 18604 5627 18656 5636
rect 18604 5593 18613 5627
rect 18613 5593 18647 5627
rect 18647 5593 18656 5627
rect 18604 5584 18656 5593
rect 19892 5584 19944 5636
rect 17868 5516 17920 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 3056 5312 3108 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 3976 5312 4028 5364
rect 5724 5312 5776 5364
rect 1492 5287 1544 5296
rect 1492 5253 1501 5287
rect 1501 5253 1535 5287
rect 1535 5253 1544 5287
rect 1492 5244 1544 5253
rect 3608 5244 3660 5296
rect 4160 5244 4212 5296
rect 2136 5219 2188 5228
rect 2136 5185 2170 5219
rect 2170 5185 2188 5219
rect 2136 5176 2188 5185
rect 2596 5176 2648 5228
rect 3056 5176 3108 5228
rect 3884 5176 3936 5228
rect 5172 5244 5224 5296
rect 6644 5312 6696 5364
rect 8116 5312 8168 5364
rect 9772 5244 9824 5296
rect 5540 5219 5592 5228
rect 5540 5185 5549 5219
rect 5549 5185 5583 5219
rect 5583 5185 5592 5219
rect 5540 5176 5592 5185
rect 5908 5176 5960 5228
rect 7656 5176 7708 5228
rect 3240 5108 3292 5160
rect 4344 5151 4396 5160
rect 4344 5117 4353 5151
rect 4353 5117 4387 5151
rect 4387 5117 4396 5151
rect 4344 5108 4396 5117
rect 4528 5151 4580 5160
rect 4528 5117 4537 5151
rect 4537 5117 4571 5151
rect 4571 5117 4580 5151
rect 4528 5108 4580 5117
rect 2136 4972 2188 5024
rect 2596 4972 2648 5024
rect 4988 5040 5040 5092
rect 6736 5108 6788 5160
rect 7932 5108 7984 5160
rect 8300 5176 8352 5228
rect 9036 5219 9088 5228
rect 9036 5185 9045 5219
rect 9045 5185 9079 5219
rect 9079 5185 9088 5219
rect 9036 5176 9088 5185
rect 10232 5176 10284 5228
rect 11060 5312 11112 5364
rect 10876 5287 10928 5296
rect 10876 5253 10885 5287
rect 10885 5253 10919 5287
rect 10919 5253 10928 5287
rect 10876 5244 10928 5253
rect 11888 5312 11940 5364
rect 12256 5312 12308 5364
rect 13636 5312 13688 5364
rect 11336 5244 11388 5296
rect 11428 5244 11480 5296
rect 11888 5176 11940 5228
rect 12532 5244 12584 5296
rect 13728 5287 13780 5296
rect 13728 5253 13746 5287
rect 13746 5253 13780 5287
rect 13728 5244 13780 5253
rect 14924 5312 14976 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 15292 5312 15344 5321
rect 17408 5312 17460 5364
rect 17868 5312 17920 5364
rect 15568 5244 15620 5296
rect 15752 5244 15804 5296
rect 12440 5176 12492 5228
rect 5632 5040 5684 5092
rect 5816 5040 5868 5092
rect 8208 5040 8260 5092
rect 4436 4972 4488 5024
rect 5908 5015 5960 5024
rect 5908 4981 5917 5015
rect 5917 4981 5951 5015
rect 5951 4981 5960 5015
rect 5908 4972 5960 4981
rect 6092 4972 6144 5024
rect 6828 4972 6880 5024
rect 7472 4972 7524 5024
rect 7840 5015 7892 5024
rect 7840 4981 7849 5015
rect 7849 4981 7883 5015
rect 7883 4981 7892 5015
rect 7840 4972 7892 4981
rect 8484 4972 8536 5024
rect 9404 4972 9456 5024
rect 9772 4972 9824 5024
rect 14280 5108 14332 5160
rect 14924 5176 14976 5228
rect 14648 5151 14700 5160
rect 14648 5117 14657 5151
rect 14657 5117 14691 5151
rect 14691 5117 14700 5151
rect 15384 5176 15436 5228
rect 17684 5176 17736 5228
rect 18236 5176 18288 5228
rect 18880 5244 18932 5296
rect 20076 5312 20128 5364
rect 20168 5355 20220 5364
rect 20168 5321 20177 5355
rect 20177 5321 20211 5355
rect 20211 5321 20220 5355
rect 20168 5312 20220 5321
rect 22560 5244 22612 5296
rect 18972 5176 19024 5228
rect 20628 5176 20680 5228
rect 21916 5176 21968 5228
rect 14648 5108 14700 5117
rect 15292 5108 15344 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16304 5108 16356 5160
rect 16488 5108 16540 5160
rect 17224 5108 17276 5160
rect 20996 5151 21048 5160
rect 15476 5040 15528 5092
rect 18144 5040 18196 5092
rect 19892 5040 19944 5092
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 21364 5040 21416 5092
rect 12532 5015 12584 5024
rect 12532 4981 12541 5015
rect 12541 4981 12575 5015
rect 12575 4981 12584 5015
rect 12532 4972 12584 4981
rect 12716 4972 12768 5024
rect 13636 4972 13688 5024
rect 15384 4972 15436 5024
rect 15660 4972 15712 5024
rect 17500 4972 17552 5024
rect 20904 4972 20956 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 1768 4768 1820 4820
rect 4620 4811 4672 4820
rect 4620 4777 4629 4811
rect 4629 4777 4663 4811
rect 4663 4777 4672 4811
rect 4620 4768 4672 4777
rect 5908 4768 5960 4820
rect 2964 4632 3016 4684
rect 4344 4675 4396 4684
rect 4344 4641 4353 4675
rect 4353 4641 4387 4675
rect 4387 4641 4396 4675
rect 4344 4632 4396 4641
rect 5448 4675 5500 4684
rect 5448 4641 5457 4675
rect 5457 4641 5491 4675
rect 5491 4641 5500 4675
rect 6092 4675 6144 4684
rect 5448 4632 5500 4641
rect 6092 4641 6101 4675
rect 6101 4641 6135 4675
rect 6135 4641 6144 4675
rect 6092 4632 6144 4641
rect 2136 4564 2188 4616
rect 3332 4564 3384 4616
rect 4528 4564 4580 4616
rect 5264 4564 5316 4616
rect 5540 4607 5592 4616
rect 5540 4573 5549 4607
rect 5549 4573 5583 4607
rect 5583 4573 5592 4607
rect 5540 4564 5592 4573
rect 6368 4607 6420 4616
rect 6368 4573 6377 4607
rect 6377 4573 6411 4607
rect 6411 4573 6420 4607
rect 6368 4564 6420 4573
rect 2964 4496 3016 4548
rect 4252 4539 4304 4548
rect 2044 4428 2096 4480
rect 4252 4505 4261 4539
rect 4261 4505 4295 4539
rect 4295 4505 4304 4539
rect 4252 4496 4304 4505
rect 4344 4496 4396 4548
rect 5356 4496 5408 4548
rect 6644 4700 6696 4752
rect 7012 4675 7064 4684
rect 7012 4641 7021 4675
rect 7021 4641 7055 4675
rect 7055 4641 7064 4675
rect 7012 4632 7064 4641
rect 8484 4700 8536 4752
rect 9312 4700 9364 4752
rect 9680 4768 9732 4820
rect 10876 4768 10928 4820
rect 11060 4768 11112 4820
rect 11428 4768 11480 4820
rect 11888 4768 11940 4820
rect 12348 4768 12400 4820
rect 12440 4768 12492 4820
rect 12808 4768 12860 4820
rect 12900 4768 12952 4820
rect 13452 4768 13504 4820
rect 6552 4564 6604 4616
rect 8208 4632 8260 4684
rect 9956 4632 10008 4684
rect 10048 4632 10100 4684
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 7932 4564 7984 4616
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 12164 4743 12216 4752
rect 12164 4709 12173 4743
rect 12173 4709 12207 4743
rect 12207 4709 12216 4743
rect 12164 4700 12216 4709
rect 14740 4700 14792 4752
rect 11612 4675 11664 4684
rect 11612 4641 11621 4675
rect 11621 4641 11655 4675
rect 11655 4641 11664 4675
rect 11612 4632 11664 4641
rect 11704 4632 11756 4684
rect 11980 4632 12032 4684
rect 12348 4564 12400 4616
rect 12532 4632 12584 4684
rect 12808 4632 12860 4684
rect 12900 4632 12952 4684
rect 13176 4632 13228 4684
rect 13636 4675 13688 4684
rect 13636 4641 13645 4675
rect 13645 4641 13679 4675
rect 13679 4641 13688 4675
rect 13636 4632 13688 4641
rect 14188 4632 14240 4684
rect 13544 4607 13596 4616
rect 13544 4573 13553 4607
rect 13553 4573 13587 4607
rect 13587 4573 13596 4607
rect 13544 4564 13596 4573
rect 14096 4564 14148 4616
rect 17224 4768 17276 4820
rect 18328 4768 18380 4820
rect 18420 4768 18472 4820
rect 15660 4700 15712 4752
rect 17408 4700 17460 4752
rect 19064 4768 19116 4820
rect 20260 4768 20312 4820
rect 22744 4768 22796 4820
rect 15108 4632 15160 4684
rect 19892 4675 19944 4684
rect 15384 4564 15436 4616
rect 16488 4564 16540 4616
rect 8576 4496 8628 4548
rect 8760 4496 8812 4548
rect 9496 4496 9548 4548
rect 9864 4496 9916 4548
rect 10232 4496 10284 4548
rect 11612 4496 11664 4548
rect 11980 4496 12032 4548
rect 19892 4641 19901 4675
rect 19901 4641 19935 4675
rect 19935 4641 19944 4675
rect 19892 4632 19944 4641
rect 20904 4675 20956 4684
rect 20904 4641 20913 4675
rect 20913 4641 20947 4675
rect 20947 4641 20956 4675
rect 20904 4632 20956 4641
rect 21548 4632 21600 4684
rect 17500 4539 17552 4548
rect 17500 4505 17509 4539
rect 17509 4505 17543 4539
rect 17543 4505 17552 4539
rect 17500 4496 17552 4505
rect 22008 4564 22060 4616
rect 17960 4539 18012 4548
rect 3792 4471 3844 4480
rect 3792 4437 3801 4471
rect 3801 4437 3835 4471
rect 3835 4437 3844 4471
rect 3792 4428 3844 4437
rect 5816 4428 5868 4480
rect 7288 4428 7340 4480
rect 7656 4428 7708 4480
rect 8300 4428 8352 4480
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 9312 4428 9364 4480
rect 9772 4428 9824 4480
rect 10600 4428 10652 4480
rect 10968 4428 11020 4480
rect 11244 4428 11296 4480
rect 12072 4471 12124 4480
rect 12072 4437 12081 4471
rect 12081 4437 12115 4471
rect 12115 4437 12124 4471
rect 12072 4428 12124 4437
rect 12164 4428 12216 4480
rect 12532 4428 12584 4480
rect 13176 4471 13228 4480
rect 13176 4437 13185 4471
rect 13185 4437 13219 4471
rect 13219 4437 13228 4471
rect 14280 4471 14332 4480
rect 13176 4428 13228 4437
rect 14280 4437 14289 4471
rect 14289 4437 14323 4471
rect 14323 4437 14332 4471
rect 14280 4428 14332 4437
rect 14556 4471 14608 4480
rect 14556 4437 14565 4471
rect 14565 4437 14599 4471
rect 14599 4437 14608 4471
rect 14556 4428 14608 4437
rect 14740 4428 14792 4480
rect 16948 4428 17000 4480
rect 17408 4471 17460 4480
rect 17408 4437 17417 4471
rect 17417 4437 17451 4471
rect 17451 4437 17460 4471
rect 17408 4428 17460 4437
rect 17960 4505 17994 4539
rect 17994 4505 18012 4539
rect 17960 4496 18012 4505
rect 18880 4496 18932 4548
rect 20996 4496 21048 4548
rect 21180 4496 21232 4548
rect 21548 4496 21600 4548
rect 18236 4428 18288 4480
rect 18972 4428 19024 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 5724 4267 5776 4276
rect 3792 4156 3844 4208
rect 3884 4156 3936 4208
rect 4252 4156 4304 4208
rect 5724 4233 5733 4267
rect 5733 4233 5767 4267
rect 5767 4233 5776 4267
rect 5724 4224 5776 4233
rect 6000 4224 6052 4276
rect 6644 4224 6696 4276
rect 8484 4224 8536 4276
rect 9496 4224 9548 4276
rect 9956 4224 10008 4276
rect 6736 4156 6788 4208
rect 204 4088 256 4140
rect 940 4088 992 4140
rect 1952 4131 2004 4140
rect 1952 4097 1961 4131
rect 1961 4097 1995 4131
rect 1995 4097 2004 4131
rect 1952 4088 2004 4097
rect 2228 4131 2280 4140
rect 2228 4097 2237 4131
rect 2237 4097 2271 4131
rect 2271 4097 2280 4131
rect 2228 4088 2280 4097
rect 2596 4131 2648 4140
rect 2596 4097 2605 4131
rect 2605 4097 2639 4131
rect 2639 4097 2648 4131
rect 2596 4088 2648 4097
rect 3424 4131 3476 4140
rect 3424 4097 3433 4131
rect 3433 4097 3467 4131
rect 3467 4097 3476 4131
rect 3424 4088 3476 4097
rect 4804 4088 4856 4140
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 1768 3952 1820 4004
rect 2320 3952 2372 4004
rect 3056 3952 3108 4004
rect 4620 4020 4672 4072
rect 5080 4063 5132 4072
rect 5080 4029 5089 4063
rect 5089 4029 5123 4063
rect 5123 4029 5132 4063
rect 5080 4020 5132 4029
rect 5264 4063 5316 4072
rect 5264 4029 5273 4063
rect 5273 4029 5307 4063
rect 5307 4029 5316 4063
rect 5264 4020 5316 4029
rect 3884 3995 3936 4004
rect 3884 3961 3893 3995
rect 3893 3961 3927 3995
rect 3927 3961 3936 3995
rect 3884 3952 3936 3961
rect 1216 3884 1268 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 4804 3952 4856 4004
rect 5356 3884 5408 3936
rect 5724 4020 5776 4072
rect 5632 3952 5684 4004
rect 7196 4156 7248 4208
rect 7380 4156 7432 4208
rect 10600 4156 10652 4208
rect 7104 4131 7156 4140
rect 7104 4097 7138 4131
rect 7138 4097 7156 4131
rect 7104 4088 7156 4097
rect 8484 4088 8536 4140
rect 8852 4088 8904 4140
rect 10232 4088 10284 4140
rect 10416 4131 10468 4140
rect 10416 4097 10425 4131
rect 10425 4097 10459 4131
rect 10459 4097 10468 4131
rect 10416 4088 10468 4097
rect 6828 4063 6880 4072
rect 6828 4029 6837 4063
rect 6837 4029 6871 4063
rect 6871 4029 6880 4063
rect 6828 4020 6880 4029
rect 8392 4063 8444 4072
rect 6736 3952 6788 4004
rect 8392 4029 8401 4063
rect 8401 4029 8435 4063
rect 8435 4029 8444 4063
rect 8392 4020 8444 4029
rect 8576 4063 8628 4072
rect 8576 4029 8585 4063
rect 8585 4029 8619 4063
rect 8619 4029 8628 4063
rect 8576 4020 8628 4029
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10416 3952 10468 4004
rect 10876 4224 10928 4276
rect 10784 4020 10836 4072
rect 11060 4088 11112 4140
rect 12072 4224 12124 4276
rect 12440 4224 12492 4276
rect 13176 4224 13228 4276
rect 13544 4224 13596 4276
rect 14280 4224 14332 4276
rect 15476 4267 15528 4276
rect 15476 4233 15485 4267
rect 15485 4233 15519 4267
rect 15519 4233 15528 4267
rect 15476 4224 15528 4233
rect 18880 4267 18932 4276
rect 18880 4233 18889 4267
rect 18889 4233 18923 4267
rect 18923 4233 18932 4267
rect 18880 4224 18932 4233
rect 19616 4224 19668 4276
rect 12900 4199 12952 4208
rect 12900 4165 12909 4199
rect 12909 4165 12943 4199
rect 12943 4165 12952 4199
rect 12900 4156 12952 4165
rect 14004 4156 14056 4208
rect 15568 4156 15620 4208
rect 11428 4088 11480 4140
rect 12164 4088 12216 4140
rect 12440 4088 12492 4140
rect 12808 4088 12860 4140
rect 11520 4020 11572 4072
rect 12256 4020 12308 4072
rect 12532 4020 12584 4072
rect 13360 4020 13412 4072
rect 13912 4088 13964 4140
rect 15476 4088 15528 4140
rect 14372 4020 14424 4072
rect 14648 4063 14700 4072
rect 14648 4029 14657 4063
rect 14657 4029 14691 4063
rect 14691 4029 14700 4063
rect 14648 4020 14700 4029
rect 15292 4063 15344 4072
rect 6460 3884 6512 3936
rect 10784 3884 10836 3936
rect 13728 3952 13780 4004
rect 14188 3952 14240 4004
rect 15292 4029 15301 4063
rect 15301 4029 15335 4063
rect 15335 4029 15344 4063
rect 17500 4156 17552 4208
rect 18052 4156 18104 4208
rect 17224 4088 17276 4140
rect 18512 4131 18564 4140
rect 15292 4020 15344 4029
rect 15108 3952 15160 4004
rect 16120 3995 16172 4004
rect 11152 3884 11204 3936
rect 11244 3884 11296 3936
rect 11704 3884 11756 3936
rect 13820 3884 13872 3936
rect 14464 3884 14516 3936
rect 15844 3927 15896 3936
rect 15844 3893 15853 3927
rect 15853 3893 15887 3927
rect 15887 3893 15896 3927
rect 15844 3884 15896 3893
rect 16120 3961 16129 3995
rect 16129 3961 16163 3995
rect 16163 3961 16172 3995
rect 16120 3952 16172 3961
rect 16580 3952 16632 4004
rect 18512 4097 18521 4131
rect 18521 4097 18555 4131
rect 18555 4097 18564 4131
rect 18512 4088 18564 4097
rect 20720 4224 20772 4276
rect 20168 4088 20220 4140
rect 21640 4088 21692 4140
rect 18788 4020 18840 4072
rect 18972 4020 19024 4072
rect 17040 3884 17092 3936
rect 18236 3884 18288 3936
rect 18972 3884 19024 3936
rect 19064 3884 19116 3936
rect 19340 4020 19392 4072
rect 19616 4020 19668 4072
rect 20260 4063 20312 4072
rect 20260 4029 20269 4063
rect 20269 4029 20303 4063
rect 20303 4029 20312 4063
rect 20260 4020 20312 4029
rect 20352 4063 20404 4072
rect 20352 4029 20361 4063
rect 20361 4029 20395 4063
rect 20395 4029 20404 4063
rect 20352 4020 20404 4029
rect 21824 4020 21876 4072
rect 20720 3884 20772 3936
rect 21732 3884 21784 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2964 3680 3016 3732
rect 5172 3680 5224 3732
rect 5724 3680 5776 3732
rect 2780 3612 2832 3664
rect 6000 3612 6052 3664
rect 2688 3544 2740 3596
rect 4160 3587 4212 3596
rect 4160 3553 4169 3587
rect 4169 3553 4203 3587
rect 4203 3553 4212 3587
rect 4160 3544 4212 3553
rect 4620 3544 4672 3596
rect 5448 3587 5500 3596
rect 5448 3553 5457 3587
rect 5457 3553 5491 3587
rect 5491 3553 5500 3587
rect 5448 3544 5500 3553
rect 5724 3544 5776 3596
rect 6092 3587 6144 3596
rect 6092 3553 6101 3587
rect 6101 3553 6135 3587
rect 6135 3553 6144 3587
rect 6092 3544 6144 3553
rect 6276 3587 6328 3596
rect 6276 3553 6285 3587
rect 6285 3553 6319 3587
rect 6319 3553 6328 3587
rect 6276 3544 6328 3553
rect 6828 3680 6880 3732
rect 7104 3680 7156 3732
rect 8576 3680 8628 3732
rect 9864 3680 9916 3732
rect 10508 3680 10560 3732
rect 10784 3680 10836 3732
rect 12256 3680 12308 3732
rect 13360 3723 13412 3732
rect 7932 3612 7984 3664
rect 10140 3612 10192 3664
rect 11796 3612 11848 3664
rect 13360 3689 13369 3723
rect 13369 3689 13403 3723
rect 13403 3689 13412 3723
rect 13360 3680 13412 3689
rect 13452 3680 13504 3732
rect 15476 3680 15528 3732
rect 18788 3723 18840 3732
rect 14832 3612 14884 3664
rect 17960 3655 18012 3664
rect 17960 3621 17969 3655
rect 17969 3621 18003 3655
rect 18003 3621 18012 3655
rect 17960 3612 18012 3621
rect 8300 3587 8352 3596
rect 8300 3553 8309 3587
rect 8309 3553 8343 3587
rect 8343 3553 8352 3587
rect 8300 3544 8352 3553
rect 940 3476 992 3528
rect 2872 3519 2924 3528
rect 2872 3485 2881 3519
rect 2881 3485 2915 3519
rect 2915 3485 2924 3519
rect 2872 3476 2924 3485
rect 1032 3408 1084 3460
rect 4528 3476 4580 3528
rect 4712 3476 4764 3528
rect 9312 3544 9364 3596
rect 8944 3476 8996 3528
rect 11612 3544 11664 3596
rect 11888 3544 11940 3596
rect 4252 3408 4304 3460
rect 3976 3340 4028 3392
rect 4712 3383 4764 3392
rect 4712 3349 4721 3383
rect 4721 3349 4755 3383
rect 4755 3349 4764 3383
rect 4712 3340 4764 3349
rect 6460 3408 6512 3460
rect 7748 3408 7800 3460
rect 8208 3408 8260 3460
rect 5172 3383 5224 3392
rect 5172 3349 5181 3383
rect 5181 3349 5215 3383
rect 5215 3349 5224 3383
rect 5172 3340 5224 3349
rect 5448 3340 5500 3392
rect 5816 3340 5868 3392
rect 6644 3340 6696 3392
rect 6828 3340 6880 3392
rect 9128 3408 9180 3460
rect 13544 3544 13596 3596
rect 14648 3587 14700 3596
rect 14648 3553 14657 3587
rect 14657 3553 14691 3587
rect 14691 3553 14700 3587
rect 14648 3544 14700 3553
rect 15292 3544 15344 3596
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 18788 3689 18797 3723
rect 18797 3689 18831 3723
rect 18831 3689 18840 3723
rect 18788 3680 18840 3689
rect 19064 3680 19116 3732
rect 19616 3680 19668 3732
rect 22836 3680 22888 3732
rect 19524 3612 19576 3664
rect 20076 3612 20128 3664
rect 20260 3612 20312 3664
rect 19708 3587 19760 3596
rect 9680 3408 9732 3460
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 9404 3383 9456 3392
rect 9404 3349 9413 3383
rect 9413 3349 9447 3383
rect 9447 3349 9456 3383
rect 9772 3383 9824 3392
rect 9404 3340 9456 3349
rect 9772 3349 9781 3383
rect 9781 3349 9815 3383
rect 9815 3349 9824 3383
rect 9772 3340 9824 3349
rect 9956 3408 10008 3460
rect 11060 3408 11112 3460
rect 12716 3476 12768 3528
rect 13728 3519 13780 3528
rect 12440 3408 12492 3460
rect 13728 3485 13737 3519
rect 13737 3485 13771 3519
rect 13771 3485 13780 3519
rect 13728 3476 13780 3485
rect 14464 3519 14516 3528
rect 14464 3485 14473 3519
rect 14473 3485 14507 3519
rect 14507 3485 14516 3519
rect 14464 3476 14516 3485
rect 15476 3476 15528 3528
rect 15936 3476 15988 3528
rect 13728 3340 13780 3392
rect 13820 3340 13872 3392
rect 14924 3408 14976 3460
rect 16028 3451 16080 3460
rect 16028 3417 16037 3451
rect 16037 3417 16071 3451
rect 16071 3417 16080 3451
rect 16028 3408 16080 3417
rect 17408 3476 17460 3528
rect 17776 3476 17828 3528
rect 19708 3553 19717 3587
rect 19717 3553 19751 3587
rect 19751 3553 19760 3587
rect 19708 3544 19760 3553
rect 18604 3476 18656 3528
rect 19156 3476 19208 3528
rect 20352 3544 20404 3596
rect 20076 3519 20128 3528
rect 20076 3485 20085 3519
rect 20085 3485 20119 3519
rect 20119 3485 20128 3519
rect 20076 3476 20128 3485
rect 20444 3519 20496 3528
rect 20444 3485 20453 3519
rect 20453 3485 20487 3519
rect 20487 3485 20496 3519
rect 20444 3476 20496 3485
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 22008 3476 22060 3528
rect 17960 3408 18012 3460
rect 19524 3408 19576 3460
rect 15936 3383 15988 3392
rect 15936 3349 15945 3383
rect 15945 3349 15979 3383
rect 15979 3349 15988 3383
rect 15936 3340 15988 3349
rect 16304 3383 16356 3392
rect 16304 3349 16313 3383
rect 16313 3349 16347 3383
rect 16347 3349 16356 3383
rect 16304 3340 16356 3349
rect 18420 3383 18472 3392
rect 18420 3349 18429 3383
rect 18429 3349 18463 3383
rect 18463 3349 18472 3383
rect 18420 3340 18472 3349
rect 18788 3340 18840 3392
rect 19616 3383 19668 3392
rect 19616 3349 19625 3383
rect 19625 3349 19659 3383
rect 19659 3349 19668 3383
rect 19616 3340 19668 3349
rect 19800 3340 19852 3392
rect 21364 3383 21416 3392
rect 21364 3349 21373 3383
rect 21373 3349 21407 3383
rect 21407 3349 21416 3383
rect 21364 3340 21416 3349
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 5816 3136 5868 3188
rect 6552 3136 6604 3188
rect 6736 3136 6788 3188
rect 7840 3136 7892 3188
rect 8208 3136 8260 3188
rect 8944 3136 8996 3188
rect 9036 3136 9088 3188
rect 9496 3136 9548 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 10140 3136 10192 3188
rect 10784 3136 10836 3188
rect 11244 3136 11296 3188
rect 14924 3179 14976 3188
rect 2596 3111 2648 3120
rect 2596 3077 2605 3111
rect 2605 3077 2639 3111
rect 2639 3077 2648 3111
rect 2596 3068 2648 3077
rect 3056 3068 3108 3120
rect 8300 3068 8352 3120
rect 9772 3111 9824 3120
rect 9772 3077 9781 3111
rect 9781 3077 9815 3111
rect 9815 3077 9824 3111
rect 9772 3068 9824 3077
rect 11336 3068 11388 3120
rect 11796 3068 11848 3120
rect 12348 3068 12400 3120
rect 572 3000 624 3052
rect 2412 3000 2464 3052
rect 4160 3000 4212 3052
rect 4436 3000 4488 3052
rect 4804 3043 4856 3052
rect 4804 3009 4838 3043
rect 4838 3009 4856 3043
rect 4804 3000 4856 3009
rect 5356 3000 5408 3052
rect 1952 2975 2004 2984
rect 1952 2941 1961 2975
rect 1961 2941 1995 2975
rect 1995 2941 2004 2975
rect 1952 2932 2004 2941
rect 2964 2864 3016 2916
rect 4068 2796 4120 2848
rect 6092 3000 6144 3052
rect 7656 3000 7708 3052
rect 7932 3000 7984 3052
rect 9128 3043 9180 3052
rect 9128 3009 9137 3043
rect 9137 3009 9171 3043
rect 9171 3009 9180 3043
rect 9128 3000 9180 3009
rect 5632 2932 5684 2984
rect 6828 2932 6880 2984
rect 7104 2975 7156 2984
rect 7104 2941 7113 2975
rect 7113 2941 7147 2975
rect 7147 2941 7156 2975
rect 7104 2932 7156 2941
rect 8024 2932 8076 2984
rect 6552 2864 6604 2916
rect 11336 2975 11388 2984
rect 11336 2941 11345 2975
rect 11345 2941 11379 2975
rect 11379 2941 11388 2975
rect 11336 2932 11388 2941
rect 5908 2839 5960 2848
rect 5908 2805 5917 2839
rect 5917 2805 5951 2839
rect 5951 2805 5960 2839
rect 5908 2796 5960 2805
rect 6000 2796 6052 2848
rect 7012 2796 7064 2848
rect 7748 2839 7800 2848
rect 7748 2805 7757 2839
rect 7757 2805 7791 2839
rect 7791 2805 7800 2839
rect 7748 2796 7800 2805
rect 9864 2864 9916 2916
rect 11520 3000 11572 3052
rect 11796 2932 11848 2984
rect 13360 3068 13412 3120
rect 12716 3043 12768 3052
rect 12716 3009 12725 3043
rect 12725 3009 12759 3043
rect 12759 3009 12768 3043
rect 12716 3000 12768 3009
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 15200 3136 15252 3188
rect 18512 3179 18564 3188
rect 15016 3068 15068 3120
rect 12624 2932 12676 2984
rect 13728 2932 13780 2984
rect 14832 3000 14884 3052
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15752 3043 15804 3052
rect 15752 3009 15761 3043
rect 15761 3009 15795 3043
rect 15795 3009 15804 3043
rect 15752 3000 15804 3009
rect 16212 3043 16264 3052
rect 16212 3009 16221 3043
rect 16221 3009 16255 3043
rect 16255 3009 16264 3043
rect 16212 3000 16264 3009
rect 16028 2932 16080 2984
rect 16948 3043 17000 3052
rect 16948 3009 16957 3043
rect 16957 3009 16991 3043
rect 16991 3009 17000 3043
rect 17316 3043 17368 3052
rect 16948 3000 17000 3009
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 17592 3000 17644 3052
rect 18052 3111 18104 3120
rect 18052 3077 18061 3111
rect 18061 3077 18095 3111
rect 18095 3077 18104 3111
rect 18052 3068 18104 3077
rect 17776 2975 17828 2984
rect 17776 2941 17785 2975
rect 17785 2941 17819 2975
rect 17819 2941 17828 2975
rect 17776 2932 17828 2941
rect 18236 3000 18288 3052
rect 8484 2796 8536 2848
rect 10048 2796 10100 2848
rect 10140 2796 10192 2848
rect 11428 2796 11480 2848
rect 11704 2796 11756 2848
rect 12440 2796 12492 2848
rect 14648 2864 14700 2916
rect 15200 2907 15252 2916
rect 15200 2873 15209 2907
rect 15209 2873 15243 2907
rect 15243 2873 15252 2907
rect 15200 2864 15252 2873
rect 15568 2907 15620 2916
rect 15568 2873 15577 2907
rect 15577 2873 15611 2907
rect 15611 2873 15620 2907
rect 15568 2864 15620 2873
rect 14280 2796 14332 2848
rect 14464 2839 14516 2848
rect 14464 2805 14473 2839
rect 14473 2805 14507 2839
rect 14507 2805 14516 2839
rect 14464 2796 14516 2805
rect 16672 2839 16724 2848
rect 16672 2805 16681 2839
rect 16681 2805 16715 2839
rect 16715 2805 16724 2839
rect 16672 2796 16724 2805
rect 17224 2796 17276 2848
rect 17316 2796 17368 2848
rect 18512 3145 18521 3179
rect 18521 3145 18555 3179
rect 18555 3145 18564 3179
rect 18512 3136 18564 3145
rect 18880 3136 18932 3188
rect 21088 3136 21140 3188
rect 19800 3068 19852 3120
rect 20628 3111 20680 3120
rect 20628 3077 20637 3111
rect 20637 3077 20671 3111
rect 20671 3077 20680 3111
rect 20628 3068 20680 3077
rect 18972 3000 19024 3052
rect 19156 2975 19208 2984
rect 19156 2941 19165 2975
rect 19165 2941 19199 2975
rect 19199 2941 19208 2975
rect 19156 2932 19208 2941
rect 19708 2932 19760 2984
rect 19984 3000 20036 3052
rect 20720 3043 20772 3052
rect 20720 3009 20729 3043
rect 20729 3009 20763 3043
rect 20763 3009 20772 3043
rect 20720 3000 20772 3009
rect 20536 2932 20588 2984
rect 19064 2864 19116 2916
rect 20628 2864 20680 2916
rect 18512 2796 18564 2848
rect 18604 2796 18656 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 5724 2592 5776 2644
rect 6092 2592 6144 2644
rect 6920 2592 6972 2644
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 7564 2524 7616 2576
rect 7656 2524 7708 2576
rect 12716 2592 12768 2644
rect 9312 2524 9364 2576
rect 10692 2524 10744 2576
rect 12072 2524 12124 2576
rect 2228 2456 2280 2508
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 2780 2456 2832 2508
rect 5816 2499 5868 2508
rect 5816 2465 5825 2499
rect 5825 2465 5859 2499
rect 5859 2465 5868 2499
rect 5816 2456 5868 2465
rect 7012 2456 7064 2508
rect 8116 2456 8168 2508
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 2412 2431 2464 2440
rect 2412 2397 2421 2431
rect 2421 2397 2455 2431
rect 2455 2397 2464 2431
rect 2412 2388 2464 2397
rect 3884 2388 3936 2440
rect 4804 2388 4856 2440
rect 7196 2431 7248 2440
rect 7196 2397 7205 2431
rect 7205 2397 7239 2431
rect 7239 2397 7248 2431
rect 7196 2388 7248 2397
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 4436 2320 4488 2372
rect 7288 2320 7340 2372
rect 8760 2388 8812 2440
rect 9496 2388 9548 2440
rect 9772 2456 9824 2508
rect 10784 2499 10836 2508
rect 10784 2465 10793 2499
rect 10793 2465 10827 2499
rect 10827 2465 10836 2499
rect 10784 2456 10836 2465
rect 10876 2456 10928 2508
rect 11704 2456 11756 2508
rect 13084 2524 13136 2576
rect 9588 2320 9640 2372
rect 10508 2388 10560 2440
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 11152 2388 11204 2440
rect 11888 2431 11940 2440
rect 11888 2397 11897 2431
rect 11897 2397 11931 2431
rect 11931 2397 11940 2431
rect 11888 2388 11940 2397
rect 12532 2456 12584 2508
rect 14280 2592 14332 2644
rect 15936 2592 15988 2644
rect 13820 2524 13872 2576
rect 14004 2524 14056 2576
rect 14832 2524 14884 2576
rect 16028 2524 16080 2576
rect 16948 2524 17000 2576
rect 14740 2431 14792 2440
rect 14740 2397 14749 2431
rect 14749 2397 14783 2431
rect 14783 2397 14792 2431
rect 14740 2388 14792 2397
rect 16672 2456 16724 2508
rect 14464 2320 14516 2372
rect 14556 2320 14608 2372
rect 15936 2431 15988 2440
rect 15936 2397 15945 2431
rect 15945 2397 15979 2431
rect 15979 2397 15988 2431
rect 15936 2388 15988 2397
rect 16212 2388 16264 2440
rect 18420 2592 18472 2644
rect 19892 2592 19944 2644
rect 18236 2456 18288 2508
rect 18328 2499 18380 2508
rect 18328 2465 18337 2499
rect 18337 2465 18371 2499
rect 18371 2465 18380 2499
rect 20996 2524 21048 2576
rect 21732 2524 21784 2576
rect 22652 2524 22704 2576
rect 18328 2456 18380 2465
rect 18420 2431 18472 2440
rect 3884 2252 3936 2304
rect 4068 2252 4120 2304
rect 7472 2252 7524 2304
rect 8208 2252 8260 2304
rect 8576 2295 8628 2304
rect 8576 2261 8585 2295
rect 8585 2261 8619 2295
rect 8619 2261 8628 2295
rect 8576 2252 8628 2261
rect 9312 2252 9364 2304
rect 9772 2295 9824 2304
rect 9772 2261 9781 2295
rect 9781 2261 9815 2295
rect 9815 2261 9824 2295
rect 9772 2252 9824 2261
rect 12164 2252 12216 2304
rect 12440 2252 12492 2304
rect 13544 2252 13596 2304
rect 14372 2252 14424 2304
rect 15200 2252 15252 2304
rect 15752 2252 15804 2304
rect 16396 2320 16448 2372
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 22192 2456 22244 2508
rect 19064 2431 19116 2440
rect 18420 2388 18472 2397
rect 19064 2397 19073 2431
rect 19073 2397 19107 2431
rect 19107 2397 19116 2431
rect 19064 2388 19116 2397
rect 19248 2431 19300 2440
rect 19248 2397 19257 2431
rect 19257 2397 19291 2431
rect 19291 2397 19300 2431
rect 19248 2388 19300 2397
rect 20352 2431 20404 2440
rect 20352 2397 20361 2431
rect 20361 2397 20395 2431
rect 20395 2397 20404 2431
rect 20352 2388 20404 2397
rect 20720 2431 20772 2440
rect 20720 2397 20729 2431
rect 20729 2397 20763 2431
rect 20763 2397 20772 2431
rect 20720 2388 20772 2397
rect 22560 2388 22612 2440
rect 18696 2252 18748 2304
rect 21824 2320 21876 2372
rect 18972 2252 19024 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 6000 2048 6052 2100
rect 11704 2048 11756 2100
rect 12440 2048 12492 2100
rect 16304 2048 16356 2100
rect 19248 2048 19300 2100
rect 2412 1980 2464 2032
rect 7104 1980 7156 2032
rect 8208 1980 8260 2032
rect 9220 1980 9272 2032
rect 17776 1980 17828 2032
rect 20352 1980 20404 2032
rect 848 1912 900 1964
rect 4804 1912 4856 1964
rect 8300 1912 8352 1964
rect 11888 1912 11940 1964
rect 12624 1912 12676 1964
rect 1952 1844 2004 1896
rect 5908 1844 5960 1896
rect 10876 1844 10928 1896
rect 16120 1844 16172 1896
rect 19248 1844 19300 1896
rect 21824 1844 21876 1896
rect 22376 1844 22428 1896
rect 2872 1776 2924 1828
rect 10692 1776 10744 1828
rect 15016 1776 15068 1828
rect 19064 1776 19116 1828
rect 3976 1708 4028 1760
rect 11060 1708 11112 1760
rect 9772 1640 9824 1692
rect 10508 1640 10560 1692
rect 11980 1640 12032 1692
rect 17224 1436 17276 1488
rect 18144 1436 18196 1488
rect 17684 1368 17736 1420
rect 18972 1368 19024 1420
rect 22008 1368 22060 1420
rect 22744 1368 22796 1420
rect 3240 1300 3292 1352
rect 10324 1300 10376 1352
rect 17132 1300 17184 1352
rect 18696 1300 18748 1352
rect 3516 1232 3568 1284
rect 5724 1232 5776 1284
rect 13176 1232 13228 1284
rect 18512 1232 18564 1284
rect 20260 1232 20312 1284
rect 3240 1164 3292 1216
rect 4528 1164 4580 1216
rect 1032 1028 1084 1080
rect 12808 1028 12860 1080
rect 7840 960 7892 1012
rect 17960 960 18012 1012
rect 6644 892 6696 944
rect 14648 892 14700 944
rect 21364 892 21416 944
<< metal2 >>
rect 202 22200 258 23000
rect 294 22944 350 22953
rect 294 22879 350 22888
rect 20 21684 72 21690
rect 20 21626 72 21632
rect 32 7886 60 21626
rect 216 17864 244 22200
rect 124 17836 244 17864
rect 124 14482 152 17836
rect 112 14476 164 14482
rect 112 14418 164 14424
rect 20 7880 72 7886
rect 20 7822 72 7828
rect 308 6914 336 22879
rect 570 22200 626 23000
rect 938 22200 994 23000
rect 1030 22536 1086 22545
rect 1030 22471 1086 22480
rect 584 18154 612 22200
rect 848 22092 900 22098
rect 848 22034 900 22040
rect 860 18902 888 22034
rect 952 20806 980 22200
rect 1044 22098 1072 22471
rect 1122 22400 1178 22409
rect 1122 22335 1178 22344
rect 1032 22092 1084 22098
rect 1032 22034 1084 22040
rect 1030 21992 1086 22001
rect 1030 21927 1086 21936
rect 940 20800 992 20806
rect 940 20742 992 20748
rect 1044 19156 1072 21927
rect 952 19128 1072 19156
rect 848 18896 900 18902
rect 848 18838 900 18844
rect 572 18148 624 18154
rect 572 18090 624 18096
rect 846 14070 902 14079
rect 846 14005 902 14014
rect 388 10804 440 10810
rect 388 10746 440 10752
rect 216 6886 336 6914
rect 216 4146 244 6886
rect 294 6760 350 6769
rect 294 6695 350 6704
rect 204 4140 256 4146
rect 204 4082 256 4088
rect 308 3482 336 6695
rect 400 6390 428 10746
rect 860 9518 888 14005
rect 848 9512 900 9518
rect 848 9454 900 9460
rect 756 7540 808 7546
rect 756 7482 808 7488
rect 388 6384 440 6390
rect 388 6326 440 6332
rect 216 3454 336 3482
rect 216 800 244 3454
rect 572 3052 624 3058
rect 572 2994 624 3000
rect 584 800 612 2994
rect 202 0 258 800
rect 570 0 626 800
rect 768 354 796 7482
rect 952 6914 980 19128
rect 1136 18986 1164 22335
rect 1306 22200 1362 23000
rect 1674 22200 1730 23000
rect 2042 22200 2098 23000
rect 2410 22672 2466 22681
rect 2410 22607 2466 22616
rect 1214 20904 1270 20913
rect 1214 20839 1270 20848
rect 1044 18958 1164 18986
rect 1044 10985 1072 18958
rect 1124 18896 1176 18902
rect 1124 18838 1176 18844
rect 1030 10976 1086 10985
rect 1030 10911 1086 10920
rect 1032 9512 1084 9518
rect 1030 9480 1032 9489
rect 1084 9480 1086 9489
rect 1030 9415 1086 9424
rect 1032 7880 1084 7886
rect 1030 7848 1032 7857
rect 1084 7848 1086 7857
rect 1030 7783 1086 7792
rect 1030 7712 1086 7721
rect 1030 7647 1086 7656
rect 860 6886 980 6914
rect 860 1970 888 6886
rect 1044 6866 1072 7647
rect 1032 6860 1084 6866
rect 1032 6802 1084 6808
rect 940 6384 992 6390
rect 940 6326 992 6332
rect 952 6089 980 6326
rect 938 6080 994 6089
rect 938 6015 994 6024
rect 1136 4593 1164 18838
rect 1122 4584 1178 4593
rect 1122 4519 1178 4528
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 4049 980 4082
rect 938 4040 994 4049
rect 938 3975 994 3984
rect 952 3534 980 3975
rect 1228 3942 1256 20839
rect 1320 20466 1348 22200
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1308 20460 1360 20466
rect 1308 20402 1360 20408
rect 1320 19009 1348 20402
rect 1306 19000 1362 19009
rect 1306 18935 1362 18944
rect 1412 14890 1440 21490
rect 1582 20224 1638 20233
rect 1582 20159 1638 20168
rect 1596 20058 1624 20159
rect 1584 20052 1636 20058
rect 1584 19994 1636 20000
rect 1492 19848 1544 19854
rect 1490 19816 1492 19825
rect 1544 19816 1546 19825
rect 1688 19802 1716 22200
rect 1766 21040 1822 21049
rect 1766 20975 1822 20984
rect 1490 19751 1546 19760
rect 1596 19774 1716 19802
rect 1492 19712 1544 19718
rect 1490 19680 1492 19689
rect 1544 19680 1546 19689
rect 1490 19615 1546 19624
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1490 18864 1546 18873
rect 1490 18799 1546 18808
rect 1596 18737 1624 19774
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 18766 1716 19654
rect 1780 18970 1808 20975
rect 2056 20482 2084 22200
rect 2226 21856 2282 21865
rect 2226 21791 2282 21800
rect 1872 20454 2084 20482
rect 1872 19496 1900 20454
rect 1952 20392 2004 20398
rect 1952 20334 2004 20340
rect 2042 20360 2098 20369
rect 1964 19689 1992 20334
rect 2042 20295 2098 20304
rect 2056 19854 2084 20295
rect 2044 19848 2096 19854
rect 2044 19790 2096 19796
rect 1950 19680 2006 19689
rect 1950 19615 2006 19624
rect 1872 19468 2176 19496
rect 1950 19408 2006 19417
rect 1950 19343 1952 19352
rect 2004 19343 2006 19352
rect 2044 19372 2096 19378
rect 1952 19314 2004 19320
rect 2044 19314 2096 19320
rect 1858 19272 1914 19281
rect 1858 19207 1860 19216
rect 1912 19207 1914 19216
rect 1860 19178 1912 19184
rect 1768 18964 1820 18970
rect 1768 18906 1820 18912
rect 1676 18760 1728 18766
rect 1582 18728 1638 18737
rect 1676 18702 1728 18708
rect 1582 18663 1638 18672
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1676 18284 1728 18290
rect 1676 18226 1728 18232
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17649 1532 18022
rect 1688 17882 1716 18226
rect 1860 18080 1912 18086
rect 1858 18048 1860 18057
rect 1912 18048 1914 18057
rect 1858 17983 1914 17992
rect 2056 17882 2084 19314
rect 2148 18578 2176 19468
rect 2240 18970 2268 21791
rect 2318 21720 2374 21729
rect 2318 21655 2374 21664
rect 2332 19378 2360 21655
rect 2320 19372 2372 19378
rect 2320 19314 2372 19320
rect 2318 19272 2374 19281
rect 2318 19207 2374 19216
rect 2228 18964 2280 18970
rect 2228 18906 2280 18912
rect 2332 18766 2360 19207
rect 2424 18970 2452 22607
rect 2502 22200 2558 23000
rect 2870 22200 2926 23000
rect 3238 22200 3294 23000
rect 3606 22200 3662 23000
rect 3974 22200 4030 23000
rect 4158 22264 4214 22273
rect 2516 21554 2544 22200
rect 2504 21548 2556 21554
rect 2504 21490 2556 21496
rect 2596 21480 2648 21486
rect 2502 21448 2558 21457
rect 2596 21422 2648 21428
rect 2502 21383 2558 21392
rect 2516 19378 2544 21383
rect 2608 19836 2636 21422
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2688 21072 2740 21078
rect 2688 21014 2740 21020
rect 2700 19990 2728 21014
rect 2688 19984 2740 19990
rect 2688 19926 2740 19932
rect 2608 19808 2728 19836
rect 2596 19508 2648 19514
rect 2596 19450 2648 19456
rect 2504 19372 2556 19378
rect 2504 19314 2556 19320
rect 2412 18964 2464 18970
rect 2412 18906 2464 18912
rect 2320 18760 2372 18766
rect 2320 18702 2372 18708
rect 2148 18550 2268 18578
rect 2134 18456 2190 18465
rect 2134 18391 2190 18400
rect 2148 18086 2176 18391
rect 2136 18080 2188 18086
rect 2134 18048 2136 18057
rect 2188 18048 2190 18057
rect 2134 17983 2190 17992
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 2044 17876 2096 17882
rect 2044 17818 2096 17824
rect 1950 17776 2006 17785
rect 1768 17740 1820 17746
rect 1950 17711 2006 17720
rect 1768 17682 1820 17688
rect 1490 17640 1546 17649
rect 1490 17575 1546 17584
rect 1492 17536 1544 17542
rect 1492 17478 1544 17484
rect 1504 17241 1532 17478
rect 1780 17338 1808 17682
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1490 17232 1546 17241
rect 1490 17167 1546 17176
rect 1676 17196 1728 17202
rect 1676 17138 1728 17144
rect 1492 16992 1544 16998
rect 1492 16934 1544 16940
rect 1504 16833 1532 16934
rect 1490 16824 1546 16833
rect 1688 16794 1716 17138
rect 1490 16759 1546 16768
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1780 16726 1808 17274
rect 1860 17196 1912 17202
rect 1860 17138 1912 17144
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1504 16289 1532 16390
rect 1490 16280 1546 16289
rect 1490 16215 1546 16224
rect 1688 16114 1716 16390
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1780 16046 1808 16662
rect 1872 16574 1900 17138
rect 1964 17066 1992 17711
rect 2044 17604 2096 17610
rect 2044 17546 2096 17552
rect 1952 17060 2004 17066
rect 1952 17002 2004 17008
rect 1872 16546 1992 16574
rect 1768 16040 1820 16046
rect 1768 15982 1820 15988
rect 1492 15904 1544 15910
rect 1490 15872 1492 15881
rect 1544 15872 1546 15881
rect 1490 15807 1546 15816
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1858 15464 1914 15473
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15065 1532 15302
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1584 14952 1636 14958
rect 1584 14894 1636 14900
rect 1400 14884 1452 14890
rect 1400 14826 1452 14832
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14657 1532 14758
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1596 14362 1624 14894
rect 1688 14890 1716 15438
rect 1858 15399 1914 15408
rect 1872 15366 1900 15399
rect 1860 15360 1912 15366
rect 1860 15302 1912 15308
rect 1676 14884 1728 14890
rect 1676 14826 1728 14832
rect 1674 14512 1730 14521
rect 1674 14447 1730 14456
rect 1412 14334 1624 14362
rect 1308 12232 1360 12238
rect 1412 12209 1440 14334
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1492 13728 1544 13734
rect 1492 13670 1544 13676
rect 1504 13433 1532 13670
rect 1490 13424 1546 13433
rect 1688 13410 1716 14447
rect 1964 14362 1992 16546
rect 2056 16522 2084 17546
rect 2240 17377 2268 18550
rect 2608 18426 2636 19450
rect 2700 18766 2728 19808
rect 2792 19378 2820 21286
rect 2884 20754 2912 22200
rect 3148 20936 3200 20942
rect 3148 20878 3200 20884
rect 3056 20800 3108 20806
rect 2884 20726 3004 20754
rect 3056 20742 3108 20748
rect 2870 20632 2926 20641
rect 2870 20567 2926 20576
rect 2884 19446 2912 20567
rect 2872 19440 2924 19446
rect 2872 19382 2924 19388
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2872 19304 2924 19310
rect 2872 19246 2924 19252
rect 2688 18760 2740 18766
rect 2688 18702 2740 18708
rect 2884 18601 2912 19246
rect 2976 19242 3004 20726
rect 3068 19281 3096 20742
rect 3054 19272 3110 19281
rect 2964 19236 3016 19242
rect 3054 19207 3110 19216
rect 2964 19178 3016 19184
rect 2870 18592 2926 18601
rect 2870 18527 2926 18536
rect 2596 18420 2648 18426
rect 2596 18362 2648 18368
rect 2872 18352 2924 18358
rect 2872 18294 2924 18300
rect 2504 18216 2556 18222
rect 2504 18158 2556 18164
rect 2320 18080 2372 18086
rect 2320 18022 2372 18028
rect 2332 17678 2360 18022
rect 2320 17672 2372 17678
rect 2320 17614 2372 17620
rect 2226 17368 2282 17377
rect 2226 17303 2282 17312
rect 2410 17232 2466 17241
rect 2410 17167 2412 17176
rect 2464 17167 2466 17176
rect 2412 17138 2464 17144
rect 2136 16992 2188 16998
rect 2136 16934 2188 16940
rect 2228 16992 2280 16998
rect 2228 16934 2280 16940
rect 2148 16561 2176 16934
rect 2240 16590 2268 16934
rect 2228 16584 2280 16590
rect 2134 16552 2190 16561
rect 2044 16516 2096 16522
rect 2516 16574 2544 18158
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2688 17740 2740 17746
rect 2688 17682 2740 17688
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2228 16526 2280 16532
rect 2424 16546 2544 16574
rect 2134 16487 2190 16496
rect 2044 16458 2096 16464
rect 2424 16182 2452 16546
rect 2502 16280 2558 16289
rect 2502 16215 2558 16224
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 2412 16176 2464 16182
rect 2412 16118 2464 16124
rect 2240 15706 2268 16118
rect 2516 15910 2544 16215
rect 2504 15904 2556 15910
rect 2504 15846 2556 15852
rect 2228 15700 2280 15706
rect 2228 15642 2280 15648
rect 2044 15496 2096 15502
rect 2044 15438 2096 15444
rect 2056 15162 2084 15438
rect 2608 15162 2636 17478
rect 2700 16425 2728 17682
rect 2792 17610 2820 18022
rect 2884 17814 2912 18294
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2780 17604 2832 17610
rect 2780 17546 2832 17552
rect 3160 17320 3188 20878
rect 3252 19854 3280 22200
rect 3620 21214 3648 22200
rect 3608 21208 3660 21214
rect 3422 21176 3478 21185
rect 3608 21150 3660 21156
rect 3422 21111 3478 21120
rect 3332 21004 3384 21010
rect 3332 20946 3384 20952
rect 3344 20466 3372 20946
rect 3332 20460 3384 20466
rect 3332 20402 3384 20408
rect 3240 19848 3292 19854
rect 3344 19825 3372 20402
rect 3240 19790 3292 19796
rect 3330 19816 3386 19825
rect 3330 19751 3386 19760
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3240 19372 3292 19378
rect 3240 19314 3292 19320
rect 3252 17513 3280 19314
rect 3344 18193 3372 19654
rect 3436 18970 3464 21111
rect 3620 20466 3648 21150
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3884 20256 3936 20262
rect 3884 20198 3936 20204
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 3608 19984 3660 19990
rect 3608 19926 3660 19932
rect 3792 19984 3844 19990
rect 3792 19926 3844 19932
rect 3620 19334 3648 19926
rect 3700 19848 3752 19854
rect 3700 19790 3752 19796
rect 3712 19378 3740 19790
rect 3804 19718 3832 19926
rect 3792 19712 3844 19718
rect 3792 19654 3844 19660
rect 3528 19310 3648 19334
rect 3700 19372 3752 19378
rect 3700 19314 3752 19320
rect 3516 19306 3648 19310
rect 3516 19304 3568 19306
rect 3516 19246 3568 19252
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 3424 18964 3476 18970
rect 3424 18906 3476 18912
rect 3700 18896 3752 18902
rect 3896 18850 3924 20198
rect 3988 19990 4016 22200
rect 4158 22199 4214 22208
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5170 22200 5226 23000
rect 5538 22200 5594 23000
rect 5906 22200 5962 23000
rect 6012 22222 6224 22250
rect 4068 21276 4120 21282
rect 4068 21218 4120 21224
rect 3976 19984 4028 19990
rect 3976 19926 4028 19932
rect 4080 19922 4108 21218
rect 4068 19916 4120 19922
rect 4068 19858 4120 19864
rect 3976 19440 4028 19446
rect 4172 19417 4200 22199
rect 4252 20800 4304 20806
rect 4252 20742 4304 20748
rect 3976 19382 4028 19388
rect 4158 19408 4214 19417
rect 3988 19174 4016 19382
rect 4158 19343 4214 19352
rect 4068 19304 4120 19310
rect 4068 19246 4120 19252
rect 3976 19168 4028 19174
rect 3976 19110 4028 19116
rect 3700 18838 3752 18844
rect 3712 18766 3740 18838
rect 3804 18822 3924 18850
rect 3700 18760 3752 18766
rect 3700 18702 3752 18708
rect 3608 18624 3660 18630
rect 3804 18601 3832 18822
rect 3988 18766 4016 19110
rect 3884 18760 3936 18766
rect 3884 18702 3936 18708
rect 3976 18760 4028 18766
rect 3976 18702 4028 18708
rect 3608 18566 3660 18572
rect 3790 18592 3846 18601
rect 3620 18426 3648 18566
rect 3790 18527 3846 18536
rect 3608 18420 3660 18426
rect 3608 18362 3660 18368
rect 3330 18184 3386 18193
rect 3330 18119 3386 18128
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3896 17882 3924 18702
rect 3332 17876 3384 17882
rect 3332 17818 3384 17824
rect 3884 17876 3936 17882
rect 3884 17818 3936 17824
rect 3344 17678 3372 17818
rect 3988 17746 4016 18702
rect 4080 18426 4108 19246
rect 4160 19236 4212 19242
rect 4160 19178 4212 19184
rect 4172 19009 4200 19178
rect 4158 19000 4214 19009
rect 4264 18970 4292 20742
rect 4356 20330 4384 22200
rect 4712 21548 4764 21554
rect 4712 21490 4764 21496
rect 4436 21140 4488 21146
rect 4436 21082 4488 21088
rect 4344 20324 4396 20330
rect 4344 20266 4396 20272
rect 4448 20040 4476 21082
rect 4620 20392 4672 20398
rect 4620 20334 4672 20340
rect 4356 20012 4476 20040
rect 4158 18935 4214 18944
rect 4252 18964 4304 18970
rect 4252 18906 4304 18912
rect 4160 18624 4212 18630
rect 4160 18566 4212 18572
rect 4068 18420 4120 18426
rect 4068 18362 4120 18368
rect 4068 18284 4120 18290
rect 4068 18226 4120 18232
rect 4080 17882 4108 18226
rect 4172 17921 4200 18566
rect 4158 17912 4214 17921
rect 4068 17876 4120 17882
rect 4356 17898 4384 20012
rect 4434 19952 4490 19961
rect 4434 19887 4490 19896
rect 4448 19689 4476 19887
rect 4434 19680 4490 19689
rect 4434 19615 4490 19624
rect 4448 18358 4476 19615
rect 4528 18828 4580 18834
rect 4528 18770 4580 18776
rect 4436 18352 4488 18358
rect 4436 18294 4488 18300
rect 4158 17847 4214 17856
rect 4264 17870 4384 17898
rect 4068 17818 4120 17824
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3332 17672 3384 17678
rect 4172 17649 4200 17847
rect 3332 17614 3384 17620
rect 4158 17640 4214 17649
rect 4158 17575 4214 17584
rect 3976 17536 4028 17542
rect 3238 17504 3294 17513
rect 3976 17478 4028 17484
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 3238 17439 3294 17448
rect 3160 17292 3372 17320
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3252 16658 3280 17138
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 2964 16516 3016 16522
rect 2964 16458 3016 16464
rect 2686 16416 2742 16425
rect 2686 16351 2742 16360
rect 2976 16250 3004 16458
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 2596 15156 2648 15162
rect 2596 15098 2648 15104
rect 2320 15020 2372 15026
rect 2320 14962 2372 14968
rect 2596 15020 2648 15026
rect 2596 14962 2648 14968
rect 2228 14408 2280 14414
rect 1964 14334 2176 14362
rect 2228 14350 2280 14356
rect 2044 14272 2096 14278
rect 2044 14214 2096 14220
rect 2056 13938 2084 14214
rect 2044 13932 2096 13938
rect 2044 13874 2096 13880
rect 1858 13832 1914 13841
rect 1858 13767 1860 13776
rect 1912 13767 1914 13776
rect 2042 13832 2098 13841
rect 2042 13767 2098 13776
rect 1860 13738 1912 13744
rect 1490 13359 1546 13368
rect 1596 13382 1716 13410
rect 1950 13424 2006 13433
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 12889 1532 13126
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12481 1532 12582
rect 1490 12472 1546 12481
rect 1490 12407 1546 12416
rect 1308 12174 1360 12180
rect 1398 12200 1454 12209
rect 1320 9654 1348 12174
rect 1398 12135 1454 12144
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11393 1532 12038
rect 1490 11384 1546 11393
rect 1490 11319 1546 11328
rect 1490 10840 1546 10849
rect 1490 10775 1546 10784
rect 1504 10742 1532 10775
rect 1492 10736 1544 10742
rect 1492 10678 1544 10684
rect 1596 10112 1624 13382
rect 1950 13359 2006 13368
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1688 12986 1716 13262
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1676 12980 1728 12986
rect 1676 12922 1728 12928
rect 1676 12844 1728 12850
rect 1676 12786 1728 12792
rect 1768 12844 1820 12850
rect 1768 12786 1820 12792
rect 1688 12102 1716 12786
rect 1780 12442 1808 12786
rect 1768 12436 1820 12442
rect 1768 12378 1820 12384
rect 1676 12096 1728 12102
rect 1676 12038 1728 12044
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1688 11218 1716 11834
rect 1780 11286 1808 12378
rect 1872 12073 1900 13126
rect 1858 12064 1914 12073
rect 1858 11999 1914 12008
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1768 11280 1820 11286
rect 1872 11257 1900 11698
rect 1768 11222 1820 11228
rect 1858 11248 1914 11257
rect 1676 11212 1728 11218
rect 1858 11183 1914 11192
rect 1676 11154 1728 11160
rect 1768 11008 1820 11014
rect 1768 10950 1820 10956
rect 1780 10266 1808 10950
rect 1860 10668 1912 10674
rect 1860 10610 1912 10616
rect 1768 10260 1820 10266
rect 1768 10202 1820 10208
rect 1596 10084 1808 10112
rect 1674 10024 1730 10033
rect 1674 9959 1676 9968
rect 1728 9959 1730 9968
rect 1676 9930 1728 9936
rect 1582 9752 1638 9761
rect 1582 9687 1638 9696
rect 1308 9648 1360 9654
rect 1308 9590 1360 9596
rect 1320 9081 1348 9590
rect 1400 9376 1452 9382
rect 1400 9318 1452 9324
rect 1306 9072 1362 9081
rect 1306 9007 1362 9016
rect 1306 8256 1362 8265
rect 1306 8191 1362 8200
rect 1320 7041 1348 8191
rect 1306 7032 1362 7041
rect 1306 6967 1362 6976
rect 1320 6798 1348 6967
rect 1308 6792 1360 6798
rect 1308 6734 1360 6740
rect 1412 6633 1440 9318
rect 1596 8974 1624 9687
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1504 8673 1532 8910
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1490 8664 1546 8673
rect 1490 8599 1546 8608
rect 1596 8537 1624 8774
rect 1582 8528 1638 8537
rect 1582 8463 1638 8472
rect 1688 8430 1716 9590
rect 1780 9330 1808 10084
rect 1872 9518 1900 10610
rect 1964 10470 1992 13359
rect 2056 12918 2084 13767
rect 2044 12912 2096 12918
rect 2044 12854 2096 12860
rect 2148 11880 2176 14334
rect 2240 13870 2268 14350
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2332 13784 2360 14962
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2424 14006 2452 14214
rect 2608 14074 2636 14962
rect 2700 14414 2728 15302
rect 2976 15162 3004 16050
rect 3056 16040 3108 16046
rect 3056 15982 3108 15988
rect 3146 16008 3202 16017
rect 2964 15156 3016 15162
rect 2964 15098 3016 15104
rect 3068 14618 3096 15982
rect 3146 15943 3202 15952
rect 3056 14612 3108 14618
rect 3056 14554 3108 14560
rect 2964 14544 3016 14550
rect 2964 14486 3016 14492
rect 2688 14408 2740 14414
rect 2740 14368 2820 14396
rect 2688 14350 2740 14356
rect 2686 14240 2742 14249
rect 2686 14175 2742 14184
rect 2596 14068 2648 14074
rect 2596 14010 2648 14016
rect 2412 14000 2464 14006
rect 2412 13942 2464 13948
rect 2700 13938 2728 14175
rect 2688 13932 2740 13938
rect 2688 13874 2740 13880
rect 2332 13756 2452 13784
rect 2320 13252 2372 13258
rect 2320 13194 2372 13200
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2056 11852 2176 11880
rect 1952 10464 2004 10470
rect 1952 10406 2004 10412
rect 2056 9625 2084 11852
rect 2136 11756 2188 11762
rect 2136 11698 2188 11704
rect 2148 11665 2176 11698
rect 2134 11656 2190 11665
rect 2134 11591 2190 11600
rect 2240 11218 2268 12582
rect 2228 11212 2280 11218
rect 2228 11154 2280 11160
rect 2240 10742 2268 11154
rect 2228 10736 2280 10742
rect 2228 10678 2280 10684
rect 2332 10554 2360 13194
rect 2424 12170 2452 13756
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2700 12646 2728 13670
rect 2792 13297 2820 14368
rect 2976 13569 3004 14486
rect 3160 14362 3188 15943
rect 3252 15706 3280 16594
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 14952 3292 14958
rect 3238 14920 3240 14929
rect 3292 14920 3294 14929
rect 3238 14855 3294 14864
rect 3068 14334 3188 14362
rect 2962 13560 3018 13569
rect 2962 13495 3018 13504
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2780 12912 2832 12918
rect 2780 12854 2832 12860
rect 2688 12640 2740 12646
rect 2688 12582 2740 12588
rect 2700 12442 2728 12582
rect 2688 12436 2740 12442
rect 2688 12378 2740 12384
rect 2686 12200 2742 12209
rect 2412 12164 2464 12170
rect 2412 12106 2464 12112
rect 2504 12164 2556 12170
rect 2686 12135 2742 12144
rect 2504 12106 2556 12112
rect 2410 11656 2466 11665
rect 2410 11591 2466 11600
rect 2424 11558 2452 11591
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2148 10526 2360 10554
rect 2042 9616 2098 9625
rect 2042 9551 2098 9560
rect 1860 9512 1912 9518
rect 1860 9454 1912 9460
rect 1950 9480 2006 9489
rect 1950 9415 1952 9424
rect 2004 9415 2006 9424
rect 1952 9386 2004 9392
rect 2148 9382 2176 10526
rect 2516 10470 2544 12106
rect 2594 12064 2650 12073
rect 2594 11999 2650 12008
rect 2504 10464 2556 10470
rect 2504 10406 2556 10412
rect 2516 10130 2544 10406
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2228 9920 2280 9926
rect 2228 9862 2280 9868
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2502 9888 2558 9897
rect 2136 9376 2188 9382
rect 1780 9302 2084 9330
rect 2136 9318 2188 9324
rect 1766 9072 1822 9081
rect 1766 9007 1822 9016
rect 1676 8424 1728 8430
rect 1676 8366 1728 8372
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1492 7472 1544 7478
rect 1490 7440 1492 7449
rect 1544 7440 1546 7449
rect 1490 7375 1546 7384
rect 1596 7206 1624 7822
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 1688 7313 1716 7754
rect 1674 7304 1730 7313
rect 1674 7239 1730 7248
rect 1584 7200 1636 7206
rect 1584 7142 1636 7148
rect 1596 6905 1624 7142
rect 1780 6914 1808 9007
rect 1858 8936 1914 8945
rect 1858 8871 1914 8880
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1688 6886 1808 6914
rect 1398 6624 1454 6633
rect 1398 6559 1454 6568
rect 1412 6458 1440 6559
rect 1400 6452 1452 6458
rect 1400 6394 1452 6400
rect 1306 5944 1362 5953
rect 1306 5879 1362 5888
rect 1216 3936 1268 3942
rect 1216 3878 1268 3884
rect 940 3528 992 3534
rect 940 3470 992 3476
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 848 1964 900 1970
rect 848 1906 900 1912
rect 1044 1086 1072 3402
rect 1320 2009 1348 5879
rect 1596 5778 1624 6831
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 1490 5536 1546 5545
rect 1490 5471 1546 5480
rect 1504 5302 1532 5471
rect 1492 5296 1544 5302
rect 1492 5238 1544 5244
rect 1306 2000 1362 2009
rect 1306 1935 1362 1944
rect 1032 1080 1084 1086
rect 1032 1022 1084 1028
rect 1044 800 1072 1022
rect 1412 870 1532 898
rect 1412 800 1440 870
rect 768 326 980 354
rect 952 241 980 326
rect 938 232 994 241
rect 938 167 994 176
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1504 762 1532 870
rect 1688 762 1716 6886
rect 1872 6662 1900 8871
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1964 8090 1992 8434
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1964 6866 1992 8026
rect 1952 6860 2004 6866
rect 1952 6802 2004 6808
rect 2056 6730 2084 9302
rect 2240 9178 2268 9862
rect 2332 9722 2360 9862
rect 2502 9823 2558 9832
rect 2320 9716 2372 9722
rect 2320 9658 2372 9664
rect 2320 9444 2372 9450
rect 2320 9386 2372 9392
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2228 9172 2280 9178
rect 2228 9114 2280 9120
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 7721 2268 8366
rect 2226 7712 2282 7721
rect 2226 7647 2282 7656
rect 2044 6724 2096 6730
rect 2044 6666 2096 6672
rect 1860 6656 1912 6662
rect 1860 6598 1912 6604
rect 2136 6656 2188 6662
rect 2136 6598 2188 6604
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1964 5778 1992 6054
rect 2148 5914 2176 6598
rect 2240 6458 2268 7647
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 6118 2360 9386
rect 2424 9178 2452 9386
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 2516 9110 2544 9823
rect 2504 9104 2556 9110
rect 2504 9046 2556 9052
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2424 8090 2452 8774
rect 2516 8634 2544 8774
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2502 8392 2558 8401
rect 2502 8327 2558 8336
rect 2412 8084 2464 8090
rect 2412 8026 2464 8032
rect 2410 7984 2466 7993
rect 2410 7919 2466 7928
rect 2424 6254 2452 7919
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2320 6112 2372 6118
rect 2320 6054 2372 6060
rect 2516 5930 2544 8327
rect 2608 7585 2636 11999
rect 2700 11121 2728 12135
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2700 10742 2728 11047
rect 2688 10736 2740 10742
rect 2688 10678 2740 10684
rect 2792 10441 2820 12854
rect 2962 12608 3018 12617
rect 2962 12543 3018 12552
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11354 2912 12174
rect 2976 11778 3004 12543
rect 3068 12481 3096 14334
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3160 13190 3188 14214
rect 3344 14056 3372 17292
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 3988 16833 4016 17478
rect 3974 16824 4030 16833
rect 3974 16759 4030 16768
rect 3976 16584 4028 16590
rect 3976 16526 4028 16532
rect 3988 15978 4016 16526
rect 4172 16289 4200 17478
rect 4264 16674 4292 17870
rect 4436 17740 4488 17746
rect 4436 17682 4488 17688
rect 4448 17270 4476 17682
rect 4436 17264 4488 17270
rect 4436 17206 4488 17212
rect 4436 16992 4488 16998
rect 4540 16969 4568 18770
rect 4632 18057 4660 20334
rect 4724 18358 4752 21490
rect 4816 21418 4844 22200
rect 4804 21412 4856 21418
rect 4804 21354 4856 21360
rect 5080 21412 5132 21418
rect 5080 21354 5132 21360
rect 4988 20392 5040 20398
rect 4988 20334 5040 20340
rect 4896 20256 4948 20262
rect 4802 20224 4858 20233
rect 4896 20198 4948 20204
rect 4802 20159 4858 20168
rect 4816 18714 4844 20159
rect 4908 19802 4936 20198
rect 5000 20097 5028 20334
rect 4986 20088 5042 20097
rect 4986 20023 5042 20032
rect 4908 19774 5028 19802
rect 4896 19712 4948 19718
rect 4896 19654 4948 19660
rect 4908 19446 4936 19654
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 4908 18834 4936 19382
rect 4896 18828 4948 18834
rect 4896 18770 4948 18776
rect 4816 18686 4936 18714
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4712 18352 4764 18358
rect 4710 18320 4712 18329
rect 4764 18320 4766 18329
rect 4710 18255 4766 18264
rect 4816 18222 4844 18566
rect 4908 18222 4936 18686
rect 4804 18216 4856 18222
rect 4804 18158 4856 18164
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 4712 18148 4764 18154
rect 4712 18090 4764 18096
rect 4618 18048 4674 18057
rect 4618 17983 4674 17992
rect 4620 17672 4672 17678
rect 4620 17614 4672 17620
rect 4632 17105 4660 17614
rect 4618 17096 4674 17105
rect 4618 17031 4674 17040
rect 4436 16934 4488 16940
rect 4526 16960 4582 16969
rect 4264 16646 4384 16674
rect 4448 16658 4476 16934
rect 4526 16895 4582 16904
rect 4250 16552 4306 16561
rect 4250 16487 4306 16496
rect 4264 16454 4292 16487
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4158 16280 4214 16289
rect 4158 16215 4214 16224
rect 4356 16114 4384 16646
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 4540 16454 4568 16895
rect 4724 16590 4752 18090
rect 4712 16584 4764 16590
rect 4712 16526 4764 16532
rect 4528 16448 4580 16454
rect 4528 16390 4580 16396
rect 4344 16108 4396 16114
rect 4344 16050 4396 16056
rect 4068 16040 4120 16046
rect 4068 15982 4120 15988
rect 3976 15972 4028 15978
rect 3976 15914 4028 15920
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 4080 15162 4108 15982
rect 4356 15910 4384 16050
rect 4344 15904 4396 15910
rect 4344 15846 4396 15852
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 4264 15094 4292 15438
rect 4252 15088 4304 15094
rect 4252 15030 4304 15036
rect 4160 14884 4212 14890
rect 4160 14826 4212 14832
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 4172 14482 4200 14826
rect 4540 14618 4568 16390
rect 4816 15978 4844 18158
rect 4896 18080 4948 18086
rect 4896 18022 4948 18028
rect 4908 16250 4936 18022
rect 4896 16244 4948 16250
rect 4896 16186 4948 16192
rect 4896 16040 4948 16046
rect 4896 15982 4948 15988
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4816 15638 4844 15914
rect 4804 15632 4856 15638
rect 4804 15574 4856 15580
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4632 14958 4660 15438
rect 4712 15360 4764 15366
rect 4712 15302 4764 15308
rect 4620 14952 4672 14958
rect 4620 14894 4672 14900
rect 4528 14612 4580 14618
rect 4528 14554 4580 14560
rect 4160 14476 4212 14482
rect 4160 14418 4212 14424
rect 3884 14408 3936 14414
rect 3884 14350 3936 14356
rect 3516 14272 3568 14278
rect 3516 14214 3568 14220
rect 3252 14028 3372 14056
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3252 13002 3280 14028
rect 3528 13977 3556 14214
rect 3514 13968 3570 13977
rect 3332 13932 3384 13938
rect 3514 13903 3570 13912
rect 3332 13874 3384 13880
rect 3344 13530 3372 13874
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 3896 13530 3924 14350
rect 4068 14272 4120 14278
rect 4066 14240 4068 14249
rect 4436 14272 4488 14278
rect 4120 14240 4122 14249
rect 4436 14214 4488 14220
rect 4528 14272 4580 14278
rect 4528 14214 4580 14220
rect 4066 14175 4122 14184
rect 4068 13864 4120 13870
rect 3988 13824 4068 13852
rect 3332 13524 3384 13530
rect 3332 13466 3384 13472
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3332 13252 3384 13258
rect 3436 13240 3464 13466
rect 3882 13424 3938 13433
rect 3882 13359 3938 13368
rect 3384 13212 3464 13240
rect 3332 13194 3384 13200
rect 3160 12974 3280 13002
rect 3054 12472 3110 12481
rect 3054 12407 3110 12416
rect 3056 12368 3108 12374
rect 3056 12310 3108 12316
rect 3068 11898 3096 12310
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2976 11750 3096 11778
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2964 11008 3016 11014
rect 2964 10950 3016 10956
rect 2778 10432 2834 10441
rect 2778 10367 2834 10376
rect 2792 10062 2820 10367
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2976 9926 3004 10950
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2780 9920 2832 9926
rect 2780 9862 2832 9868
rect 2964 9920 3016 9926
rect 2964 9862 3016 9868
rect 2700 9722 2728 9862
rect 2688 9716 2740 9722
rect 2688 9658 2740 9664
rect 2688 9512 2740 9518
rect 2688 9454 2740 9460
rect 2700 9042 2728 9454
rect 2792 9058 2820 9862
rect 2964 9716 3016 9722
rect 2964 9658 3016 9664
rect 2872 9580 2924 9586
rect 2872 9522 2924 9528
rect 2884 9178 2912 9522
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2688 9036 2740 9042
rect 2792 9030 2912 9058
rect 2688 8978 2740 8984
rect 2780 8968 2832 8974
rect 2780 8910 2832 8916
rect 2686 7848 2742 7857
rect 2686 7783 2742 7792
rect 2594 7576 2650 7585
rect 2594 7511 2650 7520
rect 2596 6860 2648 6866
rect 2596 6802 2648 6808
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 2424 5902 2544 5930
rect 1952 5772 2004 5778
rect 1952 5714 2004 5720
rect 1768 5568 1820 5574
rect 1768 5510 1820 5516
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 1780 4826 1808 5510
rect 2136 5228 2188 5234
rect 2056 5188 2136 5216
rect 1768 4820 1820 4826
rect 1768 4762 1820 4768
rect 2056 4486 2084 5188
rect 2136 5170 2188 5176
rect 2136 5024 2188 5030
rect 2136 4966 2188 4972
rect 2148 4622 2176 4966
rect 2226 4856 2282 4865
rect 2226 4791 2282 4800
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 2044 4480 2096 4486
rect 2044 4422 2096 4428
rect 1950 4176 2006 4185
rect 2240 4146 2268 4791
rect 1950 4111 1952 4120
rect 2004 4111 2006 4120
rect 2228 4140 2280 4146
rect 1952 4082 2004 4088
rect 2228 4082 2280 4088
rect 2332 4010 2360 5510
rect 1768 4004 1820 4010
rect 1768 3946 1820 3952
rect 2320 4004 2372 4010
rect 2320 3946 2372 3952
rect 1780 2446 1808 3946
rect 1858 3632 1914 3641
rect 1858 3567 1914 3576
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 1872 800 1900 3567
rect 2424 3058 2452 5902
rect 2504 5636 2556 5642
rect 2504 5578 2556 5584
rect 2516 4078 2544 5578
rect 2608 5234 2636 6802
rect 2596 5228 2648 5234
rect 2596 5170 2648 5176
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2608 4146 2636 4966
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2700 3602 2728 7783
rect 2792 6662 2820 8910
rect 2884 8906 2912 9030
rect 2872 8900 2924 8906
rect 2872 8842 2924 8848
rect 2870 8800 2926 8809
rect 2870 8735 2926 8744
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2780 6112 2832 6118
rect 2780 6054 2832 6060
rect 2792 3670 2820 6054
rect 2884 5137 2912 8735
rect 2976 7546 3004 9658
rect 3068 8265 3096 11750
rect 3160 10810 3188 12974
rect 3240 12844 3292 12850
rect 3240 12786 3292 12792
rect 3252 12442 3280 12786
rect 3344 12714 3372 13194
rect 3516 13184 3568 13190
rect 3516 13126 3568 13132
rect 3528 12918 3556 13126
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3896 12782 3924 13359
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3988 12646 4016 13824
rect 4068 13806 4120 13812
rect 4344 13728 4396 13734
rect 4344 13670 4396 13676
rect 4356 13433 4384 13670
rect 4342 13424 4398 13433
rect 4068 13388 4120 13394
rect 4342 13359 4344 13368
rect 4068 13330 4120 13336
rect 4396 13359 4398 13368
rect 4344 13330 4396 13336
rect 4080 13138 4108 13330
rect 4356 13299 4384 13330
rect 4252 13184 4304 13190
rect 4080 13110 4200 13138
rect 4252 13126 4304 13132
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3976 12640 4028 12646
rect 3976 12582 4028 12588
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3988 12306 4016 12582
rect 4080 12442 4108 12786
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 3976 12300 4028 12306
rect 3976 12242 4028 12248
rect 3884 12232 3936 12238
rect 3884 12174 3936 12180
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3344 10470 3372 11630
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3792 11144 3844 11150
rect 3790 11112 3792 11121
rect 3844 11112 3846 11121
rect 3424 11076 3476 11082
rect 3790 11047 3846 11056
rect 3424 11018 3476 11024
rect 3332 10464 3384 10470
rect 3332 10406 3384 10412
rect 3436 10130 3464 11018
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3790 10160 3846 10169
rect 3424 10124 3476 10130
rect 3476 10084 3740 10112
rect 3790 10095 3846 10104
rect 3424 10066 3476 10072
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 2964 7540 3016 7546
rect 2964 7482 3016 7488
rect 2964 7404 3016 7410
rect 2964 7346 3016 7352
rect 2976 6254 3004 7346
rect 3160 6914 3188 9998
rect 3608 9988 3660 9994
rect 3528 9948 3608 9976
rect 3332 9920 3384 9926
rect 3332 9862 3384 9868
rect 3240 9376 3292 9382
rect 3344 9353 3372 9862
rect 3528 9432 3556 9948
rect 3608 9930 3660 9936
rect 3712 9654 3740 10084
rect 3804 10062 3832 10095
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9722 3832 9998
rect 3792 9716 3844 9722
rect 3792 9658 3844 9664
rect 3700 9648 3752 9654
rect 3700 9590 3752 9596
rect 3712 9450 3740 9590
rect 3436 9404 3556 9432
rect 3700 9444 3752 9450
rect 3240 9318 3292 9324
rect 3330 9344 3386 9353
rect 3252 8838 3280 9318
rect 3330 9279 3386 9288
rect 3436 9042 3464 9404
rect 3700 9386 3752 9392
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3896 9178 3924 12174
rect 4172 11898 4200 13110
rect 4264 12238 4292 13126
rect 4448 12986 4476 14214
rect 4540 13530 4568 14214
rect 4620 14000 4672 14006
rect 4724 13988 4752 15302
rect 4804 14884 4856 14890
rect 4804 14826 4856 14832
rect 4816 14618 4844 14826
rect 4804 14612 4856 14618
rect 4804 14554 4856 14560
rect 4672 13960 4752 13988
rect 4620 13942 4672 13948
rect 4724 13734 4752 13960
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4528 13524 4580 13530
rect 4528 13466 4580 13472
rect 4526 13424 4582 13433
rect 4526 13359 4582 13368
rect 4436 12980 4488 12986
rect 4436 12922 4488 12928
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 11892 4212 11898
rect 4160 11834 4212 11840
rect 3988 11750 4200 11778
rect 3988 11354 4016 11750
rect 4172 11694 4200 11750
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4068 11688 4120 11694
rect 4068 11630 4120 11636
rect 4160 11688 4212 11694
rect 4160 11630 4212 11636
rect 4080 11354 4108 11630
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3988 10742 4016 11290
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 4080 10810 4108 11154
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3974 10432 4030 10441
rect 3974 10367 4030 10376
rect 3988 10266 4016 10367
rect 3976 10260 4028 10266
rect 3976 10202 4028 10208
rect 3974 10024 4030 10033
rect 3974 9959 4030 9968
rect 3884 9172 3936 9178
rect 3884 9114 3936 9120
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3068 6886 3188 6914
rect 3068 6390 3096 6886
rect 3252 6798 3280 7958
rect 3332 7336 3384 7342
rect 3332 7278 3384 7284
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3056 6384 3108 6390
rect 3056 6326 3108 6332
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 2870 5128 2926 5137
rect 2870 5063 2926 5072
rect 2976 4690 3004 6190
rect 3240 6112 3292 6118
rect 3240 6054 3292 6060
rect 3054 5672 3110 5681
rect 3054 5607 3110 5616
rect 3068 5370 3096 5607
rect 3252 5370 3280 6054
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2964 4548 3016 4554
rect 2964 4490 3016 4496
rect 2976 3738 3004 4490
rect 3068 4457 3096 5170
rect 3240 5160 3292 5166
rect 3240 5102 3292 5108
rect 3054 4448 3110 4457
rect 3054 4383 3110 4392
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2780 3664 2832 3670
rect 2780 3606 2832 3612
rect 2688 3596 2740 3602
rect 2688 3538 2740 3544
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 2594 3224 2650 3233
rect 2594 3159 2650 3168
rect 2608 3126 2636 3159
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1952 2984 2004 2990
rect 1952 2926 2004 2932
rect 2778 2952 2834 2961
rect 1964 1902 1992 2926
rect 2778 2887 2834 2896
rect 2686 2816 2742 2825
rect 2686 2751 2742 2760
rect 2700 2514 2728 2751
rect 2792 2514 2820 2887
rect 2228 2508 2280 2514
rect 2228 2450 2280 2456
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2780 2508 2832 2514
rect 2780 2450 2832 2456
rect 1952 1896 2004 1902
rect 1952 1838 2004 1844
rect 2240 800 2268 2450
rect 2412 2440 2464 2446
rect 2792 2394 2820 2450
rect 2412 2382 2464 2388
rect 2424 2038 2452 2382
rect 2700 2366 2820 2394
rect 2412 2032 2464 2038
rect 2412 1974 2464 1980
rect 2700 800 2728 2366
rect 2884 1834 2912 3470
rect 2976 2922 3004 3674
rect 3068 3126 3096 3946
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2872 1828 2924 1834
rect 2872 1770 2924 1776
rect 3252 1358 3280 5102
rect 3344 4622 3372 7278
rect 3436 6458 3464 8978
rect 3528 8809 3556 8978
rect 3514 8800 3570 8809
rect 3514 8735 3570 8744
rect 3988 8673 4016 9959
rect 4080 9926 4108 10746
rect 4068 9920 4120 9926
rect 4172 9897 4200 11018
rect 4264 10538 4292 11698
rect 4356 10674 4384 12786
rect 4434 12744 4490 12753
rect 4434 12679 4490 12688
rect 4344 10668 4396 10674
rect 4344 10610 4396 10616
rect 4252 10532 4304 10538
rect 4252 10474 4304 10480
rect 4356 10441 4384 10610
rect 4342 10432 4398 10441
rect 4342 10367 4398 10376
rect 4250 10296 4306 10305
rect 4250 10231 4306 10240
rect 4264 10062 4292 10231
rect 4252 10056 4304 10062
rect 4252 9998 4304 10004
rect 4068 9862 4120 9868
rect 4158 9888 4214 9897
rect 4158 9823 4214 9832
rect 4264 9738 4292 9998
rect 4080 9710 4292 9738
rect 4344 9716 4396 9722
rect 4080 9178 4108 9710
rect 4344 9658 4396 9664
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 4264 9489 4292 9522
rect 4250 9480 4306 9489
rect 4250 9415 4306 9424
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4158 9208 4214 9217
rect 4068 9172 4120 9178
rect 4158 9143 4214 9152
rect 4068 9114 4120 9120
rect 4066 9072 4122 9081
rect 4066 9007 4122 9016
rect 4080 8974 4108 9007
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3974 8664 4030 8673
rect 3974 8599 4030 8608
rect 3882 8528 3938 8537
rect 3882 8463 3938 8472
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 3896 8072 3924 8463
rect 3976 8288 4028 8294
rect 4080 8265 4108 8774
rect 3976 8230 4028 8236
rect 4066 8256 4122 8265
rect 3804 8044 3924 8072
rect 3514 7984 3570 7993
rect 3514 7919 3570 7928
rect 3528 7886 3556 7919
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3606 7440 3662 7449
rect 3712 7410 3740 7754
rect 3804 7721 3832 8044
rect 3882 7984 3938 7993
rect 3988 7954 4016 8230
rect 4066 8191 4122 8200
rect 4066 8120 4122 8129
rect 4066 8055 4122 8064
rect 3882 7919 3938 7928
rect 3976 7948 4028 7954
rect 3790 7712 3846 7721
rect 3790 7647 3846 7656
rect 3606 7375 3662 7384
rect 3700 7404 3752 7410
rect 3620 7342 3648 7375
rect 3700 7346 3752 7352
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3514 6896 3570 6905
rect 3514 6831 3516 6840
rect 3568 6831 3570 6840
rect 3698 6896 3754 6905
rect 3698 6831 3754 6840
rect 3516 6802 3568 6808
rect 3424 6452 3476 6458
rect 3424 6394 3476 6400
rect 3712 6322 3740 6831
rect 3896 6610 3924 7919
rect 3976 7890 4028 7896
rect 4080 7750 4108 8055
rect 4172 7886 4200 9143
rect 4264 7954 4292 9318
rect 4356 9217 4384 9658
rect 4448 9586 4476 12679
rect 4540 12170 4568 13359
rect 4724 13326 4752 13670
rect 4712 13320 4764 13326
rect 4712 13262 4764 13268
rect 4816 13172 4844 14554
rect 4908 14346 4936 15982
rect 4896 14340 4948 14346
rect 4896 14282 4948 14288
rect 5000 13530 5028 19774
rect 5092 18358 5120 21354
rect 5184 20602 5212 22200
rect 5172 20596 5224 20602
rect 5552 20584 5580 22200
rect 5552 20556 5764 20584
rect 5172 20538 5224 20544
rect 5080 18352 5132 18358
rect 5184 18329 5212 20538
rect 5632 20460 5684 20466
rect 5632 20402 5684 20408
rect 5540 20392 5592 20398
rect 5540 20334 5592 20340
rect 5356 20256 5408 20262
rect 5356 20198 5408 20204
rect 5368 19258 5396 20198
rect 5552 19922 5580 20334
rect 5540 19916 5592 19922
rect 5540 19858 5592 19864
rect 5448 19848 5500 19854
rect 5448 19790 5500 19796
rect 5460 19378 5488 19790
rect 5540 19780 5592 19786
rect 5540 19722 5592 19728
rect 5448 19372 5500 19378
rect 5448 19314 5500 19320
rect 5276 19230 5396 19258
rect 5080 18294 5132 18300
rect 5170 18320 5226 18329
rect 5170 18255 5226 18264
rect 5276 18222 5304 19230
rect 5356 18896 5408 18902
rect 5356 18838 5408 18844
rect 5172 18216 5224 18222
rect 5172 18158 5224 18164
rect 5264 18216 5316 18222
rect 5264 18158 5316 18164
rect 5078 17776 5134 17785
rect 5078 17711 5134 17720
rect 5092 17678 5120 17711
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 5080 17536 5132 17542
rect 5080 17478 5132 17484
rect 5092 17270 5120 17478
rect 5080 17264 5132 17270
rect 5080 17206 5132 17212
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5092 15366 5120 16390
rect 5080 15360 5132 15366
rect 5080 15302 5132 15308
rect 5184 15314 5212 18158
rect 5262 18048 5318 18057
rect 5262 17983 5318 17992
rect 5276 16402 5304 17983
rect 5368 17882 5396 18838
rect 5448 18692 5500 18698
rect 5448 18634 5500 18640
rect 5460 18601 5488 18634
rect 5446 18592 5502 18601
rect 5446 18527 5502 18536
rect 5448 18284 5500 18290
rect 5448 18226 5500 18232
rect 5460 18086 5488 18226
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5356 17876 5408 17882
rect 5356 17818 5408 17824
rect 5356 17740 5408 17746
rect 5356 17682 5408 17688
rect 5368 16794 5396 17682
rect 5460 17678 5488 18022
rect 5448 17672 5500 17678
rect 5448 17614 5500 17620
rect 5552 17134 5580 19722
rect 5644 19514 5672 20402
rect 5632 19508 5684 19514
rect 5632 19450 5684 19456
rect 5736 19394 5764 20556
rect 5920 20482 5948 22200
rect 6012 20534 6040 22222
rect 6196 22114 6224 22222
rect 6274 22200 6330 23000
rect 6642 22200 6698 23000
rect 7102 22200 7158 23000
rect 7470 22200 7526 23000
rect 7746 22808 7802 22817
rect 7746 22743 7802 22752
rect 6288 22114 6316 22200
rect 6196 22086 6316 22114
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 6550 20632 6606 20641
rect 6288 20576 6550 20584
rect 6288 20567 6606 20576
rect 6288 20556 6592 20567
rect 5828 20454 5948 20482
rect 6000 20528 6052 20534
rect 6000 20470 6052 20476
rect 5828 20330 5856 20454
rect 5816 20324 5868 20330
rect 5816 20266 5868 20272
rect 5644 19366 5764 19394
rect 5644 18601 5672 19366
rect 5828 19145 5856 20266
rect 6012 19496 6040 20470
rect 6288 20233 6316 20556
rect 6550 20496 6606 20505
rect 6550 20431 6606 20440
rect 6460 20256 6512 20262
rect 6274 20224 6330 20233
rect 6274 20159 6330 20168
rect 6458 20224 6460 20233
rect 6512 20224 6514 20233
rect 6458 20159 6514 20168
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 6012 19468 6224 19496
rect 5908 19440 5960 19446
rect 5960 19388 6040 19394
rect 5908 19382 6040 19388
rect 5920 19366 6040 19382
rect 5908 19304 5960 19310
rect 5908 19246 5960 19252
rect 5814 19136 5870 19145
rect 5814 19071 5870 19080
rect 5724 18692 5776 18698
rect 5724 18634 5776 18640
rect 5630 18592 5686 18601
rect 5630 18527 5686 18536
rect 5630 18456 5686 18465
rect 5630 18391 5686 18400
rect 5644 18057 5672 18391
rect 5736 18306 5764 18634
rect 5816 18624 5868 18630
rect 5816 18566 5868 18572
rect 5828 18426 5856 18566
rect 5920 18426 5948 19246
rect 5816 18420 5868 18426
rect 5816 18362 5868 18368
rect 5908 18420 5960 18426
rect 5908 18362 5960 18368
rect 5736 18278 5856 18306
rect 5724 18216 5776 18222
rect 5724 18158 5776 18164
rect 5630 18048 5686 18057
rect 5630 17983 5686 17992
rect 5632 17672 5684 17678
rect 5736 17649 5764 18158
rect 5632 17614 5684 17620
rect 5722 17640 5778 17649
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5644 16969 5672 17614
rect 5722 17575 5778 17584
rect 5724 17536 5776 17542
rect 5722 17504 5724 17513
rect 5776 17504 5778 17513
rect 5722 17439 5778 17448
rect 5736 17338 5764 17439
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5724 17196 5776 17202
rect 5724 17138 5776 17144
rect 5630 16960 5686 16969
rect 5630 16895 5686 16904
rect 5356 16788 5408 16794
rect 5356 16730 5408 16736
rect 5632 16720 5684 16726
rect 5632 16662 5684 16668
rect 5538 16552 5594 16561
rect 5460 16522 5538 16538
rect 5448 16516 5538 16522
rect 5500 16510 5538 16516
rect 5538 16487 5594 16496
rect 5448 16458 5500 16464
rect 5540 16448 5592 16454
rect 5276 16374 5488 16402
rect 5540 16390 5592 16396
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5276 16114 5304 16186
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5356 16040 5408 16046
rect 5356 15982 5408 15988
rect 5184 15286 5304 15314
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 5078 14920 5134 14929
rect 5078 14855 5134 14864
rect 5092 14113 5120 14855
rect 5184 14414 5212 15098
rect 5276 14618 5304 15286
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5172 14408 5224 14414
rect 5172 14350 5224 14356
rect 5264 14408 5316 14414
rect 5264 14350 5316 14356
rect 5078 14104 5134 14113
rect 5078 14039 5134 14048
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4724 13144 4844 13172
rect 4988 13184 5040 13190
rect 4620 12368 4672 12374
rect 4620 12310 4672 12316
rect 4528 12164 4580 12170
rect 4528 12106 4580 12112
rect 4632 12102 4660 12310
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 10538 4568 11494
rect 4528 10532 4580 10538
rect 4528 10474 4580 10480
rect 4528 9920 4580 9926
rect 4528 9862 4580 9868
rect 4436 9580 4488 9586
rect 4436 9522 4488 9528
rect 4436 9444 4488 9450
rect 4436 9386 4488 9392
rect 4342 9208 4398 9217
rect 4342 9143 4398 9152
rect 4344 9104 4396 9110
rect 4448 9092 4476 9386
rect 4396 9064 4476 9092
rect 4344 9046 4396 9052
rect 4344 8968 4396 8974
rect 4344 8910 4396 8916
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4356 8838 4384 8910
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8498 4384 8774
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 7744 4120 7750
rect 4068 7686 4120 7692
rect 4344 7744 4396 7750
rect 4344 7686 4396 7692
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6798 4016 7142
rect 4080 7002 4108 7346
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 4264 6798 4292 7346
rect 4356 7206 4384 7686
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3804 6582 3924 6610
rect 3804 6497 3832 6582
rect 3790 6488 3846 6497
rect 3790 6423 3846 6432
rect 3884 6452 3936 6458
rect 3884 6394 3936 6400
rect 3700 6316 3752 6322
rect 3700 6258 3752 6264
rect 3424 6180 3476 6186
rect 3424 6122 3476 6128
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3436 4146 3464 6122
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3608 5840 3660 5846
rect 3606 5808 3608 5817
rect 3660 5808 3662 5817
rect 3606 5743 3662 5752
rect 3790 5808 3846 5817
rect 3790 5743 3846 5752
rect 3804 5710 3832 5743
rect 3608 5704 3660 5710
rect 3608 5646 3660 5652
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3620 5302 3648 5646
rect 3608 5296 3660 5302
rect 3804 5273 3832 5646
rect 3608 5238 3660 5244
rect 3790 5264 3846 5273
rect 3896 5234 3924 6394
rect 3988 5642 4016 6734
rect 4080 6254 4108 6734
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4068 6248 4120 6254
rect 4068 6190 4120 6196
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 3976 5364 4028 5370
rect 3976 5306 4028 5312
rect 3790 5199 3846 5208
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3882 4584 3938 4593
rect 3882 4519 3938 4528
rect 3792 4480 3844 4486
rect 3792 4422 3844 4428
rect 3804 4214 3832 4422
rect 3896 4214 3924 4519
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3884 4208 3936 4214
rect 3884 4150 3936 4156
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3422 4040 3478 4049
rect 3422 3975 3478 3984
rect 3882 4040 3938 4049
rect 3882 3975 3884 3984
rect 3240 1352 3292 1358
rect 3240 1294 3292 1300
rect 3240 1216 3292 1222
rect 3240 1158 3292 1164
rect 3252 921 3280 1158
rect 3238 912 3294 921
rect 3068 870 3188 898
rect 3068 800 3096 870
rect 1504 734 1716 762
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3160 762 3188 870
rect 3238 847 3294 856
rect 3436 762 3464 3975
rect 3936 3975 3938 3984
rect 3884 3946 3936 3952
rect 3988 3890 4016 5306
rect 4080 4865 4108 5782
rect 4172 5302 4200 6598
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 4264 5914 4292 6190
rect 4252 5908 4304 5914
rect 4252 5850 4304 5856
rect 4356 5794 4384 7142
rect 4264 5766 4384 5794
rect 4160 5296 4212 5302
rect 4160 5238 4212 5244
rect 4158 5128 4214 5137
rect 4158 5063 4214 5072
rect 4066 4856 4122 4865
rect 4066 4791 4122 4800
rect 3896 3862 4016 3890
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 3896 2446 3924 3862
rect 4172 3754 4200 5063
rect 4264 4554 4292 5766
rect 4344 5704 4396 5710
rect 4344 5646 4396 5652
rect 4356 5166 4384 5646
rect 4344 5160 4396 5166
rect 4448 5137 4476 8910
rect 4540 6905 4568 9862
rect 4526 6896 4582 6905
rect 4526 6831 4582 6840
rect 4528 6792 4580 6798
rect 4528 6734 4580 6740
rect 4540 6390 4568 6734
rect 4528 6384 4580 6390
rect 4528 6326 4580 6332
rect 4528 5160 4580 5166
rect 4344 5102 4396 5108
rect 4434 5128 4490 5137
rect 4356 4690 4384 5102
rect 4528 5102 4580 5108
rect 4434 5063 4490 5072
rect 4436 5024 4488 5030
rect 4436 4966 4488 4972
rect 4344 4684 4396 4690
rect 4344 4626 4396 4632
rect 4342 4584 4398 4593
rect 4252 4548 4304 4554
rect 4342 4519 4344 4528
rect 4252 4490 4304 4496
rect 4396 4519 4398 4528
rect 4344 4490 4396 4496
rect 4342 4312 4398 4321
rect 4342 4247 4398 4256
rect 4252 4208 4304 4214
rect 4252 4150 4304 4156
rect 4080 3726 4200 3754
rect 3976 3392 4028 3398
rect 3976 3334 4028 3340
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3516 1284 3568 1290
rect 3516 1226 3568 1232
rect 3528 800 3556 1226
rect 3896 800 3924 2246
rect 3988 1766 4016 3334
rect 4080 2938 4108 3726
rect 4264 3641 4292 4150
rect 4250 3632 4306 3641
rect 4160 3596 4212 3602
rect 4250 3567 4306 3576
rect 4160 3538 4212 3544
rect 4172 3058 4200 3538
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 4080 2910 4200 2938
rect 4068 2848 4120 2854
rect 4172 2825 4200 2910
rect 4068 2790 4120 2796
rect 4158 2816 4214 2825
rect 4080 2310 4108 2790
rect 4158 2751 4214 2760
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4264 1873 4292 3402
rect 4250 1864 4306 1873
rect 4250 1799 4306 1808
rect 3976 1760 4028 1766
rect 3976 1702 4028 1708
rect 4356 800 4384 4247
rect 4448 3058 4476 4966
rect 4540 4622 4568 5102
rect 4632 4826 4660 11698
rect 4724 11558 4752 13144
rect 4988 13126 5040 13132
rect 4896 12980 4948 12986
rect 4896 12922 4948 12928
rect 4908 12288 4936 12922
rect 5000 12714 5028 13126
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 4988 12708 5040 12714
rect 4988 12650 5040 12656
rect 5092 12442 5120 12786
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 4816 12260 5028 12288
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4724 11218 4752 11494
rect 4712 11212 4764 11218
rect 4712 11154 4764 11160
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 4724 10198 4752 10542
rect 4712 10192 4764 10198
rect 4712 10134 4764 10140
rect 4712 9920 4764 9926
rect 4712 9862 4764 9868
rect 4724 9722 4752 9862
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4712 9512 4764 9518
rect 4712 9454 4764 9460
rect 4724 9353 4752 9454
rect 4710 9344 4766 9353
rect 4710 9279 4766 9288
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4724 7857 4752 9114
rect 4710 7848 4766 7857
rect 4710 7783 4766 7792
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 4528 4616 4580 4622
rect 4528 4558 4580 4564
rect 4618 4448 4674 4457
rect 4618 4383 4674 4392
rect 4632 4078 4660 4383
rect 4620 4072 4672 4078
rect 4620 4014 4672 4020
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4526 3768 4582 3777
rect 4526 3703 4582 3712
rect 4540 3534 4568 3703
rect 4632 3602 4660 3878
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4724 3534 4752 6598
rect 4816 4146 4844 12260
rect 4894 12200 4950 12209
rect 5000 12170 5028 12260
rect 4894 12135 4950 12144
rect 4988 12164 5040 12170
rect 4908 12102 4936 12135
rect 4988 12106 5040 12112
rect 4896 12096 4948 12102
rect 4896 12038 4948 12044
rect 4988 11688 5040 11694
rect 4988 11630 5040 11636
rect 4896 11212 4948 11218
rect 4896 11154 4948 11160
rect 4908 10606 4936 11154
rect 5000 11150 5028 11630
rect 5080 11552 5132 11558
rect 5078 11520 5080 11529
rect 5132 11520 5134 11529
rect 5078 11455 5134 11464
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5000 10849 5028 11086
rect 5092 11082 5120 11455
rect 5184 11257 5212 14350
rect 5276 14278 5304 14350
rect 5264 14272 5316 14278
rect 5264 14214 5316 14220
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5276 11898 5304 14010
rect 5368 12866 5396 15982
rect 5460 13569 5488 16374
rect 5552 16046 5580 16390
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5552 15706 5580 15982
rect 5644 15706 5672 16662
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 5630 15464 5686 15473
rect 5630 15399 5686 15408
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 14793 5580 15302
rect 5538 14784 5594 14793
rect 5538 14719 5594 14728
rect 5540 14272 5592 14278
rect 5540 14214 5592 14220
rect 5552 13841 5580 14214
rect 5538 13832 5594 13841
rect 5538 13767 5594 13776
rect 5446 13560 5502 13569
rect 5446 13495 5502 13504
rect 5448 13184 5500 13190
rect 5448 13126 5500 13132
rect 5460 12986 5488 13126
rect 5448 12980 5500 12986
rect 5448 12922 5500 12928
rect 5368 12838 5488 12866
rect 5354 12608 5410 12617
rect 5354 12543 5410 12552
rect 5368 12442 5396 12543
rect 5356 12436 5408 12442
rect 5356 12378 5408 12384
rect 5356 12096 5408 12102
rect 5356 12038 5408 12044
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5368 11801 5396 12038
rect 5354 11792 5410 11801
rect 5264 11756 5316 11762
rect 5354 11727 5410 11736
rect 5264 11698 5316 11704
rect 5170 11248 5226 11257
rect 5276 11218 5304 11698
rect 5170 11183 5226 11192
rect 5264 11212 5316 11218
rect 5264 11154 5316 11160
rect 5368 11098 5396 11727
rect 5080 11076 5132 11082
rect 5080 11018 5132 11024
rect 5184 11070 5396 11098
rect 4986 10840 5042 10849
rect 5184 10826 5212 11070
rect 5264 11008 5316 11014
rect 5316 10968 5396 10996
rect 5264 10950 5316 10956
rect 5184 10798 5304 10826
rect 4986 10775 5042 10784
rect 4988 10736 5040 10742
rect 4988 10678 5040 10684
rect 4896 10600 4948 10606
rect 4896 10542 4948 10548
rect 4908 10470 4936 10542
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4908 10130 4936 10406
rect 5000 10266 5028 10678
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5184 10266 5212 10542
rect 5276 10470 5304 10798
rect 5264 10464 5316 10470
rect 5264 10406 5316 10412
rect 5262 10296 5318 10305
rect 4988 10260 5040 10266
rect 4988 10202 5040 10208
rect 5172 10260 5224 10266
rect 5262 10231 5264 10240
rect 5172 10202 5224 10208
rect 5316 10231 5318 10240
rect 5264 10202 5316 10208
rect 4896 10124 4948 10130
rect 5368 10112 5396 10968
rect 5460 10198 5488 12838
rect 5540 12640 5592 12646
rect 5540 12582 5592 12588
rect 5552 11694 5580 12582
rect 5540 11688 5592 11694
rect 5540 11630 5592 11636
rect 5644 11506 5672 15399
rect 5736 15065 5764 17138
rect 5828 15586 5856 18278
rect 6012 18154 6040 19366
rect 6092 19304 6144 19310
rect 6092 19246 6144 19252
rect 6104 18970 6132 19246
rect 6092 18964 6144 18970
rect 6092 18906 6144 18912
rect 6196 18698 6224 19468
rect 6460 19372 6512 19378
rect 6460 19314 6512 19320
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6184 18692 6236 18698
rect 6184 18634 6236 18640
rect 6380 18612 6408 19178
rect 6472 18766 6500 19314
rect 6564 19174 6592 20431
rect 6656 19378 6684 22200
rect 6920 20596 6972 20602
rect 6920 20538 6972 20544
rect 6932 20482 6960 20538
rect 6840 20466 6960 20482
rect 6828 20460 6960 20466
rect 6880 20454 6960 20460
rect 6828 20402 6880 20408
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 6736 20324 6788 20330
rect 6736 20266 6788 20272
rect 6748 19854 6776 20266
rect 6828 20256 6880 20262
rect 6828 20198 6880 20204
rect 6840 19922 6868 20198
rect 6828 19916 6880 19922
rect 6828 19858 6880 19864
rect 6736 19848 6788 19854
rect 6736 19790 6788 19796
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6748 19310 6776 19790
rect 6828 19780 6880 19786
rect 6828 19722 6880 19728
rect 6736 19304 6788 19310
rect 6736 19246 6788 19252
rect 6840 19174 6868 19722
rect 6932 19718 6960 20334
rect 7012 20256 7064 20262
rect 7012 20198 7064 20204
rect 6920 19712 6972 19718
rect 6920 19654 6972 19660
rect 7024 19446 7052 20198
rect 7116 19990 7144 22200
rect 7484 22114 7512 22200
rect 7760 22137 7788 22743
rect 7838 22200 7894 23000
rect 8206 22200 8262 23000
rect 8574 22200 8630 23000
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9770 22200 9826 23000
rect 10138 22200 10194 23000
rect 10506 22200 10562 23000
rect 10874 22200 10930 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12070 22200 12126 23000
rect 12438 22200 12494 23000
rect 12806 22200 12862 23000
rect 13174 22200 13230 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14370 22200 14426 23000
rect 14738 22200 14794 23000
rect 15106 22200 15162 23000
rect 15474 22200 15530 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16670 22200 16726 23000
rect 16776 22222 16988 22250
rect 7392 22086 7512 22114
rect 7746 22128 7802 22137
rect 7392 20602 7420 22086
rect 7746 22063 7802 22072
rect 7470 21992 7526 22001
rect 7470 21927 7526 21936
rect 7484 21729 7512 21927
rect 7470 21720 7526 21729
rect 7470 21655 7526 21664
rect 7564 21616 7616 21622
rect 7564 21558 7616 21564
rect 7576 21078 7604 21558
rect 7564 21072 7616 21078
rect 7564 21014 7616 21020
rect 7380 20596 7432 20602
rect 7380 20538 7432 20544
rect 7852 20466 7880 22200
rect 8220 21026 8248 22200
rect 8128 20998 8248 21026
rect 7472 20460 7524 20466
rect 7472 20402 7524 20408
rect 7840 20460 7892 20466
rect 8128 20448 8156 20998
rect 8208 20868 8260 20874
rect 8208 20810 8260 20816
rect 8220 20602 8248 20810
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8208 20460 8260 20466
rect 8128 20420 8208 20448
rect 7840 20402 7892 20408
rect 8208 20402 8260 20408
rect 8484 20460 8536 20466
rect 8588 20448 8616 22200
rect 8668 20596 8720 20602
rect 8668 20538 8720 20544
rect 8536 20420 8616 20448
rect 8484 20402 8536 20408
rect 7380 20256 7432 20262
rect 7380 20198 7432 20204
rect 7104 19984 7156 19990
rect 7104 19926 7156 19932
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7194 19816 7250 19825
rect 7116 19689 7144 19790
rect 7194 19751 7250 19760
rect 7102 19680 7158 19689
rect 7102 19615 7158 19624
rect 7102 19544 7158 19553
rect 7102 19479 7158 19488
rect 7012 19440 7064 19446
rect 7012 19382 7064 19388
rect 7012 19304 7064 19310
rect 6918 19272 6974 19281
rect 7012 19246 7064 19252
rect 6918 19207 6974 19216
rect 6932 19174 6960 19207
rect 6552 19168 6604 19174
rect 6552 19110 6604 19116
rect 6828 19168 6880 19174
rect 6828 19110 6880 19116
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6736 18964 6788 18970
rect 6656 18924 6736 18952
rect 6460 18760 6512 18766
rect 6460 18702 6512 18708
rect 6380 18584 6592 18612
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 6000 18148 6052 18154
rect 6000 18090 6052 18096
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6288 17610 6316 17818
rect 6276 17604 6328 17610
rect 6276 17546 6328 17552
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 6000 17536 6052 17542
rect 6564 17513 6592 18584
rect 6000 17478 6052 17484
rect 6550 17504 6606 17513
rect 5920 16590 5948 17478
rect 6012 16726 6040 17478
rect 6148 17436 6456 17456
rect 6550 17439 6606 17448
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6552 17332 6604 17338
rect 6552 17274 6604 17280
rect 6184 17264 6236 17270
rect 6184 17206 6236 17212
rect 6196 17105 6224 17206
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6182 17096 6238 17105
rect 6182 17031 6238 17040
rect 6196 16726 6224 17031
rect 6274 16824 6330 16833
rect 6274 16759 6330 16768
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6184 16720 6236 16726
rect 6184 16662 6236 16668
rect 6288 16590 6316 16759
rect 6380 16590 6408 17138
rect 6460 17128 6512 17134
rect 6460 17070 6512 17076
rect 6472 16794 6500 17070
rect 6460 16788 6512 16794
rect 6460 16730 6512 16736
rect 5908 16584 5960 16590
rect 5908 16526 5960 16532
rect 6000 16584 6052 16590
rect 6000 16526 6052 16532
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5920 16250 5948 16390
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5908 16108 5960 16114
rect 5908 16050 5960 16056
rect 5920 15978 5948 16050
rect 5908 15972 5960 15978
rect 5908 15914 5960 15920
rect 5828 15558 5948 15586
rect 5816 15496 5868 15502
rect 5816 15438 5868 15444
rect 5722 15056 5778 15065
rect 5722 14991 5778 15000
rect 5736 14618 5764 14991
rect 5724 14612 5776 14618
rect 5724 14554 5776 14560
rect 5736 13394 5764 14554
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5828 12646 5856 15438
rect 5920 14600 5948 15558
rect 6012 14822 6040 16526
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 6092 16176 6144 16182
rect 6564 16130 6592 17274
rect 6092 16118 6144 16124
rect 6104 15910 6132 16118
rect 6288 16102 6592 16130
rect 6184 16040 6236 16046
rect 6184 15982 6236 15988
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 6196 15706 6224 15982
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6288 15502 6316 16102
rect 6552 16040 6604 16046
rect 6552 15982 6604 15988
rect 6460 15972 6512 15978
rect 6460 15914 6512 15920
rect 6276 15496 6328 15502
rect 6276 15438 6328 15444
rect 6472 15434 6500 15914
rect 6564 15502 6592 15982
rect 6656 15910 6684 18924
rect 6736 18906 6788 18912
rect 6840 18698 6868 19110
rect 6736 18692 6788 18698
rect 6736 18634 6788 18640
rect 6828 18692 6880 18698
rect 6828 18634 6880 18640
rect 6748 18601 6776 18634
rect 6734 18592 6790 18601
rect 6734 18527 6790 18536
rect 6734 18456 6790 18465
rect 6734 18391 6790 18400
rect 6748 18290 6776 18391
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 6748 18057 6776 18226
rect 6840 18222 6868 18634
rect 7024 18465 7052 19246
rect 7010 18456 7066 18465
rect 7010 18391 7066 18400
rect 6920 18352 6972 18358
rect 6920 18294 6972 18300
rect 6828 18216 6880 18222
rect 6828 18158 6880 18164
rect 6734 18048 6790 18057
rect 6734 17983 6790 17992
rect 6932 17882 6960 18294
rect 7012 18284 7064 18290
rect 7012 18226 7064 18232
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6828 17740 6880 17746
rect 6828 17682 6880 17688
rect 6736 17128 6788 17134
rect 6736 17070 6788 17076
rect 6748 16250 6776 17070
rect 6840 16726 6868 17682
rect 7024 17678 7052 18226
rect 7012 17672 7064 17678
rect 7012 17614 7064 17620
rect 7116 17338 7144 19479
rect 7208 18426 7236 19751
rect 7288 19712 7340 19718
rect 7288 19654 7340 19660
rect 7300 19514 7328 19654
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7392 19334 7420 20198
rect 7300 19306 7420 19334
rect 7300 19224 7328 19306
rect 7300 19196 7420 19224
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 7300 18426 7328 18906
rect 7392 18766 7420 19196
rect 7484 18970 7512 20402
rect 7564 20052 7616 20058
rect 7564 19994 7616 20000
rect 7576 19334 7604 19994
rect 7748 19848 7800 19854
rect 7748 19790 7800 19796
rect 7760 19334 7788 19790
rect 7545 19306 7604 19334
rect 7668 19306 7788 19334
rect 7545 19258 7573 19306
rect 7545 19230 7604 19258
rect 7472 18964 7524 18970
rect 7472 18906 7524 18912
rect 7380 18760 7432 18766
rect 7380 18702 7432 18708
rect 7470 18456 7526 18465
rect 7196 18420 7248 18426
rect 7196 18362 7248 18368
rect 7288 18420 7340 18426
rect 7470 18391 7526 18400
rect 7288 18362 7340 18368
rect 7484 18290 7512 18391
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7286 17912 7342 17921
rect 7286 17847 7342 17856
rect 7300 17678 7328 17847
rect 7288 17672 7340 17678
rect 7288 17614 7340 17620
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7104 17332 7156 17338
rect 7104 17274 7156 17280
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 6828 16720 6880 16726
rect 6828 16662 6880 16668
rect 6736 16244 6788 16250
rect 6736 16186 6788 16192
rect 6736 15972 6788 15978
rect 6736 15914 6788 15920
rect 6644 15904 6696 15910
rect 6644 15846 6696 15852
rect 6552 15496 6604 15502
rect 6552 15438 6604 15444
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6564 15162 6592 15438
rect 6748 15178 6776 15914
rect 6552 15156 6604 15162
rect 6552 15098 6604 15104
rect 6656 15150 6776 15178
rect 6092 14884 6144 14890
rect 6092 14826 6144 14832
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 5920 14572 6040 14600
rect 5908 14476 5960 14482
rect 5908 14418 5960 14424
rect 5920 14074 5948 14418
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6012 14006 6040 14572
rect 6104 14414 6132 14826
rect 6564 14482 6592 15098
rect 6656 14822 6684 15150
rect 6736 15020 6788 15026
rect 6840 15008 6868 16662
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6920 15972 6972 15978
rect 7024 15960 7052 16526
rect 6972 15932 7052 15960
rect 6920 15914 6972 15920
rect 7010 15192 7066 15201
rect 7010 15127 7066 15136
rect 6788 14980 6868 15008
rect 6736 14962 6788 14968
rect 6644 14816 6696 14822
rect 6644 14758 6696 14764
rect 6656 14618 6684 14758
rect 6644 14612 6696 14618
rect 6644 14554 6696 14560
rect 6748 14482 6776 14962
rect 7024 14890 7052 15127
rect 7116 15026 7144 16934
rect 7194 16824 7250 16833
rect 7194 16759 7250 16768
rect 7208 16425 7236 16759
rect 7300 16590 7328 17478
rect 7470 17368 7526 17377
rect 7470 17303 7526 17312
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7288 16584 7340 16590
rect 7288 16526 7340 16532
rect 7194 16416 7250 16425
rect 7194 16351 7250 16360
rect 7208 16250 7236 16351
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7392 15978 7420 17138
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7104 15020 7156 15026
rect 7156 14980 7236 15008
rect 7104 14962 7156 14968
rect 7012 14884 7064 14890
rect 7012 14826 7064 14832
rect 7208 14822 7236 14980
rect 7196 14816 7248 14822
rect 7196 14758 7248 14764
rect 6826 14648 6882 14657
rect 6826 14583 6882 14592
rect 6840 14550 6868 14583
rect 6828 14544 6880 14550
rect 6828 14486 6880 14492
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6092 14408 6144 14414
rect 6092 14350 6144 14356
rect 6734 14376 6790 14385
rect 7300 14362 7328 15302
rect 6734 14311 6736 14320
rect 6788 14311 6790 14320
rect 7208 14334 7328 14362
rect 6736 14282 6788 14288
rect 7208 14278 7236 14334
rect 6552 14272 6604 14278
rect 6550 14240 6552 14249
rect 7196 14272 7248 14278
rect 6604 14240 6606 14249
rect 6148 14172 6456 14192
rect 7288 14272 7340 14278
rect 7196 14214 7248 14220
rect 7286 14240 7288 14249
rect 7340 14240 7342 14249
rect 6550 14175 6606 14184
rect 7286 14175 7342 14184
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 6000 14000 6052 14006
rect 6000 13942 6052 13948
rect 5908 13864 5960 13870
rect 5908 13806 5960 13812
rect 6460 13864 6512 13870
rect 6564 13852 6592 14175
rect 6826 14104 6882 14113
rect 6826 14039 6882 14048
rect 7104 14068 7156 14074
rect 6840 14006 6868 14039
rect 7156 14028 7236 14056
rect 7104 14010 7156 14016
rect 6644 14000 6696 14006
rect 6644 13942 6696 13948
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 6512 13824 6592 13852
rect 6460 13806 6512 13812
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5920 12322 5948 13806
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6380 13394 6408 13738
rect 6552 13728 6604 13734
rect 6552 13670 6604 13676
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6564 13326 6592 13670
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6000 13184 6052 13190
rect 6000 13126 6052 13132
rect 6012 12986 6040 13126
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6460 12912 6512 12918
rect 5998 12880 6054 12889
rect 6460 12854 6512 12860
rect 5998 12815 6054 12824
rect 5724 12300 5776 12306
rect 5724 12242 5776 12248
rect 5828 12294 5948 12322
rect 6012 12306 6040 12815
rect 6472 12714 6500 12854
rect 6460 12708 6512 12714
rect 6460 12650 6512 12656
rect 6564 12646 6592 13262
rect 6552 12640 6604 12646
rect 6552 12582 6604 12588
rect 6000 12300 6052 12306
rect 5552 11478 5672 11506
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 4896 10066 4948 10072
rect 5276 10084 5396 10112
rect 5172 9920 5224 9926
rect 5170 9888 5172 9897
rect 5224 9888 5226 9897
rect 5170 9823 5226 9832
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4988 9716 5040 9722
rect 4988 9658 5040 9664
rect 4908 9489 4936 9658
rect 4894 9480 4950 9489
rect 4894 9415 4950 9424
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4908 8294 4936 9318
rect 5000 8634 5028 9658
rect 5170 9616 5226 9625
rect 5170 9551 5226 9560
rect 5080 9512 5132 9518
rect 5080 9454 5132 9460
rect 5092 9024 5120 9454
rect 5184 9450 5212 9551
rect 5172 9444 5224 9450
rect 5172 9386 5224 9392
rect 5276 9024 5304 10084
rect 5552 10033 5580 11478
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10810 5672 10950
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5632 10464 5684 10470
rect 5632 10406 5684 10412
rect 5538 10024 5594 10033
rect 5356 9988 5408 9994
rect 5538 9959 5594 9968
rect 5356 9930 5408 9936
rect 5368 9722 5396 9930
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5356 9716 5408 9722
rect 5356 9658 5408 9664
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5092 8996 5212 9024
rect 5276 8996 5396 9024
rect 5184 8956 5212 8996
rect 5184 8928 5304 8956
rect 5170 8800 5226 8809
rect 5170 8735 5226 8744
rect 5184 8634 5212 8735
rect 5276 8634 5304 8928
rect 4988 8628 5040 8634
rect 4988 8570 5040 8576
rect 5172 8628 5224 8634
rect 5172 8570 5224 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5262 8528 5318 8537
rect 5262 8463 5264 8472
rect 5316 8463 5318 8472
rect 5264 8434 5316 8440
rect 4908 8266 5028 8294
rect 4896 8016 4948 8022
rect 4896 7958 4948 7964
rect 4908 6934 4936 7958
rect 5000 7410 5028 8266
rect 5172 7948 5224 7954
rect 5172 7890 5224 7896
rect 5080 7744 5132 7750
rect 5080 7686 5132 7692
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4896 6928 4948 6934
rect 4896 6870 4948 6876
rect 4896 6792 4948 6798
rect 4896 6734 4948 6740
rect 4908 6474 4936 6734
rect 5000 6730 5028 7210
rect 4988 6724 5040 6730
rect 4988 6666 5040 6672
rect 4908 6446 5028 6474
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4908 5914 4936 6258
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4804 4140 4856 4146
rect 4804 4082 4856 4088
rect 4804 4004 4856 4010
rect 4804 3946 4856 3952
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4448 2378 4476 2994
rect 4526 2816 4582 2825
rect 4526 2751 4582 2760
rect 4436 2372 4488 2378
rect 4436 2314 4488 2320
rect 4540 1222 4568 2751
rect 4724 2689 4752 3334
rect 4816 3058 4844 3946
rect 4908 3505 4936 5510
rect 5000 5216 5028 6446
rect 5092 6118 5120 7686
rect 5184 7546 5212 7890
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5172 7540 5224 7546
rect 5172 7482 5224 7488
rect 5184 7410 5212 7482
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 5172 6792 5224 6798
rect 5170 6760 5172 6769
rect 5224 6760 5226 6769
rect 5170 6695 5226 6704
rect 5172 6316 5224 6322
rect 5172 6258 5224 6264
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5184 5302 5212 6258
rect 5172 5296 5224 5302
rect 5172 5238 5224 5244
rect 5000 5188 5120 5216
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4894 3496 4950 3505
rect 4894 3431 4950 3440
rect 4804 3052 4856 3058
rect 4804 2994 4856 3000
rect 4710 2680 4766 2689
rect 4710 2615 4766 2624
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4816 1970 4844 2382
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4528 1216 4580 1222
rect 4528 1158 4580 1164
rect 4816 800 4844 1906
rect 4908 1057 4936 3431
rect 5000 2417 5028 5034
rect 5092 4185 5120 5188
rect 5276 4622 5304 7822
rect 5368 7585 5396 8996
rect 5460 8090 5488 9522
rect 5448 8084 5500 8090
rect 5448 8026 5500 8032
rect 5552 7732 5580 9862
rect 5644 9761 5672 10406
rect 5630 9752 5686 9761
rect 5630 9687 5686 9696
rect 5736 9602 5764 12242
rect 5828 11937 5856 12294
rect 6000 12242 6052 12248
rect 5908 12232 5960 12238
rect 5908 12174 5960 12180
rect 5814 11928 5870 11937
rect 5814 11863 5870 11872
rect 5920 11830 5948 12174
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 6012 11762 6040 12038
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 6368 11824 6420 11830
rect 6368 11766 6420 11772
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 5828 11286 5856 11698
rect 5908 11688 5960 11694
rect 5908 11630 5960 11636
rect 5816 11280 5868 11286
rect 5816 11222 5868 11228
rect 5816 11144 5868 11150
rect 5816 11086 5868 11092
rect 5828 10742 5856 11086
rect 5816 10736 5868 10742
rect 5816 10678 5868 10684
rect 5920 10033 5948 11630
rect 6012 11218 6040 11698
rect 6380 11558 6408 11766
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6380 11218 6408 11494
rect 6564 11393 6592 12582
rect 6656 12345 6684 13942
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6748 12918 6776 13466
rect 6736 12912 6788 12918
rect 6736 12854 6788 12860
rect 6840 12782 6868 13738
rect 6920 13728 6972 13734
rect 6920 13670 6972 13676
rect 6932 13462 6960 13670
rect 7024 13530 7052 13874
rect 7012 13524 7064 13530
rect 7012 13466 7064 13472
rect 6920 13456 6972 13462
rect 6920 13398 6972 13404
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6920 12708 6972 12714
rect 6920 12650 6972 12656
rect 6828 12640 6880 12646
rect 6828 12582 6880 12588
rect 6642 12336 6698 12345
rect 6642 12271 6698 12280
rect 6736 12232 6788 12238
rect 6736 12174 6788 12180
rect 6642 11928 6698 11937
rect 6642 11863 6698 11872
rect 6656 11762 6684 11863
rect 6748 11830 6776 12174
rect 6840 12170 6868 12582
rect 6828 12164 6880 12170
rect 6828 12106 6880 12112
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6932 11393 6960 12650
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6550 11384 6606 11393
rect 6550 11319 6606 11328
rect 6918 11384 6974 11393
rect 6918 11319 6974 11328
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6368 11212 6420 11218
rect 6368 11154 6420 11160
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6288 10996 6316 11086
rect 6012 10968 6316 10996
rect 6564 10996 6592 11319
rect 6736 11144 6788 11150
rect 6788 11092 6960 11098
rect 6736 11086 6960 11092
rect 6748 11070 6960 11086
rect 6564 10968 6776 10996
rect 6012 10538 6040 10968
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6550 10432 6606 10441
rect 6550 10367 6606 10376
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5906 10024 5962 10033
rect 5906 9959 5962 9968
rect 5908 9920 5960 9926
rect 5908 9862 5960 9868
rect 5920 9722 5948 9862
rect 5816 9716 5868 9722
rect 5816 9658 5868 9664
rect 5908 9716 5960 9722
rect 5908 9658 5960 9664
rect 5644 9574 5764 9602
rect 5644 9081 5672 9574
rect 5724 9444 5776 9450
rect 5724 9386 5776 9392
rect 5630 9072 5686 9081
rect 5630 9007 5686 9016
rect 5632 8900 5684 8906
rect 5632 8842 5684 8848
rect 5644 8022 5672 8842
rect 5736 8838 5764 9386
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5736 8378 5764 8774
rect 5828 8634 5856 9658
rect 6012 9450 6040 10066
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6458 9616 6514 9625
rect 6458 9551 6460 9560
rect 6512 9551 6514 9560
rect 6460 9522 6512 9528
rect 6000 9444 6052 9450
rect 6000 9386 6052 9392
rect 6564 9353 6592 10367
rect 6644 10056 6696 10062
rect 6642 10024 6644 10033
rect 6696 10024 6698 10033
rect 6642 9959 6698 9968
rect 6644 9920 6696 9926
rect 6644 9862 6696 9868
rect 6550 9344 6606 9353
rect 6550 9279 6606 9288
rect 5998 9072 6054 9081
rect 5998 9007 6054 9016
rect 5908 8900 5960 8906
rect 5908 8842 5960 8848
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5920 8566 5948 8842
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5736 8350 5856 8378
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5632 8016 5684 8022
rect 5632 7958 5684 7964
rect 5736 7954 5764 8230
rect 5724 7948 5776 7954
rect 5724 7890 5776 7896
rect 5724 7744 5776 7750
rect 5552 7704 5724 7732
rect 5724 7686 5776 7692
rect 5354 7576 5410 7585
rect 5354 7511 5410 7520
rect 5630 7576 5686 7585
rect 5828 7562 5856 8350
rect 6012 7993 6040 9007
rect 6564 8820 6592 9279
rect 6656 8974 6684 9862
rect 6644 8968 6696 8974
rect 6644 8910 6696 8916
rect 6748 8820 6776 10968
rect 6826 10976 6882 10985
rect 6826 10911 6882 10920
rect 6840 8888 6868 10911
rect 6932 10266 6960 11070
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6932 10062 6960 10202
rect 6920 10056 6972 10062
rect 6920 9998 6972 10004
rect 6920 9512 6972 9518
rect 7024 9500 7052 12378
rect 7116 12238 7144 13330
rect 7208 13326 7236 14028
rect 7196 13320 7248 13326
rect 7196 13262 7248 13268
rect 7392 12986 7420 15302
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 7196 12844 7248 12850
rect 7196 12786 7248 12792
rect 7208 12442 7236 12786
rect 7288 12776 7340 12782
rect 7288 12718 7340 12724
rect 7380 12776 7432 12782
rect 7380 12718 7432 12724
rect 7300 12442 7328 12718
rect 7196 12436 7248 12442
rect 7196 12378 7248 12384
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7116 11830 7144 12174
rect 7104 11824 7156 11830
rect 7104 11766 7156 11772
rect 7208 11762 7236 12242
rect 7392 12186 7420 12718
rect 7300 12158 7420 12186
rect 7300 11898 7328 12158
rect 7380 12096 7432 12102
rect 7378 12064 7380 12073
rect 7432 12064 7434 12073
rect 7378 11999 7434 12008
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7392 11801 7420 11999
rect 7378 11792 7434 11801
rect 7196 11756 7248 11762
rect 7378 11727 7434 11736
rect 7196 11698 7248 11704
rect 7208 10742 7236 11698
rect 7286 11112 7342 11121
rect 7286 11047 7342 11056
rect 7380 11076 7432 11082
rect 7300 10810 7328 11047
rect 7380 11018 7432 11024
rect 7288 10804 7340 10810
rect 7288 10746 7340 10752
rect 7196 10736 7248 10742
rect 7196 10678 7248 10684
rect 7196 10600 7248 10606
rect 7196 10542 7248 10548
rect 7286 10568 7342 10577
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 7116 9926 7144 10066
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 6972 9472 7052 9500
rect 6920 9454 6972 9460
rect 6932 9110 6960 9454
rect 7012 9376 7064 9382
rect 7012 9318 7064 9324
rect 6920 9104 6972 9110
rect 6920 9046 6972 9052
rect 6840 8860 6960 8888
rect 6564 8792 6684 8820
rect 6748 8792 6868 8820
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6092 8492 6144 8498
rect 6092 8434 6144 8440
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6104 8265 6132 8434
rect 6090 8256 6146 8265
rect 6090 8191 6146 8200
rect 6380 8022 6408 8434
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6368 8016 6420 8022
rect 5998 7984 6054 7993
rect 6472 7993 6500 8366
rect 6552 8356 6604 8362
rect 6552 8298 6604 8304
rect 6368 7958 6420 7964
rect 6458 7984 6514 7993
rect 5998 7919 6054 7928
rect 6458 7919 6514 7928
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 5630 7511 5686 7520
rect 5736 7534 5856 7562
rect 5368 6390 5396 7511
rect 5644 6882 5672 7511
rect 5552 6854 5672 6882
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 5356 6384 5408 6390
rect 5356 6326 5408 6332
rect 5460 5574 5488 6734
rect 5552 5624 5580 6854
rect 5736 6780 5764 7534
rect 6012 6848 6040 7754
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6184 7472 6236 7478
rect 6184 7414 6236 7420
rect 6460 7472 6512 7478
rect 6460 7414 6512 7420
rect 6196 6848 6224 7414
rect 6472 7041 6500 7414
rect 6564 7177 6592 8298
rect 6656 8106 6684 8792
rect 6734 8664 6790 8673
rect 6734 8599 6790 8608
rect 6748 8430 6776 8599
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6656 8078 6776 8106
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6656 7478 6684 7822
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 6644 7336 6696 7342
rect 6644 7278 6696 7284
rect 6550 7168 6606 7177
rect 6550 7103 6606 7112
rect 6458 7032 6514 7041
rect 6458 6967 6514 6976
rect 5920 6820 6040 6848
rect 6104 6820 6224 6848
rect 6656 6848 6684 7278
rect 6748 7041 6776 8078
rect 6840 7818 6868 8792
rect 6932 8378 6960 8860
rect 7024 8673 7052 9318
rect 7010 8664 7066 8673
rect 7010 8599 7066 8608
rect 7208 8514 7236 10542
rect 7286 10503 7342 10512
rect 7300 9897 7328 10503
rect 7392 10198 7420 11018
rect 7484 10538 7512 17303
rect 7576 13190 7604 19230
rect 7668 18426 7696 19306
rect 7852 19258 7880 20402
rect 8024 20392 8076 20398
rect 8024 20334 8076 20340
rect 7932 19780 7984 19786
rect 7932 19722 7984 19728
rect 7760 19230 7880 19258
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7760 18222 7788 19230
rect 7944 19174 7972 19722
rect 8036 19174 8064 20334
rect 8114 19952 8170 19961
rect 8114 19887 8170 19896
rect 8128 19718 8156 19887
rect 8116 19712 8168 19718
rect 8114 19680 8116 19689
rect 8168 19680 8170 19689
rect 8114 19615 8170 19624
rect 8220 19334 8248 20402
rect 8390 20360 8446 20369
rect 8390 20295 8446 20304
rect 8300 19916 8352 19922
rect 8300 19858 8352 19864
rect 8312 19378 8340 19858
rect 8128 19306 8248 19334
rect 8300 19372 8352 19378
rect 8300 19314 8352 19320
rect 7932 19168 7984 19174
rect 7932 19110 7984 19116
rect 8024 19168 8076 19174
rect 8128 19145 8156 19306
rect 8312 19242 8340 19314
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8208 19168 8260 19174
rect 8024 19110 8076 19116
rect 8114 19136 8170 19145
rect 8208 19110 8260 19116
rect 8114 19071 8170 19080
rect 8116 18964 8168 18970
rect 8116 18906 8168 18912
rect 8024 18760 8076 18766
rect 7944 18720 8024 18748
rect 7840 18624 7892 18630
rect 7840 18566 7892 18572
rect 7656 18216 7708 18222
rect 7656 18158 7708 18164
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7668 17610 7696 18158
rect 7852 17882 7880 18566
rect 7944 18426 7972 18720
rect 8024 18702 8076 18708
rect 8128 18630 8156 18906
rect 8024 18624 8076 18630
rect 8024 18566 8076 18572
rect 8116 18624 8168 18630
rect 8116 18566 8168 18572
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 7746 17776 7802 17785
rect 7746 17711 7748 17720
rect 7800 17711 7802 17720
rect 7932 17740 7984 17746
rect 7748 17682 7800 17688
rect 7932 17682 7984 17688
rect 7656 17604 7708 17610
rect 7656 17546 7708 17552
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7760 15881 7788 17478
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7852 16658 7880 17138
rect 7944 16726 7972 17682
rect 7932 16720 7984 16726
rect 7932 16662 7984 16668
rect 7840 16652 7892 16658
rect 7840 16594 7892 16600
rect 7746 15872 7802 15881
rect 7746 15807 7802 15816
rect 7654 15736 7710 15745
rect 7654 15671 7710 15680
rect 7668 13734 7696 15671
rect 7852 15570 7880 16594
rect 8036 16454 8064 18566
rect 8114 18456 8170 18465
rect 8114 18391 8170 18400
rect 8128 18290 8156 18391
rect 8116 18284 8168 18290
rect 8116 18226 8168 18232
rect 8116 18148 8168 18154
rect 8116 18090 8168 18096
rect 8128 17785 8156 18090
rect 8114 17776 8170 17785
rect 8114 17711 8170 17720
rect 8220 17270 8248 19110
rect 8312 18358 8340 19178
rect 8404 18902 8432 20295
rect 8496 19174 8524 20402
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8588 19961 8616 20198
rect 8574 19952 8630 19961
rect 8574 19887 8630 19896
rect 8680 19417 8708 20538
rect 8956 20466 8984 22200
rect 9312 20596 9364 20602
rect 9312 20538 9364 20544
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 9128 20392 9180 20398
rect 9128 20334 9180 20340
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 9140 19904 9168 20334
rect 9218 20088 9274 20097
rect 9218 20023 9274 20032
rect 8956 19876 9168 19904
rect 8760 19848 8812 19854
rect 8760 19790 8812 19796
rect 8666 19408 8722 19417
rect 8576 19372 8628 19378
rect 8666 19343 8722 19352
rect 8576 19314 8628 19320
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8392 18896 8444 18902
rect 8392 18838 8444 18844
rect 8496 18850 8524 18906
rect 8588 18850 8616 19314
rect 8772 19156 8800 19790
rect 8956 19553 8984 19876
rect 9128 19780 9180 19786
rect 9128 19722 9180 19728
rect 9140 19553 9168 19722
rect 9232 19718 9260 20023
rect 9220 19712 9272 19718
rect 9220 19654 9272 19660
rect 8942 19544 8998 19553
rect 8942 19479 8998 19488
rect 9126 19544 9182 19553
rect 9324 19514 9352 20538
rect 9416 20262 9444 22200
rect 9496 20528 9548 20534
rect 9496 20470 9548 20476
rect 9404 20256 9456 20262
rect 9404 20198 9456 20204
rect 9416 19786 9444 20198
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 9126 19479 9182 19488
rect 9312 19508 9364 19514
rect 9312 19450 9364 19456
rect 9508 19394 9536 20470
rect 9680 20460 9732 20466
rect 9680 20402 9732 20408
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9600 19514 9628 19790
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9128 19372 9180 19378
rect 9508 19366 9628 19394
rect 9128 19314 9180 19320
rect 8680 19128 8800 19156
rect 8680 18970 8708 19128
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 8668 18964 8720 18970
rect 8668 18906 8720 18912
rect 9140 18902 9168 19314
rect 9496 19304 9548 19310
rect 9496 19246 9548 19252
rect 9508 19009 9536 19246
rect 9494 19000 9550 19009
rect 9494 18935 9550 18944
rect 9128 18896 9180 18902
rect 8496 18822 8800 18850
rect 9128 18838 9180 18844
rect 8392 18760 8444 18766
rect 8392 18702 8444 18708
rect 8482 18728 8538 18737
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8300 18216 8352 18222
rect 8300 18158 8352 18164
rect 8320 18068 8348 18158
rect 8312 18040 8348 18068
rect 8312 17882 8340 18040
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 8404 17338 8432 18702
rect 8482 18663 8538 18672
rect 8496 18465 8524 18663
rect 8772 18578 8800 18822
rect 9600 18816 9628 19366
rect 9532 18788 9628 18816
rect 9532 18766 9560 18788
rect 9496 18760 9560 18766
rect 9548 18720 9560 18760
rect 9496 18702 9548 18708
rect 8772 18550 8984 18578
rect 8482 18456 8538 18465
rect 8482 18391 8538 18400
rect 8760 18352 8812 18358
rect 8758 18320 8760 18329
rect 8812 18320 8814 18329
rect 8668 18284 8720 18290
rect 8758 18255 8814 18264
rect 8668 18226 8720 18232
rect 8680 18136 8708 18226
rect 8760 18216 8812 18222
rect 8956 18204 8984 18550
rect 9218 18456 9274 18465
rect 9048 18414 9218 18442
rect 9048 18358 9076 18414
rect 9218 18391 9274 18400
rect 9036 18352 9088 18358
rect 9036 18294 9088 18300
rect 9218 18320 9274 18329
rect 9218 18255 9274 18264
rect 9588 18284 9640 18290
rect 9232 18204 9260 18255
rect 9588 18226 9640 18232
rect 9312 18216 9364 18222
rect 8956 18176 9168 18204
rect 9232 18176 9312 18204
rect 8760 18158 8812 18164
rect 8588 18108 8708 18136
rect 8484 17876 8536 17882
rect 8484 17818 8536 17824
rect 8496 17746 8524 17818
rect 8588 17814 8616 18108
rect 8772 18068 8800 18158
rect 8680 18040 8800 18068
rect 8576 17808 8628 17814
rect 8576 17750 8628 17756
rect 8484 17740 8536 17746
rect 8484 17682 8536 17688
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8208 17264 8260 17270
rect 8208 17206 8260 17212
rect 8300 17264 8352 17270
rect 8300 17206 8352 17212
rect 8312 16969 8340 17206
rect 8496 17066 8524 17682
rect 8680 17338 8708 18040
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 9140 17921 9168 18176
rect 9600 18193 9628 18226
rect 9312 18158 9364 18164
rect 9402 18184 9458 18193
rect 9402 18119 9458 18128
rect 9586 18184 9642 18193
rect 9586 18119 9642 18128
rect 9126 17912 9182 17921
rect 9126 17847 9182 17856
rect 8668 17332 8720 17338
rect 8668 17274 8720 17280
rect 9140 17270 9168 17847
rect 9416 17338 9444 18119
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9218 17232 9274 17241
rect 8668 17196 8720 17202
rect 9218 17167 9220 17176
rect 8668 17138 8720 17144
rect 9272 17167 9274 17176
rect 9220 17138 9272 17144
rect 8484 17060 8536 17066
rect 8484 17002 8536 17008
rect 8298 16960 8354 16969
rect 8298 16895 8354 16904
rect 8496 16810 8524 17002
rect 8576 16992 8628 16998
rect 8680 16946 8708 17138
rect 9128 17128 9180 17134
rect 8850 17096 8906 17105
rect 9128 17070 9180 17076
rect 8850 17031 8852 17040
rect 8904 17031 8906 17040
rect 8852 17002 8904 17008
rect 8628 16940 8708 16946
rect 8576 16934 8708 16940
rect 8588 16918 8708 16934
rect 8496 16782 8616 16810
rect 8588 16658 8616 16782
rect 8576 16652 8628 16658
rect 8576 16594 8628 16600
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8116 16516 8168 16522
rect 8116 16458 8168 16464
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 8022 16280 8078 16289
rect 8022 16215 8078 16224
rect 7840 15564 7892 15570
rect 7840 15506 7892 15512
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7656 13728 7708 13734
rect 7656 13670 7708 13676
rect 7760 13530 7788 15302
rect 7944 15162 7972 15438
rect 8036 15201 8064 16215
rect 8128 16114 8156 16458
rect 8220 16250 8248 16458
rect 8392 16448 8444 16454
rect 8392 16390 8444 16396
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8404 16130 8432 16390
rect 8496 16289 8524 16526
rect 8482 16280 8538 16289
rect 8482 16215 8538 16224
rect 8116 16108 8168 16114
rect 8404 16102 8524 16130
rect 8116 16050 8168 16056
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 8392 16040 8444 16046
rect 8392 15982 8444 15988
rect 8022 15192 8078 15201
rect 7932 15156 7984 15162
rect 8022 15127 8078 15136
rect 7932 15098 7984 15104
rect 8036 15042 8064 15127
rect 7944 15014 8064 15042
rect 7840 14340 7892 14346
rect 7840 14282 7892 14288
rect 7748 13524 7800 13530
rect 7748 13466 7800 13472
rect 7564 13184 7616 13190
rect 7564 13126 7616 13132
rect 7748 12912 7800 12918
rect 7748 12854 7800 12860
rect 7564 12776 7616 12782
rect 7564 12718 7616 12724
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7380 10192 7432 10198
rect 7380 10134 7432 10140
rect 7380 9988 7432 9994
rect 7380 9930 7432 9936
rect 7286 9888 7342 9897
rect 7286 9823 7342 9832
rect 7392 9330 7420 9930
rect 7472 9512 7524 9518
rect 7472 9454 7524 9460
rect 7300 9302 7420 9330
rect 7300 8922 7328 9302
rect 7378 9208 7434 9217
rect 7484 9178 7512 9454
rect 7378 9143 7434 9152
rect 7472 9172 7524 9178
rect 7392 9058 7420 9143
rect 7472 9114 7524 9120
rect 7392 9030 7512 9058
rect 7300 8894 7420 8922
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7107 8486 7236 8514
rect 6932 8350 7052 8378
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6828 7472 6880 7478
rect 6826 7440 6828 7449
rect 6880 7440 6882 7449
rect 6826 7375 6882 7384
rect 7024 7290 7052 8350
rect 7107 8106 7135 8486
rect 7196 8288 7248 8294
rect 7300 8276 7328 8774
rect 7392 8362 7420 8894
rect 7484 8673 7512 9030
rect 7470 8664 7526 8673
rect 7470 8599 7526 8608
rect 7380 8356 7432 8362
rect 7380 8298 7432 8304
rect 7248 8248 7328 8276
rect 7472 8288 7524 8294
rect 7378 8256 7434 8265
rect 7196 8230 7248 8236
rect 7472 8230 7524 8236
rect 7378 8191 7434 8200
rect 7107 8078 7236 8106
rect 6840 7262 7052 7290
rect 6734 7032 6790 7041
rect 6734 6967 6790 6976
rect 6736 6860 6788 6866
rect 6656 6820 6736 6848
rect 5816 6792 5868 6798
rect 5736 6752 5816 6780
rect 5816 6734 5868 6740
rect 5920 6662 5948 6820
rect 5632 6656 5684 6662
rect 5908 6656 5960 6662
rect 5632 6598 5684 6604
rect 5722 6624 5778 6633
rect 5644 5692 5672 6598
rect 6104 6644 6132 6820
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 5908 6598 5960 6604
rect 6012 6616 6132 6644
rect 5722 6559 5778 6568
rect 5736 6458 5764 6559
rect 5814 6488 5870 6497
rect 5724 6452 5776 6458
rect 6012 6458 6040 6616
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 5814 6423 5816 6432
rect 5724 6394 5776 6400
rect 5868 6423 5870 6432
rect 6000 6452 6052 6458
rect 5816 6394 5868 6400
rect 6000 6394 6052 6400
rect 6196 6412 6408 6440
rect 5736 6310 6040 6338
rect 6196 6322 6224 6412
rect 6380 6372 6408 6412
rect 6573 6372 6601 6666
rect 6656 6633 6684 6820
rect 6736 6802 6788 6808
rect 6642 6624 6698 6633
rect 6840 6610 6868 7262
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6932 6746 6960 7142
rect 7104 6928 7156 6934
rect 7104 6870 7156 6876
rect 6932 6718 7052 6746
rect 6642 6559 6698 6568
rect 6748 6582 6868 6610
rect 6918 6624 6974 6633
rect 6748 6474 6776 6582
rect 6918 6559 6974 6568
rect 6274 6352 6330 6361
rect 5736 6254 5764 6310
rect 5724 6248 5776 6254
rect 5724 6190 5776 6196
rect 5814 6216 5870 6225
rect 6012 6186 6040 6310
rect 6184 6316 6236 6322
rect 6380 6344 6601 6372
rect 6656 6446 6776 6474
rect 6828 6452 6880 6458
rect 6274 6287 6330 6296
rect 6184 6258 6236 6264
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 5814 6151 5870 6160
rect 6000 6180 6052 6186
rect 5724 5704 5776 5710
rect 5644 5664 5724 5692
rect 5724 5646 5776 5652
rect 5552 5596 5672 5624
rect 5448 5568 5500 5574
rect 5448 5510 5500 5516
rect 5644 5250 5672 5596
rect 5724 5568 5776 5574
rect 5724 5510 5776 5516
rect 5736 5370 5764 5510
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5540 5228 5592 5234
rect 5644 5222 5764 5250
rect 5540 5170 5592 5176
rect 5552 5137 5580 5170
rect 5538 5128 5594 5137
rect 5538 5063 5594 5072
rect 5632 5092 5684 5098
rect 5632 5034 5684 5040
rect 5448 4684 5500 4690
rect 5448 4626 5500 4632
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5262 4448 5318 4457
rect 5262 4383 5318 4392
rect 5078 4176 5134 4185
rect 5078 4111 5134 4120
rect 5276 4078 5304 4383
rect 5080 4072 5132 4078
rect 5264 4072 5316 4078
rect 5080 4014 5132 4020
rect 5170 4040 5226 4049
rect 4986 2408 5042 2417
rect 4986 2343 5042 2352
rect 4894 1048 4950 1057
rect 4894 983 4950 992
rect 5092 921 5120 4014
rect 5264 4014 5316 4020
rect 5170 3975 5226 3984
rect 5184 3738 5212 3975
rect 5368 3942 5396 4490
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5184 1329 5212 3334
rect 5262 3224 5318 3233
rect 5262 3159 5318 3168
rect 5170 1320 5226 1329
rect 5170 1255 5226 1264
rect 5276 1170 5304 3159
rect 5368 3058 5396 3878
rect 5460 3602 5488 4626
rect 5540 4616 5592 4622
rect 5644 4593 5672 5034
rect 5540 4558 5592 4564
rect 5630 4584 5686 4593
rect 5552 4185 5580 4558
rect 5630 4519 5686 4528
rect 5736 4468 5764 5222
rect 5828 5098 5856 6151
rect 6000 6122 6052 6128
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5920 5545 5948 5646
rect 5906 5536 5962 5545
rect 5906 5471 5962 5480
rect 5906 5264 5962 5273
rect 5906 5199 5908 5208
rect 5960 5199 5962 5208
rect 5908 5170 5960 5176
rect 5816 5092 5868 5098
rect 5816 5034 5868 5040
rect 5908 5024 5960 5030
rect 5908 4966 5960 4972
rect 5920 4826 5948 4966
rect 5908 4820 5960 4826
rect 5908 4762 5960 4768
rect 6012 4706 6040 5782
rect 6104 5778 6132 6190
rect 6092 5772 6144 5778
rect 6092 5714 6144 5720
rect 6288 5710 6316 6287
rect 6368 6248 6420 6254
rect 6366 6216 6368 6225
rect 6460 6248 6512 6254
rect 6420 6216 6422 6225
rect 6460 6190 6512 6196
rect 6550 6216 6606 6225
rect 6366 6151 6422 6160
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6472 5556 6500 6190
rect 6550 6151 6606 6160
rect 6564 5914 6592 6151
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6472 5528 6592 5556
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 5920 4678 6040 4706
rect 6104 4690 6132 4966
rect 6564 4842 6592 5528
rect 6656 5370 6684 6446
rect 6828 6394 6880 6400
rect 6727 6316 6779 6322
rect 6727 6258 6779 6264
rect 6739 6202 6767 6258
rect 6739 6174 6776 6202
rect 6748 5681 6776 6174
rect 6734 5672 6790 5681
rect 6734 5607 6790 5616
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6734 5264 6790 5273
rect 6734 5199 6790 5208
rect 6748 5166 6776 5199
rect 6736 5160 6788 5166
rect 6736 5102 6788 5108
rect 6840 5030 6868 6394
rect 6932 6186 6960 6559
rect 7024 6458 7052 6718
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 6920 6180 6972 6186
rect 6920 6122 6972 6128
rect 7010 5944 7066 5953
rect 7010 5879 7012 5888
rect 7064 5879 7066 5888
rect 7012 5850 7064 5856
rect 7116 5778 7144 6870
rect 7208 6322 7236 8078
rect 7392 8022 7420 8191
rect 7380 8016 7432 8022
rect 7380 7958 7432 7964
rect 7484 7834 7512 8230
rect 7300 7806 7512 7834
rect 7300 7546 7328 7806
rect 7380 7744 7432 7750
rect 7380 7686 7432 7692
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7208 5817 7236 6258
rect 7300 6225 7328 6938
rect 7286 6216 7342 6225
rect 7286 6151 7342 6160
rect 7286 5944 7342 5953
rect 7286 5879 7342 5888
rect 7194 5808 7250 5817
rect 7104 5772 7156 5778
rect 7300 5778 7328 5879
rect 7194 5743 7250 5752
rect 7288 5772 7340 5778
rect 7104 5714 7156 5720
rect 7288 5714 7340 5720
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6828 5024 6880 5030
rect 6828 4966 6880 4972
rect 6564 4814 6776 4842
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6092 4684 6144 4690
rect 5644 4440 5764 4468
rect 5816 4480 5868 4486
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5644 4010 5672 4440
rect 5816 4422 5868 4428
rect 5722 4312 5778 4321
rect 5722 4247 5724 4256
rect 5776 4247 5778 4256
rect 5724 4218 5776 4224
rect 5724 4072 5776 4078
rect 5724 4014 5776 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 5736 3738 5764 4014
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5630 3632 5686 3641
rect 5448 3596 5500 3602
rect 5630 3567 5686 3576
rect 5724 3596 5776 3602
rect 5448 3538 5500 3544
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3097 5488 3334
rect 5446 3088 5502 3097
rect 5356 3052 5408 3058
rect 5446 3023 5502 3032
rect 5356 2994 5408 3000
rect 5644 2990 5672 3567
rect 5724 3538 5776 3544
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5736 2650 5764 3538
rect 5828 3398 5856 4422
rect 5816 3392 5868 3398
rect 5816 3334 5868 3340
rect 5814 3224 5870 3233
rect 5814 3159 5816 3168
rect 5868 3159 5870 3168
rect 5816 3130 5868 3136
rect 5920 2961 5948 4678
rect 6092 4626 6144 4632
rect 6368 4616 6420 4622
rect 6366 4584 6368 4593
rect 6552 4616 6604 4622
rect 6420 4584 6422 4593
rect 6552 4558 6604 4564
rect 6366 4519 6422 4528
rect 6148 4380 6456 4400
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 5998 4312 6054 4321
rect 6148 4304 6456 4324
rect 5998 4247 6000 4256
rect 6052 4247 6054 4256
rect 6000 4218 6052 4224
rect 6564 4162 6592 4558
rect 6656 4282 6684 4694
rect 6644 4276 6696 4282
rect 6644 4218 6696 4224
rect 6748 4214 6776 4814
rect 6932 4808 6960 5646
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7116 5409 7144 5510
rect 7102 5400 7158 5409
rect 7102 5335 7158 5344
rect 6840 4780 6960 4808
rect 6380 4134 6592 4162
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6840 4162 6868 4780
rect 7010 4720 7066 4729
rect 7010 4655 7012 4664
rect 7064 4655 7066 4664
rect 7012 4626 7064 4632
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7194 4312 7250 4321
rect 7194 4247 7250 4256
rect 7208 4214 7236 4247
rect 7196 4208 7248 4214
rect 6840 4134 6960 4162
rect 7196 4150 7248 4156
rect 6000 3664 6052 3670
rect 6000 3606 6052 3612
rect 6090 3632 6146 3641
rect 6012 3505 6040 3606
rect 6090 3567 6092 3576
rect 6144 3567 6146 3576
rect 6276 3596 6328 3602
rect 6092 3538 6144 3544
rect 6380 3584 6408 4134
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6460 3936 6512 3942
rect 6460 3878 6512 3884
rect 6328 3556 6408 3584
rect 6276 3538 6328 3544
rect 5998 3496 6054 3505
rect 6472 3466 6500 3878
rect 5998 3431 6054 3440
rect 6460 3460 6512 3466
rect 5906 2952 5962 2961
rect 5906 2887 5962 2896
rect 6012 2854 6040 3431
rect 6460 3402 6512 3408
rect 6644 3392 6696 3398
rect 6550 3360 6606 3369
rect 6148 3292 6456 3312
rect 6644 3334 6696 3340
rect 6550 3295 6606 3304
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 6564 3194 6592 3295
rect 6552 3188 6604 3194
rect 6552 3130 6604 3136
rect 6092 3052 6144 3058
rect 6092 2994 6144 3000
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 5814 2680 5870 2689
rect 5724 2644 5776 2650
rect 5814 2615 5870 2624
rect 5724 2586 5776 2592
rect 5828 2514 5856 2615
rect 5816 2508 5868 2514
rect 5816 2450 5868 2456
rect 5722 2272 5778 2281
rect 5722 2207 5778 2216
rect 5630 1592 5686 1601
rect 5630 1527 5686 1536
rect 5184 1142 5304 1170
rect 5078 912 5134 921
rect 5078 847 5134 856
rect 5184 800 5212 1142
rect 5644 800 5672 1527
rect 5736 1290 5764 2207
rect 5920 1902 5948 2790
rect 6104 2650 6132 2994
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6092 2644 6144 2650
rect 6092 2586 6144 2592
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 5998 2136 6054 2145
rect 6148 2128 6456 2148
rect 5998 2071 6000 2080
rect 6052 2071 6054 2080
rect 6000 2042 6052 2048
rect 5908 1896 5960 1902
rect 5908 1838 5960 1844
rect 5998 1864 6054 1873
rect 5998 1799 6054 1808
rect 5724 1284 5776 1290
rect 5724 1226 5776 1232
rect 6012 800 6040 1799
rect 6564 1442 6592 2858
rect 6472 1414 6592 1442
rect 6472 800 6500 1414
rect 6656 950 6684 3334
rect 6748 3194 6776 3946
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6840 3398 6868 3674
rect 6828 3392 6880 3398
rect 6828 3334 6880 3340
rect 6736 3188 6788 3194
rect 6932 3176 6960 4134
rect 7104 4140 7156 4146
rect 7104 4082 7156 4088
rect 7010 3768 7066 3777
rect 7116 3738 7144 4082
rect 7010 3703 7066 3712
rect 7104 3732 7156 3738
rect 6736 3130 6788 3136
rect 6840 3148 6960 3176
rect 6840 3074 6868 3148
rect 6748 3046 6868 3074
rect 6748 1737 6776 3046
rect 6828 2984 6880 2990
rect 6828 2926 6880 2932
rect 6734 1728 6790 1737
rect 6734 1663 6790 1672
rect 6644 944 6696 950
rect 6644 886 6696 892
rect 6840 800 6868 2926
rect 7024 2854 7052 3703
rect 7104 3674 7156 3680
rect 7116 2990 7144 3674
rect 7104 2984 7156 2990
rect 7104 2926 7156 2932
rect 7012 2848 7064 2854
rect 7300 2836 7328 4422
rect 7392 4321 7420 7686
rect 7484 7585 7512 7686
rect 7470 7576 7526 7585
rect 7470 7511 7526 7520
rect 7484 7410 7512 7511
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7472 6656 7524 6662
rect 7470 6624 7472 6633
rect 7524 6624 7526 6633
rect 7470 6559 7526 6568
rect 7470 6216 7526 6225
rect 7470 6151 7526 6160
rect 7484 5914 7512 6151
rect 7472 5908 7524 5914
rect 7472 5850 7524 5856
rect 7484 5642 7512 5850
rect 7576 5778 7604 12718
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7668 11898 7696 12038
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7760 11778 7788 12854
rect 7668 11750 7788 11778
rect 7668 8265 7696 11750
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10810 7788 11154
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7852 10606 7880 14282
rect 7944 14278 7972 15014
rect 8024 14952 8076 14958
rect 8024 14894 8076 14900
rect 8036 14657 8064 14894
rect 8022 14648 8078 14657
rect 8022 14583 8078 14592
rect 8220 14550 8248 15982
rect 8404 15570 8432 15982
rect 8392 15564 8444 15570
rect 8392 15506 8444 15512
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8208 14544 8260 14550
rect 8208 14486 8260 14492
rect 8024 14476 8076 14482
rect 8024 14418 8076 14424
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7932 13796 7984 13802
rect 7932 13738 7984 13744
rect 7944 13190 7972 13738
rect 8036 13530 8064 14418
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8024 13524 8076 13530
rect 8024 13466 8076 13472
rect 8022 13288 8078 13297
rect 8022 13223 8078 13232
rect 7932 13184 7984 13190
rect 7932 13126 7984 13132
rect 7944 10849 7972 13126
rect 8036 12986 8064 13223
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8128 12628 8156 14350
rect 8312 14074 8340 15302
rect 8404 15144 8432 15506
rect 8496 15337 8524 16102
rect 8576 15904 8628 15910
rect 8574 15872 8576 15881
rect 8628 15872 8630 15881
rect 8574 15807 8630 15816
rect 8680 15638 8708 16918
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 8852 16720 8904 16726
rect 8852 16662 8904 16668
rect 8864 15978 8892 16662
rect 8852 15972 8904 15978
rect 8852 15914 8904 15920
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 9140 15706 9168 17070
rect 9404 16788 9456 16794
rect 9404 16730 9456 16736
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8482 15328 8538 15337
rect 8482 15263 8538 15272
rect 8484 15156 8536 15162
rect 8404 15116 8484 15144
rect 8484 15098 8536 15104
rect 8680 15026 8708 15574
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8668 15020 8720 15026
rect 8668 14962 8720 14968
rect 8772 14804 8800 15098
rect 8574 14784 8630 14793
rect 8574 14719 8630 14728
rect 8680 14776 8800 14804
rect 9218 14784 9274 14793
rect 8484 14544 8536 14550
rect 8484 14486 8536 14492
rect 8392 14408 8444 14414
rect 8392 14350 8444 14356
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8300 13796 8352 13802
rect 8300 13738 8352 13744
rect 8208 13252 8260 13258
rect 8208 13194 8260 13200
rect 8220 12782 8248 13194
rect 8208 12776 8260 12782
rect 8312 12753 8340 13738
rect 8208 12718 8260 12724
rect 8298 12744 8354 12753
rect 8298 12679 8354 12688
rect 8128 12600 8248 12628
rect 8114 12472 8170 12481
rect 8114 12407 8116 12416
rect 8168 12407 8170 12416
rect 8116 12378 8168 12384
rect 8022 11384 8078 11393
rect 8022 11319 8078 11328
rect 7930 10840 7986 10849
rect 8036 10810 8064 11319
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7930 10775 7986 10784
rect 8024 10804 8076 10810
rect 8024 10746 8076 10752
rect 8128 10606 8156 10950
rect 7840 10600 7892 10606
rect 7840 10542 7892 10548
rect 8116 10600 8168 10606
rect 8116 10542 8168 10548
rect 8024 10532 8076 10538
rect 8024 10474 8076 10480
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7852 9722 7880 10406
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7840 9716 7892 9722
rect 7840 9658 7892 9664
rect 7944 9518 7972 9862
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 8974 7788 9114
rect 7748 8968 7800 8974
rect 7748 8910 7800 8916
rect 7654 8256 7710 8265
rect 7654 8191 7710 8200
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7668 7886 7696 8026
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7668 7546 7696 7822
rect 7656 7540 7708 7546
rect 7656 7482 7708 7488
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7668 6934 7696 7142
rect 7656 6928 7708 6934
rect 7656 6870 7708 6876
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7472 5636 7524 5642
rect 7472 5578 7524 5584
rect 7472 5024 7524 5030
rect 7472 4966 7524 4972
rect 7378 4312 7434 4321
rect 7378 4247 7434 4256
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7012 2790 7064 2796
rect 7116 2808 7328 2836
rect 7010 2680 7066 2689
rect 6920 2644 6972 2650
rect 7010 2615 7066 2624
rect 6920 2586 6972 2592
rect 6932 1737 6960 2586
rect 7024 2514 7052 2615
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7116 2038 7144 2808
rect 7196 2440 7248 2446
rect 7196 2382 7248 2388
rect 7208 2281 7236 2382
rect 7288 2372 7340 2378
rect 7288 2314 7340 2320
rect 7194 2272 7250 2281
rect 7194 2207 7250 2216
rect 7104 2032 7156 2038
rect 7104 1974 7156 1980
rect 6918 1728 6974 1737
rect 6918 1663 6974 1672
rect 7208 1601 7236 2207
rect 7300 2009 7328 2314
rect 7286 2000 7342 2009
rect 7286 1935 7342 1944
rect 7194 1592 7250 1601
rect 7194 1527 7250 1536
rect 7300 800 7328 1935
rect 3160 734 3464 762
rect 3514 0 3570 800
rect 3882 0 3938 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7392 762 7420 4150
rect 7484 2310 7512 4966
rect 7576 2582 7604 5714
rect 7668 5234 7696 6870
rect 7760 5710 7788 8910
rect 7852 8634 7880 9318
rect 7944 8974 7972 9454
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 7840 8492 7892 8498
rect 7840 8434 7892 8440
rect 7852 8106 7880 8434
rect 7944 8430 7972 8910
rect 8036 8498 8064 10474
rect 8128 10062 8156 10542
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8128 9518 8156 9998
rect 8116 9512 8168 9518
rect 8116 9454 8168 9460
rect 8128 9042 8156 9454
rect 8116 9036 8168 9042
rect 8116 8978 8168 8984
rect 8114 8936 8170 8945
rect 8114 8871 8170 8880
rect 8128 8838 8156 8871
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 7932 8424 7984 8430
rect 7932 8366 7984 8372
rect 8114 8392 8170 8401
rect 8024 8356 8076 8362
rect 8114 8327 8170 8336
rect 8024 8298 8076 8304
rect 7852 8078 7972 8106
rect 7944 7834 7972 8078
rect 7852 7806 7972 7834
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 7852 5534 7880 7806
rect 8036 6882 8064 8298
rect 8128 7993 8156 8327
rect 8114 7984 8170 7993
rect 8114 7919 8170 7928
rect 8220 7002 8248 12600
rect 8298 12336 8354 12345
rect 8298 12271 8354 12280
rect 8312 10062 8340 12271
rect 8404 12209 8432 14350
rect 8496 14113 8524 14486
rect 8482 14104 8538 14113
rect 8482 14039 8538 14048
rect 8496 14006 8524 14039
rect 8588 14006 8616 14719
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8576 13864 8628 13870
rect 8576 13806 8628 13812
rect 8484 13728 8536 13734
rect 8484 13670 8536 13676
rect 8496 12782 8524 13670
rect 8484 12776 8536 12782
rect 8484 12718 8536 12724
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12306 8524 12582
rect 8484 12300 8536 12306
rect 8484 12242 8536 12248
rect 8390 12200 8446 12209
rect 8390 12135 8446 12144
rect 8404 11914 8432 12135
rect 8588 12084 8616 13806
rect 8680 13274 8708 14776
rect 8747 14716 9055 14736
rect 9218 14719 9274 14728
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 9126 14648 9182 14657
rect 9126 14583 9182 14592
rect 8760 14476 8812 14482
rect 8760 14418 8812 14424
rect 8772 13870 8800 14418
rect 9140 14414 9168 14583
rect 9232 14482 9260 14719
rect 9416 14498 9444 16730
rect 9508 16658 9536 17614
rect 9692 16969 9720 20402
rect 9784 19786 9812 22200
rect 9862 20632 9918 20641
rect 9862 20567 9918 20576
rect 9876 20369 9904 20567
rect 9862 20360 9918 20369
rect 9862 20295 9918 20304
rect 10152 20097 10180 22200
rect 10520 20466 10548 22200
rect 10692 20800 10744 20806
rect 10692 20742 10744 20748
rect 10704 20466 10732 20742
rect 10888 20602 10916 22200
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10508 20460 10560 20466
rect 10508 20402 10560 20408
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10784 20392 10836 20398
rect 10784 20334 10836 20340
rect 10876 20392 10928 20398
rect 10876 20334 10928 20340
rect 10508 20256 10560 20262
rect 10508 20198 10560 20204
rect 10692 20256 10744 20262
rect 10692 20198 10744 20204
rect 10138 20088 10194 20097
rect 10138 20023 10194 20032
rect 10152 19786 10180 20023
rect 9772 19780 9824 19786
rect 9772 19722 9824 19728
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 9784 18850 9812 19722
rect 9956 19712 10008 19718
rect 9956 19654 10008 19660
rect 10324 19712 10376 19718
rect 10324 19654 10376 19660
rect 9864 19508 9916 19514
rect 9864 19450 9916 19456
rect 9876 19292 9904 19450
rect 9968 19417 9996 19654
rect 10140 19440 10192 19446
rect 9954 19408 10010 19417
rect 9954 19343 10010 19352
rect 10060 19388 10140 19394
rect 10336 19417 10364 19654
rect 10060 19382 10192 19388
rect 10322 19408 10378 19417
rect 10060 19366 10180 19382
rect 10232 19372 10284 19378
rect 9876 19264 9996 19292
rect 9862 19000 9918 19009
rect 9862 18935 9864 18944
rect 9916 18935 9918 18944
rect 9864 18906 9916 18912
rect 9784 18822 9904 18850
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 9784 17649 9812 18702
rect 9876 18306 9904 18822
rect 9968 18426 9996 19264
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9876 18278 9996 18306
rect 9864 18080 9916 18086
rect 9864 18022 9916 18028
rect 9876 17882 9904 18022
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9968 17746 9996 18278
rect 10060 17882 10088 19366
rect 10322 19343 10378 19352
rect 10232 19314 10284 19320
rect 10138 19272 10194 19281
rect 10138 19207 10194 19216
rect 10152 18737 10180 19207
rect 10244 18970 10272 19314
rect 10414 19272 10470 19281
rect 10324 19236 10376 19242
rect 10414 19207 10470 19216
rect 10324 19178 10376 19184
rect 10336 19009 10364 19178
rect 10322 19000 10378 19009
rect 10232 18964 10284 18970
rect 10322 18935 10378 18944
rect 10232 18906 10284 18912
rect 10324 18760 10376 18766
rect 10138 18728 10194 18737
rect 10324 18702 10376 18708
rect 10138 18663 10194 18672
rect 10140 18624 10192 18630
rect 10140 18566 10192 18572
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 10152 17814 10180 18566
rect 10336 18222 10364 18702
rect 10324 18216 10376 18222
rect 10324 18158 10376 18164
rect 10140 17808 10192 17814
rect 10140 17750 10192 17756
rect 9956 17740 10008 17746
rect 9956 17682 10008 17688
rect 10336 17678 10364 18158
rect 10428 18057 10456 19207
rect 10520 18970 10548 20198
rect 10704 20058 10732 20198
rect 10692 20052 10744 20058
rect 10692 19994 10744 20000
rect 10796 19825 10824 20334
rect 10888 20058 10916 20334
rect 10966 20224 11022 20233
rect 10966 20159 11022 20168
rect 10876 20052 10928 20058
rect 10876 19994 10928 20000
rect 10980 19854 11008 20159
rect 11256 19990 11284 22200
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 11716 20584 11744 22200
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11796 20596 11848 20602
rect 11716 20556 11796 20584
rect 11796 20538 11848 20544
rect 11992 20482 12020 20878
rect 12084 20602 12112 22200
rect 12164 21276 12216 21282
rect 12164 21218 12216 21224
rect 12176 20942 12204 21218
rect 12164 20936 12216 20942
rect 12164 20878 12216 20884
rect 12452 20602 12480 22200
rect 12820 20602 12848 22200
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 12440 20596 12492 20602
rect 12440 20538 12492 20544
rect 12808 20596 12860 20602
rect 12808 20538 12860 20544
rect 11888 20460 11940 20466
rect 11992 20454 12112 20482
rect 11888 20402 11940 20408
rect 11900 20058 11928 20402
rect 11978 20088 12034 20097
rect 11888 20052 11940 20058
rect 11978 20023 12034 20032
rect 11888 19994 11940 20000
rect 11244 19984 11296 19990
rect 11244 19926 11296 19932
rect 11704 19916 11756 19922
rect 11704 19858 11756 19864
rect 10968 19848 11020 19854
rect 10598 19816 10654 19825
rect 10782 19816 10838 19825
rect 10654 19774 10732 19802
rect 10598 19751 10654 19760
rect 10704 19530 10732 19774
rect 10968 19790 11020 19796
rect 11060 19848 11112 19854
rect 11060 19790 11112 19796
rect 10782 19751 10838 19760
rect 10704 19502 11008 19530
rect 11072 19514 11100 19790
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11150 19680 11206 19689
rect 11150 19615 11206 19624
rect 10784 19440 10836 19446
rect 10784 19382 10836 19388
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10692 18624 10744 18630
rect 10692 18566 10744 18572
rect 10508 18420 10560 18426
rect 10560 18380 10640 18408
rect 10508 18362 10560 18368
rect 10508 18216 10560 18222
rect 10508 18158 10560 18164
rect 10414 18048 10470 18057
rect 10414 17983 10470 17992
rect 10520 17785 10548 18158
rect 10506 17776 10562 17785
rect 10506 17711 10562 17720
rect 10324 17672 10376 17678
rect 9770 17640 9826 17649
rect 10324 17614 10376 17620
rect 9770 17575 9826 17584
rect 10336 17542 10364 17614
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 9678 16960 9734 16969
rect 9678 16895 9734 16904
rect 9496 16652 9548 16658
rect 9496 16594 9548 16600
rect 9508 16182 9536 16594
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9508 15706 9536 16118
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9600 15706 9628 16050
rect 9678 15736 9734 15745
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9588 15700 9640 15706
rect 9784 15706 9812 17138
rect 9678 15671 9734 15680
rect 9772 15700 9824 15706
rect 9588 15642 9640 15648
rect 9588 15564 9640 15570
rect 9588 15506 9640 15512
rect 9600 15094 9628 15506
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9220 14476 9272 14482
rect 9416 14470 9536 14498
rect 9600 14482 9628 15030
rect 9220 14418 9272 14424
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 9312 14408 9364 14414
rect 9312 14350 9364 14356
rect 9140 13977 9168 14350
rect 9220 14272 9272 14278
rect 9220 14214 9272 14220
rect 9126 13968 9182 13977
rect 9126 13903 9182 13912
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 9128 13456 9180 13462
rect 9128 13398 9180 13404
rect 9034 13288 9090 13297
rect 8680 13246 8892 13274
rect 8668 13184 8720 13190
rect 8668 13126 8720 13132
rect 8760 13184 8812 13190
rect 8760 13126 8812 13132
rect 8680 12986 8708 13126
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8680 12152 8708 12922
rect 8772 12918 8800 13126
rect 8760 12912 8812 12918
rect 8760 12854 8812 12860
rect 8864 12714 8892 13246
rect 9034 13223 9090 13232
rect 9048 12918 9076 13223
rect 9036 12912 9088 12918
rect 9036 12854 9088 12860
rect 9140 12782 9168 13398
rect 9232 12832 9260 14214
rect 9324 13938 9352 14350
rect 9404 14340 9456 14346
rect 9404 14282 9456 14288
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9232 12804 9352 12832
rect 9128 12776 9180 12782
rect 9128 12718 9180 12724
rect 8852 12708 8904 12714
rect 8852 12650 8904 12656
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 9140 12170 9168 12718
rect 9220 12708 9272 12714
rect 9220 12650 9272 12656
rect 9232 12442 9260 12650
rect 9220 12436 9272 12442
rect 9220 12378 9272 12384
rect 9128 12164 9180 12170
rect 8680 12124 8800 12152
rect 8588 12056 8708 12084
rect 8404 11886 8616 11914
rect 8390 11792 8446 11801
rect 8390 11727 8392 11736
rect 8444 11727 8446 11736
rect 8392 11698 8444 11704
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8392 9988 8444 9994
rect 8392 9930 8444 9936
rect 8404 9761 8432 9930
rect 8390 9752 8446 9761
rect 8390 9687 8446 9696
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 8300 9444 8352 9450
rect 8300 9386 8352 9392
rect 8312 8566 8340 9386
rect 8404 9217 8432 9590
rect 8390 9208 8446 9217
rect 8390 9143 8446 9152
rect 8404 9042 8432 9143
rect 8496 9110 8524 10950
rect 8588 10742 8616 11886
rect 8680 11830 8708 12056
rect 8772 11830 8800 12124
rect 9128 12106 9180 12112
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8864 11898 8892 12038
rect 8852 11892 8904 11898
rect 8852 11834 8904 11840
rect 8668 11824 8720 11830
rect 8668 11766 8720 11772
rect 8760 11824 8812 11830
rect 8760 11766 8812 11772
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 11540 9076 11698
rect 9140 11694 9168 12106
rect 9128 11688 9180 11694
rect 9128 11630 9180 11636
rect 9048 11512 9168 11540
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8576 10736 8628 10742
rect 8576 10678 8628 10684
rect 8574 10432 8630 10441
rect 8574 10367 8630 10376
rect 8588 9926 8616 10367
rect 8576 9920 8628 9926
rect 8576 9862 8628 9868
rect 8680 9489 8708 11290
rect 9140 11082 9168 11512
rect 9220 11144 9272 11150
rect 9218 11112 9220 11121
rect 9272 11112 9274 11121
rect 9128 11076 9180 11082
rect 9218 11047 9274 11056
rect 9128 11018 9180 11024
rect 9324 11014 9352 12804
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9220 10600 9272 10606
rect 9220 10542 9272 10548
rect 9128 10464 9180 10470
rect 9128 10406 9180 10412
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 9140 10266 9168 10406
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 8852 10192 8904 10198
rect 8852 10134 8904 10140
rect 8864 9586 8892 10134
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 8944 9920 8996 9926
rect 8996 9880 9076 9908
rect 8944 9862 8996 9868
rect 9048 9625 9076 9880
rect 9034 9616 9090 9625
rect 8852 9580 8904 9586
rect 9034 9551 9090 9560
rect 8852 9522 8904 9528
rect 8666 9480 8722 9489
rect 8666 9415 8722 9424
rect 9140 9382 9168 9930
rect 8668 9376 8720 9382
rect 8574 9344 8630 9353
rect 8668 9318 8720 9324
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 8574 9279 8630 9288
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8588 8945 8616 9279
rect 8680 9110 8708 9318
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 9036 8968 9088 8974
rect 8390 8936 8446 8945
rect 8574 8936 8630 8945
rect 8446 8894 8524 8922
rect 8390 8871 8446 8880
rect 8392 8832 8444 8838
rect 8496 8820 8524 8894
rect 9036 8910 9088 8916
rect 8574 8871 8630 8880
rect 8668 8832 8720 8838
rect 8496 8792 8668 8820
rect 8392 8774 8444 8780
rect 8668 8774 8720 8780
rect 8300 8560 8352 8566
rect 8300 8502 8352 8508
rect 8300 8356 8352 8362
rect 8300 8298 8352 8304
rect 8312 7954 8340 8298
rect 8300 7948 8352 7954
rect 8300 7890 8352 7896
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7002 8340 7686
rect 8404 7546 8432 8774
rect 8484 8424 8536 8430
rect 8484 8366 8536 8372
rect 8496 7546 8524 8366
rect 9048 8294 9076 8910
rect 9140 8430 9168 9318
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 9048 8266 9168 8294
rect 8574 8256 8630 8265
rect 8574 8191 8630 8200
rect 8588 8022 8616 8191
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8588 7750 8616 7958
rect 8576 7744 8628 7750
rect 8576 7686 8628 7692
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8392 7404 8444 7410
rect 8392 7346 8444 7352
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8300 6996 8352 7002
rect 8300 6938 8352 6944
rect 8036 6866 8340 6882
rect 8036 6860 8352 6866
rect 8036 6854 8300 6860
rect 8300 6802 8352 6808
rect 8116 6792 8168 6798
rect 8022 6760 8078 6769
rect 8168 6752 8248 6780
rect 8116 6734 8168 6740
rect 8022 6695 8078 6704
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6202 7972 6598
rect 8036 6440 8064 6695
rect 8116 6452 8168 6458
rect 8036 6412 8116 6440
rect 8116 6394 8168 6400
rect 8128 6225 8156 6394
rect 8220 6322 8248 6752
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 8300 6248 8352 6254
rect 8114 6216 8170 6225
rect 7944 6186 8064 6202
rect 7944 6180 8076 6186
rect 7944 6174 8024 6180
rect 8300 6190 8352 6196
rect 8114 6151 8170 6160
rect 8208 6180 8260 6186
rect 8024 6122 8076 6128
rect 8208 6122 8260 6128
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7944 5914 7972 6054
rect 8128 5953 8156 6054
rect 8114 5944 8170 5953
rect 7932 5908 7984 5914
rect 8114 5879 8170 5888
rect 7932 5850 7984 5856
rect 8116 5704 8168 5710
rect 8114 5672 8116 5681
rect 8168 5672 8170 5681
rect 8220 5658 8248 6122
rect 8312 5778 8340 6190
rect 8404 5953 8432 7346
rect 8680 6984 8708 8026
rect 9036 7880 9088 7886
rect 9140 7868 9168 8266
rect 9088 7840 9168 7868
rect 9036 7822 9088 7828
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 8747 7100 9055 7120
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 8680 6956 8800 6984
rect 8668 6860 8720 6866
rect 8668 6802 8720 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8390 5944 8446 5953
rect 8390 5879 8446 5888
rect 8496 5778 8524 6734
rect 8300 5772 8352 5778
rect 8300 5714 8352 5720
rect 8484 5772 8536 5778
rect 8484 5714 8536 5720
rect 8220 5630 8524 5658
rect 8114 5607 8170 5616
rect 8300 5568 8352 5574
rect 7852 5506 7972 5534
rect 7944 5250 7972 5506
rect 8266 5516 8300 5534
rect 8266 5510 8352 5516
rect 8266 5506 8340 5510
rect 8266 5386 8294 5506
rect 8128 5370 8294 5386
rect 8116 5364 8294 5370
rect 8168 5358 8294 5364
rect 8116 5306 8168 5312
rect 7656 5228 7708 5234
rect 7944 5222 8156 5250
rect 7656 5170 7708 5176
rect 7932 5160 7984 5166
rect 7932 5102 7984 5108
rect 7840 5024 7892 5030
rect 7746 4992 7802 5001
rect 7944 5001 7972 5102
rect 7840 4966 7892 4972
rect 7930 4992 7986 5001
rect 7746 4927 7802 4936
rect 7656 4480 7708 4486
rect 7654 4448 7656 4457
rect 7708 4448 7710 4457
rect 7654 4383 7710 4392
rect 7760 4321 7788 4927
rect 7746 4312 7802 4321
rect 7746 4247 7802 4256
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7668 3058 7696 3703
rect 7748 3460 7800 3466
rect 7748 3402 7800 3408
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7760 2854 7788 3402
rect 7852 3194 7880 4966
rect 7930 4927 7986 4936
rect 8022 4856 8078 4865
rect 8022 4791 8078 4800
rect 7932 4616 7984 4622
rect 7932 4558 7984 4564
rect 7944 3670 7972 4558
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7944 3058 7972 3606
rect 8036 3097 8064 4791
rect 8022 3088 8078 3097
rect 7932 3052 7984 3058
rect 8022 3023 8078 3032
rect 7932 2994 7984 3000
rect 8024 2984 8076 2990
rect 8024 2926 8076 2932
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7838 2816 7894 2825
rect 7838 2751 7894 2760
rect 7654 2680 7710 2689
rect 7654 2615 7710 2624
rect 7668 2582 7696 2615
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7656 2576 7708 2582
rect 7656 2518 7708 2524
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7484 1193 7512 2246
rect 7470 1184 7526 1193
rect 7470 1119 7526 1128
rect 7852 1018 7880 2751
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 7944 1465 7972 2382
rect 8036 2292 8064 2926
rect 8128 2514 8156 5222
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8208 5092 8260 5098
rect 8208 5034 8260 5040
rect 8220 4690 8248 5034
rect 8312 4865 8340 5170
rect 8496 5114 8524 5630
rect 8680 5574 8708 6802
rect 8772 6769 8800 6956
rect 8942 6896 8998 6905
rect 8942 6831 8998 6840
rect 8758 6760 8814 6769
rect 8758 6695 8814 6704
rect 8956 6458 8984 6831
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8747 6012 9055 6032
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 9140 5846 9168 7346
rect 9232 6798 9260 10542
rect 9324 9178 9352 10950
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9324 8838 9352 9114
rect 9312 8832 9364 8838
rect 9416 8809 9444 14282
rect 9508 14278 9536 14470
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9496 14272 9548 14278
rect 9496 14214 9548 14220
rect 9496 13932 9548 13938
rect 9496 13874 9548 13880
rect 9508 13258 9536 13874
rect 9600 13870 9628 14418
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9692 13705 9720 15671
rect 9772 15642 9824 15648
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 15360 9824 15366
rect 9876 15337 9904 15438
rect 9772 15302 9824 15308
rect 9862 15328 9918 15337
rect 9784 14804 9812 15302
rect 9862 15263 9918 15272
rect 9876 14958 9904 15263
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9784 14776 9904 14804
rect 9678 13696 9734 13705
rect 9678 13631 9734 13640
rect 9678 13560 9734 13569
rect 9678 13495 9734 13504
rect 9692 13394 9720 13495
rect 9680 13388 9732 13394
rect 9680 13330 9732 13336
rect 9496 13252 9548 13258
rect 9496 13194 9548 13200
rect 9508 9897 9536 13194
rect 9692 12481 9720 13330
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9784 12782 9812 12922
rect 9772 12776 9824 12782
rect 9876 12753 9904 14776
rect 9968 13326 9996 17274
rect 10336 17134 10364 17478
rect 10520 17338 10548 17478
rect 10508 17332 10560 17338
rect 10508 17274 10560 17280
rect 10048 17128 10100 17134
rect 10048 17070 10100 17076
rect 10324 17128 10376 17134
rect 10324 17070 10376 17076
rect 10506 17096 10562 17105
rect 10060 16522 10088 17070
rect 10506 17031 10562 17040
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10048 16516 10100 16522
rect 10048 16458 10100 16464
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10060 15162 10088 15302
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 10046 15056 10102 15065
rect 10046 14991 10102 15000
rect 10060 14958 10088 14991
rect 10048 14952 10100 14958
rect 10048 14894 10100 14900
rect 10152 14521 10180 16934
rect 10520 16590 10548 17031
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10336 16250 10364 16458
rect 10612 16250 10640 18380
rect 10704 18057 10732 18566
rect 10690 18048 10746 18057
rect 10690 17983 10746 17992
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10704 17649 10732 17818
rect 10690 17640 10746 17649
rect 10690 17575 10746 17584
rect 10692 17536 10744 17542
rect 10692 17478 10744 17484
rect 10704 17377 10732 17478
rect 10690 17368 10746 17377
rect 10796 17338 10824 19382
rect 10876 19372 10928 19378
rect 10980 19360 11008 19502
rect 11060 19508 11112 19514
rect 11060 19450 11112 19456
rect 11164 19446 11192 19615
rect 11256 19514 11284 19722
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 11716 19514 11744 19858
rect 11888 19780 11940 19786
rect 11992 19768 12020 20023
rect 11940 19740 12020 19768
rect 11888 19722 11940 19728
rect 12084 19700 12112 20454
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12624 20324 12676 20330
rect 12624 20266 12676 20272
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 12268 19972 12296 20198
rect 12438 20088 12494 20097
rect 12438 20023 12440 20032
rect 12492 20023 12494 20032
rect 12440 19994 12492 20000
rect 12348 19984 12400 19990
rect 12268 19944 12348 19972
rect 12348 19926 12400 19932
rect 12452 19854 12480 19994
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12348 19780 12400 19786
rect 12348 19722 12400 19728
rect 11992 19672 12112 19700
rect 12164 19712 12216 19718
rect 11244 19508 11296 19514
rect 11244 19450 11296 19456
rect 11704 19508 11756 19514
rect 11704 19450 11756 19456
rect 11152 19440 11204 19446
rect 11152 19382 11204 19388
rect 11888 19440 11940 19446
rect 11888 19382 11940 19388
rect 10980 19332 11100 19360
rect 10876 19314 10928 19320
rect 10888 18426 10916 19314
rect 10966 19136 11022 19145
rect 10966 19071 11022 19080
rect 10980 18698 11008 19071
rect 10968 18692 11020 18698
rect 10968 18634 11020 18640
rect 11072 18601 11100 19332
rect 11520 19304 11572 19310
rect 11520 19246 11572 19252
rect 11150 19000 11206 19009
rect 11150 18935 11206 18944
rect 11058 18592 11114 18601
rect 11058 18527 11114 18536
rect 11164 18465 11192 18935
rect 11532 18748 11560 19246
rect 11612 18760 11664 18766
rect 11532 18720 11612 18748
rect 11664 18720 11744 18748
rect 11612 18702 11664 18708
rect 11244 18624 11296 18630
rect 11244 18566 11296 18572
rect 11150 18456 11206 18465
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 10968 18420 11020 18426
rect 11020 18380 11100 18408
rect 11150 18391 11206 18400
rect 10968 18362 11020 18368
rect 11072 18340 11100 18380
rect 11256 18340 11284 18566
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 11072 18312 11284 18340
rect 11428 18352 11480 18358
rect 11428 18294 11480 18300
rect 11060 18216 11112 18222
rect 11112 18176 11192 18204
rect 11060 18158 11112 18164
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 10874 17776 10930 17785
rect 10874 17711 10876 17720
rect 10928 17711 10930 17720
rect 10876 17682 10928 17688
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10690 17303 10746 17312
rect 10784 17332 10836 17338
rect 10784 17274 10836 17280
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 10704 16998 10732 17138
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10888 16794 10916 17546
rect 10980 17202 11008 18022
rect 11072 17746 11100 18022
rect 11060 17740 11112 17746
rect 11060 17682 11112 17688
rect 11164 17354 11192 18176
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 11256 17678 11284 18090
rect 11440 18057 11468 18294
rect 11426 18048 11482 18057
rect 11426 17983 11482 17992
rect 11716 17814 11744 18720
rect 11794 18048 11850 18057
rect 11794 17983 11850 17992
rect 11704 17808 11756 17814
rect 11704 17750 11756 17756
rect 11244 17672 11296 17678
rect 11244 17614 11296 17620
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11440 17524 11468 17614
rect 11256 17496 11468 17524
rect 11256 17354 11284 17496
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11072 17326 11284 17354
rect 10968 17196 11020 17202
rect 10968 17138 11020 17144
rect 10876 16788 10928 16794
rect 10876 16730 10928 16736
rect 10782 16552 10838 16561
rect 10782 16487 10784 16496
rect 10836 16487 10838 16496
rect 10784 16458 10836 16464
rect 10692 16448 10744 16454
rect 10692 16390 10744 16396
rect 10324 16244 10376 16250
rect 10324 16186 10376 16192
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10232 15904 10284 15910
rect 10232 15846 10284 15852
rect 10138 14512 10194 14521
rect 10138 14447 10194 14456
rect 10048 14272 10100 14278
rect 10048 14214 10100 14220
rect 10060 14074 10088 14214
rect 10048 14068 10100 14074
rect 10048 14010 10100 14016
rect 10152 13954 10180 14447
rect 10060 13926 10180 13954
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9772 12718 9824 12724
rect 9862 12744 9918 12753
rect 9784 12628 9812 12718
rect 9862 12679 9918 12688
rect 9784 12600 9904 12628
rect 9678 12472 9734 12481
rect 9678 12407 9734 12416
rect 9678 12336 9734 12345
rect 9678 12271 9734 12280
rect 9692 11937 9720 12271
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9678 11928 9734 11937
rect 9678 11863 9734 11872
rect 9680 10600 9732 10606
rect 9680 10542 9732 10548
rect 9586 10296 9642 10305
rect 9586 10231 9642 10240
rect 9600 9926 9628 10231
rect 9692 10062 9720 10542
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9588 9920 9640 9926
rect 9494 9888 9550 9897
rect 9588 9862 9640 9868
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9494 9823 9550 9832
rect 9600 9761 9628 9862
rect 9586 9752 9642 9761
rect 9496 9716 9548 9722
rect 9586 9687 9642 9696
rect 9496 9658 9548 9664
rect 9508 9217 9536 9658
rect 9494 9208 9550 9217
rect 9494 9143 9550 9152
rect 9588 8900 9640 8906
rect 9588 8842 9640 8848
rect 9312 8774 9364 8780
rect 9402 8800 9458 8809
rect 9402 8735 9458 8744
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9312 8424 9364 8430
rect 9312 8366 9364 8372
rect 9324 8090 9352 8366
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9310 7984 9366 7993
rect 9310 7919 9366 7928
rect 9324 7750 9352 7919
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 9324 7206 9352 7414
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 9324 7041 9352 7142
rect 9310 7032 9366 7041
rect 9416 7002 9444 8434
rect 9508 7750 9536 8502
rect 9600 8401 9628 8842
rect 9586 8392 9642 8401
rect 9586 8327 9642 8336
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9600 7342 9628 7754
rect 9692 7721 9720 9862
rect 9678 7712 9734 7721
rect 9678 7647 9734 7656
rect 9588 7336 9640 7342
rect 9508 7296 9588 7324
rect 9310 6967 9366 6976
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9310 6896 9366 6905
rect 9310 6831 9366 6840
rect 9324 6798 9352 6831
rect 9220 6792 9272 6798
rect 9220 6734 9272 6740
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9220 6656 9272 6662
rect 9312 6656 9364 6662
rect 9220 6598 9272 6604
rect 9310 6624 9312 6633
rect 9364 6624 9366 6633
rect 9128 5840 9180 5846
rect 9128 5782 9180 5788
rect 8852 5704 8904 5710
rect 8850 5672 8852 5681
rect 8904 5672 8906 5681
rect 8850 5607 8906 5616
rect 9034 5672 9090 5681
rect 9034 5607 9090 5616
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 9048 5386 9076 5607
rect 8956 5358 9076 5386
rect 8496 5086 8616 5114
rect 8484 5024 8536 5030
rect 8390 4992 8446 5001
rect 8484 4966 8536 4972
rect 8390 4927 8446 4936
rect 8298 4856 8354 4865
rect 8298 4791 8354 4800
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8220 3466 8248 4626
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8312 3602 8340 4422
rect 8404 4078 8432 4927
rect 8496 4758 8524 4966
rect 8484 4752 8536 4758
rect 8484 4694 8536 4700
rect 8588 4554 8616 5086
rect 8956 5012 8984 5358
rect 9036 5228 9088 5234
rect 9140 5216 9168 5782
rect 9088 5188 9168 5216
rect 9036 5170 9088 5176
rect 8956 4984 9168 5012
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 8850 4584 8906 4593
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8760 4548 8812 4554
rect 8850 4519 8906 4528
rect 8760 4490 8812 4496
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8496 4282 8524 4422
rect 8484 4276 8536 4282
rect 8484 4218 8536 4224
rect 8772 4162 8800 4490
rect 8484 4140 8536 4146
rect 8484 4082 8536 4088
rect 8680 4134 8800 4162
rect 8864 4146 8892 4519
rect 8852 4140 8904 4146
rect 8392 4072 8444 4078
rect 8392 4014 8444 4020
rect 8300 3596 8352 3602
rect 8300 3538 8352 3544
rect 8208 3460 8260 3466
rect 8208 3402 8260 3408
rect 8220 3194 8248 3402
rect 8208 3188 8260 3194
rect 8208 3130 8260 3136
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 8208 2304 8260 2310
rect 8036 2264 8156 2292
rect 7930 1456 7986 1465
rect 7930 1391 7986 1400
rect 7840 1012 7892 1018
rect 7840 954 7892 960
rect 7576 870 7696 898
rect 7576 762 7604 870
rect 7668 800 7696 870
rect 8128 800 8156 2264
rect 8208 2246 8260 2252
rect 8220 2038 8248 2246
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8312 1970 8340 3062
rect 8496 2854 8524 4082
rect 8576 4072 8628 4078
rect 8576 4014 8628 4020
rect 8588 3738 8616 4014
rect 8576 3732 8628 3738
rect 8576 3674 8628 3680
rect 8574 3224 8630 3233
rect 8574 3159 8630 3168
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8588 2553 8616 3159
rect 8574 2544 8630 2553
rect 8574 2479 8630 2488
rect 8576 2304 8628 2310
rect 8576 2246 8628 2252
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8588 1601 8616 2246
rect 8574 1592 8630 1601
rect 8574 1527 8630 1536
rect 8680 1442 8708 4134
rect 8852 4082 8904 4088
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 9140 3584 9168 4984
rect 9048 3556 9168 3584
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8956 3194 8984 3470
rect 9048 3194 9076 3556
rect 9128 3460 9180 3466
rect 9128 3402 9180 3408
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 9140 3058 9168 3402
rect 9128 3052 9180 3058
rect 9128 2994 9180 3000
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 9126 2680 9182 2689
rect 9126 2615 9128 2624
rect 9180 2615 9182 2624
rect 9128 2586 9180 2592
rect 8758 2544 8814 2553
rect 8758 2479 8814 2488
rect 9126 2544 9182 2553
rect 9126 2479 9182 2488
rect 8772 2446 8800 2479
rect 8760 2440 8812 2446
rect 8760 2382 8812 2388
rect 8942 1728 8998 1737
rect 8942 1663 8998 1672
rect 8496 1414 8708 1442
rect 8496 800 8524 1414
rect 8956 800 8984 1663
rect 7392 734 7604 762
rect 7654 0 7710 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8942 0 8998 800
rect 9140 762 9168 2479
rect 9232 2038 9260 6598
rect 9310 6559 9366 6568
rect 9312 6384 9364 6390
rect 9312 6326 9364 6332
rect 9324 5574 9352 6326
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9310 5400 9366 5409
rect 9310 5335 9366 5344
rect 9324 4758 9352 5335
rect 9416 5030 9444 6938
rect 9508 6866 9536 7296
rect 9588 7278 9640 7284
rect 9496 6860 9548 6866
rect 9496 6802 9548 6808
rect 9784 6746 9812 12174
rect 9876 11354 9904 12600
rect 9968 12102 9996 13126
rect 10060 12986 10088 13926
rect 10140 13796 10192 13802
rect 10140 13738 10192 13744
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10152 12918 10180 13738
rect 10140 12912 10192 12918
rect 10140 12854 10192 12860
rect 10048 12640 10100 12646
rect 10046 12608 10048 12617
rect 10100 12608 10102 12617
rect 10046 12543 10102 12552
rect 10046 12200 10102 12209
rect 10046 12135 10102 12144
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 10060 11830 10088 12135
rect 10048 11824 10100 11830
rect 9968 11784 10048 11812
rect 9864 11348 9916 11354
rect 9864 11290 9916 11296
rect 9968 11286 9996 11784
rect 10048 11766 10100 11772
rect 10244 11694 10272 15846
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10324 15360 10376 15366
rect 10324 15302 10376 15308
rect 10336 14074 10364 15302
rect 10416 15156 10468 15162
rect 10416 15098 10468 15104
rect 10428 15065 10456 15098
rect 10414 15056 10470 15065
rect 10414 14991 10470 15000
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10416 13864 10468 13870
rect 10520 13852 10548 15438
rect 10598 15328 10654 15337
rect 10598 15263 10654 15272
rect 10612 15162 10640 15263
rect 10600 15156 10652 15162
rect 10600 15098 10652 15104
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10612 14482 10640 14758
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10704 13954 10732 16390
rect 10796 15910 10824 16458
rect 10888 16046 10916 16730
rect 10968 16108 11020 16114
rect 10968 16050 11020 16056
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10784 15904 10836 15910
rect 10980 15881 11008 16050
rect 10784 15846 10836 15852
rect 10966 15872 11022 15881
rect 10966 15807 11022 15816
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14006 10824 14758
rect 10888 14618 10916 15302
rect 11072 15094 11100 17326
rect 11244 17060 11296 17066
rect 11244 17002 11296 17008
rect 11256 16969 11284 17002
rect 11242 16960 11298 16969
rect 11242 16895 11298 16904
rect 11518 16824 11574 16833
rect 11518 16759 11574 16768
rect 11532 16658 11560 16759
rect 11716 16658 11744 17750
rect 11808 17592 11836 17983
rect 11900 17882 11928 19382
rect 11992 18465 12020 19672
rect 12164 19654 12216 19660
rect 12176 19378 12204 19654
rect 12256 19440 12308 19446
rect 12256 19382 12308 19388
rect 12164 19372 12216 19378
rect 12164 19314 12216 19320
rect 12268 19174 12296 19382
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12360 18601 12388 19722
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12452 19174 12480 19450
rect 12530 19408 12586 19417
rect 12530 19343 12586 19352
rect 12544 19310 12572 19343
rect 12636 19334 12664 20266
rect 12820 20058 12848 20402
rect 12808 20052 12860 20058
rect 12808 19994 12860 20000
rect 12532 19304 12584 19310
rect 12636 19306 12756 19334
rect 12532 19246 12584 19252
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12624 19168 12676 19174
rect 12624 19110 12676 19116
rect 12636 18884 12664 19110
rect 12544 18856 12664 18884
rect 12544 18766 12572 18856
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12728 18680 12756 19306
rect 12808 18828 12860 18834
rect 12808 18770 12860 18776
rect 12636 18652 12756 18680
rect 12440 18624 12492 18630
rect 12346 18592 12402 18601
rect 12440 18566 12492 18572
rect 12346 18527 12402 18536
rect 11978 18456 12034 18465
rect 12452 18426 12480 18566
rect 11978 18391 12034 18400
rect 12440 18420 12492 18426
rect 12440 18362 12492 18368
rect 12532 18352 12584 18358
rect 12530 18320 12532 18329
rect 12584 18320 12586 18329
rect 12530 18255 12586 18264
rect 11980 18216 12032 18222
rect 11980 18158 12032 18164
rect 11992 18086 12020 18158
rect 12348 18148 12400 18154
rect 12348 18090 12400 18096
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11808 17564 11928 17592
rect 11794 17504 11850 17513
rect 11794 17439 11850 17448
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11520 16652 11572 16658
rect 11520 16594 11572 16600
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11164 15201 11192 16594
rect 11244 16584 11296 16590
rect 11244 16526 11296 16532
rect 11256 16250 11284 16526
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11336 16108 11388 16114
rect 11336 16050 11388 16056
rect 11348 15910 11376 16050
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 11704 15904 11756 15910
rect 11704 15846 11756 15852
rect 11716 15609 11744 15846
rect 11702 15600 11758 15609
rect 11702 15535 11758 15544
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11150 15192 11206 15201
rect 11346 15184 11654 15204
rect 11150 15127 11206 15136
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10980 14822 11008 14962
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10876 14612 10928 14618
rect 10876 14554 10928 14560
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 14074 10916 14214
rect 10876 14068 10928 14074
rect 10876 14010 10928 14016
rect 10468 13824 10548 13852
rect 10612 13926 10732 13954
rect 10784 14000 10836 14006
rect 10784 13942 10836 13948
rect 10416 13806 10468 13812
rect 10428 13297 10456 13806
rect 10414 13288 10470 13297
rect 10414 13223 10470 13232
rect 10324 13184 10376 13190
rect 10376 13144 10456 13172
rect 10324 13126 10376 13132
rect 10324 12436 10376 12442
rect 10324 12378 10376 12384
rect 10336 11898 10364 12378
rect 10428 12306 10456 13144
rect 10508 12640 10560 12646
rect 10508 12582 10560 12588
rect 10416 12300 10468 12306
rect 10416 12242 10468 12248
rect 10324 11892 10376 11898
rect 10324 11834 10376 11840
rect 10232 11688 10284 11694
rect 10046 11656 10102 11665
rect 10232 11630 10284 11636
rect 10046 11591 10102 11600
rect 9956 11280 10008 11286
rect 9956 11222 10008 11228
rect 9968 11082 9996 11222
rect 10060 11218 10088 11591
rect 10140 11552 10192 11558
rect 10140 11494 10192 11500
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 9956 11076 10008 11082
rect 9956 11018 10008 11024
rect 9954 10840 10010 10849
rect 9954 10775 10010 10784
rect 9864 10532 9916 10538
rect 9864 10474 9916 10480
rect 9876 10062 9904 10474
rect 9864 10056 9916 10062
rect 9864 9998 9916 10004
rect 9968 9654 9996 10775
rect 10152 10282 10180 11494
rect 10230 11112 10286 11121
rect 10230 11047 10286 11056
rect 10244 10810 10272 11047
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10336 10742 10364 11834
rect 10428 11762 10456 12242
rect 10520 12238 10548 12582
rect 10508 12232 10560 12238
rect 10508 12174 10560 12180
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10520 11642 10548 12038
rect 10428 11614 10548 11642
rect 10324 10736 10376 10742
rect 10324 10678 10376 10684
rect 10230 10568 10286 10577
rect 10230 10503 10286 10512
rect 10060 10254 10180 10282
rect 10060 10169 10088 10254
rect 10046 10160 10102 10169
rect 10046 10095 10102 10104
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10048 9920 10100 9926
rect 10048 9862 10100 9868
rect 9956 9648 10008 9654
rect 9956 9590 10008 9596
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9876 7818 9904 9386
rect 9968 8673 9996 9590
rect 9954 8664 10010 8673
rect 9954 8599 9956 8608
rect 10008 8599 10010 8608
rect 9956 8570 10008 8576
rect 10060 8514 10088 9862
rect 10152 9586 10180 10066
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10152 9042 10180 9522
rect 10140 9036 10192 9042
rect 10140 8978 10192 8984
rect 9968 8486 10088 8514
rect 9864 7812 9916 7818
rect 9864 7754 9916 7760
rect 9862 7032 9918 7041
rect 9862 6967 9918 6976
rect 9508 6718 9812 6746
rect 9404 5024 9456 5030
rect 9404 4966 9456 4972
rect 9312 4752 9364 4758
rect 9312 4694 9364 4700
rect 9508 4554 9536 6718
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9586 6488 9642 6497
rect 9784 6458 9812 6598
rect 9586 6423 9588 6432
rect 9640 6423 9642 6432
rect 9772 6452 9824 6458
rect 9588 6394 9640 6400
rect 9772 6394 9824 6400
rect 9680 6248 9732 6254
rect 9680 6190 9732 6196
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 9496 4548 9548 4554
rect 9496 4490 9548 4496
rect 9312 4480 9364 4486
rect 9312 4422 9364 4428
rect 9324 3602 9352 4422
rect 9494 4312 9550 4321
rect 9494 4247 9496 4256
rect 9548 4247 9550 4256
rect 9496 4218 9548 4224
rect 9600 4060 9628 6054
rect 9692 4826 9720 6190
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9784 5302 9812 6122
rect 9876 5681 9904 6967
rect 9968 6322 9996 8486
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10060 7313 10088 8366
rect 10152 8362 10180 8978
rect 10140 8356 10192 8362
rect 10140 8298 10192 8304
rect 10152 8090 10180 8298
rect 10140 8084 10192 8090
rect 10140 8026 10192 8032
rect 10140 7812 10192 7818
rect 10140 7754 10192 7760
rect 10046 7304 10102 7313
rect 10046 7239 10102 7248
rect 10060 6882 10088 7239
rect 10152 7206 10180 7754
rect 10244 7546 10272 10503
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 8906 10364 10406
rect 10428 9722 10456 11614
rect 10612 11286 10640 13926
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10600 11280 10652 11286
rect 10600 11222 10652 11228
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10612 10674 10640 10950
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10520 10266 10548 10610
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10416 9716 10468 9722
rect 10416 9658 10468 9664
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 9382 10456 9454
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10520 9042 10548 10202
rect 10600 10192 10652 10198
rect 10600 10134 10652 10140
rect 10612 9722 10640 10134
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10600 9512 10652 9518
rect 10600 9454 10652 9460
rect 10612 9178 10640 9454
rect 10600 9172 10652 9178
rect 10600 9114 10652 9120
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10704 8922 10732 13806
rect 10980 13569 11008 14758
rect 11072 14074 11100 15030
rect 11164 14521 11192 15127
rect 11426 15056 11482 15065
rect 11426 14991 11482 15000
rect 11440 14822 11468 14991
rect 11520 14952 11572 14958
rect 11520 14894 11572 14900
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11150 14512 11206 14521
rect 11150 14447 11206 14456
rect 11440 14414 11468 14758
rect 11532 14550 11560 14894
rect 11808 14618 11836 17439
rect 11900 16454 11928 17564
rect 11888 16448 11940 16454
rect 11888 16390 11940 16396
rect 11888 15904 11940 15910
rect 11888 15846 11940 15852
rect 11900 15473 11928 15846
rect 11886 15464 11942 15473
rect 11886 15399 11942 15408
rect 11992 14793 12020 18022
rect 12254 17776 12310 17785
rect 12360 17762 12388 18090
rect 12438 17912 12494 17921
rect 12438 17847 12494 17856
rect 12310 17734 12388 17762
rect 12254 17711 12310 17720
rect 12348 17604 12400 17610
rect 12348 17546 12400 17552
rect 12164 17536 12216 17542
rect 12164 17478 12216 17484
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 12084 16998 12112 17206
rect 12072 16992 12124 16998
rect 12072 16934 12124 16940
rect 12176 16574 12204 17478
rect 12360 17338 12388 17546
rect 12452 17338 12480 17847
rect 12532 17536 12584 17542
rect 12532 17478 12584 17484
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12348 16992 12400 16998
rect 12348 16934 12400 16940
rect 12084 16546 12204 16574
rect 11978 14784 12034 14793
rect 11978 14719 12034 14728
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11164 13954 11192 14350
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 11888 14272 11940 14278
rect 12084 14249 12112 16546
rect 12162 16280 12218 16289
rect 12162 16215 12218 16224
rect 12176 16182 12204 16215
rect 12164 16176 12216 16182
rect 12164 16118 12216 16124
rect 12164 15904 12216 15910
rect 12164 15846 12216 15852
rect 12176 15502 12204 15846
rect 12268 15570 12296 16934
rect 12360 16794 12388 16934
rect 12544 16810 12572 17478
rect 12452 16794 12572 16810
rect 12348 16788 12400 16794
rect 12348 16730 12400 16736
rect 12440 16788 12572 16794
rect 12492 16782 12572 16788
rect 12440 16730 12492 16736
rect 12636 16640 12664 18652
rect 12714 18592 12770 18601
rect 12714 18527 12770 18536
rect 12728 18426 12756 18527
rect 12716 18420 12768 18426
rect 12716 18362 12768 18368
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 12544 16612 12664 16640
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12348 16176 12400 16182
rect 12348 16118 12400 16124
rect 12360 15706 12388 16118
rect 12348 15700 12400 15706
rect 12348 15642 12400 15648
rect 12452 15638 12480 16458
rect 12440 15632 12492 15638
rect 12440 15574 12492 15580
rect 12256 15564 12308 15570
rect 12256 15506 12308 15512
rect 12164 15496 12216 15502
rect 12164 15438 12216 15444
rect 12452 14822 12480 15574
rect 12440 14816 12492 14822
rect 12440 14758 12492 14764
rect 12164 14612 12216 14618
rect 12348 14612 12400 14618
rect 12216 14572 12296 14600
rect 12164 14554 12216 14560
rect 11888 14214 11940 14220
rect 12070 14240 12126 14249
rect 11072 13926 11192 13954
rect 10966 13560 11022 13569
rect 10966 13495 11022 13504
rect 10876 13252 10928 13258
rect 10876 13194 10928 13200
rect 10888 12782 10916 13194
rect 11072 13190 11100 13926
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 10966 13016 11022 13025
rect 10966 12951 10968 12960
rect 11020 12951 11022 12960
rect 10968 12922 11020 12928
rect 10876 12776 10928 12782
rect 10876 12718 10928 12724
rect 11164 12288 11192 13806
rect 11256 12986 11284 14214
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11716 14074 11744 14214
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 11796 14068 11848 14074
rect 11796 14010 11848 14016
rect 11610 13968 11666 13977
rect 11336 13932 11388 13938
rect 11808 13938 11836 14010
rect 11610 13903 11666 13912
rect 11796 13932 11848 13938
rect 11336 13874 11388 13880
rect 11348 13530 11376 13874
rect 11624 13870 11652 13903
rect 11796 13874 11848 13880
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11520 13728 11572 13734
rect 11520 13670 11572 13676
rect 11532 13530 11560 13670
rect 11336 13524 11388 13530
rect 11336 13466 11388 13472
rect 11520 13524 11572 13530
rect 11520 13466 11572 13472
rect 11612 13388 11664 13394
rect 11612 13330 11664 13336
rect 11624 13240 11652 13330
rect 11624 13212 11744 13240
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11244 12980 11296 12986
rect 11716 12968 11744 13212
rect 11244 12922 11296 12928
rect 11624 12940 11744 12968
rect 11244 12708 11296 12714
rect 11244 12650 11296 12656
rect 11072 12260 11192 12288
rect 10968 12232 11020 12238
rect 10888 12192 10968 12220
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 10796 10266 10824 11222
rect 10888 10588 10916 12192
rect 10968 12174 11020 12180
rect 10966 11248 11022 11257
rect 10966 11183 11022 11192
rect 10980 11150 11008 11183
rect 10968 11144 11020 11150
rect 10968 11086 11020 11092
rect 10968 10600 11020 10606
rect 10888 10560 10968 10588
rect 10968 10542 11020 10548
rect 10784 10260 10836 10266
rect 10784 10202 10836 10208
rect 10796 9926 10824 10202
rect 10876 9988 10928 9994
rect 10980 9976 11008 10542
rect 11072 10010 11100 12260
rect 11152 12164 11204 12170
rect 11152 12106 11204 12112
rect 11164 11626 11192 12106
rect 11256 12102 11284 12650
rect 11624 12170 11652 12940
rect 11716 12782 11744 12813
rect 11704 12776 11756 12782
rect 11808 12730 11836 13738
rect 11756 12724 11836 12730
rect 11704 12718 11836 12724
rect 11716 12702 11836 12718
rect 11716 12442 11744 12702
rect 11796 12640 11848 12646
rect 11796 12582 11848 12588
rect 11704 12436 11756 12442
rect 11704 12378 11756 12384
rect 11808 12306 11836 12582
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11900 12238 11928 14214
rect 12070 14175 12126 14184
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11992 13258 12020 14010
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 12084 12434 12112 13942
rect 12162 13696 12218 13705
rect 12162 13631 12218 13640
rect 12176 13025 12204 13631
rect 12268 13410 12296 14572
rect 12348 14554 12400 14560
rect 12360 14362 12388 14554
rect 12452 14482 12480 14758
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12360 14334 12480 14362
rect 12346 14104 12402 14113
rect 12346 14039 12402 14048
rect 12360 13841 12388 14039
rect 12346 13832 12402 13841
rect 12346 13767 12402 13776
rect 12268 13382 12388 13410
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12162 13016 12218 13025
rect 12162 12951 12218 12960
rect 12164 12776 12216 12782
rect 12164 12718 12216 12724
rect 12176 12442 12204 12718
rect 11992 12406 12112 12434
rect 12164 12436 12216 12442
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11612 12164 11664 12170
rect 11612 12106 11664 12112
rect 11244 12096 11296 12102
rect 11244 12038 11296 12044
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11704 11688 11756 11694
rect 11704 11630 11756 11636
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11218 11192 11562
rect 11716 11354 11744 11630
rect 11244 11348 11296 11354
rect 11244 11290 11296 11296
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11164 10810 11192 11154
rect 11256 11014 11284 11290
rect 11900 11218 11928 11698
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 11796 11076 11848 11082
rect 11796 11018 11848 11024
rect 11888 11076 11940 11082
rect 11888 11018 11940 11024
rect 11244 11008 11296 11014
rect 11808 10985 11836 11018
rect 11244 10950 11296 10956
rect 11794 10976 11850 10985
rect 11346 10908 11654 10928
rect 11794 10911 11850 10920
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11900 10810 11928 11018
rect 11152 10804 11204 10810
rect 11152 10746 11204 10752
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11888 10532 11940 10538
rect 11888 10474 11940 10480
rect 11796 10192 11848 10198
rect 11702 10160 11758 10169
rect 11796 10134 11848 10140
rect 11702 10095 11758 10104
rect 11072 9982 11192 10010
rect 10928 9948 11008 9976
rect 10876 9930 10928 9936
rect 10784 9920 10836 9926
rect 11060 9920 11112 9926
rect 10784 9862 10836 9868
rect 11058 9888 11060 9897
rect 11112 9888 11114 9897
rect 11058 9823 11114 9832
rect 11164 9466 11192 9982
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11334 9616 11390 9625
rect 11334 9551 11390 9560
rect 10888 9438 11192 9466
rect 10784 9376 10836 9382
rect 10784 9318 10836 9324
rect 10796 8974 10824 9318
rect 10888 9178 10916 9438
rect 11152 9376 11204 9382
rect 11072 9336 11152 9364
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10520 8894 10732 8922
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10336 8537 10364 8842
rect 10416 8832 10468 8838
rect 10414 8800 10416 8809
rect 10468 8800 10470 8809
rect 10414 8735 10470 8744
rect 10322 8528 10378 8537
rect 10322 8463 10378 8472
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10324 8356 10376 8362
rect 10324 8298 10376 8304
rect 10336 7993 10364 8298
rect 10322 7984 10378 7993
rect 10322 7919 10378 7928
rect 10428 7868 10456 8434
rect 10336 7840 10456 7868
rect 10336 7721 10364 7840
rect 10416 7744 10468 7750
rect 10322 7712 10378 7721
rect 10416 7686 10468 7692
rect 10322 7647 10378 7656
rect 10322 7576 10378 7585
rect 10232 7540 10284 7546
rect 10322 7511 10378 7520
rect 10232 7482 10284 7488
rect 10232 7336 10284 7342
rect 10336 7313 10364 7511
rect 10232 7278 10284 7284
rect 10322 7304 10378 7313
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10060 6854 10180 6882
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9956 6316 10008 6322
rect 9956 6258 10008 6264
rect 9862 5672 9918 5681
rect 9862 5607 9918 5616
rect 9956 5636 10008 5642
rect 9956 5578 10008 5584
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 9772 5296 9824 5302
rect 9772 5238 9824 5244
rect 9772 5024 9824 5030
rect 9772 4966 9824 4972
rect 9680 4820 9732 4826
rect 9680 4762 9732 4768
rect 9784 4486 9812 4966
rect 9876 4554 9904 5510
rect 9968 4690 9996 5578
rect 10060 4690 10088 6734
rect 10152 6662 10180 6854
rect 10244 6798 10272 7278
rect 10322 7239 10378 7248
rect 10322 6896 10378 6905
rect 10322 6831 10378 6840
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10140 6656 10192 6662
rect 10140 6598 10192 6604
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 10152 5001 10180 6258
rect 10336 5930 10364 6831
rect 10244 5902 10364 5930
rect 10244 5234 10272 5902
rect 10324 5840 10376 5846
rect 10324 5782 10376 5788
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10138 4992 10194 5001
rect 10138 4927 10194 4936
rect 9956 4684 10008 4690
rect 9956 4626 10008 4632
rect 10048 4684 10100 4690
rect 10048 4626 10100 4632
rect 9864 4548 9916 4554
rect 9864 4490 9916 4496
rect 9772 4480 9824 4486
rect 9772 4422 9824 4428
rect 9956 4276 10008 4282
rect 9956 4218 10008 4224
rect 9772 4072 9824 4078
rect 9600 4032 9772 4060
rect 9494 3904 9550 3913
rect 9494 3839 9550 3848
rect 9312 3596 9364 3602
rect 9312 3538 9364 3544
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9404 3392 9456 3398
rect 9508 3369 9536 3839
rect 9600 3448 9628 4032
rect 9772 4014 9824 4020
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9680 3460 9732 3466
rect 9600 3420 9680 3448
rect 9680 3402 9732 3408
rect 9404 3334 9456 3340
rect 9494 3360 9550 3369
rect 9324 2582 9352 3334
rect 9312 2576 9364 2582
rect 9312 2518 9364 2524
rect 9416 2428 9444 3334
rect 9494 3295 9550 3304
rect 9692 3194 9720 3402
rect 9772 3392 9824 3398
rect 9772 3334 9824 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9508 2774 9536 3130
rect 9784 3126 9812 3334
rect 9772 3120 9824 3126
rect 9772 3062 9824 3068
rect 9678 2952 9734 2961
rect 9678 2887 9734 2896
rect 9508 2746 9628 2774
rect 9324 2400 9444 2428
rect 9496 2440 9548 2446
rect 9324 2310 9352 2400
rect 9496 2382 9548 2388
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9508 2258 9536 2382
rect 9600 2378 9628 2746
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 9692 2258 9720 2887
rect 9784 2514 9812 3062
rect 9876 2922 9904 3674
rect 9968 3466 9996 4218
rect 10152 3754 10180 4927
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10244 4554 10272 4626
rect 10232 4548 10284 4554
rect 10232 4490 10284 4496
rect 10232 4140 10284 4146
rect 10232 4082 10284 4088
rect 10060 3726 10180 3754
rect 9956 3460 10008 3466
rect 9956 3402 10008 3408
rect 9968 3194 9996 3402
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 9508 2230 9720 2258
rect 9772 2304 9824 2310
rect 9772 2246 9824 2252
rect 9220 2032 9272 2038
rect 9220 1974 9272 1980
rect 9784 1698 9812 2246
rect 9772 1692 9824 1698
rect 9772 1634 9824 1640
rect 9876 1170 9904 2858
rect 10060 2854 10088 3726
rect 10140 3664 10192 3670
rect 10140 3606 10192 3612
rect 10152 3194 10180 3606
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10244 3074 10272 4082
rect 10152 3046 10272 3074
rect 10152 2854 10180 3046
rect 10230 2952 10286 2961
rect 10230 2887 10286 2896
rect 10048 2848 10100 2854
rect 10048 2790 10100 2796
rect 10140 2848 10192 2854
rect 10140 2790 10192 2796
rect 9784 1142 9904 1170
rect 9324 870 9444 898
rect 9324 762 9352 870
rect 9416 800 9444 870
rect 9784 800 9812 1142
rect 10244 800 10272 2887
rect 10336 1358 10364 5782
rect 10428 5574 10456 7686
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10414 4856 10470 4865
rect 10414 4791 10470 4800
rect 10428 4146 10456 4791
rect 10416 4140 10468 4146
rect 10416 4082 10468 4088
rect 10416 4004 10468 4010
rect 10416 3946 10468 3952
rect 10428 3641 10456 3946
rect 10520 3738 10548 8894
rect 10692 8832 10744 8838
rect 10888 8786 10916 9114
rect 10692 8774 10744 8780
rect 10704 8634 10732 8774
rect 10796 8758 10916 8786
rect 10968 8832 11020 8838
rect 10968 8774 11020 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10600 8560 10652 8566
rect 10600 8502 10652 8508
rect 10690 8528 10746 8537
rect 10612 7478 10640 8502
rect 10690 8463 10746 8472
rect 10704 8294 10732 8463
rect 10692 8288 10744 8294
rect 10692 8230 10744 8236
rect 10796 8090 10824 8758
rect 10874 8664 10930 8673
rect 10874 8599 10876 8608
rect 10928 8599 10930 8608
rect 10876 8570 10928 8576
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10888 8090 10916 8298
rect 10784 8084 10836 8090
rect 10784 8026 10836 8032
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10692 7812 10744 7818
rect 10692 7754 10744 7760
rect 10600 7472 10652 7478
rect 10600 7414 10652 7420
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 6934 10640 7142
rect 10600 6928 10652 6934
rect 10600 6870 10652 6876
rect 10704 6186 10732 7754
rect 10796 7154 10824 8026
rect 10876 7744 10928 7750
rect 10876 7686 10928 7692
rect 10888 7274 10916 7686
rect 10876 7268 10928 7274
rect 10876 7210 10928 7216
rect 10796 7126 10916 7154
rect 10888 6662 10916 7126
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10600 6180 10652 6186
rect 10600 6122 10652 6128
rect 10692 6180 10744 6186
rect 10692 6122 10744 6128
rect 10612 5914 10640 6122
rect 10600 5908 10652 5914
rect 10600 5850 10652 5856
rect 10600 5568 10652 5574
rect 10600 5510 10652 5516
rect 10612 4865 10640 5510
rect 10598 4856 10654 4865
rect 10598 4791 10654 4800
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10612 4214 10640 4422
rect 10600 4208 10652 4214
rect 10600 4150 10652 4156
rect 10508 3732 10560 3738
rect 10508 3674 10560 3680
rect 10414 3632 10470 3641
rect 10414 3567 10470 3576
rect 10428 2009 10456 3567
rect 10704 2802 10732 6122
rect 10796 5914 10824 6258
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10888 5302 10916 6054
rect 10876 5296 10928 5302
rect 10876 5238 10928 5244
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10888 4282 10916 4762
rect 10980 4622 11008 8774
rect 11072 8362 11100 9336
rect 11152 9318 11204 9324
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11164 8566 11192 8978
rect 11348 8945 11376 9551
rect 11716 9432 11744 10095
rect 11808 9926 11836 10134
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11532 9404 11744 9432
rect 11532 8974 11560 9404
rect 11610 9344 11666 9353
rect 11610 9279 11666 9288
rect 11624 9110 11652 9279
rect 11702 9208 11758 9217
rect 11702 9143 11758 9152
rect 11796 9172 11848 9178
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11520 8968 11572 8974
rect 11334 8936 11390 8945
rect 11716 8945 11744 9143
rect 11796 9114 11848 9120
rect 11520 8910 11572 8916
rect 11702 8936 11758 8945
rect 11334 8871 11390 8880
rect 11808 8906 11836 9114
rect 11702 8871 11758 8880
rect 11796 8900 11848 8906
rect 11796 8842 11848 8848
rect 11244 8832 11296 8838
rect 11244 8774 11296 8780
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11247 8634 11275 8774
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8560 11204 8566
rect 11204 8508 11284 8514
rect 11152 8502 11284 8508
rect 11164 8486 11284 8502
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7936 11192 8298
rect 11072 7908 11192 7936
rect 11072 6866 11100 7908
rect 11256 7886 11284 8486
rect 11336 8288 11388 8294
rect 11336 8230 11388 8236
rect 11244 7880 11296 7886
rect 11348 7857 11376 8230
rect 11612 8084 11664 8090
rect 11440 8044 11612 8072
rect 11244 7822 11296 7828
rect 11334 7848 11390 7857
rect 11334 7783 11390 7792
rect 11440 7732 11468 8044
rect 11612 8026 11664 8032
rect 11256 7704 11468 7732
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11060 6112 11112 6118
rect 11060 6054 11112 6060
rect 11072 5370 11100 6054
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 11164 5148 11192 7142
rect 11256 6866 11284 7704
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11256 6390 11284 6666
rect 11716 6662 11744 8774
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11808 7426 11836 8230
rect 11900 7750 11928 10474
rect 11992 10266 12020 12406
rect 12164 12378 12216 12384
rect 12268 12374 12296 13126
rect 12360 12986 12388 13382
rect 12348 12980 12400 12986
rect 12348 12922 12400 12928
rect 12072 12368 12124 12374
rect 12072 12310 12124 12316
rect 12256 12368 12308 12374
rect 12256 12310 12308 12316
rect 12084 11762 12112 12310
rect 12164 12300 12216 12306
rect 12164 12242 12216 12248
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 12070 11384 12126 11393
rect 12070 11319 12126 11328
rect 12084 10810 12112 11319
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 12176 10470 12204 12242
rect 12254 12200 12310 12209
rect 12254 12135 12310 12144
rect 12268 11370 12296 12135
rect 12348 12096 12400 12102
rect 12348 12038 12400 12044
rect 12360 11898 12388 12038
rect 12348 11892 12400 11898
rect 12348 11834 12400 11840
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 12360 11626 12388 11698
rect 12348 11620 12400 11626
rect 12348 11562 12400 11568
rect 12268 11354 12388 11370
rect 12268 11348 12400 11354
rect 12268 11342 12348 11348
rect 12348 11290 12400 11296
rect 12256 11280 12308 11286
rect 12256 11222 12308 11228
rect 12072 10464 12124 10470
rect 12072 10406 12124 10412
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11992 9722 12020 10202
rect 11980 9716 12032 9722
rect 11980 9658 12032 9664
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11992 9024 12020 9114
rect 11983 8996 12020 9024
rect 11983 8820 12011 8996
rect 11983 8792 12020 8820
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11992 7546 12020 8792
rect 11980 7540 12032 7546
rect 11980 7482 12032 7488
rect 11808 7398 11928 7426
rect 11796 7336 11848 7342
rect 11796 7278 11848 7284
rect 11808 6662 11836 7278
rect 11704 6656 11756 6662
rect 11704 6598 11756 6604
rect 11796 6656 11848 6662
rect 11796 6598 11848 6604
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 11900 6474 11928 7398
rect 12084 7041 12112 10406
rect 12176 10169 12204 10406
rect 12162 10160 12218 10169
rect 12268 10130 12296 11222
rect 12452 10996 12480 14334
rect 12544 14006 12572 16612
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12636 16250 12664 16458
rect 12624 16244 12676 16250
rect 12624 16186 12676 16192
rect 12728 16046 12756 17138
rect 12820 16454 12848 18770
rect 12912 18426 12940 21354
rect 13084 21072 13136 21078
rect 13084 21014 13136 21020
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 13004 18902 13032 20810
rect 12992 18896 13044 18902
rect 12992 18838 13044 18844
rect 12900 18420 12952 18426
rect 12900 18362 12952 18368
rect 13096 17921 13124 21014
rect 13188 20602 13216 22200
rect 13268 21208 13320 21214
rect 13268 21150 13320 21156
rect 13176 20596 13228 20602
rect 13176 20538 13228 20544
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13188 20058 13216 20402
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 13176 19848 13228 19854
rect 13176 19790 13228 19796
rect 13188 19514 13216 19790
rect 13176 19508 13228 19514
rect 13176 19450 13228 19456
rect 13174 19136 13230 19145
rect 13174 19071 13230 19080
rect 13188 18834 13216 19071
rect 13176 18828 13228 18834
rect 13176 18770 13228 18776
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 13082 17912 13138 17921
rect 13082 17847 13138 17856
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 13004 17270 13032 17750
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 12992 17264 13044 17270
rect 12992 17206 13044 17212
rect 12992 16584 13044 16590
rect 12992 16526 13044 16532
rect 12808 16448 12860 16454
rect 12808 16390 12860 16396
rect 12820 16114 12848 16390
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12716 16040 12768 16046
rect 12716 15982 12768 15988
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 15162 12664 15302
rect 12624 15156 12676 15162
rect 12624 15098 12676 15104
rect 12728 15094 12756 15982
rect 13004 15348 13032 16526
rect 13096 16250 13124 17478
rect 13188 17202 13216 18566
rect 13280 18426 13308 21150
rect 13556 20602 13584 22200
rect 14016 20602 14044 22200
rect 14280 21684 14332 21690
rect 14280 21626 14332 21632
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 14004 20596 14056 20602
rect 14004 20538 14056 20544
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 20058 13492 20334
rect 13542 20224 13598 20233
rect 13542 20159 13598 20168
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13556 19938 13584 20159
rect 13740 20058 13768 20402
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 13728 20052 13780 20058
rect 13728 19994 13780 20000
rect 13360 19916 13412 19922
rect 13360 19858 13412 19864
rect 13464 19910 13584 19938
rect 13372 19174 13400 19858
rect 13464 19174 13492 19910
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13544 19236 13596 19242
rect 13544 19178 13596 19184
rect 13360 19168 13412 19174
rect 13360 19110 13412 19116
rect 13452 19168 13504 19174
rect 13452 19110 13504 19116
rect 13268 18420 13320 18426
rect 13268 18362 13320 18368
rect 13372 18034 13400 19110
rect 13464 18154 13492 19110
rect 13556 18426 13584 19178
rect 13544 18420 13596 18426
rect 13544 18362 13596 18368
rect 13544 18284 13596 18290
rect 13544 18226 13596 18232
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13372 18006 13492 18034
rect 13360 17876 13412 17882
rect 13360 17818 13412 17824
rect 13268 17536 13320 17542
rect 13268 17478 13320 17484
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13084 16244 13136 16250
rect 13084 16186 13136 16192
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13084 15972 13136 15978
rect 13084 15914 13136 15920
rect 12820 15320 13032 15348
rect 12716 15088 12768 15094
rect 12716 15030 12768 15036
rect 12714 14648 12770 14657
rect 12624 14612 12676 14618
rect 12714 14583 12770 14592
rect 12624 14554 12676 14560
rect 12636 14482 12664 14554
rect 12624 14476 12676 14482
rect 12624 14418 12676 14424
rect 12728 14249 12756 14583
rect 12714 14240 12770 14249
rect 12714 14175 12770 14184
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12624 13728 12676 13734
rect 12624 13670 12676 13676
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12544 12850 12572 13194
rect 12636 12889 12664 13670
rect 12622 12880 12678 12889
rect 12532 12844 12584 12850
rect 12622 12815 12678 12824
rect 12532 12786 12584 12792
rect 12530 12744 12586 12753
rect 12530 12679 12586 12688
rect 12544 12345 12572 12679
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12530 12336 12586 12345
rect 12530 12271 12586 12280
rect 12532 12232 12584 12238
rect 12530 12200 12532 12209
rect 12584 12200 12586 12209
rect 12530 12135 12586 12144
rect 12530 12064 12586 12073
rect 12530 11999 12586 12008
rect 12360 10968 12480 10996
rect 12162 10095 12218 10104
rect 12256 10124 12308 10130
rect 12256 10066 12308 10072
rect 12162 9888 12218 9897
rect 12162 9823 12218 9832
rect 12070 7032 12126 7041
rect 11980 6996 12032 7002
rect 12070 6967 12126 6976
rect 11980 6938 12032 6944
rect 11716 6446 11928 6474
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11428 6248 11480 6254
rect 11428 6190 11480 6196
rect 11336 6112 11388 6118
rect 11336 6054 11388 6060
rect 11348 5914 11376 6054
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11348 5817 11376 5850
rect 11334 5808 11390 5817
rect 11440 5778 11468 6190
rect 11334 5743 11390 5752
rect 11428 5772 11480 5778
rect 11428 5714 11480 5720
rect 11440 5642 11468 5714
rect 11428 5636 11480 5642
rect 11428 5578 11480 5584
rect 11716 5574 11744 6446
rect 11886 6352 11942 6361
rect 11886 6287 11888 6296
rect 11940 6287 11942 6296
rect 11888 6258 11940 6264
rect 11992 6254 12020 6938
rect 12070 6896 12126 6905
rect 12070 6831 12126 6840
rect 12084 6730 12112 6831
rect 12072 6724 12124 6730
rect 12072 6666 12124 6672
rect 12070 6624 12126 6633
rect 12070 6559 12126 6568
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11796 6180 11848 6186
rect 11796 6122 11848 6128
rect 11808 5681 11836 6122
rect 12084 6066 12112 6559
rect 12176 6186 12204 9823
rect 12268 9586 12296 10066
rect 12256 9580 12308 9586
rect 12256 9522 12308 9528
rect 12268 9382 12296 9522
rect 12256 9376 12308 9382
rect 12256 9318 12308 9324
rect 12268 8566 12296 9318
rect 12256 8560 12308 8566
rect 12256 8502 12308 8508
rect 12360 7834 12388 10968
rect 12544 10674 12572 11999
rect 12636 11082 12664 12582
rect 12728 11257 12756 13670
rect 12820 12889 12848 15320
rect 12990 15056 13046 15065
rect 12990 14991 13046 15000
rect 12900 14340 12952 14346
rect 12900 14282 12952 14288
rect 12806 12880 12862 12889
rect 12806 12815 12862 12824
rect 12806 11928 12862 11937
rect 12806 11863 12808 11872
rect 12860 11863 12862 11872
rect 12808 11834 12860 11840
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 11558 12848 11698
rect 12808 11552 12860 11558
rect 12806 11520 12808 11529
rect 12860 11520 12862 11529
rect 12806 11455 12862 11464
rect 12808 11348 12860 11354
rect 12808 11290 12860 11296
rect 12714 11248 12770 11257
rect 12714 11183 12770 11192
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12532 10668 12584 10674
rect 12532 10610 12584 10616
rect 12440 8968 12492 8974
rect 12438 8936 12440 8945
rect 12492 8936 12494 8945
rect 12438 8871 12494 8880
rect 12532 8832 12584 8838
rect 12532 8774 12584 8780
rect 12544 8673 12572 8774
rect 12530 8664 12586 8673
rect 12530 8599 12586 8608
rect 12636 8378 12664 11018
rect 12820 10606 12848 11290
rect 12808 10600 12860 10606
rect 12808 10542 12860 10548
rect 12716 9716 12768 9722
rect 12716 9658 12768 9664
rect 12544 8350 12664 8378
rect 12544 8294 12572 8350
rect 12532 8288 12584 8294
rect 12532 8230 12584 8236
rect 12624 8288 12676 8294
rect 12624 8230 12676 8236
rect 12728 8242 12756 9658
rect 12912 9178 12940 14282
rect 13004 14074 13032 14991
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12992 13864 13044 13870
rect 12990 13832 12992 13841
rect 13044 13832 13046 13841
rect 12990 13767 13046 13776
rect 13096 13462 13124 15914
rect 13188 15706 13216 16050
rect 13280 15745 13308 17478
rect 13372 17270 13400 17818
rect 13464 17660 13492 18006
rect 13556 17882 13584 18226
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13648 17785 13676 19314
rect 13728 19236 13780 19242
rect 13728 19178 13780 19184
rect 13740 19009 13768 19178
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13726 19000 13782 19009
rect 13832 18970 13860 19110
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 13726 18935 13782 18944
rect 13820 18964 13872 18970
rect 13820 18906 13872 18912
rect 13728 18896 13780 18902
rect 13728 18838 13780 18844
rect 13740 18057 13768 18838
rect 13818 18728 13874 18737
rect 13818 18663 13820 18672
rect 13872 18663 13874 18672
rect 13820 18634 13872 18640
rect 14292 18358 14320 21626
rect 14384 20602 14412 22200
rect 14554 21584 14610 21593
rect 14554 21519 14610 21528
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14464 20460 14516 20466
rect 14464 20402 14516 20408
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18873 14412 19110
rect 14476 18970 14504 20402
rect 14568 19904 14596 21519
rect 14752 20602 14780 22200
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14740 20596 14792 20602
rect 14740 20538 14792 20544
rect 14648 20460 14700 20466
rect 14648 20402 14700 20408
rect 14660 20058 14688 20402
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14568 19876 14688 19904
rect 14556 19780 14608 19786
rect 14556 19722 14608 19728
rect 14464 18964 14516 18970
rect 14464 18906 14516 18912
rect 14370 18864 14426 18873
rect 14568 18850 14596 19722
rect 14370 18799 14426 18808
rect 14476 18822 14596 18850
rect 14370 18728 14426 18737
rect 14370 18663 14426 18672
rect 14384 18358 14412 18663
rect 14280 18352 14332 18358
rect 14280 18294 14332 18300
rect 14372 18352 14424 18358
rect 14372 18294 14424 18300
rect 14280 18080 14332 18086
rect 13726 18048 13782 18057
rect 14280 18022 14332 18028
rect 13726 17983 13782 17992
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 13820 17808 13872 17814
rect 13634 17776 13690 17785
rect 13634 17711 13690 17720
rect 13818 17776 13820 17785
rect 13872 17776 13874 17785
rect 13818 17711 13874 17720
rect 13728 17672 13780 17678
rect 13464 17632 13676 17660
rect 13360 17264 13412 17270
rect 13360 17206 13412 17212
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13464 16674 13492 17138
rect 13542 16960 13598 16969
rect 13542 16895 13598 16904
rect 13556 16794 13584 16895
rect 13544 16788 13596 16794
rect 13544 16730 13596 16736
rect 13464 16658 13584 16674
rect 13464 16652 13596 16658
rect 13464 16646 13544 16652
rect 13544 16594 13596 16600
rect 13556 16046 13584 16594
rect 13648 16590 13676 17632
rect 13728 17614 13780 17620
rect 13740 17202 13768 17614
rect 13820 17604 13872 17610
rect 13820 17546 13872 17552
rect 13728 17196 13780 17202
rect 13728 17138 13780 17144
rect 13636 16584 13688 16590
rect 13636 16526 13688 16532
rect 13728 16448 13780 16454
rect 13728 16390 13780 16396
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13452 16040 13504 16046
rect 13452 15982 13504 15988
rect 13544 16040 13596 16046
rect 13544 15982 13596 15988
rect 13266 15736 13322 15745
rect 13176 15700 13228 15706
rect 13266 15671 13322 15680
rect 13176 15642 13228 15648
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 15162 13400 15302
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14952 13320 14958
rect 13268 14894 13320 14900
rect 13176 13864 13228 13870
rect 13176 13806 13228 13812
rect 13084 13456 13136 13462
rect 13188 13433 13216 13806
rect 13084 13398 13136 13404
rect 13174 13424 13230 13433
rect 13174 13359 13230 13368
rect 13280 13308 13308 14894
rect 13372 14822 13400 14962
rect 13360 14816 13412 14822
rect 13360 14758 13412 14764
rect 13464 14618 13492 15982
rect 13648 15638 13676 16050
rect 13636 15632 13688 15638
rect 13636 15574 13688 15580
rect 13740 15194 13768 16390
rect 13832 16250 13860 17546
rect 14292 17513 14320 18022
rect 14278 17504 14334 17513
rect 14278 17439 14334 17448
rect 14280 17060 14332 17066
rect 14280 17002 14332 17008
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 14292 16658 14320 17002
rect 14280 16652 14332 16658
rect 14280 16594 14332 16600
rect 13912 16448 13964 16454
rect 13912 16390 13964 16396
rect 14372 16448 14424 16454
rect 14372 16390 14424 16396
rect 13924 16250 13952 16390
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13912 16244 13964 16250
rect 13912 16186 13964 16192
rect 13924 15892 13952 16186
rect 14384 16182 14412 16390
rect 14372 16176 14424 16182
rect 14372 16118 14424 16124
rect 13832 15864 13952 15892
rect 13832 15201 13860 15864
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 14384 15502 14412 16118
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14280 15428 14332 15434
rect 14280 15370 14332 15376
rect 13648 15166 13768 15194
rect 13818 15192 13874 15201
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13360 14544 13412 14550
rect 13360 14486 13412 14492
rect 13372 14278 13400 14486
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13464 14006 13492 14350
rect 13544 14272 13596 14278
rect 13544 14214 13596 14220
rect 13452 14000 13504 14006
rect 13452 13942 13504 13948
rect 13360 13456 13412 13462
rect 13360 13398 13412 13404
rect 13450 13424 13506 13433
rect 13188 13280 13308 13308
rect 12992 13184 13044 13190
rect 12992 13126 13044 13132
rect 13084 13184 13136 13190
rect 13084 13126 13136 13132
rect 13004 12918 13032 13126
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12992 12368 13044 12374
rect 12990 12336 12992 12345
rect 13044 12336 13046 12345
rect 12990 12271 13046 12280
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13004 11150 13032 12174
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 12992 10736 13044 10742
rect 13096 10713 13124 13126
rect 13188 12628 13216 13280
rect 13372 13258 13400 13398
rect 13450 13359 13506 13368
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 13280 12753 13308 12922
rect 13266 12744 13322 12753
rect 13266 12679 13322 12688
rect 13188 12600 13308 12628
rect 13280 12345 13308 12600
rect 13266 12336 13322 12345
rect 13266 12271 13322 12280
rect 13174 11520 13230 11529
rect 13174 11455 13230 11464
rect 13188 11354 13216 11455
rect 13176 11348 13228 11354
rect 13176 11290 13228 11296
rect 12992 10678 13044 10684
rect 13082 10704 13138 10713
rect 13004 9761 13032 10678
rect 13280 10674 13308 12271
rect 13372 11370 13400 13194
rect 13464 12617 13492 13359
rect 13556 12850 13584 14214
rect 13544 12844 13596 12850
rect 13544 12786 13596 12792
rect 13450 12608 13506 12617
rect 13450 12543 13506 12552
rect 13648 12374 13676 15166
rect 13818 15127 13874 15136
rect 13728 14816 13780 14822
rect 13728 14758 13780 14764
rect 13740 13190 13768 14758
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 14004 14544 14056 14550
rect 14004 14486 14056 14492
rect 14016 13938 14044 14486
rect 14292 14482 14320 15370
rect 14476 14958 14504 18822
rect 14556 18760 14608 18766
rect 14556 18702 14608 18708
rect 14568 18426 14596 18702
rect 14660 18426 14688 19876
rect 14832 19848 14884 19854
rect 14832 19790 14884 19796
rect 14740 19304 14792 19310
rect 14738 19272 14740 19281
rect 14792 19272 14794 19281
rect 14738 19207 14794 19216
rect 14738 19136 14794 19145
rect 14738 19071 14794 19080
rect 14556 18420 14608 18426
rect 14556 18362 14608 18368
rect 14648 18420 14700 18426
rect 14648 18362 14700 18368
rect 14752 18358 14780 19071
rect 14740 18352 14792 18358
rect 14740 18294 14792 18300
rect 14556 18216 14608 18222
rect 14556 18158 14608 18164
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14464 14816 14516 14822
rect 14462 14784 14464 14793
rect 14516 14784 14518 14793
rect 14462 14719 14518 14728
rect 14280 14476 14332 14482
rect 14280 14418 14332 14424
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13818 13560 13874 13569
rect 13945 13552 14253 13572
rect 14370 13560 14426 13569
rect 13818 13495 13874 13504
rect 14370 13495 14426 13504
rect 13832 13462 13860 13495
rect 14384 13462 14412 13495
rect 13820 13456 13872 13462
rect 13820 13398 13872 13404
rect 14372 13456 14424 13462
rect 14372 13398 14424 13404
rect 13818 13288 13874 13297
rect 13818 13223 13820 13232
rect 13872 13223 13874 13232
rect 13820 13194 13872 13200
rect 13728 13184 13780 13190
rect 13728 13126 13780 13132
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13740 12306 13768 12786
rect 14280 12708 14332 12714
rect 14280 12650 14332 12656
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13544 12096 13596 12102
rect 13544 12038 13596 12044
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 13556 11762 13584 12038
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13452 11688 13504 11694
rect 13450 11656 13452 11665
rect 14108 11665 14136 12038
rect 13504 11656 13506 11665
rect 14094 11656 14150 11665
rect 13450 11591 13506 11600
rect 13636 11620 13688 11626
rect 14094 11591 14150 11600
rect 13636 11562 13688 11568
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13372 11342 13492 11370
rect 13556 11354 13584 11494
rect 13360 11280 13412 11286
rect 13360 11222 13412 11228
rect 13082 10639 13138 10648
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13268 10464 13320 10470
rect 13268 10406 13320 10412
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 12990 9752 13046 9761
rect 12990 9687 13046 9696
rect 13188 9518 13216 9862
rect 13280 9586 13308 10406
rect 13372 10130 13400 11222
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13176 9512 13228 9518
rect 13464 9466 13492 11342
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13544 11212 13596 11218
rect 13544 11154 13596 11160
rect 13556 10742 13584 11154
rect 13648 10996 13676 11562
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13818 11520 13874 11529
rect 13740 11150 13768 11494
rect 13818 11455 13874 11464
rect 13832 11218 13860 11455
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13912 11212 13964 11218
rect 13912 11154 13964 11160
rect 13728 11144 13780 11150
rect 13924 11098 13952 11154
rect 13728 11086 13780 11092
rect 13832 11070 13952 11098
rect 13832 10996 13860 11070
rect 13648 10968 13860 10996
rect 13912 11008 13964 11014
rect 13740 10742 13768 10968
rect 13912 10950 13964 10956
rect 13544 10736 13596 10742
rect 13728 10736 13780 10742
rect 13544 10678 13596 10684
rect 13634 10704 13690 10713
rect 13556 10441 13584 10678
rect 13728 10678 13780 10684
rect 13634 10639 13690 10648
rect 13542 10432 13598 10441
rect 13542 10367 13598 10376
rect 13556 10062 13584 10367
rect 13648 10266 13676 10639
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 13740 10130 13768 10678
rect 13924 10606 13952 10950
rect 13912 10600 13964 10606
rect 13912 10542 13964 10548
rect 14004 10600 14056 10606
rect 14004 10542 14056 10548
rect 14016 10452 14044 10542
rect 13832 10441 14044 10452
rect 13818 10432 14044 10441
rect 13874 10424 14044 10432
rect 13818 10367 13874 10376
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 13820 10192 13872 10198
rect 13820 10134 13872 10140
rect 14188 10192 14240 10198
rect 14188 10134 14240 10140
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 13648 9704 13676 10066
rect 13556 9676 13676 9704
rect 13556 9586 13584 9676
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 13636 9580 13688 9586
rect 13636 9522 13688 9528
rect 13176 9454 13228 9460
rect 12992 9444 13044 9450
rect 12992 9386 13044 9392
rect 13280 9438 13492 9466
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 13004 9110 13032 9386
rect 13082 9208 13138 9217
rect 13082 9143 13138 9152
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12820 8634 12848 8978
rect 13096 8838 13124 9143
rect 13176 8968 13228 8974
rect 13176 8910 13228 8916
rect 13084 8832 13136 8838
rect 13084 8774 13136 8780
rect 12898 8664 12954 8673
rect 12808 8628 12860 8634
rect 12898 8599 12954 8608
rect 12808 8570 12860 8576
rect 12438 8120 12494 8129
rect 12438 8055 12440 8064
rect 12492 8055 12494 8064
rect 12440 8026 12492 8032
rect 12532 7948 12584 7954
rect 12532 7890 12584 7896
rect 12256 7812 12308 7818
rect 12360 7806 12480 7834
rect 12256 7754 12308 7760
rect 12268 7546 12296 7754
rect 12348 7744 12400 7750
rect 12348 7686 12400 7692
rect 12256 7540 12308 7546
rect 12256 7482 12308 7488
rect 12360 7342 12388 7686
rect 12348 7336 12400 7342
rect 12268 7296 12348 7324
rect 12268 6905 12296 7296
rect 12348 7278 12400 7284
rect 12452 7154 12480 7806
rect 12544 7342 12572 7890
rect 12636 7818 12664 8230
rect 12728 8214 12848 8242
rect 12820 8090 12848 8214
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12808 8084 12860 8090
rect 12808 8026 12860 8032
rect 12624 7812 12676 7818
rect 12624 7754 12676 7760
rect 12728 7546 12756 8026
rect 12806 7984 12862 7993
rect 12806 7919 12862 7928
rect 12820 7886 12848 7919
rect 12808 7880 12860 7886
rect 12808 7822 12860 7828
rect 12820 7585 12848 7822
rect 12806 7576 12862 7585
rect 12716 7540 12768 7546
rect 12806 7511 12862 7520
rect 12716 7482 12768 7488
rect 12912 7410 12940 8599
rect 13096 7993 13124 8774
rect 13188 8294 13216 8910
rect 13280 8362 13308 9438
rect 13360 9376 13412 9382
rect 13360 9318 13412 9324
rect 13268 8356 13320 8362
rect 13268 8298 13320 8304
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13082 7984 13138 7993
rect 13082 7919 13138 7928
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13096 7546 13124 7754
rect 13188 7546 13216 7754
rect 13084 7540 13136 7546
rect 13084 7482 13136 7488
rect 13176 7540 13228 7546
rect 13176 7482 13228 7488
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12532 7336 12584 7342
rect 12532 7278 12584 7284
rect 12716 7268 12768 7274
rect 12716 7210 12768 7216
rect 12360 7126 12480 7154
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12254 6896 12310 6905
rect 12254 6831 12310 6840
rect 12360 6746 12388 7126
rect 12544 6914 12572 7142
rect 12544 6886 12664 6914
rect 12440 6792 12492 6798
rect 12268 6718 12388 6746
rect 12438 6760 12440 6769
rect 12492 6760 12494 6769
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12084 6038 12204 6066
rect 11794 5672 11850 5681
rect 11794 5607 11850 5616
rect 11978 5672 12034 5681
rect 11978 5607 11980 5616
rect 12032 5607 12034 5616
rect 11980 5578 12032 5584
rect 11244 5568 11296 5574
rect 11244 5510 11296 5516
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11072 5120 11192 5148
rect 11072 4826 11100 5120
rect 11060 4820 11112 4826
rect 11060 4762 11112 4768
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 11256 4486 11284 5510
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 11794 5400 11850 5409
rect 11794 5335 11850 5344
rect 11888 5364 11940 5370
rect 11336 5296 11388 5302
rect 11336 5238 11388 5244
rect 11428 5296 11480 5302
rect 11808 5284 11836 5335
rect 11940 5324 12020 5352
rect 11888 5306 11940 5312
rect 11428 5238 11480 5244
rect 11692 5256 11836 5284
rect 11348 4593 11376 5238
rect 11440 4826 11468 5238
rect 11692 5148 11720 5256
rect 11888 5228 11940 5234
rect 11888 5170 11940 5176
rect 11692 5120 11836 5148
rect 11610 4856 11666 4865
rect 11428 4820 11480 4826
rect 11610 4791 11666 4800
rect 11428 4762 11480 4768
rect 11624 4690 11652 4791
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11704 4684 11756 4690
rect 11704 4626 11756 4632
rect 11334 4584 11390 4593
rect 11624 4554 11652 4626
rect 11334 4519 11390 4528
rect 11612 4548 11664 4554
rect 11612 4490 11664 4496
rect 10968 4480 11020 4486
rect 11244 4480 11296 4486
rect 10968 4422 11020 4428
rect 11150 4448 11206 4457
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10784 4072 10836 4078
rect 10980 4060 11008 4422
rect 11206 4428 11244 4434
rect 11206 4422 11296 4428
rect 11206 4406 11284 4422
rect 11150 4383 11206 4392
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11150 4312 11206 4321
rect 11346 4304 11654 4324
rect 11150 4247 11206 4256
rect 11060 4140 11112 4146
rect 11164 4128 11192 4247
rect 11428 4140 11480 4146
rect 11164 4100 11428 4128
rect 11060 4082 11112 4088
rect 11428 4082 11480 4088
rect 10784 4014 10836 4020
rect 10888 4032 11008 4060
rect 10796 3942 10824 4014
rect 10784 3936 10836 3942
rect 10784 3878 10836 3884
rect 10784 3732 10836 3738
rect 10784 3674 10836 3680
rect 10796 3194 10824 3674
rect 10784 3188 10836 3194
rect 10784 3130 10836 3136
rect 10612 2774 10732 2802
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10414 2000 10470 2009
rect 10414 1935 10470 1944
rect 10520 1698 10548 2382
rect 10508 1692 10560 1698
rect 10508 1634 10560 1640
rect 10324 1352 10376 1358
rect 10324 1294 10376 1300
rect 10612 800 10640 2774
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10704 2446 10732 2518
rect 10796 2514 10824 3130
rect 10888 2514 10916 4032
rect 11072 3584 11100 4082
rect 11520 4072 11572 4078
rect 11164 4020 11520 4026
rect 11716 4026 11744 4626
rect 11164 4014 11572 4020
rect 11164 3998 11560 4014
rect 11624 3998 11744 4026
rect 11164 3942 11192 3998
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 11244 3936 11296 3942
rect 11244 3878 11296 3884
rect 10980 3556 11100 3584
rect 10980 3233 11008 3556
rect 11060 3460 11112 3466
rect 11060 3402 11112 3408
rect 10966 3224 11022 3233
rect 10966 3159 11022 3168
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10704 1834 10732 2382
rect 10888 1902 10916 2450
rect 10876 1896 10928 1902
rect 10876 1838 10928 1844
rect 10692 1828 10744 1834
rect 10692 1770 10744 1776
rect 11072 1766 11100 3402
rect 11150 3224 11206 3233
rect 11256 3194 11284 3878
rect 11624 3602 11652 3998
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3596 11664 3602
rect 11612 3538 11664 3544
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 11150 3159 11206 3168
rect 11244 3188 11296 3194
rect 11164 2446 11192 3159
rect 11244 3130 11296 3136
rect 11336 3120 11388 3126
rect 11716 3108 11744 3878
rect 11808 3670 11836 5120
rect 11900 4826 11928 5170
rect 11888 4820 11940 4826
rect 11888 4762 11940 4768
rect 11796 3664 11848 3670
rect 11796 3606 11848 3612
rect 11900 3602 11928 4762
rect 11992 4690 12020 5324
rect 12176 5284 12204 6038
rect 12268 5370 12296 6718
rect 12438 6695 12494 6704
rect 12348 6656 12400 6662
rect 12348 6598 12400 6604
rect 12360 6390 12388 6598
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12636 5914 12664 6886
rect 12728 6361 12756 7210
rect 12992 7200 13044 7206
rect 12992 7142 13044 7148
rect 13004 7002 13032 7142
rect 12992 6996 13044 7002
rect 12898 6930 12954 6939
rect 12992 6938 13044 6944
rect 13096 6905 13124 7346
rect 13372 7342 13400 9318
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13452 8832 13504 8838
rect 13450 8800 13452 8809
rect 13504 8800 13506 8809
rect 13450 8735 13506 8744
rect 13556 8514 13584 9114
rect 13648 8906 13676 9522
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13728 8560 13780 8566
rect 13556 8486 13676 8514
rect 13728 8502 13780 8508
rect 13544 8424 13596 8430
rect 13544 8366 13596 8372
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13464 7585 13492 8298
rect 13556 7954 13584 8366
rect 13544 7948 13596 7954
rect 13648 7936 13676 8486
rect 13740 8090 13768 8502
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13648 7908 13768 7936
rect 13544 7890 13596 7896
rect 13634 7848 13690 7857
rect 13634 7783 13690 7792
rect 13544 7744 13596 7750
rect 13544 7686 13596 7692
rect 13450 7576 13506 7585
rect 13450 7511 13506 7520
rect 13360 7336 13412 7342
rect 13360 7278 13412 7284
rect 13176 7200 13228 7206
rect 13176 7142 13228 7148
rect 13360 7200 13412 7206
rect 13360 7142 13412 7148
rect 12898 6865 12954 6874
rect 13082 6896 13138 6905
rect 12714 6352 12770 6361
rect 12714 6287 12770 6296
rect 12624 5908 12676 5914
rect 12624 5850 12676 5856
rect 12912 5778 12940 6865
rect 13082 6831 13138 6840
rect 13188 6798 13216 7142
rect 13176 6792 13228 6798
rect 13176 6734 13228 6740
rect 13266 6624 13322 6633
rect 13266 6559 13322 6568
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12716 5772 12768 5778
rect 12716 5714 12768 5720
rect 12900 5772 12952 5778
rect 12900 5714 12952 5720
rect 12440 5636 12492 5642
rect 12360 5596 12440 5624
rect 12256 5364 12308 5370
rect 12256 5306 12308 5312
rect 12084 5256 12204 5284
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 12084 4604 12112 5256
rect 12162 5128 12218 5137
rect 12162 5063 12218 5072
rect 12176 4758 12204 5063
rect 12268 4865 12296 5306
rect 12254 4856 12310 4865
rect 12360 4826 12388 5596
rect 12440 5578 12492 5584
rect 12544 5302 12572 5714
rect 12622 5672 12678 5681
rect 12622 5607 12678 5616
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12440 5228 12492 5234
rect 12440 5170 12492 5176
rect 12452 5001 12480 5170
rect 12532 5024 12584 5030
rect 12438 4992 12494 5001
rect 12532 4966 12584 4972
rect 12438 4927 12494 4936
rect 12254 4791 12310 4800
rect 12348 4820 12400 4826
rect 12348 4762 12400 4768
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12164 4752 12216 4758
rect 12164 4694 12216 4700
rect 12348 4616 12400 4622
rect 12084 4576 12296 4604
rect 11980 4548 12032 4554
rect 11980 4490 12032 4496
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11900 3448 11928 3538
rect 11808 3420 11928 3448
rect 11808 3126 11836 3420
rect 11886 3360 11942 3369
rect 11886 3295 11942 3304
rect 11336 3062 11388 3068
rect 11624 3080 11744 3108
rect 11796 3120 11848 3126
rect 11348 2990 11376 3062
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11336 2984 11388 2990
rect 11336 2926 11388 2932
rect 11428 2848 11480 2854
rect 11532 2836 11560 2994
rect 11480 2808 11560 2836
rect 11428 2790 11480 2796
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 11072 800 11100 1702
rect 9140 734 9352 762
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10598 0 10654 800
rect 11058 0 11114 800
rect 11164 762 11192 2382
rect 11624 2292 11652 3080
rect 11796 3062 11848 3068
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 11704 2848 11756 2854
rect 11808 2825 11836 2926
rect 11704 2790 11756 2796
rect 11794 2816 11850 2825
rect 11716 2514 11744 2790
rect 11794 2751 11850 2760
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11900 2446 11928 3295
rect 11888 2440 11940 2446
rect 11888 2382 11940 2388
rect 11624 2264 11744 2292
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 11716 2106 11744 2264
rect 11704 2100 11756 2106
rect 11704 2042 11756 2048
rect 11888 1964 11940 1970
rect 11888 1906 11940 1912
rect 11348 870 11468 898
rect 11348 762 11376 870
rect 11440 800 11468 870
rect 11900 800 11928 1906
rect 11992 1698 12020 4490
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12164 4480 12216 4486
rect 12164 4422 12216 4428
rect 12084 4282 12112 4422
rect 12072 4276 12124 4282
rect 12072 4218 12124 4224
rect 12176 4146 12204 4422
rect 12268 4154 12296 4576
rect 12348 4558 12400 4564
rect 12360 4457 12388 4558
rect 12346 4448 12402 4457
rect 12346 4383 12402 4392
rect 12452 4282 12480 4762
rect 12544 4690 12572 4966
rect 12532 4684 12584 4690
rect 12532 4626 12584 4632
rect 12530 4584 12586 4593
rect 12530 4519 12586 4528
rect 12544 4486 12572 4519
rect 12532 4480 12584 4486
rect 12532 4422 12584 4428
rect 12440 4276 12492 4282
rect 12440 4218 12492 4224
rect 12164 4140 12216 4146
rect 12268 4126 12388 4154
rect 12164 4082 12216 4088
rect 12256 4072 12308 4078
rect 12254 4040 12256 4049
rect 12308 4040 12310 4049
rect 12254 3975 12310 3984
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 12162 3632 12218 3641
rect 12162 3567 12218 3576
rect 12070 3224 12126 3233
rect 12070 3159 12126 3168
rect 12084 2582 12112 3159
rect 12072 2576 12124 2582
rect 12072 2518 12124 2524
rect 12176 2310 12204 3567
rect 12164 2304 12216 2310
rect 12164 2246 12216 2252
rect 11980 1692 12032 1698
rect 11980 1634 12032 1640
rect 12268 800 12296 3674
rect 12360 3126 12388 4126
rect 12440 4140 12492 4146
rect 12440 4082 12492 4088
rect 12452 3466 12480 4082
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 12438 3360 12494 3369
rect 12438 3295 12494 3304
rect 12348 3120 12400 3126
rect 12348 3062 12400 3068
rect 12452 2854 12480 3295
rect 12440 2848 12492 2854
rect 12440 2790 12492 2796
rect 12544 2514 12572 4014
rect 12636 3641 12664 5607
rect 12728 5030 12756 5714
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12716 5024 12768 5030
rect 12716 4966 12768 4972
rect 12728 4672 12756 4966
rect 12820 4826 12848 5510
rect 12898 4856 12954 4865
rect 12808 4820 12860 4826
rect 12898 4791 12900 4800
rect 12808 4762 12860 4768
rect 12952 4791 12954 4800
rect 12900 4762 12952 4768
rect 12808 4684 12860 4690
rect 12728 4644 12808 4672
rect 12808 4626 12860 4632
rect 12900 4684 12952 4690
rect 12900 4626 12952 4632
rect 12714 4584 12770 4593
rect 12714 4519 12770 4528
rect 12622 3632 12678 3641
rect 12728 3618 12756 4519
rect 12820 4146 12848 4626
rect 12912 4214 12940 4626
rect 12900 4208 12952 4214
rect 12900 4150 12952 4156
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 13004 3777 13032 6326
rect 13174 5944 13230 5953
rect 13174 5879 13230 5888
rect 13188 5681 13216 5879
rect 13174 5672 13230 5681
rect 13174 5607 13230 5616
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13082 5264 13138 5273
rect 13082 5199 13138 5208
rect 12990 3768 13046 3777
rect 12990 3703 13046 3712
rect 13096 3641 13124 5199
rect 13188 4690 13216 5510
rect 13176 4684 13228 4690
rect 13176 4626 13228 4632
rect 13176 4480 13228 4486
rect 13176 4422 13228 4428
rect 13188 4282 13216 4422
rect 13176 4276 13228 4282
rect 13176 4218 13228 4224
rect 13082 3632 13138 3641
rect 12728 3590 12940 3618
rect 12622 3567 12678 3576
rect 12716 3528 12768 3534
rect 12716 3470 12768 3476
rect 12728 3058 12756 3470
rect 12716 3052 12768 3058
rect 12716 2994 12768 3000
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12452 2106 12480 2246
rect 12440 2100 12492 2106
rect 12440 2042 12492 2048
rect 12636 1970 12664 2926
rect 12912 2774 12940 3590
rect 13082 3567 13138 3576
rect 13280 2774 13308 6559
rect 13372 4162 13400 7142
rect 13464 6746 13492 7511
rect 13556 6866 13584 7686
rect 13648 7546 13676 7783
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13740 7426 13768 7908
rect 13832 7546 13860 10134
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 14016 9518 14044 9998
rect 14200 9926 14228 10134
rect 14188 9920 14240 9926
rect 14188 9862 14240 9868
rect 14004 9512 14056 9518
rect 14004 9454 14056 9460
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 14292 9081 14320 12650
rect 14464 12640 14516 12646
rect 14462 12608 14464 12617
rect 14516 12608 14518 12617
rect 14462 12543 14518 12552
rect 14370 12472 14426 12481
rect 14370 12407 14372 12416
rect 14424 12407 14426 12416
rect 14372 12378 14424 12384
rect 14372 12232 14424 12238
rect 14372 12174 14424 12180
rect 14384 11286 14412 12174
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14372 10668 14424 10674
rect 14372 10610 14424 10616
rect 14384 10266 14412 10610
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 14370 9208 14426 9217
rect 14370 9143 14372 9152
rect 14424 9143 14426 9152
rect 14372 9114 14424 9120
rect 14278 9072 14334 9081
rect 14188 9036 14240 9042
rect 14278 9007 14334 9016
rect 14188 8978 14240 8984
rect 14200 8673 14228 8978
rect 14476 8922 14504 12038
rect 14568 10198 14596 18158
rect 14648 17264 14700 17270
rect 14648 17206 14700 17212
rect 14660 16998 14688 17206
rect 14648 16992 14700 16998
rect 14648 16934 14700 16940
rect 14740 16448 14792 16454
rect 14740 16390 14792 16396
rect 14648 15904 14700 15910
rect 14648 15846 14700 15852
rect 14660 15706 14688 15846
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14660 15366 14688 15642
rect 14648 15360 14700 15366
rect 14752 15348 14780 16390
rect 14844 16182 14872 19790
rect 14936 18426 14964 20878
rect 15120 20584 15148 22200
rect 15382 20632 15438 20641
rect 15200 20596 15252 20602
rect 15120 20556 15200 20584
rect 15488 20602 15516 22200
rect 15660 21548 15712 21554
rect 15660 21490 15712 21496
rect 15382 20567 15438 20576
rect 15476 20596 15528 20602
rect 15200 20538 15252 20544
rect 15290 20496 15346 20505
rect 15016 20460 15068 20466
rect 15290 20431 15346 20440
rect 15016 20402 15068 20408
rect 15028 20058 15056 20402
rect 15016 20052 15068 20058
rect 15016 19994 15068 20000
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15212 19360 15240 19790
rect 15120 19332 15240 19360
rect 15120 19258 15148 19332
rect 15304 19310 15332 20431
rect 15396 19360 15424 20567
rect 15476 20538 15528 20544
rect 15568 20460 15620 20466
rect 15568 20402 15620 20408
rect 15396 19332 15516 19360
rect 15292 19304 15344 19310
rect 15028 19230 15148 19258
rect 15198 19272 15254 19281
rect 15028 19174 15056 19230
rect 15292 19246 15344 19252
rect 15382 19272 15438 19281
rect 15198 19207 15254 19216
rect 15382 19207 15438 19216
rect 15016 19168 15068 19174
rect 15016 19110 15068 19116
rect 14924 18420 14976 18426
rect 14924 18362 14976 18368
rect 15028 18086 15056 19110
rect 15212 18426 15240 19207
rect 15292 19168 15344 19174
rect 15292 19110 15344 19116
rect 15304 18902 15332 19110
rect 15292 18896 15344 18902
rect 15292 18838 15344 18844
rect 15290 18592 15346 18601
rect 15290 18527 15346 18536
rect 15304 18426 15332 18527
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15396 18358 15424 19207
rect 15384 18352 15436 18358
rect 15384 18294 15436 18300
rect 15016 18080 15068 18086
rect 15016 18022 15068 18028
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15016 17128 15068 17134
rect 15120 17082 15148 17478
rect 15200 17196 15252 17202
rect 15200 17138 15252 17144
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15068 17076 15148 17082
rect 15016 17070 15148 17076
rect 15028 17054 15148 17070
rect 14924 16992 14976 16998
rect 14924 16934 14976 16940
rect 14832 16176 14884 16182
rect 14832 16118 14884 16124
rect 14936 15502 14964 16934
rect 15120 16522 15148 17054
rect 15212 16522 15240 17138
rect 15292 17128 15344 17134
rect 15292 17070 15344 17076
rect 15108 16516 15160 16522
rect 15108 16458 15160 16464
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15120 16046 15148 16458
rect 15304 16250 15332 17070
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15570 15148 15982
rect 15396 15706 15424 17138
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 14924 15496 14976 15502
rect 14924 15438 14976 15444
rect 14832 15360 14884 15366
rect 14752 15320 14832 15348
rect 14648 15302 14700 15308
rect 14832 15302 14884 15308
rect 15200 15360 15252 15366
rect 15200 15302 15252 15308
rect 14660 13190 14688 15302
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14752 13870 14780 14894
rect 14844 14822 14872 15302
rect 15212 15094 15240 15302
rect 15200 15088 15252 15094
rect 15200 15030 15252 15036
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 15014 14376 15070 14385
rect 15014 14311 15070 14320
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14556 10192 14608 10198
rect 14556 10134 14608 10140
rect 14556 9920 14608 9926
rect 14556 9862 14608 9868
rect 14568 9722 14596 9862
rect 14556 9716 14608 9722
rect 14556 9658 14608 9664
rect 14660 9489 14688 12582
rect 14752 12170 14780 13806
rect 14844 13734 14872 14214
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14740 12164 14792 12170
rect 14740 12106 14792 12112
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14646 9480 14702 9489
rect 14556 9444 14608 9450
rect 14646 9415 14702 9424
rect 14556 9386 14608 9392
rect 14292 8894 14504 8922
rect 14186 8664 14242 8673
rect 14186 8599 14188 8608
rect 14240 8599 14242 8608
rect 14188 8570 14240 8576
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 13912 7948 13964 7954
rect 13912 7890 13964 7896
rect 13820 7540 13872 7546
rect 13820 7482 13872 7488
rect 13636 7404 13688 7410
rect 13740 7398 13860 7426
rect 13636 7346 13688 7352
rect 13544 6860 13596 6866
rect 13544 6802 13596 6808
rect 13464 6718 13584 6746
rect 13450 6080 13506 6089
rect 13450 6015 13506 6024
rect 13464 4826 13492 6015
rect 13556 5930 13584 6718
rect 13648 6390 13676 7346
rect 13728 7268 13780 7274
rect 13728 7210 13780 7216
rect 13740 7177 13768 7210
rect 13726 7168 13782 7177
rect 13726 7103 13782 7112
rect 13832 6882 13860 7398
rect 13924 7342 13952 7890
rect 14292 7426 14320 8894
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14384 8430 14412 8774
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 14384 7954 14412 8366
rect 14476 8242 14504 8774
rect 14568 8430 14596 9386
rect 14648 9376 14700 9382
rect 14646 9344 14648 9353
rect 14700 9344 14702 9353
rect 14646 9279 14702 9288
rect 14660 8537 14688 9279
rect 14646 8528 14702 8537
rect 14646 8463 14702 8472
rect 14556 8424 14608 8430
rect 14554 8392 14556 8401
rect 14608 8392 14610 8401
rect 14554 8327 14610 8336
rect 14476 8214 14596 8242
rect 14568 8090 14596 8214
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14464 8016 14516 8022
rect 14464 7958 14516 7964
rect 14372 7948 14424 7954
rect 14372 7890 14424 7896
rect 14292 7398 14412 7426
rect 14476 7410 14504 7958
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 13945 7100 14253 7120
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 13832 6854 13952 6882
rect 13728 6724 13780 6730
rect 13728 6666 13780 6672
rect 13740 6458 13768 6666
rect 13924 6662 13952 6854
rect 13912 6656 13964 6662
rect 13912 6598 13964 6604
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 14292 6322 14320 7210
rect 14280 6316 14332 6322
rect 14280 6258 14332 6264
rect 13728 6180 13780 6186
rect 13728 6122 13780 6128
rect 13556 5902 13676 5930
rect 13544 5840 13596 5846
rect 13544 5782 13596 5788
rect 13452 4820 13504 4826
rect 13452 4762 13504 4768
rect 13556 4622 13584 5782
rect 13648 5574 13676 5902
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 13636 5364 13688 5370
rect 13636 5306 13688 5312
rect 13648 5114 13676 5306
rect 13740 5302 13768 6122
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5710 13860 6054
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 13820 5704 13872 5710
rect 13820 5646 13872 5652
rect 13728 5296 13780 5302
rect 13728 5238 13780 5244
rect 13648 5086 13768 5114
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4690 13676 4966
rect 13636 4684 13688 4690
rect 13636 4626 13688 4632
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13740 4321 13768 5086
rect 13726 4312 13782 4321
rect 13544 4276 13596 4282
rect 13726 4247 13782 4256
rect 13544 4218 13596 4224
rect 13372 4134 13492 4162
rect 13360 4072 13412 4078
rect 13360 4014 13412 4020
rect 13372 3738 13400 4014
rect 13464 3738 13492 4134
rect 13360 3732 13412 3738
rect 13360 3674 13412 3680
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13372 3126 13400 3674
rect 13556 3602 13584 4218
rect 13728 4004 13780 4010
rect 13728 3946 13780 3952
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13740 3534 13768 3946
rect 13832 3942 13860 5646
rect 14292 5642 14320 6258
rect 14280 5636 14332 5642
rect 14280 5578 14332 5584
rect 14292 5166 14320 5578
rect 14280 5160 14332 5166
rect 14280 5102 14332 5108
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 14002 4720 14058 4729
rect 14002 4655 14058 4664
rect 14188 4684 14240 4690
rect 14016 4214 14044 4655
rect 14188 4626 14240 4632
rect 14096 4616 14148 4622
rect 14096 4558 14148 4564
rect 14108 4457 14136 4558
rect 14094 4448 14150 4457
rect 14094 4383 14150 4392
rect 14004 4208 14056 4214
rect 14004 4150 14056 4156
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13924 4049 13952 4082
rect 13910 4040 13966 4049
rect 14200 4010 14228 4626
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 14292 4282 14320 4422
rect 14280 4276 14332 4282
rect 14280 4218 14332 4224
rect 14384 4162 14412 7398
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14476 6866 14504 7346
rect 14464 6860 14516 6866
rect 14464 6802 14516 6808
rect 14660 6746 14688 8463
rect 14752 7290 14780 11222
rect 14844 9450 14872 13670
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14936 11762 14964 12922
rect 15028 12646 15056 14311
rect 15212 14074 15240 14894
rect 15304 14346 15332 15506
rect 15488 14929 15516 19332
rect 15580 18970 15608 20402
rect 15568 18964 15620 18970
rect 15568 18906 15620 18912
rect 15672 17864 15700 21490
rect 15856 20602 15884 22200
rect 16212 21616 16264 21622
rect 16212 21558 16264 21564
rect 16120 21480 16172 21486
rect 16120 21422 16172 21428
rect 16028 21140 16080 21146
rect 16028 21082 16080 21088
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15936 20460 15988 20466
rect 15936 20402 15988 20408
rect 15948 20058 15976 20402
rect 16040 20262 16068 21082
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16132 20058 16160 21422
rect 15936 20052 15988 20058
rect 15936 19994 15988 20000
rect 16120 20052 16172 20058
rect 16120 19994 16172 20000
rect 15844 19984 15896 19990
rect 15844 19926 15896 19932
rect 15752 19168 15804 19174
rect 15752 19110 15804 19116
rect 15764 18193 15792 19110
rect 15750 18184 15806 18193
rect 15750 18119 15806 18128
rect 15672 17836 15792 17864
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15580 17338 15608 17478
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15672 16726 15700 17002
rect 15660 16720 15712 16726
rect 15660 16662 15712 16668
rect 15658 16280 15714 16289
rect 15658 16215 15660 16224
rect 15712 16215 15714 16224
rect 15660 16186 15712 16192
rect 15660 15496 15712 15502
rect 15660 15438 15712 15444
rect 15672 15366 15700 15438
rect 15660 15360 15712 15366
rect 15660 15302 15712 15308
rect 15764 15201 15792 17836
rect 15750 15192 15806 15201
rect 15750 15127 15806 15136
rect 15752 15020 15804 15026
rect 15752 14962 15804 14968
rect 15474 14920 15530 14929
rect 15474 14855 15530 14864
rect 15476 14408 15528 14414
rect 15476 14350 15528 14356
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15108 13932 15160 13938
rect 15108 13874 15160 13880
rect 15120 13530 15148 13874
rect 15108 13524 15160 13530
rect 15108 13466 15160 13472
rect 15304 13394 15332 14282
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15200 13320 15252 13326
rect 15200 13262 15252 13268
rect 15108 13252 15160 13258
rect 15108 13194 15160 13200
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15120 11914 15148 13194
rect 15028 11886 15148 11914
rect 15212 11898 15240 13262
rect 15292 13184 15344 13190
rect 15292 13126 15344 13132
rect 15304 12986 15332 13126
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15396 12458 15424 14214
rect 15488 14074 15516 14350
rect 15658 14104 15714 14113
rect 15476 14068 15528 14074
rect 15658 14039 15714 14048
rect 15476 14010 15528 14016
rect 15672 14006 15700 14039
rect 15660 14000 15712 14006
rect 15660 13942 15712 13948
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 12850 15516 13262
rect 15568 13184 15620 13190
rect 15566 13152 15568 13161
rect 15620 13152 15622 13161
rect 15566 13087 15622 13096
rect 15672 12986 15700 13806
rect 15764 13530 15792 14962
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15660 12980 15712 12986
rect 15660 12922 15712 12928
rect 15476 12844 15528 12850
rect 15476 12786 15528 12792
rect 15568 12708 15620 12714
rect 15568 12650 15620 12656
rect 15396 12430 15516 12458
rect 15384 12232 15436 12238
rect 15384 12174 15436 12180
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15200 11892 15252 11898
rect 14924 11756 14976 11762
rect 14924 11698 14976 11704
rect 15028 11354 15056 11886
rect 15200 11834 15252 11840
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15016 11348 15068 11354
rect 15016 11290 15068 11296
rect 14924 11212 14976 11218
rect 14924 11154 14976 11160
rect 14936 10690 14964 11154
rect 15028 11082 15056 11290
rect 15016 11076 15068 11082
rect 15016 11018 15068 11024
rect 14936 10662 15056 10690
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10266 14964 10542
rect 14924 10260 14976 10266
rect 14924 10202 14976 10208
rect 14924 9920 14976 9926
rect 14924 9862 14976 9868
rect 14936 9761 14964 9862
rect 14922 9752 14978 9761
rect 15028 9722 15056 10662
rect 15120 10470 15148 11698
rect 15200 11348 15252 11354
rect 15200 11290 15252 11296
rect 15212 11257 15240 11290
rect 15304 11286 15332 12038
rect 15396 11762 15424 12174
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15292 11280 15344 11286
rect 15198 11248 15254 11257
rect 15292 11222 15344 11228
rect 15198 11183 15254 11192
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10130 15148 10406
rect 15212 10169 15240 11086
rect 15304 11014 15332 11222
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15292 10736 15344 10742
rect 15292 10678 15344 10684
rect 15198 10160 15254 10169
rect 15108 10124 15160 10130
rect 15198 10095 15254 10104
rect 15108 10066 15160 10072
rect 15304 9926 15332 10678
rect 15384 10600 15436 10606
rect 15384 10542 15436 10548
rect 15396 10198 15424 10542
rect 15384 10192 15436 10198
rect 15384 10134 15436 10140
rect 15396 10062 15424 10093
rect 15384 10056 15436 10062
rect 15382 10024 15384 10033
rect 15436 10024 15438 10033
rect 15382 9959 15438 9968
rect 15292 9920 15344 9926
rect 15292 9862 15344 9868
rect 15396 9722 15424 9959
rect 14922 9687 14978 9696
rect 15016 9716 15068 9722
rect 14832 9444 14884 9450
rect 14832 9386 14884 9392
rect 14936 9382 14964 9687
rect 15016 9658 15068 9664
rect 15384 9716 15436 9722
rect 15384 9658 15436 9664
rect 15028 9518 15056 9658
rect 15488 9654 15516 12430
rect 15580 10742 15608 12650
rect 15856 12594 15884 19926
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 15948 19242 15976 19790
rect 16224 19334 16252 21558
rect 16316 20346 16344 22200
rect 16684 22114 16712 22200
rect 16776 22114 16804 22222
rect 16684 22086 16804 22114
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 16672 20460 16724 20466
rect 16672 20402 16724 20408
rect 16316 20330 16620 20346
rect 16316 20324 16632 20330
rect 16316 20318 16580 20324
rect 16580 20266 16632 20272
rect 16396 20256 16448 20262
rect 16396 20198 16448 20204
rect 16408 19854 16436 20198
rect 16684 19854 16712 20402
rect 16960 19990 16988 22222
rect 17038 22200 17094 23000
rect 17406 22200 17462 23000
rect 17774 22200 17830 23000
rect 17958 22264 18014 22273
rect 17052 20058 17080 22200
rect 17314 20904 17370 20913
rect 17314 20839 17370 20848
rect 17132 20460 17184 20466
rect 17132 20402 17184 20408
rect 17040 20052 17092 20058
rect 17040 19994 17092 20000
rect 16948 19984 17000 19990
rect 16948 19926 17000 19932
rect 16396 19848 16448 19854
rect 16396 19790 16448 19796
rect 16672 19848 16724 19854
rect 16672 19790 16724 19796
rect 16948 19848 17000 19854
rect 17000 19796 17080 19802
rect 16948 19790 17080 19796
rect 16132 19306 16252 19334
rect 15936 19236 15988 19242
rect 15936 19178 15988 19184
rect 15936 18760 15988 18766
rect 15936 18702 15988 18708
rect 15948 18426 15976 18702
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16028 17740 16080 17746
rect 16028 17682 16080 17688
rect 15936 17536 15988 17542
rect 15936 17478 15988 17484
rect 15948 16250 15976 17478
rect 16040 16590 16068 17682
rect 16132 17218 16160 19306
rect 16304 19304 16356 19310
rect 16304 19246 16356 19252
rect 16316 18306 16344 19246
rect 16408 19174 16436 19790
rect 16960 19774 17080 19790
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 17052 19174 17080 19774
rect 17144 19718 17172 20402
rect 17224 20256 17276 20262
rect 17224 20198 17276 20204
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 16396 19168 16448 19174
rect 16396 19110 16448 19116
rect 17040 19168 17092 19174
rect 17040 19110 17092 19116
rect 16408 18426 16436 19110
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 17052 18442 17080 19110
rect 17236 18766 17264 20198
rect 17328 19514 17356 20839
rect 17420 19990 17448 22200
rect 17500 20528 17552 20534
rect 17500 20470 17552 20476
rect 17408 19984 17460 19990
rect 17408 19926 17460 19932
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17328 18902 17356 19178
rect 17420 18970 17448 19790
rect 17512 18970 17540 20470
rect 17788 20058 17816 22200
rect 17958 22199 18014 22208
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 18970 22200 19026 23000
rect 19338 22200 19394 23000
rect 19706 22200 19762 23000
rect 20074 22200 20130 23000
rect 20442 22200 20498 23000
rect 20534 22672 20590 22681
rect 20534 22607 20590 22616
rect 17868 21344 17920 21350
rect 17868 21286 17920 21292
rect 17776 20052 17828 20058
rect 17776 19994 17828 20000
rect 17592 19848 17644 19854
rect 17592 19790 17644 19796
rect 17604 19514 17632 19790
rect 17880 19514 17908 21286
rect 17972 20602 18000 22199
rect 18156 20602 18184 22200
rect 17960 20596 18012 20602
rect 17960 20538 18012 20544
rect 18144 20596 18196 20602
rect 18144 20538 18196 20544
rect 18616 20330 18644 22200
rect 18984 20534 19012 22200
rect 18972 20528 19024 20534
rect 18972 20470 19024 20476
rect 18878 20360 18934 20369
rect 18604 20324 18656 20330
rect 18878 20295 18934 20304
rect 18604 20266 18656 20272
rect 18892 20058 18920 20295
rect 19352 20244 19380 22200
rect 19720 21978 19748 22200
rect 19720 21950 19932 21978
rect 19706 21856 19762 21865
rect 19706 21791 19762 21800
rect 19524 20596 19576 20602
rect 19524 20538 19576 20544
rect 19430 20496 19486 20505
rect 19536 20466 19564 20538
rect 19430 20431 19486 20440
rect 19524 20460 19576 20466
rect 19444 20398 19472 20431
rect 19524 20402 19576 20408
rect 19432 20392 19484 20398
rect 19432 20334 19484 20340
rect 19616 20256 19668 20262
rect 19352 20216 19564 20244
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 18696 20052 18748 20058
rect 18696 19994 18748 20000
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18604 19780 18656 19786
rect 18604 19722 18656 19728
rect 18512 19712 18564 19718
rect 18512 19654 18564 19660
rect 18050 19544 18106 19553
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17868 19508 17920 19514
rect 18050 19479 18106 19488
rect 18156 19502 18460 19530
rect 18524 19514 18552 19654
rect 17868 19450 17920 19456
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 17592 19304 17644 19310
rect 17592 19246 17644 19252
rect 17408 18964 17460 18970
rect 17408 18906 17460 18912
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17316 18896 17368 18902
rect 17316 18838 17368 18844
rect 17224 18760 17276 18766
rect 17224 18702 17276 18708
rect 17408 18624 17460 18630
rect 17406 18592 17408 18601
rect 17604 18612 17632 19246
rect 17972 18902 18000 19314
rect 18064 18970 18092 19479
rect 18156 19446 18184 19502
rect 18144 19440 18196 19446
rect 18144 19382 18196 19388
rect 18432 19378 18460 19502
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18510 19408 18566 19417
rect 18236 19372 18288 19378
rect 18420 19372 18472 19378
rect 18288 19332 18368 19360
rect 18236 19314 18288 19320
rect 18234 19000 18290 19009
rect 18052 18964 18104 18970
rect 18234 18935 18236 18944
rect 18052 18906 18104 18912
rect 18288 18935 18290 18944
rect 18236 18906 18288 18912
rect 17960 18896 18012 18902
rect 17960 18838 18012 18844
rect 18236 18760 18288 18766
rect 18236 18702 18288 18708
rect 17460 18592 17632 18612
rect 17462 18584 17632 18592
rect 17406 18527 17462 18536
rect 16396 18420 16448 18426
rect 17052 18414 17172 18442
rect 18248 18426 18276 18702
rect 18340 18630 18368 19332
rect 18510 19343 18566 19352
rect 18420 19314 18472 19320
rect 18524 19258 18552 19343
rect 18432 19230 18552 19258
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 16396 18362 16448 18368
rect 16316 18278 16620 18306
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16224 17338 16252 17546
rect 16304 17536 16356 17542
rect 16304 17478 16356 17484
rect 16316 17338 16344 17478
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16132 17190 16252 17218
rect 16408 17202 16436 18090
rect 16592 17785 16620 18278
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16854 17912 16910 17921
rect 16854 17847 16910 17856
rect 16578 17776 16634 17785
rect 16868 17746 16896 17847
rect 16578 17711 16634 17720
rect 16856 17740 16908 17746
rect 16856 17682 16908 17688
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 16028 16040 16080 16046
rect 16028 15982 16080 15988
rect 15936 14952 15988 14958
rect 15936 14894 15988 14900
rect 15948 14618 15976 14894
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15948 13870 15976 14554
rect 15936 13864 15988 13870
rect 15936 13806 15988 13812
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15948 12986 15976 13194
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15934 12880 15990 12889
rect 15934 12815 15936 12824
rect 15988 12815 15990 12824
rect 15936 12786 15988 12792
rect 15672 12566 15884 12594
rect 15672 12102 15700 12566
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15764 11898 15792 12378
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 15672 11121 15700 11698
rect 15764 11218 15792 11834
rect 15856 11694 15884 12378
rect 15936 11824 15988 11830
rect 15936 11766 15988 11772
rect 15844 11688 15896 11694
rect 15844 11630 15896 11636
rect 15844 11280 15896 11286
rect 15948 11257 15976 11766
rect 15844 11222 15896 11228
rect 15934 11248 15990 11257
rect 15752 11212 15804 11218
rect 15752 11154 15804 11160
rect 15658 11112 15714 11121
rect 15658 11047 15714 11056
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15568 10736 15620 10742
rect 15568 10678 15620 10684
rect 15566 10160 15622 10169
rect 15566 10095 15622 10104
rect 15580 9926 15608 10095
rect 15672 9926 15700 10950
rect 15764 10742 15792 10950
rect 15752 10736 15804 10742
rect 15752 10678 15804 10684
rect 15764 10577 15792 10678
rect 15750 10568 15806 10577
rect 15750 10503 15806 10512
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15764 9994 15792 10202
rect 15752 9988 15804 9994
rect 15752 9930 15804 9936
rect 15568 9920 15620 9926
rect 15568 9862 15620 9868
rect 15660 9920 15712 9926
rect 15660 9862 15712 9868
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15474 9480 15530 9489
rect 15474 9415 15530 9424
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14830 9208 14886 9217
rect 14830 9143 14886 9152
rect 14844 8974 14872 9143
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14844 8634 14872 8910
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14832 8356 14884 8362
rect 14832 8298 14884 8304
rect 14844 8022 14872 8298
rect 14832 8016 14884 8022
rect 14832 7958 14884 7964
rect 14832 7744 14884 7750
rect 14830 7712 14832 7721
rect 14884 7712 14886 7721
rect 14830 7647 14886 7656
rect 14844 7410 14872 7647
rect 14832 7404 14884 7410
rect 14832 7346 14884 7352
rect 14752 7262 14872 7290
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14292 4134 14412 4162
rect 14476 6718 14688 6746
rect 13910 3975 13966 3984
rect 14188 4004 14240 4010
rect 14188 3946 14240 3952
rect 13820 3936 13872 3942
rect 13820 3878 13872 3884
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 13728 3528 13780 3534
rect 13728 3470 13780 3476
rect 13728 3392 13780 3398
rect 13728 3334 13780 3340
rect 13820 3392 13872 3398
rect 13820 3334 13872 3340
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13740 2990 13768 3334
rect 13728 2984 13780 2990
rect 13728 2926 13780 2932
rect 12820 2746 12940 2774
rect 13188 2746 13308 2774
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 12624 1964 12676 1970
rect 12624 1906 12676 1912
rect 12728 800 12756 2586
rect 12820 1086 12848 2746
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 12808 1080 12860 1086
rect 12808 1022 12860 1028
rect 13096 800 13124 2518
rect 13188 1290 13216 2746
rect 13832 2582 13860 3334
rect 14292 2961 14320 4134
rect 14372 4072 14424 4078
rect 14476 4049 14504 6718
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14568 5574 14596 6598
rect 14648 6384 14700 6390
rect 14648 6326 14700 6332
rect 14660 5778 14688 6326
rect 14752 5778 14780 7142
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14740 5772 14792 5778
rect 14740 5714 14792 5720
rect 14556 5568 14608 5574
rect 14556 5510 14608 5516
rect 14660 5166 14688 5714
rect 14738 5536 14794 5545
rect 14738 5471 14794 5480
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14752 4758 14780 5471
rect 14740 4752 14792 4758
rect 14738 4720 14740 4729
rect 14792 4720 14794 4729
rect 14738 4655 14794 4664
rect 14556 4480 14608 4486
rect 14556 4422 14608 4428
rect 14740 4480 14792 4486
rect 14740 4422 14792 4428
rect 14372 4014 14424 4020
rect 14462 4040 14518 4049
rect 14384 3505 14412 4014
rect 14462 3975 14518 3984
rect 14464 3936 14516 3942
rect 14464 3878 14516 3884
rect 14476 3534 14504 3878
rect 14464 3528 14516 3534
rect 14370 3496 14426 3505
rect 14464 3470 14516 3476
rect 14370 3431 14426 3440
rect 14278 2952 14334 2961
rect 14278 2887 14334 2896
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14464 2848 14516 2854
rect 14464 2790 14516 2796
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 14292 2650 14320 2790
rect 14280 2644 14332 2650
rect 14280 2586 14332 2592
rect 13820 2576 13872 2582
rect 13820 2518 13872 2524
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13176 1284 13228 1290
rect 13176 1226 13228 1232
rect 13556 800 13584 2246
rect 14016 800 14044 2518
rect 14476 2378 14504 2790
rect 14568 2378 14596 4422
rect 14648 4072 14700 4078
rect 14648 4014 14700 4020
rect 14660 3913 14688 4014
rect 14646 3904 14702 3913
rect 14646 3839 14702 3848
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14660 2922 14688 3538
rect 14648 2916 14700 2922
rect 14648 2858 14700 2864
rect 14646 2680 14702 2689
rect 14646 2615 14702 2624
rect 14464 2372 14516 2378
rect 14464 2314 14516 2320
rect 14556 2372 14608 2378
rect 14556 2314 14608 2320
rect 14372 2304 14424 2310
rect 14372 2246 14424 2252
rect 14384 800 14412 2246
rect 14660 950 14688 2615
rect 14752 2446 14780 4422
rect 14844 3670 14872 7262
rect 14936 6118 14964 9318
rect 15382 9208 15438 9217
rect 15108 9172 15160 9178
rect 15382 9143 15438 9152
rect 15108 9114 15160 9120
rect 15016 8832 15068 8838
rect 15016 8774 15068 8780
rect 15028 8430 15056 8774
rect 15016 8424 15068 8430
rect 15016 8366 15068 8372
rect 15016 8084 15068 8090
rect 15016 8026 15068 8032
rect 14924 6112 14976 6118
rect 14924 6054 14976 6060
rect 14922 5944 14978 5953
rect 15028 5930 15056 8026
rect 15120 7546 15148 9114
rect 15396 8673 15424 9143
rect 15382 8664 15438 8673
rect 15488 8634 15516 9415
rect 15580 9353 15608 9862
rect 15672 9761 15700 9862
rect 15658 9752 15714 9761
rect 15658 9687 15660 9696
rect 15712 9687 15714 9696
rect 15660 9658 15712 9664
rect 15672 9627 15700 9658
rect 15660 9512 15712 9518
rect 15660 9454 15712 9460
rect 15566 9344 15622 9353
rect 15566 9279 15622 9288
rect 15568 9036 15620 9042
rect 15568 8978 15620 8984
rect 15382 8599 15438 8608
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15384 8288 15436 8294
rect 15198 8256 15254 8265
rect 15384 8230 15436 8236
rect 15198 8191 15254 8200
rect 15212 7585 15240 8191
rect 15396 7886 15424 8230
rect 15580 8090 15608 8978
rect 15568 8084 15620 8090
rect 15568 8026 15620 8032
rect 15384 7880 15436 7886
rect 15384 7822 15436 7828
rect 15476 7744 15528 7750
rect 15476 7686 15528 7692
rect 15672 7698 15700 9454
rect 15752 9376 15804 9382
rect 15752 9318 15804 9324
rect 15764 7818 15792 9318
rect 15856 8974 15884 11222
rect 15934 11183 15990 11192
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 15948 10810 15976 10950
rect 15936 10804 15988 10810
rect 15936 10746 15988 10752
rect 15948 10266 15976 10746
rect 16040 10538 16068 15982
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 16132 15162 16160 15302
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16132 13394 16160 14214
rect 16224 13734 16252 17190
rect 16396 17196 16448 17202
rect 16396 17138 16448 17144
rect 16960 17066 16988 18226
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 16948 17060 17000 17066
rect 16948 17002 17000 17008
rect 16396 16992 16448 16998
rect 16396 16934 16448 16940
rect 16408 15502 16436 16934
rect 16948 16516 17000 16522
rect 16948 16458 17000 16464
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 16960 16130 16988 16458
rect 16776 16114 16988 16130
rect 16764 16108 16988 16114
rect 16816 16102 16988 16108
rect 16764 16050 16816 16056
rect 16776 15706 16804 16050
rect 16764 15700 16816 15706
rect 16764 15642 16816 15648
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16304 15360 16356 15366
rect 16304 15302 16356 15308
rect 16316 14414 16344 15302
rect 16408 15065 16436 15438
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 16394 15056 16450 15065
rect 16394 14991 16450 15000
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16316 13938 16344 14350
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16132 12782 16160 13330
rect 16212 13320 16264 13326
rect 16212 13262 16264 13268
rect 16224 13190 16252 13262
rect 16212 13184 16264 13190
rect 16212 13126 16264 13132
rect 16120 12776 16172 12782
rect 16120 12718 16172 12724
rect 16212 12776 16264 12782
rect 16212 12718 16264 12724
rect 16120 12640 16172 12646
rect 16224 12617 16252 12718
rect 16120 12582 16172 12588
rect 16210 12608 16266 12617
rect 16132 12374 16160 12582
rect 16210 12543 16266 12552
rect 16120 12368 16172 12374
rect 16120 12310 16172 12316
rect 16132 11354 16160 12310
rect 16316 12238 16344 13874
rect 16408 13326 16436 14894
rect 16948 14816 17000 14822
rect 16948 14758 17000 14764
rect 16960 14278 16988 14758
rect 16948 14272 17000 14278
rect 16948 14214 17000 14220
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 16580 13864 16632 13870
rect 16580 13806 16632 13812
rect 16592 13705 16620 13806
rect 16672 13728 16724 13734
rect 16578 13696 16634 13705
rect 16672 13670 16724 13676
rect 16578 13631 16634 13640
rect 16396 13320 16448 13326
rect 16684 13297 16712 13670
rect 16396 13262 16448 13268
rect 16670 13288 16726 13297
rect 16670 13223 16726 13232
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16408 12850 16436 13126
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16960 12850 16988 14214
rect 17052 13682 17080 17614
rect 17144 16998 17172 18414
rect 17592 18420 17644 18426
rect 17592 18362 17644 18368
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 17314 18320 17370 18329
rect 17314 18255 17370 18264
rect 17408 18284 17460 18290
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17236 16794 17264 17070
rect 17328 16794 17356 18255
rect 17408 18226 17460 18232
rect 17420 17882 17448 18226
rect 17408 17876 17460 17882
rect 17408 17818 17460 17824
rect 17224 16788 17276 16794
rect 17224 16730 17276 16736
rect 17316 16788 17368 16794
rect 17316 16730 17368 16736
rect 17236 16250 17264 16730
rect 17500 16720 17552 16726
rect 17500 16662 17552 16668
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17224 16244 17276 16250
rect 17224 16186 17276 16192
rect 17130 16008 17186 16017
rect 17130 15943 17186 15952
rect 17144 14074 17172 15943
rect 17222 14512 17278 14521
rect 17222 14447 17278 14456
rect 17236 14278 17264 14447
rect 17224 14272 17276 14278
rect 17222 14240 17224 14249
rect 17276 14240 17278 14249
rect 17222 14175 17278 14184
rect 17222 14104 17278 14113
rect 17132 14068 17184 14074
rect 17222 14039 17278 14048
rect 17132 14010 17184 14016
rect 17236 13938 17264 14039
rect 17224 13932 17276 13938
rect 17224 13874 17276 13880
rect 17132 13864 17184 13870
rect 17130 13832 17132 13841
rect 17184 13832 17186 13841
rect 17130 13767 17186 13776
rect 17224 13796 17276 13802
rect 17224 13738 17276 13744
rect 17052 13654 17172 13682
rect 17038 13288 17094 13297
rect 17038 13223 17094 13232
rect 16396 12844 16448 12850
rect 16396 12786 16448 12792
rect 16948 12844 17000 12850
rect 16948 12786 17000 12792
rect 16408 12442 16436 12786
rect 17052 12782 17080 13223
rect 17040 12776 17092 12782
rect 17040 12718 17092 12724
rect 16762 12608 16818 12617
rect 16762 12543 16818 12552
rect 16396 12436 16448 12442
rect 16396 12378 16448 12384
rect 16580 12300 16632 12306
rect 16776 12288 16804 12543
rect 16946 12472 17002 12481
rect 16946 12407 17002 12416
rect 16580 12242 16632 12248
rect 16684 12260 16804 12288
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16396 12232 16448 12238
rect 16592 12209 16620 12242
rect 16396 12174 16448 12180
rect 16578 12200 16634 12209
rect 16212 12096 16264 12102
rect 16212 12038 16264 12044
rect 16302 12064 16358 12073
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16132 10810 16160 11086
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 16028 10532 16080 10538
rect 16028 10474 16080 10480
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15936 10124 15988 10130
rect 15936 10066 15988 10072
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15856 8090 15884 8910
rect 15948 8566 15976 10066
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15948 8294 15976 8502
rect 15936 8288 15988 8294
rect 15936 8230 15988 8236
rect 15844 8084 15896 8090
rect 15844 8026 15896 8032
rect 15842 7984 15898 7993
rect 15842 7919 15844 7928
rect 15896 7919 15898 7928
rect 15844 7890 15896 7896
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15198 7576 15254 7585
rect 15108 7540 15160 7546
rect 15198 7511 15254 7520
rect 15108 7482 15160 7488
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15200 7404 15252 7410
rect 15200 7346 15252 7352
rect 15108 7200 15160 7206
rect 15108 7142 15160 7148
rect 15120 6254 15148 7142
rect 15108 6248 15160 6254
rect 15108 6190 15160 6196
rect 15120 6089 15148 6190
rect 15106 6080 15162 6089
rect 15106 6015 15162 6024
rect 14978 5902 15056 5930
rect 14922 5879 14978 5888
rect 14936 5681 14964 5879
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 14922 5672 14978 5681
rect 14922 5607 14978 5616
rect 15016 5636 15068 5642
rect 14936 5370 14964 5607
rect 15016 5578 15068 5584
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 3058 14872 3606
rect 14936 3466 14964 5170
rect 14924 3460 14976 3466
rect 14924 3402 14976 3408
rect 14936 3369 14964 3402
rect 14922 3360 14978 3369
rect 14922 3295 14978 3304
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14832 2576 14884 2582
rect 14832 2518 14884 2524
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14648 944 14700 950
rect 14648 886 14700 892
rect 14844 800 14872 2518
rect 14936 1329 14964 3130
rect 15028 3126 15056 5578
rect 15120 4690 15148 5714
rect 15108 4684 15160 4690
rect 15108 4626 15160 4632
rect 15120 4010 15148 4626
rect 15108 4004 15160 4010
rect 15108 3946 15160 3952
rect 15106 3768 15162 3777
rect 15106 3703 15162 3712
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 15120 2774 15148 3703
rect 15212 3194 15240 7346
rect 15292 6724 15344 6730
rect 15292 6666 15344 6672
rect 15304 6186 15332 6666
rect 15292 6180 15344 6186
rect 15292 6122 15344 6128
rect 15304 5930 15332 6122
rect 15396 6066 15424 7414
rect 15488 6390 15516 7686
rect 15672 7670 15792 7698
rect 15764 7410 15792 7670
rect 15752 7404 15804 7410
rect 15752 7346 15804 7352
rect 15566 7168 15622 7177
rect 15566 7103 15622 7112
rect 15580 6662 15608 7103
rect 15658 7032 15714 7041
rect 15764 7002 15792 7346
rect 15948 7342 15976 8230
rect 16040 7546 16068 10474
rect 16120 10260 16172 10266
rect 16120 10202 16172 10208
rect 16132 9160 16160 10202
rect 16224 10130 16252 12038
rect 16302 11999 16358 12008
rect 16316 11830 16344 11999
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16316 11529 16344 11766
rect 16302 11520 16358 11529
rect 16302 11455 16358 11464
rect 16408 11082 16436 12174
rect 16684 12170 16712 12260
rect 16762 12200 16818 12209
rect 16578 12135 16634 12144
rect 16672 12164 16724 12170
rect 16960 12170 16988 12407
rect 17040 12300 17092 12306
rect 17040 12242 17092 12248
rect 16762 12135 16764 12144
rect 16672 12106 16724 12112
rect 16816 12135 16818 12144
rect 16948 12164 17000 12170
rect 16764 12106 16816 12112
rect 16948 12106 17000 12112
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 17052 11937 17080 12242
rect 17038 11928 17094 11937
rect 17038 11863 17094 11872
rect 16488 11756 16540 11762
rect 16672 11756 16724 11762
rect 16540 11716 16620 11744
rect 16488 11698 16540 11704
rect 16592 11234 16620 11716
rect 16672 11698 16724 11704
rect 16684 11354 16712 11698
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16592 11206 17080 11234
rect 16396 11076 16448 11082
rect 16396 11018 16448 11024
rect 16948 11076 17000 11082
rect 16948 11018 17000 11024
rect 16212 10124 16264 10130
rect 16212 10066 16264 10072
rect 16408 10062 16436 11018
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16960 10606 16988 11018
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 16960 10198 16988 10542
rect 16948 10192 17000 10198
rect 16948 10134 17000 10140
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 16212 9988 16264 9994
rect 16212 9930 16264 9936
rect 16304 9988 16356 9994
rect 16304 9930 16356 9936
rect 16224 9722 16252 9930
rect 16212 9716 16264 9722
rect 16212 9658 16264 9664
rect 16316 9654 16344 9930
rect 16396 9920 16448 9926
rect 16396 9862 16448 9868
rect 16304 9648 16356 9654
rect 16210 9616 16266 9625
rect 16304 9590 16356 9596
rect 16210 9551 16212 9560
rect 16264 9551 16266 9560
rect 16212 9522 16264 9528
rect 16132 9132 16344 9160
rect 16212 9036 16264 9042
rect 16212 8978 16264 8984
rect 16120 8832 16172 8838
rect 16120 8774 16172 8780
rect 16132 8634 16160 8774
rect 16120 8628 16172 8634
rect 16120 8570 16172 8576
rect 16118 8392 16174 8401
rect 16118 8327 16174 8336
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16132 7426 16160 8327
rect 16224 7970 16252 8978
rect 16316 8412 16344 9132
rect 16408 8616 16436 9862
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 16960 9722 16988 9998
rect 16948 9716 17000 9722
rect 16948 9658 17000 9664
rect 16488 9648 16540 9654
rect 16488 9590 16540 9596
rect 16946 9616 17002 9625
rect 16500 9042 16528 9590
rect 16946 9551 17002 9560
rect 16488 9036 16540 9042
rect 16488 8978 16540 8984
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16408 8588 16620 8616
rect 16592 8548 16620 8588
rect 16764 8560 16816 8566
rect 16592 8520 16764 8548
rect 16764 8502 16816 8508
rect 16856 8424 16908 8430
rect 16316 8384 16436 8412
rect 16224 7942 16344 7970
rect 16212 7880 16264 7886
rect 16212 7822 16264 7828
rect 16224 7750 16252 7822
rect 16212 7744 16264 7750
rect 16212 7686 16264 7692
rect 16040 7398 16160 7426
rect 16224 7410 16252 7686
rect 16316 7546 16344 7942
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16212 7404 16264 7410
rect 15936 7336 15988 7342
rect 15936 7278 15988 7284
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15658 6967 15660 6976
rect 15712 6967 15714 6976
rect 15752 6996 15804 7002
rect 15660 6938 15712 6944
rect 15752 6938 15804 6944
rect 15948 6934 15976 7142
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 15936 6792 15988 6798
rect 15658 6760 15714 6769
rect 15936 6734 15988 6740
rect 15658 6695 15714 6704
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15488 6202 15516 6326
rect 15672 6322 15700 6695
rect 15856 6662 15884 6693
rect 15844 6656 15896 6662
rect 15842 6624 15844 6633
rect 15896 6624 15898 6633
rect 15842 6559 15898 6568
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15488 6174 15700 6202
rect 15396 6038 15516 6066
rect 15304 5902 15424 5930
rect 15488 5914 15516 6038
rect 15290 5808 15346 5817
rect 15290 5743 15346 5752
rect 15304 5370 15332 5743
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15396 5234 15424 5902
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15672 5817 15700 6174
rect 15658 5808 15714 5817
rect 15658 5743 15714 5752
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15384 5228 15436 5234
rect 15384 5170 15436 5176
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15304 4185 15332 5102
rect 15476 5092 15528 5098
rect 15476 5034 15528 5040
rect 15384 5024 15436 5030
rect 15384 4966 15436 4972
rect 15396 4622 15424 4966
rect 15384 4616 15436 4622
rect 15384 4558 15436 4564
rect 15396 4321 15424 4558
rect 15382 4312 15438 4321
rect 15488 4282 15516 5034
rect 15382 4247 15438 4256
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15580 4214 15608 5238
rect 15672 5030 15700 5743
rect 15856 5710 15884 6559
rect 15948 6118 15976 6734
rect 16040 6497 16068 7398
rect 16212 7346 16264 7352
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16224 6914 16252 7210
rect 16224 6886 16344 6914
rect 16120 6792 16172 6798
rect 16316 6746 16344 6886
rect 16120 6734 16172 6740
rect 16132 6633 16160 6734
rect 16224 6718 16344 6746
rect 16118 6624 16174 6633
rect 16118 6559 16174 6568
rect 16026 6488 16082 6497
rect 16026 6423 16082 6432
rect 16120 6316 16172 6322
rect 16120 6258 16172 6264
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15844 5704 15896 5710
rect 15844 5646 15896 5652
rect 15750 5400 15806 5409
rect 15750 5335 15806 5344
rect 15764 5302 15792 5335
rect 15752 5296 15804 5302
rect 15752 5238 15804 5244
rect 15856 5166 15884 5646
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15660 5024 15712 5030
rect 15660 4966 15712 4972
rect 15660 4752 15712 4758
rect 15660 4694 15712 4700
rect 15568 4208 15620 4214
rect 15290 4176 15346 4185
rect 15568 4150 15620 4156
rect 15290 4111 15346 4120
rect 15476 4140 15528 4146
rect 15476 4082 15528 4088
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 15382 4040 15438 4049
rect 15304 3602 15332 4014
rect 15382 3975 15438 3984
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15200 3188 15252 3194
rect 15200 3130 15252 3136
rect 15198 3088 15254 3097
rect 15396 3058 15424 3975
rect 15488 3738 15516 4082
rect 15476 3732 15528 3738
rect 15476 3674 15528 3680
rect 15474 3632 15530 3641
rect 15474 3567 15530 3576
rect 15488 3534 15516 3567
rect 15476 3528 15528 3534
rect 15476 3470 15528 3476
rect 15198 3023 15254 3032
rect 15384 3052 15436 3058
rect 15212 2922 15240 3023
rect 15384 2994 15436 3000
rect 15566 2952 15622 2961
rect 15200 2916 15252 2922
rect 15566 2887 15568 2896
rect 15200 2858 15252 2864
rect 15620 2887 15622 2896
rect 15568 2858 15620 2864
rect 15028 2746 15148 2774
rect 15028 1834 15056 2746
rect 15672 2530 15700 4694
rect 15750 4040 15806 4049
rect 15750 3975 15806 3984
rect 15764 3058 15792 3975
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15948 3890 15976 6054
rect 16132 4010 16160 6258
rect 16120 4004 16172 4010
rect 16120 3946 16172 3952
rect 15856 3641 15884 3878
rect 15948 3862 16160 3890
rect 15934 3768 15990 3777
rect 15934 3703 15990 3712
rect 15842 3632 15898 3641
rect 15842 3567 15898 3576
rect 15948 3534 15976 3703
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 15936 3392 15988 3398
rect 15936 3334 15988 3340
rect 15752 3052 15804 3058
rect 15752 2994 15804 3000
rect 15948 2650 15976 3334
rect 16040 2990 16068 3402
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16028 2576 16080 2582
rect 15672 2502 15976 2530
rect 16028 2518 16080 2524
rect 15948 2446 15976 2502
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15200 2304 15252 2310
rect 15200 2246 15252 2252
rect 15752 2304 15804 2310
rect 15752 2246 15804 2252
rect 15016 1828 15068 1834
rect 15016 1770 15068 1776
rect 14922 1320 14978 1329
rect 14922 1255 14978 1264
rect 15212 800 15240 2246
rect 15764 1170 15792 2246
rect 15672 1142 15792 1170
rect 15672 800 15700 1142
rect 16040 800 16068 2518
rect 16132 1902 16160 3862
rect 16224 3058 16252 6718
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16316 6458 16344 6598
rect 16304 6452 16356 6458
rect 16304 6394 16356 6400
rect 16408 6372 16436 8384
rect 16960 8401 16988 9551
rect 17052 9110 17080 11206
rect 17144 9178 17172 13654
rect 17236 12442 17264 13738
rect 17328 13433 17356 16594
rect 17512 16454 17540 16662
rect 17500 16448 17552 16454
rect 17500 16390 17552 16396
rect 17512 15858 17540 16390
rect 17420 15830 17540 15858
rect 17420 15706 17448 15830
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17500 15700 17552 15706
rect 17500 15642 17552 15648
rect 17408 15564 17460 15570
rect 17408 15506 17460 15512
rect 17420 14822 17448 15506
rect 17512 15502 17540 15642
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17408 14816 17460 14822
rect 17408 14758 17460 14764
rect 17512 14482 17540 15438
rect 17604 15348 17632 18362
rect 17958 17912 18014 17921
rect 17958 17847 18014 17856
rect 17774 17096 17830 17105
rect 17774 17031 17830 17040
rect 17788 16726 17816 17031
rect 17972 16726 18000 17847
rect 18052 17808 18104 17814
rect 18052 17750 18104 17756
rect 17776 16720 17828 16726
rect 17960 16720 18012 16726
rect 17776 16662 17828 16668
rect 17866 16688 17922 16697
rect 17960 16662 18012 16668
rect 17866 16623 17868 16632
rect 17920 16623 17922 16632
rect 17868 16594 17920 16600
rect 18064 16522 18092 17750
rect 18144 17536 18196 17542
rect 18144 17478 18196 17484
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 18064 16250 18092 16458
rect 18052 16244 18104 16250
rect 18052 16186 18104 16192
rect 17960 15904 18012 15910
rect 17960 15846 18012 15852
rect 17868 15564 17920 15570
rect 17868 15506 17920 15512
rect 17880 15366 17908 15506
rect 17776 15360 17828 15366
rect 17604 15320 17724 15348
rect 17592 15156 17644 15162
rect 17592 15098 17644 15104
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17314 13424 17370 13433
rect 17314 13359 17370 13368
rect 17224 12436 17276 12442
rect 17224 12378 17276 12384
rect 17316 12368 17368 12374
rect 17316 12310 17368 12316
rect 17224 12096 17276 12102
rect 17328 12073 17356 12310
rect 17420 12306 17448 14214
rect 17604 13870 17632 15098
rect 17592 13864 17644 13870
rect 17592 13806 17644 13812
rect 17696 13682 17724 15320
rect 17776 15302 17828 15308
rect 17868 15360 17920 15366
rect 17868 15302 17920 15308
rect 17512 13654 17724 13682
rect 17408 12300 17460 12306
rect 17408 12242 17460 12248
rect 17512 12102 17540 13654
rect 17592 13184 17644 13190
rect 17590 13152 17592 13161
rect 17644 13152 17646 13161
rect 17590 13087 17646 13096
rect 17592 12980 17644 12986
rect 17592 12922 17644 12928
rect 17604 12850 17632 12922
rect 17788 12850 17816 15302
rect 17868 14340 17920 14346
rect 17868 14282 17920 14288
rect 17880 13870 17908 14282
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17592 12844 17644 12850
rect 17776 12844 17828 12850
rect 17592 12786 17644 12792
rect 17696 12804 17776 12832
rect 17500 12096 17552 12102
rect 17224 12038 17276 12044
rect 17314 12064 17370 12073
rect 17236 9738 17264 12038
rect 17500 12038 17552 12044
rect 17314 11999 17370 12008
rect 17408 11552 17460 11558
rect 17408 11494 17460 11500
rect 17316 11076 17368 11082
rect 17316 11018 17368 11024
rect 17328 10266 17356 11018
rect 17420 10305 17448 11494
rect 17512 11234 17540 12038
rect 17604 11830 17632 12786
rect 17696 12306 17724 12804
rect 17776 12786 17828 12792
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17592 11824 17644 11830
rect 17592 11766 17644 11772
rect 17512 11206 17632 11234
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17406 10296 17462 10305
rect 17316 10260 17368 10266
rect 17406 10231 17462 10240
rect 17316 10202 17368 10208
rect 17512 10130 17540 11086
rect 17500 10124 17552 10130
rect 17500 10066 17552 10072
rect 17604 9874 17632 11206
rect 17420 9846 17632 9874
rect 17236 9710 17356 9738
rect 17328 9654 17356 9710
rect 17316 9648 17368 9654
rect 17420 9625 17448 9846
rect 17696 9674 17724 12106
rect 17788 11150 17816 12582
rect 17972 12434 18000 15846
rect 18052 13932 18104 13938
rect 18052 13874 18104 13880
rect 18064 13530 18092 13874
rect 18052 13524 18104 13530
rect 18156 13512 18184 17478
rect 18432 16454 18460 19230
rect 18510 18456 18566 18465
rect 18510 18391 18512 18400
rect 18564 18391 18566 18400
rect 18512 18362 18564 18368
rect 18510 18184 18566 18193
rect 18510 18119 18566 18128
rect 18524 17066 18552 18119
rect 18512 17060 18564 17066
rect 18512 17002 18564 17008
rect 18616 16726 18644 19722
rect 18708 18873 18736 19994
rect 18788 19984 18840 19990
rect 18788 19926 18840 19932
rect 19064 19984 19116 19990
rect 19064 19926 19116 19932
rect 18800 19514 18828 19926
rect 18880 19848 18932 19854
rect 18878 19816 18880 19825
rect 18932 19816 18934 19825
rect 18878 19751 18934 19760
rect 18788 19508 18840 19514
rect 18788 19450 18840 19456
rect 18892 19417 18920 19751
rect 18878 19408 18934 19417
rect 18878 19343 18934 19352
rect 18972 19372 19024 19378
rect 18972 19314 19024 19320
rect 18788 19168 18840 19174
rect 18788 19110 18840 19116
rect 18694 18864 18750 18873
rect 18694 18799 18750 18808
rect 18800 18766 18828 19110
rect 18880 18896 18932 18902
rect 18880 18838 18932 18844
rect 18892 18766 18920 18838
rect 18788 18760 18840 18766
rect 18788 18702 18840 18708
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18984 18748 19012 19314
rect 19076 18970 19104 19926
rect 19536 19904 19564 20216
rect 19616 20198 19668 20204
rect 19628 20097 19656 20198
rect 19614 20088 19670 20097
rect 19614 20023 19670 20032
rect 19628 19922 19656 20023
rect 19352 19876 19564 19904
rect 19616 19916 19668 19922
rect 19154 19680 19210 19689
rect 19154 19615 19210 19624
rect 19168 19514 19196 19615
rect 19156 19508 19208 19514
rect 19156 19450 19208 19456
rect 19248 19508 19300 19514
rect 19248 19450 19300 19456
rect 19260 19281 19288 19450
rect 19246 19272 19302 19281
rect 19352 19242 19380 19876
rect 19616 19858 19668 19864
rect 19614 19816 19670 19825
rect 19432 19780 19484 19786
rect 19614 19751 19670 19760
rect 19432 19722 19484 19728
rect 19444 19417 19472 19722
rect 19628 19718 19656 19751
rect 19616 19712 19668 19718
rect 19616 19654 19668 19660
rect 19430 19408 19486 19417
rect 19430 19343 19486 19352
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19246 19207 19302 19216
rect 19340 19236 19392 19242
rect 19340 19178 19392 19184
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19064 18964 19116 18970
rect 19064 18906 19116 18912
rect 19430 18864 19486 18873
rect 19430 18799 19486 18808
rect 19064 18760 19116 18766
rect 18984 18720 19064 18748
rect 18696 18624 18748 18630
rect 18696 18566 18748 18572
rect 18708 18290 18736 18566
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 18708 17678 18736 18226
rect 18788 18216 18840 18222
rect 18788 18158 18840 18164
rect 18800 18086 18828 18158
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18696 17672 18748 17678
rect 18696 17614 18748 17620
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 18604 16720 18656 16726
rect 18604 16662 18656 16668
rect 18420 16448 18472 16454
rect 18420 16390 18472 16396
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18248 15502 18276 16186
rect 18328 16176 18380 16182
rect 18326 16144 18328 16153
rect 18380 16144 18382 16153
rect 18326 16079 18382 16088
rect 18328 15972 18380 15978
rect 18328 15914 18380 15920
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18236 15020 18288 15026
rect 18236 14962 18288 14968
rect 18248 14618 18276 14962
rect 18236 14612 18288 14618
rect 18236 14554 18288 14560
rect 18156 13484 18276 13512
rect 18052 13466 18104 13472
rect 18144 13388 18196 13394
rect 18144 13330 18196 13336
rect 18156 12918 18184 13330
rect 18144 12912 18196 12918
rect 18144 12854 18196 12860
rect 17972 12406 18092 12434
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17972 11218 18000 11698
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17868 10668 17920 10674
rect 17868 10610 17920 10616
rect 17880 9722 17908 10610
rect 17972 10606 18000 11154
rect 18064 11098 18092 12406
rect 18156 12102 18184 12854
rect 18248 12617 18276 13484
rect 18234 12608 18290 12617
rect 18234 12543 18290 12552
rect 18236 12164 18288 12170
rect 18236 12106 18288 12112
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18248 11898 18276 12106
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18248 11694 18276 11834
rect 18236 11688 18288 11694
rect 18236 11630 18288 11636
rect 18064 11070 18184 11098
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 10810 18092 10950
rect 18052 10804 18104 10810
rect 18052 10746 18104 10752
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17868 9716 17920 9722
rect 17696 9646 17816 9674
rect 17868 9658 17920 9664
rect 17316 9590 17368 9596
rect 17406 9616 17462 9625
rect 17224 9512 17276 9518
rect 17224 9454 17276 9460
rect 17236 9382 17264 9454
rect 17328 9450 17356 9590
rect 17788 9602 17816 9646
rect 17406 9551 17462 9560
rect 17512 9586 17724 9602
rect 17512 9580 17736 9586
rect 17512 9574 17684 9580
rect 17316 9444 17368 9450
rect 17316 9386 17368 9392
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17328 9178 17356 9386
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17316 9172 17368 9178
rect 17316 9114 17368 9120
rect 17040 9104 17092 9110
rect 17040 9046 17092 9052
rect 17328 9058 17356 9114
rect 17224 9036 17276 9042
rect 17328 9030 17448 9058
rect 17224 8978 17276 8984
rect 17040 8832 17092 8838
rect 17040 8774 17092 8780
rect 17052 8634 17080 8774
rect 17040 8628 17092 8634
rect 17040 8570 17092 8576
rect 17040 8492 17092 8498
rect 17040 8434 17092 8440
rect 16856 8366 16908 8372
rect 16946 8392 17002 8401
rect 16868 7886 16896 8366
rect 16946 8327 17002 8336
rect 16856 7880 16908 7886
rect 16856 7822 16908 7828
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 16580 7472 16632 7478
rect 16580 7414 16632 7420
rect 16960 7426 16988 7754
rect 17052 7546 17080 8434
rect 17236 8430 17264 8978
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17224 8424 17276 8430
rect 17224 8366 17276 8372
rect 17328 7954 17356 8434
rect 17316 7948 17368 7954
rect 17316 7890 17368 7896
rect 17420 7886 17448 9030
rect 17512 8838 17540 9574
rect 17788 9574 17908 9602
rect 17684 9522 17736 9528
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17592 8900 17644 8906
rect 17592 8842 17644 8848
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17408 7880 17460 7886
rect 17408 7822 17460 7828
rect 17222 7576 17278 7585
rect 17040 7540 17092 7546
rect 17222 7511 17278 7520
rect 17040 7482 17092 7488
rect 17130 7440 17186 7449
rect 16592 7206 16620 7414
rect 16672 7404 16724 7410
rect 16960 7398 17080 7426
rect 16672 7346 16724 7352
rect 16488 7200 16540 7206
rect 16488 7142 16540 7148
rect 16580 7200 16632 7206
rect 16684 7177 16712 7346
rect 16580 7142 16632 7148
rect 16670 7168 16726 7177
rect 16500 6934 16528 7142
rect 16670 7103 16726 7112
rect 16488 6928 16540 6934
rect 16488 6870 16540 6876
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16408 6344 16528 6372
rect 16500 6254 16528 6344
rect 16578 6352 16634 6361
rect 16578 6287 16580 6296
rect 16632 6287 16634 6296
rect 16580 6258 16632 6264
rect 16488 6248 16540 6254
rect 16488 6190 16540 6196
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 5568 16356 5574
rect 16304 5510 16356 5516
rect 16316 5166 16344 5510
rect 16304 5160 16356 5166
rect 16304 5102 16356 5108
rect 16302 3496 16358 3505
rect 16302 3431 16358 3440
rect 16316 3398 16344 3431
rect 16304 3392 16356 3398
rect 16304 3334 16356 3340
rect 16212 3052 16264 3058
rect 16212 2994 16264 3000
rect 16408 2496 16436 6054
rect 16960 5778 16988 6802
rect 17052 6610 17080 7398
rect 17236 7410 17264 7511
rect 17130 7375 17186 7384
rect 17224 7404 17276 7410
rect 17144 6866 17172 7375
rect 17224 7346 17276 7352
rect 17316 7268 17368 7274
rect 17316 7210 17368 7216
rect 17408 7268 17460 7274
rect 17408 7210 17460 7216
rect 17224 6928 17276 6934
rect 17224 6870 17276 6876
rect 17132 6860 17184 6866
rect 17132 6802 17184 6808
rect 17052 6582 17172 6610
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 16948 5772 17000 5778
rect 16948 5714 17000 5720
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 16488 5160 16540 5166
rect 16488 5102 16540 5108
rect 16500 4622 16528 5102
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 16580 4004 16632 4010
rect 16580 3946 16632 3952
rect 16592 3602 16620 3946
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 16960 3058 16988 4422
rect 17052 3942 17080 6258
rect 17040 3936 17092 3942
rect 17040 3878 17092 3884
rect 16948 3052 17000 3058
rect 16948 2994 17000 3000
rect 16672 2848 16724 2854
rect 16672 2790 16724 2796
rect 16684 2514 16712 2790
rect 16948 2576 17000 2582
rect 16948 2518 17000 2524
rect 16316 2468 16436 2496
rect 16672 2508 16724 2514
rect 16212 2440 16264 2446
rect 16212 2382 16264 2388
rect 16224 2009 16252 2382
rect 16316 2106 16344 2468
rect 16672 2450 16724 2456
rect 16396 2372 16448 2378
rect 16396 2314 16448 2320
rect 16304 2100 16356 2106
rect 16304 2042 16356 2048
rect 16210 2000 16266 2009
rect 16210 1935 16266 1944
rect 16120 1896 16172 1902
rect 16120 1838 16172 1844
rect 16408 1170 16436 2314
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 16960 1170 16988 2518
rect 17144 1358 17172 6582
rect 17236 6322 17264 6870
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17236 5166 17264 6258
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 17236 4146 17264 4762
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17328 3058 17356 7210
rect 17420 7041 17448 7210
rect 17406 7032 17462 7041
rect 17406 6967 17462 6976
rect 17512 6730 17540 8774
rect 17604 7410 17632 8842
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17500 6724 17552 6730
rect 17500 6666 17552 6672
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 5370 17448 6598
rect 17408 5364 17460 5370
rect 17408 5306 17460 5312
rect 17512 5030 17540 6666
rect 17500 5024 17552 5030
rect 17500 4966 17552 4972
rect 17406 4856 17462 4865
rect 17406 4791 17462 4800
rect 17420 4758 17448 4791
rect 17408 4752 17460 4758
rect 17408 4694 17460 4700
rect 17500 4548 17552 4554
rect 17500 4490 17552 4496
rect 17408 4480 17460 4486
rect 17408 4422 17460 4428
rect 17420 3534 17448 4422
rect 17512 4214 17540 4490
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17604 3058 17632 7346
rect 17696 5642 17724 9318
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17788 7478 17816 9046
rect 17880 8242 17908 9574
rect 18064 8974 18092 9998
rect 18052 8968 18104 8974
rect 18052 8910 18104 8916
rect 17960 8628 18012 8634
rect 17960 8570 18012 8576
rect 17972 8401 18000 8570
rect 17958 8392 18014 8401
rect 17958 8327 18014 8336
rect 17880 8214 18000 8242
rect 17972 7546 18000 8214
rect 18064 8090 18092 8910
rect 18052 8084 18104 8090
rect 18052 8026 18104 8032
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17788 6361 17816 7414
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 17774 6352 17830 6361
rect 17774 6287 17830 6296
rect 17776 6180 17828 6186
rect 17776 6122 17828 6128
rect 17788 5710 17816 6122
rect 17776 5704 17828 5710
rect 17880 5681 17908 7142
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17958 6896 18014 6905
rect 17958 6831 18014 6840
rect 17972 6798 18000 6831
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18064 6644 18092 6938
rect 18156 6934 18184 11070
rect 18236 10532 18288 10538
rect 18236 10474 18288 10480
rect 18248 9926 18276 10474
rect 18236 9920 18288 9926
rect 18236 9862 18288 9868
rect 18248 9518 18276 9862
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18234 9344 18290 9353
rect 18234 9279 18290 9288
rect 18248 8498 18276 9279
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 7857 18276 8434
rect 18234 7848 18290 7857
rect 18234 7783 18290 7792
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 7002 18276 7686
rect 18236 6996 18288 7002
rect 18236 6938 18288 6944
rect 18144 6928 18196 6934
rect 18144 6870 18196 6876
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 17972 6616 18092 6644
rect 18144 6656 18196 6662
rect 17776 5646 17828 5652
rect 17866 5672 17922 5681
rect 17684 5636 17736 5642
rect 17866 5607 17922 5616
rect 17684 5578 17736 5584
rect 17696 5234 17724 5578
rect 17868 5568 17920 5574
rect 17868 5510 17920 5516
rect 17972 5522 18000 6616
rect 18144 6598 18196 6604
rect 18156 6458 18184 6598
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18144 6316 18196 6322
rect 18144 6258 18196 6264
rect 18050 5808 18106 5817
rect 18050 5743 18106 5752
rect 18064 5642 18092 5743
rect 18052 5636 18104 5642
rect 18052 5578 18104 5584
rect 17880 5370 17908 5510
rect 17972 5494 18092 5522
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17592 3052 17644 3058
rect 17592 2994 17644 3000
rect 17224 2848 17276 2854
rect 17224 2790 17276 2796
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 17236 1494 17264 2790
rect 17224 1488 17276 1494
rect 17224 1430 17276 1436
rect 17132 1352 17184 1358
rect 17132 1294 17184 1300
rect 16408 1142 16528 1170
rect 16500 800 16528 1142
rect 16868 1142 16988 1170
rect 16868 800 16896 1142
rect 17328 800 17356 2790
rect 17696 2774 17724 5170
rect 17960 4548 18012 4554
rect 17960 4490 18012 4496
rect 17972 3670 18000 4490
rect 18064 4214 18092 5494
rect 18156 5098 18184 6258
rect 18248 5778 18276 6802
rect 18340 6338 18368 15914
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18420 15564 18472 15570
rect 18420 15506 18472 15512
rect 18432 15026 18460 15506
rect 18524 15337 18552 15846
rect 18708 15450 18736 16730
rect 18616 15422 18736 15450
rect 18510 15328 18566 15337
rect 18510 15263 18566 15272
rect 18420 15020 18472 15026
rect 18420 14962 18472 14968
rect 18616 14362 18644 15422
rect 18696 15360 18748 15366
rect 18696 15302 18748 15308
rect 18708 14929 18736 15302
rect 18694 14920 18750 14929
rect 18694 14855 18750 14864
rect 18800 14414 18828 18022
rect 18892 17270 18920 18702
rect 18984 18193 19012 18720
rect 19064 18702 19116 18708
rect 19064 18284 19116 18290
rect 19064 18226 19116 18232
rect 18970 18184 19026 18193
rect 18970 18119 19026 18128
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18880 17264 18932 17270
rect 18880 17206 18932 17212
rect 18878 16552 18934 16561
rect 18878 16487 18934 16496
rect 18892 16454 18920 16487
rect 18880 16448 18932 16454
rect 18880 16390 18932 16396
rect 18892 15162 18920 16390
rect 18984 15706 19012 18022
rect 19076 17882 19104 18226
rect 19444 18068 19472 18799
rect 19536 18426 19564 19314
rect 19524 18420 19576 18426
rect 19524 18362 19576 18368
rect 19524 18080 19576 18086
rect 19444 18040 19524 18068
rect 19524 18022 19576 18028
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 19064 17876 19116 17882
rect 19064 17818 19116 17824
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19076 17134 19104 17614
rect 19536 17202 19564 18022
rect 19628 17882 19656 19314
rect 19720 18902 19748 21791
rect 19800 20596 19852 20602
rect 19800 20538 19852 20544
rect 19812 19310 19840 20538
rect 19800 19304 19852 19310
rect 19800 19246 19852 19252
rect 19708 18896 19760 18902
rect 19708 18838 19760 18844
rect 19812 18358 19840 19246
rect 19904 18902 19932 21950
rect 19984 20596 20036 20602
rect 19984 20538 20036 20544
rect 19996 18970 20024 20538
rect 19984 18964 20036 18970
rect 19984 18906 20036 18912
rect 19892 18896 19944 18902
rect 19892 18838 19944 18844
rect 19892 18760 19944 18766
rect 19892 18702 19944 18708
rect 19800 18352 19852 18358
rect 19800 18294 19852 18300
rect 19616 17876 19668 17882
rect 19616 17818 19668 17824
rect 19616 17740 19668 17746
rect 19616 17682 19668 17688
rect 19628 17338 19656 17682
rect 19708 17672 19760 17678
rect 19708 17614 19760 17620
rect 19800 17672 19852 17678
rect 19800 17614 19852 17620
rect 19616 17332 19668 17338
rect 19616 17274 19668 17280
rect 19432 17196 19484 17202
rect 19432 17138 19484 17144
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 19064 17128 19116 17134
rect 19064 17070 19116 17076
rect 19444 16980 19472 17138
rect 19616 16992 19668 16998
rect 19444 16952 19564 16980
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 19154 16552 19210 16561
rect 19154 16487 19210 16496
rect 19168 16250 19196 16487
rect 19156 16244 19208 16250
rect 19156 16186 19208 16192
rect 19536 16153 19564 16952
rect 19720 16980 19748 17614
rect 19812 16998 19840 17614
rect 19904 17338 19932 18702
rect 20088 17882 20116 22200
rect 20456 21264 20484 22200
rect 20272 21236 20484 21264
rect 20168 20324 20220 20330
rect 20168 20266 20220 20272
rect 20180 19553 20208 20266
rect 20166 19544 20222 19553
rect 20166 19479 20222 19488
rect 20272 18290 20300 21236
rect 20548 21162 20576 22607
rect 20902 22200 20958 23000
rect 21270 22200 21326 23000
rect 21638 22200 21694 23000
rect 22006 22200 22062 23000
rect 22374 22200 22430 23000
rect 22742 22200 22798 23000
rect 20626 21448 20682 21457
rect 20626 21383 20682 21392
rect 20456 21134 20576 21162
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20364 20058 20392 20402
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20352 19848 20404 19854
rect 20350 19816 20352 19825
rect 20404 19816 20406 19825
rect 20350 19751 20406 19760
rect 20352 19236 20404 19242
rect 20352 19178 20404 19184
rect 20364 18766 20392 19178
rect 20456 18970 20484 21134
rect 20534 21040 20590 21049
rect 20534 20975 20590 20984
rect 20548 20602 20576 20975
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 20640 20482 20668 21383
rect 20916 20602 20944 22200
rect 20994 20632 21050 20641
rect 20904 20596 20956 20602
rect 20994 20567 21050 20576
rect 20904 20538 20956 20544
rect 20548 20454 20668 20482
rect 20810 20496 20866 20505
rect 20548 20058 20576 20454
rect 20810 20431 20866 20440
rect 20718 20088 20774 20097
rect 20536 20052 20588 20058
rect 20718 20023 20774 20032
rect 20536 19994 20588 20000
rect 20536 19916 20588 19922
rect 20536 19858 20588 19864
rect 20548 19825 20576 19858
rect 20732 19854 20760 20023
rect 20824 19922 20852 20431
rect 20812 19916 20864 19922
rect 20812 19858 20864 19864
rect 20720 19848 20772 19854
rect 20534 19816 20590 19825
rect 20720 19790 20772 19796
rect 20534 19751 20590 19760
rect 20916 19446 20944 20538
rect 21008 20330 21036 20567
rect 20996 20324 21048 20330
rect 20996 20266 21048 20272
rect 21088 20256 21140 20262
rect 21088 20198 21140 20204
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20444 18964 20496 18970
rect 20444 18906 20496 18912
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20352 18760 20404 18766
rect 20352 18702 20404 18708
rect 20260 18284 20312 18290
rect 20260 18226 20312 18232
rect 20456 17882 20484 18770
rect 20720 18760 20772 18766
rect 20720 18702 20772 18708
rect 20732 18426 20760 18702
rect 20812 18692 20864 18698
rect 20812 18634 20864 18640
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20076 17876 20128 17882
rect 20076 17818 20128 17824
rect 20444 17876 20496 17882
rect 20444 17818 20496 17824
rect 20074 17776 20130 17785
rect 20074 17711 20130 17720
rect 20088 17678 20116 17711
rect 20732 17678 20760 18362
rect 20076 17672 20128 17678
rect 19996 17620 20076 17626
rect 19996 17614 20128 17620
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20720 17672 20772 17678
rect 20720 17614 20772 17620
rect 19996 17598 20116 17614
rect 19892 17332 19944 17338
rect 19892 17274 19944 17280
rect 19668 16952 19748 16980
rect 19616 16934 19668 16940
rect 19522 16144 19578 16153
rect 19522 16079 19578 16088
rect 19062 16008 19118 16017
rect 19062 15943 19118 15952
rect 19614 16008 19670 16017
rect 19614 15943 19616 15952
rect 19076 15706 19104 15943
rect 19668 15943 19670 15952
rect 19616 15914 19668 15920
rect 19524 15904 19576 15910
rect 19524 15846 19576 15852
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 18972 15700 19024 15706
rect 18972 15642 19024 15648
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 19352 15094 19380 15438
rect 19340 15088 19392 15094
rect 19340 15030 19392 15036
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18984 14550 19012 14962
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 18972 14544 19024 14550
rect 18972 14486 19024 14492
rect 19156 14544 19208 14550
rect 19156 14486 19208 14492
rect 18524 14334 18644 14362
rect 18788 14408 18840 14414
rect 18788 14350 18840 14356
rect 18420 14000 18472 14006
rect 18420 13942 18472 13948
rect 18432 13530 18460 13942
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18524 13297 18552 14334
rect 18604 14272 18656 14278
rect 18604 14214 18656 14220
rect 18510 13288 18566 13297
rect 18510 13223 18566 13232
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18512 13184 18564 13190
rect 18512 13126 18564 13132
rect 18432 12889 18460 13126
rect 18418 12880 18474 12889
rect 18418 12815 18474 12824
rect 18524 11898 18552 13126
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18512 11756 18564 11762
rect 18512 11698 18564 11704
rect 18420 11688 18472 11694
rect 18420 11630 18472 11636
rect 18432 11354 18460 11630
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18524 10810 18552 11698
rect 18512 10804 18564 10810
rect 18512 10746 18564 10752
rect 18420 8832 18472 8838
rect 18420 8774 18472 8780
rect 18432 6866 18460 8774
rect 18512 8560 18564 8566
rect 18510 8528 18512 8537
rect 18564 8528 18566 8537
rect 18510 8463 18566 8472
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18524 7818 18552 8366
rect 18512 7812 18564 7818
rect 18512 7754 18564 7760
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18524 7177 18552 7346
rect 18510 7168 18566 7177
rect 18510 7103 18566 7112
rect 18420 6860 18472 6866
rect 18420 6802 18472 6808
rect 18512 6792 18564 6798
rect 18510 6760 18512 6769
rect 18564 6760 18566 6769
rect 18510 6695 18566 6704
rect 18512 6656 18564 6662
rect 18512 6598 18564 6604
rect 18524 6390 18552 6598
rect 18512 6384 18564 6390
rect 18340 6310 18460 6338
rect 18512 6326 18564 6332
rect 18328 6248 18380 6254
rect 18328 6190 18380 6196
rect 18236 5772 18288 5778
rect 18236 5714 18288 5720
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18144 5092 18196 5098
rect 18144 5034 18196 5040
rect 18248 4486 18276 5170
rect 18340 4826 18368 6190
rect 18432 5817 18460 6310
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18524 5914 18552 6190
rect 18616 6186 18644 14214
rect 18694 13968 18750 13977
rect 18694 13903 18750 13912
rect 18880 13932 18932 13938
rect 18708 13002 18736 13903
rect 18880 13874 18932 13880
rect 18708 12974 18828 13002
rect 18696 12912 18748 12918
rect 18696 12854 18748 12860
rect 18708 9586 18736 12854
rect 18800 11529 18828 12974
rect 18892 12442 18920 13874
rect 19168 13870 19196 14486
rect 19432 14408 19484 14414
rect 19536 14385 19564 15846
rect 19616 15564 19668 15570
rect 19616 15506 19668 15512
rect 19432 14350 19484 14356
rect 19522 14376 19578 14385
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19352 14074 19380 14282
rect 19340 14068 19392 14074
rect 19340 14010 19392 14016
rect 18972 13864 19024 13870
rect 19156 13864 19208 13870
rect 18972 13806 19024 13812
rect 19076 13824 19156 13852
rect 18984 13462 19012 13806
rect 18972 13456 19024 13462
rect 18972 13398 19024 13404
rect 19076 13394 19104 13824
rect 19156 13806 19208 13812
rect 19444 13716 19472 14350
rect 19522 14311 19578 14320
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19536 14006 19564 14214
rect 19628 14006 19656 15506
rect 19720 14482 19748 16952
rect 19800 16992 19852 16998
rect 19800 16934 19852 16940
rect 19890 16688 19946 16697
rect 19996 16658 20024 17598
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 19890 16623 19946 16632
rect 19984 16652 20036 16658
rect 19904 16590 19932 16623
rect 19984 16594 20036 16600
rect 19892 16584 19944 16590
rect 19892 16526 19944 16532
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19800 16040 19852 16046
rect 19800 15982 19852 15988
rect 19812 15570 19840 15982
rect 19904 15638 19932 16186
rect 19996 15706 20024 16594
rect 19984 15700 20036 15706
rect 19984 15642 20036 15648
rect 19892 15632 19944 15638
rect 19892 15574 19944 15580
rect 19800 15564 19852 15570
rect 19800 15506 19852 15512
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19800 14952 19852 14958
rect 19800 14894 19852 14900
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19812 14414 19840 14894
rect 19892 14816 19944 14822
rect 19892 14758 19944 14764
rect 19800 14408 19852 14414
rect 19800 14350 19852 14356
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19720 14074 19748 14214
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19524 14000 19576 14006
rect 19524 13942 19576 13948
rect 19616 14000 19668 14006
rect 19616 13942 19668 13948
rect 19904 13870 19932 14758
rect 19996 14618 20024 14962
rect 19984 14612 20036 14618
rect 19984 14554 20036 14560
rect 20088 14498 20116 16934
rect 20180 16794 20208 16934
rect 20168 16788 20220 16794
rect 20168 16730 20220 16736
rect 20260 16720 20312 16726
rect 20260 16662 20312 16668
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20180 16289 20208 16458
rect 20166 16280 20222 16289
rect 20166 16215 20222 16224
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20180 15706 20208 16050
rect 20272 15706 20300 16662
rect 20364 16250 20392 17614
rect 20536 17536 20588 17542
rect 20536 17478 20588 17484
rect 20548 17241 20576 17478
rect 20824 17338 20852 18634
rect 20904 17604 20956 17610
rect 20904 17546 20956 17552
rect 20812 17332 20864 17338
rect 20812 17274 20864 17280
rect 20534 17232 20590 17241
rect 20534 17167 20590 17176
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20352 16244 20404 16250
rect 20352 16186 20404 16192
rect 20350 16008 20406 16017
rect 20350 15943 20352 15952
rect 20404 15943 20406 15952
rect 20352 15914 20404 15920
rect 20536 15904 20588 15910
rect 20442 15872 20498 15881
rect 20536 15846 20588 15852
rect 20442 15807 20498 15816
rect 20168 15700 20220 15706
rect 20168 15642 20220 15648
rect 20260 15700 20312 15706
rect 20260 15642 20312 15648
rect 20456 15026 20484 15807
rect 20548 15502 20576 15846
rect 20536 15496 20588 15502
rect 20536 15438 20588 15444
rect 20444 15020 20496 15026
rect 19996 14470 20116 14498
rect 20364 14980 20444 15008
rect 19892 13864 19944 13870
rect 19892 13806 19944 13812
rect 19444 13688 19840 13716
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19522 13560 19578 13569
rect 19522 13495 19578 13504
rect 19536 13462 19564 13495
rect 19524 13456 19576 13462
rect 19616 13456 19668 13462
rect 19524 13398 19576 13404
rect 19614 13424 19616 13433
rect 19668 13424 19670 13433
rect 19064 13388 19116 13394
rect 19614 13359 19670 13368
rect 19064 13330 19116 13336
rect 18972 12708 19024 12714
rect 18972 12650 19024 12656
rect 18880 12436 18932 12442
rect 18880 12378 18932 12384
rect 18786 11520 18842 11529
rect 18786 11455 18842 11464
rect 18788 11008 18840 11014
rect 18788 10950 18840 10956
rect 18800 10130 18828 10950
rect 18984 10690 19012 12650
rect 19076 12646 19104 13330
rect 19524 13252 19576 13258
rect 19524 13194 19576 13200
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19536 12434 19564 13194
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19444 12406 19564 12434
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11694 19196 12038
rect 19260 11694 19288 12242
rect 19444 12073 19472 12406
rect 19614 12200 19670 12209
rect 19720 12170 19748 12582
rect 19614 12135 19616 12144
rect 19668 12135 19670 12144
rect 19708 12164 19760 12170
rect 19616 12106 19668 12112
rect 19708 12106 19760 12112
rect 19812 12073 19840 13688
rect 19892 13184 19944 13190
rect 19996 13172 20024 14470
rect 20168 14340 20220 14346
rect 20168 14282 20220 14288
rect 20076 13864 20128 13870
rect 20074 13832 20076 13841
rect 20128 13832 20130 13841
rect 20074 13767 20130 13776
rect 20076 13184 20128 13190
rect 19996 13152 20076 13172
rect 20128 13152 20130 13161
rect 19996 13144 20074 13152
rect 19892 13126 19944 13132
rect 19430 12064 19486 12073
rect 19430 11999 19486 12008
rect 19798 12064 19854 12073
rect 19798 11999 19854 12008
rect 19338 11928 19394 11937
rect 19706 11928 19762 11937
rect 19338 11863 19340 11872
rect 19392 11863 19394 11872
rect 19524 11892 19576 11898
rect 19340 11834 19392 11840
rect 19706 11863 19762 11872
rect 19524 11834 19576 11840
rect 19156 11688 19208 11694
rect 19156 11630 19208 11636
rect 19248 11688 19300 11694
rect 19248 11630 19300 11636
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19536 11370 19564 11834
rect 19527 11342 19564 11370
rect 19527 11336 19555 11342
rect 19444 11308 19555 11336
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 19352 10996 19380 11086
rect 18892 10662 19012 10690
rect 19076 10968 19380 10996
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18800 9518 18828 10066
rect 18788 9512 18840 9518
rect 18788 9454 18840 9460
rect 18696 9104 18748 9110
rect 18696 9046 18748 9052
rect 18604 6180 18656 6186
rect 18604 6122 18656 6128
rect 18602 6080 18658 6089
rect 18602 6015 18658 6024
rect 18512 5908 18564 5914
rect 18512 5850 18564 5856
rect 18418 5808 18474 5817
rect 18616 5794 18644 6015
rect 18418 5743 18474 5752
rect 18524 5766 18644 5794
rect 18432 4826 18460 5743
rect 18524 5114 18552 5766
rect 18604 5636 18656 5642
rect 18604 5578 18656 5584
rect 18616 5273 18644 5578
rect 18602 5264 18658 5273
rect 18602 5199 18658 5208
rect 18524 5086 18644 5114
rect 18328 4820 18380 4826
rect 18328 4762 18380 4768
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18326 4720 18382 4729
rect 18326 4655 18382 4664
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18052 4208 18104 4214
rect 18052 4150 18104 4156
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 17960 3664 18012 3670
rect 17960 3606 18012 3612
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 17788 2990 17816 3470
rect 17960 3460 18012 3466
rect 17960 3402 18012 3408
rect 17972 3369 18000 3402
rect 17958 3360 18014 3369
rect 17958 3295 18014 3304
rect 18052 3120 18104 3126
rect 17972 3080 18052 3108
rect 17776 2984 17828 2990
rect 17828 2944 17908 2972
rect 17776 2926 17828 2932
rect 17880 2825 17908 2944
rect 17866 2816 17922 2825
rect 17696 2746 17816 2774
rect 17866 2751 17922 2760
rect 17788 2038 17816 2746
rect 17776 2032 17828 2038
rect 17776 1974 17828 1980
rect 17684 1420 17736 1426
rect 17684 1362 17736 1368
rect 17696 800 17724 1362
rect 17972 1018 18000 3080
rect 18052 3062 18104 3068
rect 18248 3058 18276 3878
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18234 2816 18290 2825
rect 18234 2751 18290 2760
rect 18248 2514 18276 2751
rect 18340 2514 18368 4655
rect 18512 4140 18564 4146
rect 18512 4082 18564 4088
rect 18420 3392 18472 3398
rect 18420 3334 18472 3340
rect 18432 2650 18460 3334
rect 18524 3194 18552 4082
rect 18616 3534 18644 5086
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18708 3233 18736 9046
rect 18800 9042 18828 9454
rect 18788 9036 18840 9042
rect 18788 8978 18840 8984
rect 18892 7449 18920 10662
rect 18972 10600 19024 10606
rect 18972 10542 19024 10548
rect 18984 10198 19012 10542
rect 18972 10192 19024 10198
rect 18972 10134 19024 10140
rect 18984 10033 19012 10134
rect 18970 10024 19026 10033
rect 18970 9959 19026 9968
rect 19076 9874 19104 10968
rect 19444 10588 19472 11308
rect 19720 11286 19748 11863
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19524 11212 19576 11218
rect 19524 11154 19576 11160
rect 19536 10810 19564 11154
rect 19616 11008 19668 11014
rect 19616 10950 19668 10956
rect 19524 10804 19576 10810
rect 19524 10746 19576 10752
rect 19444 10560 19564 10588
rect 19628 10577 19656 10950
rect 19708 10600 19760 10606
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19432 10056 19484 10062
rect 19430 10024 19432 10033
rect 19484 10024 19486 10033
rect 19430 9959 19486 9968
rect 18984 9846 19104 9874
rect 18984 9110 19012 9846
rect 19536 9722 19564 10560
rect 19614 10568 19670 10577
rect 19708 10542 19760 10548
rect 19614 10503 19670 10512
rect 19616 10464 19668 10470
rect 19616 10406 19668 10412
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19154 9616 19210 9625
rect 19064 9580 19116 9586
rect 19154 9551 19210 9560
rect 19524 9580 19576 9586
rect 19064 9522 19116 9528
rect 19076 9489 19104 9522
rect 19062 9480 19118 9489
rect 19168 9450 19196 9551
rect 19524 9522 19576 9528
rect 19062 9415 19118 9424
rect 19156 9444 19208 9450
rect 19156 9386 19208 9392
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19536 9178 19564 9522
rect 19524 9172 19576 9178
rect 19524 9114 19576 9120
rect 18972 9104 19024 9110
rect 18972 9046 19024 9052
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 18972 8832 19024 8838
rect 19024 8792 19104 8820
rect 18972 8774 19024 8780
rect 18972 8288 19024 8294
rect 18972 8230 19024 8236
rect 18984 8129 19012 8230
rect 18970 8120 19026 8129
rect 18970 8055 19026 8064
rect 18972 7812 19024 7818
rect 18972 7754 19024 7760
rect 18878 7440 18934 7449
rect 18878 7375 18934 7384
rect 18786 7304 18842 7313
rect 18786 7239 18842 7248
rect 18800 5846 18828 7239
rect 18892 7188 18920 7375
rect 18984 7342 19012 7754
rect 19076 7478 19104 8792
rect 19260 8634 19288 9007
rect 19248 8628 19300 8634
rect 19248 8570 19300 8576
rect 19536 8566 19564 9114
rect 19628 8673 19656 10406
rect 19720 10266 19748 10542
rect 19708 10260 19760 10266
rect 19708 10202 19760 10208
rect 19812 10198 19840 11698
rect 19904 11665 19932 13126
rect 20074 13087 20130 13096
rect 20180 12356 20208 14282
rect 20260 12640 20312 12646
rect 20260 12582 20312 12588
rect 20272 12481 20300 12582
rect 20258 12472 20314 12481
rect 20258 12407 20314 12416
rect 20088 12328 20208 12356
rect 19984 12300 20036 12306
rect 19984 12242 20036 12248
rect 19890 11656 19946 11665
rect 19890 11591 19946 11600
rect 19892 11552 19944 11558
rect 19892 11494 19944 11500
rect 19800 10192 19852 10198
rect 19706 10160 19762 10169
rect 19800 10134 19852 10140
rect 19706 10095 19708 10104
rect 19760 10095 19762 10104
rect 19708 10066 19760 10072
rect 19812 9761 19840 10134
rect 19904 10033 19932 11494
rect 19890 10024 19946 10033
rect 19890 9959 19946 9968
rect 19798 9752 19854 9761
rect 19798 9687 19854 9696
rect 19996 9674 20024 12242
rect 19904 9646 20024 9674
rect 19904 9081 19932 9646
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19890 9072 19946 9081
rect 19890 9007 19946 9016
rect 19892 8968 19944 8974
rect 19892 8910 19944 8916
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19614 8664 19670 8673
rect 19614 8599 19670 8608
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19616 8492 19668 8498
rect 19616 8434 19668 8440
rect 19524 8424 19576 8430
rect 19524 8366 19576 8372
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19536 8090 19564 8366
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19156 7744 19208 7750
rect 19156 7686 19208 7692
rect 19168 7546 19196 7686
rect 19246 7576 19302 7585
rect 19156 7540 19208 7546
rect 19628 7546 19656 8434
rect 19720 7954 19748 8774
rect 19812 8022 19840 8842
rect 19800 8016 19852 8022
rect 19800 7958 19852 7964
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19246 7511 19248 7520
rect 19156 7482 19208 7488
rect 19300 7511 19302 7520
rect 19616 7540 19668 7546
rect 19248 7482 19300 7488
rect 19616 7482 19668 7488
rect 19064 7472 19116 7478
rect 19064 7414 19116 7420
rect 19812 7342 19840 7958
rect 19904 7954 19932 8910
rect 19996 8634 20024 9522
rect 20088 9364 20116 12328
rect 20364 12288 20392 14980
rect 20444 14962 20496 14968
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20548 14278 20576 14418
rect 20536 14272 20588 14278
rect 20536 14214 20588 14220
rect 20442 13968 20498 13977
rect 20442 13903 20444 13912
rect 20496 13903 20498 13912
rect 20444 13874 20496 13880
rect 20548 13870 20576 14214
rect 20536 13864 20588 13870
rect 20536 13806 20588 13812
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20548 12442 20576 13262
rect 20640 12442 20668 16934
rect 20810 16688 20866 16697
rect 20810 16623 20866 16632
rect 20824 16590 20852 16623
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20732 15162 20760 15438
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20824 15026 20852 15302
rect 20812 15020 20864 15026
rect 20812 14962 20864 14968
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13530 20760 13874
rect 20720 13524 20772 13530
rect 20720 13466 20772 13472
rect 20720 12776 20772 12782
rect 20720 12718 20772 12724
rect 20732 12594 20760 12718
rect 20724 12566 20760 12594
rect 20536 12436 20588 12442
rect 20536 12378 20588 12384
rect 20628 12436 20680 12442
rect 20628 12378 20680 12384
rect 20724 12322 20752 12566
rect 20180 12260 20392 12288
rect 20640 12294 20752 12322
rect 20812 12368 20864 12374
rect 20812 12310 20864 12316
rect 20180 11354 20208 12260
rect 20260 12164 20312 12170
rect 20260 12106 20312 12112
rect 20352 12164 20404 12170
rect 20352 12106 20404 12112
rect 20168 11348 20220 11354
rect 20168 11290 20220 11296
rect 20272 11286 20300 12106
rect 20364 11898 20392 12106
rect 20536 12096 20588 12102
rect 20536 12038 20588 12044
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20352 11756 20404 11762
rect 20352 11698 20404 11704
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20364 11354 20392 11698
rect 20352 11348 20404 11354
rect 20352 11290 20404 11296
rect 20260 11280 20312 11286
rect 20260 11222 20312 11228
rect 20168 11212 20220 11218
rect 20168 11154 20220 11160
rect 20180 11121 20208 11154
rect 20166 11112 20222 11121
rect 20166 11047 20222 11056
rect 20352 11076 20404 11082
rect 20352 11018 20404 11024
rect 20364 10810 20392 11018
rect 20352 10804 20404 10810
rect 20352 10746 20404 10752
rect 20350 10704 20406 10713
rect 20350 10639 20406 10648
rect 20258 10568 20314 10577
rect 20258 10503 20314 10512
rect 20168 9376 20220 9382
rect 20088 9336 20168 9364
rect 20168 9318 20220 9324
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 8356 20128 8362
rect 20076 8298 20128 8304
rect 19892 7948 19944 7954
rect 19892 7890 19944 7896
rect 19984 7880 20036 7886
rect 19984 7822 20036 7828
rect 18972 7336 19024 7342
rect 18972 7278 19024 7284
rect 19064 7336 19116 7342
rect 19064 7278 19116 7284
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 18892 7160 19012 7188
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 18788 5840 18840 5846
rect 18788 5782 18840 5788
rect 18892 5778 18920 6734
rect 18984 6730 19012 7160
rect 18972 6724 19024 6730
rect 18972 6666 19024 6672
rect 19076 6458 19104 7278
rect 19708 7268 19760 7274
rect 19708 7210 19760 7216
rect 19616 7200 19668 7206
rect 19616 7142 19668 7148
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 19156 6792 19208 6798
rect 19156 6734 19208 6740
rect 19064 6452 19116 6458
rect 19064 6394 19116 6400
rect 18970 6352 19026 6361
rect 18970 6287 19026 6296
rect 18984 6186 19012 6287
rect 19168 6202 19196 6734
rect 19260 6474 19288 6870
rect 19260 6446 19564 6474
rect 19628 6458 19656 7142
rect 19536 6338 19564 6446
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19432 6316 19484 6322
rect 19536 6310 19656 6338
rect 19432 6258 19484 6264
rect 19444 6225 19472 6258
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19076 6174 19196 6202
rect 19430 6216 19486 6225
rect 18880 5772 18932 5778
rect 18880 5714 18932 5720
rect 18892 5302 18920 5714
rect 18880 5296 18932 5302
rect 18880 5238 18932 5244
rect 18972 5228 19024 5234
rect 18972 5170 19024 5176
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18892 4282 18920 4490
rect 18984 4486 19012 5170
rect 19076 4826 19104 6174
rect 19430 6151 19486 6160
rect 19522 6080 19578 6089
rect 19143 6012 19451 6032
rect 19522 6015 19578 6024
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 19536 5794 19564 6015
rect 19352 5766 19564 5794
rect 19352 5710 19380 5766
rect 19340 5704 19392 5710
rect 19340 5646 19392 5652
rect 19522 5672 19578 5681
rect 19522 5607 19578 5616
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 19064 4820 19116 4826
rect 19064 4762 19116 4768
rect 19338 4720 19394 4729
rect 19338 4655 19394 4664
rect 18972 4480 19024 4486
rect 18972 4422 19024 4428
rect 18880 4276 18932 4282
rect 18880 4218 18932 4224
rect 18984 4078 19012 4422
rect 19352 4078 19380 4655
rect 18788 4072 18840 4078
rect 18788 4014 18840 4020
rect 18972 4072 19024 4078
rect 18972 4014 19024 4020
rect 19340 4072 19392 4078
rect 19340 4014 19392 4020
rect 18800 3738 18828 4014
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18788 3392 18840 3398
rect 18788 3334 18840 3340
rect 18694 3224 18750 3233
rect 18512 3188 18564 3194
rect 18694 3159 18750 3168
rect 18512 3130 18564 3136
rect 18512 2848 18564 2854
rect 18512 2790 18564 2796
rect 18604 2848 18656 2854
rect 18800 2836 18828 3334
rect 18880 3188 18932 3194
rect 18984 3176 19012 3878
rect 19076 3738 19104 3878
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19064 3732 19116 3738
rect 19064 3674 19116 3680
rect 19536 3670 19564 5607
rect 19628 5386 19656 6310
rect 19720 6202 19748 7210
rect 19812 6322 19840 7278
rect 19996 7206 20024 7822
rect 20088 7546 20116 8298
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19984 6724 20036 6730
rect 19984 6666 20036 6672
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19904 6254 19932 6666
rect 19892 6248 19944 6254
rect 19720 6174 19840 6202
rect 19892 6190 19944 6196
rect 19628 5358 19748 5386
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19628 4282 19656 4422
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19628 3738 19656 4014
rect 19720 3777 19748 5358
rect 19706 3768 19762 3777
rect 19616 3732 19668 3738
rect 19706 3703 19762 3712
rect 19616 3674 19668 3680
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19156 3528 19208 3534
rect 19156 3470 19208 3476
rect 18984 3148 19104 3176
rect 18880 3130 18932 3136
rect 18604 2790 18656 2796
rect 18708 2808 18828 2836
rect 18420 2644 18472 2650
rect 18420 2586 18472 2592
rect 18418 2544 18474 2553
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18328 2508 18380 2514
rect 18418 2479 18474 2488
rect 18328 2450 18380 2456
rect 18432 2446 18460 2479
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 18144 1488 18196 1494
rect 18144 1430 18196 1436
rect 17960 1012 18012 1018
rect 17960 954 18012 960
rect 18156 800 18184 1430
rect 18524 1290 18552 2790
rect 18512 1284 18564 1290
rect 18512 1226 18564 1232
rect 18616 800 18644 2790
rect 18708 2310 18736 2808
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 18696 1352 18748 1358
rect 18696 1294 18748 1300
rect 18892 1306 18920 3130
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 18984 2825 19012 2994
rect 19076 2922 19104 3148
rect 19168 2990 19196 3470
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19156 2984 19208 2990
rect 19156 2926 19208 2932
rect 19064 2916 19116 2922
rect 19064 2858 19116 2864
rect 18970 2816 19026 2825
rect 18970 2751 19026 2760
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19064 2440 19116 2446
rect 19064 2382 19116 2388
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 18972 2304 19024 2310
rect 18972 2246 19024 2252
rect 18984 1426 19012 2246
rect 19076 1834 19104 2382
rect 19260 2106 19288 2382
rect 19248 2100 19300 2106
rect 19248 2042 19300 2048
rect 19248 1896 19300 1902
rect 19248 1838 19300 1844
rect 19064 1828 19116 1834
rect 19064 1770 19116 1776
rect 19260 1465 19288 1838
rect 19536 1714 19564 3402
rect 19628 3398 19656 3674
rect 19706 3632 19762 3641
rect 19706 3567 19708 3576
rect 19760 3567 19762 3576
rect 19708 3538 19760 3544
rect 19812 3482 19840 6174
rect 19904 5914 19932 6190
rect 19892 5908 19944 5914
rect 19892 5850 19944 5856
rect 19892 5636 19944 5642
rect 19892 5578 19944 5584
rect 19904 5098 19932 5578
rect 19892 5092 19944 5098
rect 19892 5034 19944 5040
rect 19904 4690 19932 5034
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19890 4176 19946 4185
rect 19890 4111 19946 4120
rect 19720 3454 19840 3482
rect 19616 3392 19668 3398
rect 19616 3334 19668 3340
rect 19614 3224 19670 3233
rect 19614 3159 19670 3168
rect 19444 1686 19564 1714
rect 19246 1456 19302 1465
rect 18972 1420 19024 1426
rect 19246 1391 19302 1400
rect 18972 1362 19024 1368
rect 18708 921 18736 1294
rect 18892 1278 19012 1306
rect 18694 912 18750 921
rect 18694 847 18750 856
rect 18984 800 19012 1278
rect 19444 800 19472 1686
rect 11164 734 11376 762
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12254 0 12310 800
rect 12714 0 12770 800
rect 13082 0 13138 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14370 0 14426 800
rect 14830 0 14886 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16854 0 16910 800
rect 17314 0 17370 800
rect 17682 0 17738 800
rect 18142 0 18198 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19430 0 19486 800
rect 19628 241 19656 3159
rect 19720 2990 19748 3454
rect 19800 3392 19852 3398
rect 19800 3334 19852 3340
rect 19812 3126 19840 3334
rect 19800 3120 19852 3126
rect 19800 3062 19852 3068
rect 19708 2984 19760 2990
rect 19708 2926 19760 2932
rect 19904 2650 19932 4111
rect 19996 3058 20024 6666
rect 20088 5370 20116 7346
rect 20180 5370 20208 8366
rect 20272 7800 20300 10503
rect 20364 9926 20392 10639
rect 20352 9920 20404 9926
rect 20352 9862 20404 9868
rect 20352 9648 20404 9654
rect 20352 9590 20404 9596
rect 20364 8498 20392 9590
rect 20352 8492 20404 8498
rect 20352 8434 20404 8440
rect 20272 7772 20392 7800
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20076 5364 20128 5370
rect 20076 5306 20128 5312
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20272 4826 20300 6258
rect 20364 5273 20392 7772
rect 20456 6662 20484 11698
rect 20548 10266 20576 12038
rect 20640 11898 20668 12294
rect 20718 12064 20774 12073
rect 20718 11999 20774 12008
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20628 11620 20680 11626
rect 20628 11562 20680 11568
rect 20640 11354 20668 11562
rect 20628 11348 20680 11354
rect 20628 11290 20680 11296
rect 20732 11200 20760 11999
rect 20824 11937 20852 12310
rect 20810 11928 20866 11937
rect 20810 11863 20866 11872
rect 20810 11792 20866 11801
rect 20810 11727 20866 11736
rect 20824 11626 20852 11727
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20812 11280 20864 11286
rect 20812 11222 20864 11228
rect 20640 11172 20760 11200
rect 20640 11014 20668 11172
rect 20824 11121 20852 11222
rect 20916 11150 20944 17546
rect 21008 17202 21036 18634
rect 21100 17762 21128 20198
rect 21284 19938 21312 22200
rect 21652 20534 21680 22200
rect 21640 20528 21692 20534
rect 21640 20470 21692 20476
rect 21364 20460 21416 20466
rect 21364 20402 21416 20408
rect 21192 19910 21312 19938
rect 21192 19174 21220 19910
rect 21272 19848 21324 19854
rect 21272 19790 21324 19796
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21284 17814 21312 19790
rect 21376 18154 21404 20402
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 18873 21496 20198
rect 21638 19952 21694 19961
rect 21638 19887 21694 19896
rect 21548 19712 21600 19718
rect 21548 19654 21600 19660
rect 21454 18864 21510 18873
rect 21454 18799 21510 18808
rect 21456 18624 21508 18630
rect 21456 18566 21508 18572
rect 21364 18148 21416 18154
rect 21364 18090 21416 18096
rect 21468 18057 21496 18566
rect 21560 18465 21588 19654
rect 21546 18456 21602 18465
rect 21546 18391 21602 18400
rect 21454 18048 21510 18057
rect 21454 17983 21510 17992
rect 21272 17808 21324 17814
rect 21100 17734 21220 17762
rect 21272 17750 21324 17756
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 20996 17196 21048 17202
rect 20996 17138 21048 17144
rect 21100 16726 21128 17614
rect 21088 16720 21140 16726
rect 21088 16662 21140 16668
rect 21086 16280 21142 16289
rect 21086 16215 21142 16224
rect 21100 16182 21128 16215
rect 21088 16176 21140 16182
rect 21088 16118 21140 16124
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 21008 15434 21036 16050
rect 21086 15464 21142 15473
rect 20996 15428 21048 15434
rect 21086 15399 21142 15408
rect 20996 15370 21048 15376
rect 21100 15366 21128 15399
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21192 15178 21220 17734
rect 21454 17640 21510 17649
rect 21454 17575 21510 17584
rect 21468 17542 21496 17575
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21272 17196 21324 17202
rect 21272 17138 21324 17144
rect 21284 16794 21312 17138
rect 21456 16992 21508 16998
rect 21456 16934 21508 16940
rect 21468 16833 21496 16934
rect 21454 16824 21510 16833
rect 21272 16788 21324 16794
rect 21454 16759 21510 16768
rect 21272 16730 21324 16736
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21284 15706 21312 16526
rect 21456 16448 21508 16454
rect 21456 16390 21508 16396
rect 21468 16289 21496 16390
rect 21454 16280 21510 16289
rect 21454 16215 21510 16224
rect 21456 15904 21508 15910
rect 21454 15872 21456 15881
rect 21508 15872 21510 15881
rect 21454 15807 21510 15816
rect 21272 15700 21324 15706
rect 21272 15642 21324 15648
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21100 15150 21220 15178
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14482 21036 14758
rect 21100 14618 21128 15150
rect 21180 15020 21232 15026
rect 21180 14962 21232 14968
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 20996 14476 21048 14482
rect 20996 14418 21048 14424
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21100 13841 21128 14010
rect 21192 14006 21220 14962
rect 21284 14890 21312 15438
rect 21456 15360 21508 15366
rect 21456 15302 21508 15308
rect 21468 15065 21496 15302
rect 21454 15056 21510 15065
rect 21454 14991 21510 15000
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 21456 14816 21508 14822
rect 21456 14758 21508 14764
rect 21468 14657 21496 14758
rect 21454 14648 21510 14657
rect 21454 14583 21510 14592
rect 21456 14272 21508 14278
rect 21454 14240 21456 14249
rect 21508 14240 21510 14249
rect 21454 14175 21510 14184
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 21272 13932 21324 13938
rect 21272 13874 21324 13880
rect 21086 13832 21142 13841
rect 21086 13767 21142 13776
rect 21284 13530 21312 13874
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 21468 13433 21496 13670
rect 21652 13569 21680 19887
rect 22020 19786 22048 22200
rect 22008 19780 22060 19786
rect 22008 19722 22060 19728
rect 22388 17338 22416 22200
rect 22756 18902 22784 22200
rect 22744 18896 22796 18902
rect 22744 18838 22796 18844
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22376 17332 22428 17338
rect 22376 17274 22428 17280
rect 21732 16652 21784 16658
rect 21732 16594 21784 16600
rect 21638 13560 21694 13569
rect 21638 13495 21694 13504
rect 21454 13424 21510 13433
rect 21454 13359 21510 13368
rect 21272 13320 21324 13326
rect 21272 13262 21324 13268
rect 21180 12844 21232 12850
rect 21180 12786 21232 12792
rect 21088 12708 21140 12714
rect 21088 12650 21140 12656
rect 20996 12640 21048 12646
rect 20996 12582 21048 12588
rect 20904 11144 20956 11150
rect 20810 11112 20866 11121
rect 20904 11086 20956 11092
rect 20810 11047 20866 11056
rect 20628 11008 20680 11014
rect 20628 10950 20680 10956
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20640 10810 20668 10950
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20720 10464 20772 10470
rect 20720 10406 20772 10412
rect 20536 10260 20588 10266
rect 20536 10202 20588 10208
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20548 9722 20576 9930
rect 20732 9874 20760 10406
rect 20824 9994 20852 10950
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20812 9988 20864 9994
rect 20812 9930 20864 9936
rect 20724 9846 20760 9874
rect 20724 9738 20752 9846
rect 20536 9716 20588 9722
rect 20724 9710 20852 9738
rect 20536 9658 20588 9664
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20732 9178 20760 9454
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20534 9072 20590 9081
rect 20534 9007 20590 9016
rect 20548 7886 20576 9007
rect 20628 8968 20680 8974
rect 20628 8910 20680 8916
rect 20536 7880 20588 7886
rect 20536 7822 20588 7828
rect 20536 7472 20588 7478
rect 20536 7414 20588 7420
rect 20444 6656 20496 6662
rect 20444 6598 20496 6604
rect 20444 6112 20496 6118
rect 20444 6054 20496 6060
rect 20350 5264 20406 5273
rect 20350 5199 20406 5208
rect 20260 4820 20312 4826
rect 20260 4762 20312 4768
rect 20168 4140 20220 4146
rect 20168 4082 20220 4088
rect 20076 3664 20128 3670
rect 20076 3606 20128 3612
rect 20088 3534 20116 3606
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 20180 3233 20208 4082
rect 20260 4072 20312 4078
rect 20258 4040 20260 4049
rect 20352 4072 20404 4078
rect 20312 4040 20314 4049
rect 20352 4014 20404 4020
rect 20258 3975 20314 3984
rect 20260 3664 20312 3670
rect 20260 3606 20312 3612
rect 20166 3224 20222 3233
rect 20166 3159 20222 3168
rect 19984 3052 20036 3058
rect 19984 2994 20036 3000
rect 20272 2666 20300 3606
rect 20364 3602 20392 4014
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20456 3534 20484 6054
rect 20444 3528 20496 3534
rect 20444 3470 20496 3476
rect 20548 2990 20576 7414
rect 20640 6458 20668 8910
rect 20718 8664 20774 8673
rect 20718 8599 20774 8608
rect 20732 8566 20760 8599
rect 20720 8560 20772 8566
rect 20720 8502 20772 8508
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20732 8265 20760 8366
rect 20718 8256 20774 8265
rect 20718 8191 20774 8200
rect 20718 7848 20774 7857
rect 20718 7783 20720 7792
rect 20772 7783 20774 7792
rect 20720 7754 20772 7760
rect 20824 7546 20852 9710
rect 20916 7546 20944 10610
rect 21008 10441 21036 12582
rect 21100 12306 21128 12650
rect 21088 12300 21140 12306
rect 21088 12242 21140 12248
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 21100 11082 21128 12038
rect 21088 11076 21140 11082
rect 21088 11018 21140 11024
rect 21100 10849 21128 11018
rect 21086 10840 21142 10849
rect 21086 10775 21142 10784
rect 20994 10432 21050 10441
rect 20994 10367 21050 10376
rect 20994 10296 21050 10305
rect 20994 10231 21050 10240
rect 21008 10198 21036 10231
rect 20996 10192 21048 10198
rect 20996 10134 21048 10140
rect 21086 10160 21142 10169
rect 21192 10146 21220 12786
rect 21284 12442 21312 13262
rect 21456 13184 21508 13190
rect 21456 13126 21508 13132
rect 21468 12889 21496 13126
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21454 12880 21510 12889
rect 21454 12815 21510 12824
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21270 11928 21326 11937
rect 21270 11863 21326 11872
rect 21284 10470 21312 11863
rect 21376 11234 21404 12650
rect 21456 12640 21508 12646
rect 21456 12582 21508 12588
rect 21468 12481 21496 12582
rect 21454 12472 21510 12481
rect 21454 12407 21510 12416
rect 21454 12336 21510 12345
rect 21560 12306 21588 12922
rect 21640 12912 21692 12918
rect 21640 12854 21692 12860
rect 21454 12271 21510 12280
rect 21548 12300 21600 12306
rect 21468 12238 21496 12271
rect 21548 12242 21600 12248
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21548 12164 21600 12170
rect 21548 12106 21600 12112
rect 21456 12096 21508 12102
rect 21454 12064 21456 12073
rect 21508 12064 21510 12073
rect 21454 11999 21510 12008
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 21468 11354 21496 11766
rect 21560 11694 21588 12106
rect 21548 11688 21600 11694
rect 21546 11656 21548 11665
rect 21600 11656 21602 11665
rect 21546 11591 21602 11600
rect 21546 11384 21602 11393
rect 21456 11348 21508 11354
rect 21546 11319 21602 11328
rect 21456 11290 21508 11296
rect 21454 11248 21510 11257
rect 21376 11206 21454 11234
rect 21454 11183 21510 11192
rect 21468 11150 21496 11183
rect 21456 11144 21508 11150
rect 21456 11086 21508 11092
rect 21560 10996 21588 11319
rect 21376 10968 21588 10996
rect 21272 10464 21324 10470
rect 21272 10406 21324 10412
rect 21192 10118 21312 10146
rect 21086 10095 21088 10104
rect 21140 10095 21142 10104
rect 21088 10066 21140 10072
rect 21180 10056 21232 10062
rect 21086 10024 21142 10033
rect 21180 9998 21232 10004
rect 21086 9959 21142 9968
rect 20994 9752 21050 9761
rect 20994 9687 21050 9696
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 20904 7404 20956 7410
rect 20904 7346 20956 7352
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20720 6724 20772 6730
rect 20720 6666 20772 6672
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20626 6352 20682 6361
rect 20626 6287 20682 6296
rect 20640 5234 20668 6287
rect 20628 5228 20680 5234
rect 20628 5170 20680 5176
rect 20626 4584 20682 4593
rect 20626 4519 20682 4528
rect 20640 3126 20668 4519
rect 20732 4282 20760 6666
rect 20720 4276 20772 4282
rect 20720 4218 20772 4224
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20628 3120 20680 3126
rect 20628 3062 20680 3068
rect 20732 3058 20760 3878
rect 20824 3534 20852 7142
rect 20916 5914 20944 7346
rect 21008 6644 21036 9687
rect 21100 9674 21128 9959
rect 21192 9897 21220 9998
rect 21178 9888 21234 9897
rect 21178 9823 21234 9832
rect 21100 9646 21220 9674
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21100 7546 21128 8774
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21086 6896 21142 6905
rect 21086 6831 21088 6840
rect 21140 6831 21142 6840
rect 21088 6802 21140 6808
rect 21008 6616 21128 6644
rect 20994 6488 21050 6497
rect 20994 6423 21050 6432
rect 21008 6322 21036 6423
rect 20996 6316 21048 6322
rect 20996 6258 21048 6264
rect 20904 5908 20956 5914
rect 20904 5850 20956 5856
rect 21100 5710 21128 6616
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20994 5536 21050 5545
rect 20994 5471 21050 5480
rect 21008 5166 21036 5471
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 20904 5024 20956 5030
rect 20904 4966 20956 4972
rect 20916 4690 20944 4966
rect 20904 4684 20956 4690
rect 20904 4626 20956 4632
rect 20996 4548 21048 4554
rect 20996 4490 21048 4496
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20536 2984 20588 2990
rect 20536 2926 20588 2932
rect 20628 2916 20680 2922
rect 20628 2858 20680 2864
rect 19892 2644 19944 2650
rect 19892 2586 19944 2592
rect 20180 2638 20300 2666
rect 19812 870 19932 898
rect 19812 800 19840 870
rect 19614 232 19670 241
rect 19614 167 19670 176
rect 19798 0 19854 800
rect 19904 762 19932 870
rect 20180 762 20208 2638
rect 20352 2440 20404 2446
rect 20352 2382 20404 2388
rect 20364 2038 20392 2382
rect 20352 2032 20404 2038
rect 20352 1974 20404 1980
rect 20260 1284 20312 1290
rect 20260 1226 20312 1232
rect 20272 800 20300 1226
rect 20640 800 20668 2858
rect 20732 2689 20760 2994
rect 20718 2680 20774 2689
rect 20718 2615 20774 2624
rect 21008 2582 21036 4490
rect 21100 3194 21128 5646
rect 21192 4554 21220 9646
rect 21284 8673 21312 10118
rect 21376 9874 21404 10968
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21454 10432 21510 10441
rect 21454 10367 21510 10376
rect 21468 10062 21496 10367
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21376 9846 21496 9874
rect 21270 8664 21326 8673
rect 21270 8599 21326 8608
rect 21272 8492 21324 8498
rect 21272 8434 21324 8440
rect 21180 4548 21232 4554
rect 21180 4490 21232 4496
rect 21088 3188 21140 3194
rect 21088 3130 21140 3136
rect 20996 2576 21048 2582
rect 20996 2518 21048 2524
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20732 1057 20760 2382
rect 21284 2122 21312 8434
rect 21362 8120 21418 8129
rect 21362 8055 21364 8064
rect 21416 8055 21418 8064
rect 21364 8026 21416 8032
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 21376 7546 21404 7890
rect 21364 7540 21416 7546
rect 21364 7482 21416 7488
rect 21376 5098 21404 7482
rect 21468 6662 21496 9846
rect 21560 7410 21588 10542
rect 21652 8265 21680 12854
rect 21638 8256 21694 8265
rect 21638 8191 21694 8200
rect 21548 7404 21600 7410
rect 21548 7346 21600 7352
rect 21560 7002 21588 7346
rect 21744 7290 21772 16594
rect 22282 16552 22338 16561
rect 22282 16487 22338 16496
rect 21916 15972 21968 15978
rect 21916 15914 21968 15920
rect 21822 14376 21878 14385
rect 21822 14311 21878 14320
rect 21836 14278 21864 14311
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21824 13252 21876 13258
rect 21824 13194 21876 13200
rect 21836 7857 21864 13194
rect 21822 7848 21878 7857
rect 21822 7783 21878 7792
rect 21652 7262 21772 7290
rect 21548 6996 21600 7002
rect 21548 6938 21600 6944
rect 21456 6656 21508 6662
rect 21456 6598 21508 6604
rect 21454 6488 21510 6497
rect 21454 6423 21510 6432
rect 21468 6254 21496 6423
rect 21456 6248 21508 6254
rect 21456 6190 21508 6196
rect 21560 5778 21588 6938
rect 21548 5772 21600 5778
rect 21548 5714 21600 5720
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21560 4690 21588 5714
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21548 4548 21600 4554
rect 21548 4490 21600 4496
rect 21454 3496 21510 3505
rect 21454 3431 21510 3440
rect 21364 3392 21416 3398
rect 21364 3334 21416 3340
rect 21100 2094 21312 2122
rect 20718 1048 20774 1057
rect 20718 983 20774 992
rect 21100 800 21128 2094
rect 21376 950 21404 3334
rect 21364 944 21416 950
rect 21364 886 21416 892
rect 21468 800 21496 3431
rect 21560 2281 21588 4490
rect 21652 4146 21680 7262
rect 21732 7200 21784 7206
rect 21732 7142 21784 7148
rect 21640 4140 21692 4146
rect 21640 4082 21692 4088
rect 21652 4049 21680 4082
rect 21638 4040 21694 4049
rect 21638 3975 21694 3984
rect 21744 3942 21772 7142
rect 21836 6798 21864 7783
rect 21824 6792 21876 6798
rect 21824 6734 21876 6740
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 21836 4078 21864 6598
rect 21928 5234 21956 15914
rect 22008 15564 22060 15570
rect 22008 15506 22060 15512
rect 22020 7206 22048 15506
rect 22192 15428 22244 15434
rect 22192 15370 22244 15376
rect 22204 12434 22232 15370
rect 22112 12406 22232 12434
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22008 7064 22060 7070
rect 22006 7032 22008 7041
rect 22060 7032 22062 7041
rect 22006 6967 22062 6976
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21928 4865 21956 5170
rect 21914 4856 21970 4865
rect 21914 4791 21970 4800
rect 22020 4622 22048 6967
rect 22008 4616 22060 4622
rect 22008 4558 22060 4564
rect 22006 4448 22062 4457
rect 22112 4434 22140 12406
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 22204 10674 22232 12242
rect 22192 10668 22244 10674
rect 22192 10610 22244 10616
rect 22296 7562 22324 16487
rect 22376 15632 22428 15638
rect 22376 15574 22428 15580
rect 22062 4406 22140 4434
rect 22204 7534 22324 7562
rect 22006 4383 22062 4392
rect 21824 4072 21876 4078
rect 21824 4014 21876 4020
rect 21732 3936 21784 3942
rect 21732 3878 21784 3884
rect 22020 3534 22048 4383
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22006 3088 22062 3097
rect 22006 3023 22062 3032
rect 21914 2952 21970 2961
rect 21914 2887 21970 2896
rect 21732 2576 21784 2582
rect 21732 2518 21784 2524
rect 21744 2417 21772 2518
rect 21730 2408 21786 2417
rect 21730 2343 21786 2352
rect 21824 2372 21876 2378
rect 21824 2314 21876 2320
rect 21546 2272 21602 2281
rect 21546 2207 21602 2216
rect 21836 1902 21864 2314
rect 21824 1896 21876 1902
rect 21822 1864 21824 1873
rect 21876 1864 21878 1873
rect 21822 1799 21878 1808
rect 21928 800 21956 2887
rect 22020 1426 22048 3023
rect 22204 2514 22232 7534
rect 22388 7070 22416 15574
rect 22468 14272 22520 14278
rect 22468 14214 22520 14220
rect 22376 7064 22428 7070
rect 22376 7006 22428 7012
rect 22282 3360 22338 3369
rect 22282 3295 22338 3304
rect 22192 2508 22244 2514
rect 22192 2450 22244 2456
rect 22008 1420 22060 1426
rect 22008 1362 22060 1368
rect 22296 800 22324 3295
rect 22480 2774 22508 14214
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22572 5302 22600 10610
rect 22560 5296 22612 5302
rect 22560 5238 22612 5244
rect 22388 2746 22508 2774
rect 22388 1902 22416 2746
rect 22572 2446 22600 5238
rect 22664 2582 22692 17546
rect 22744 14952 22796 14958
rect 22744 14894 22796 14900
rect 22756 12434 22784 14894
rect 22928 13456 22980 13462
rect 22928 13398 22980 13404
rect 22756 12406 22876 12434
rect 22744 11620 22796 11626
rect 22744 11562 22796 11568
rect 22756 4826 22784 11562
rect 22744 4820 22796 4826
rect 22744 4762 22796 4768
rect 22848 3738 22876 12406
rect 22940 6390 22968 13398
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 22836 3732 22888 3738
rect 22836 3674 22888 3680
rect 22652 2576 22704 2582
rect 22652 2518 22704 2524
rect 22560 2440 22612 2446
rect 22560 2382 22612 2388
rect 22376 1896 22428 1902
rect 22376 1838 22428 1844
rect 22744 1420 22796 1426
rect 22744 1362 22796 1368
rect 22756 800 22784 1362
rect 19904 734 20208 762
rect 20258 0 20314 800
rect 20626 0 20682 800
rect 21086 0 21142 800
rect 21454 0 21510 800
rect 21914 0 21970 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 294 22888 350 22944
rect 1030 22480 1086 22536
rect 1122 22344 1178 22400
rect 1030 21936 1086 21992
rect 846 14014 902 14070
rect 294 6704 350 6760
rect 2410 22616 2466 22672
rect 1214 20848 1270 20904
rect 1030 10920 1086 10976
rect 1030 9460 1032 9480
rect 1032 9460 1084 9480
rect 1084 9460 1086 9480
rect 1030 9424 1086 9460
rect 1030 7828 1032 7848
rect 1032 7828 1084 7848
rect 1084 7828 1086 7848
rect 1030 7792 1086 7828
rect 1030 7656 1086 7712
rect 938 6024 994 6080
rect 1122 4528 1178 4584
rect 938 3984 994 4040
rect 1306 18944 1362 19000
rect 1582 20168 1638 20224
rect 1490 19796 1492 19816
rect 1492 19796 1544 19816
rect 1544 19796 1546 19816
rect 1766 20984 1822 21040
rect 1490 19760 1546 19796
rect 1490 19660 1492 19680
rect 1492 19660 1544 19680
rect 1544 19660 1546 19680
rect 1490 19624 1546 19660
rect 1490 18808 1546 18864
rect 2226 21800 2282 21856
rect 2042 20304 2098 20360
rect 1950 19624 2006 19680
rect 1950 19372 2006 19408
rect 1950 19352 1952 19372
rect 1952 19352 2004 19372
rect 2004 19352 2006 19372
rect 1858 19236 1914 19272
rect 1858 19216 1860 19236
rect 1860 19216 1912 19236
rect 1912 19216 1914 19236
rect 1582 18672 1638 18728
rect 1490 18400 1546 18456
rect 1858 18028 1860 18048
rect 1860 18028 1912 18048
rect 1912 18028 1914 18048
rect 1858 17992 1914 18028
rect 2318 21664 2374 21720
rect 2318 19216 2374 19272
rect 4158 22208 4214 22264
rect 2502 21392 2558 21448
rect 2134 18400 2190 18456
rect 2134 18028 2136 18048
rect 2136 18028 2188 18048
rect 2188 18028 2190 18048
rect 2134 17992 2190 18028
rect 1950 17720 2006 17776
rect 1490 17584 1546 17640
rect 1490 17176 1546 17232
rect 1490 16768 1546 16824
rect 1490 16224 1546 16280
rect 1490 15852 1492 15872
rect 1492 15852 1544 15872
rect 1544 15852 1546 15872
rect 1490 15816 1546 15852
rect 1490 15000 1546 15056
rect 1490 14592 1546 14648
rect 1858 15408 1914 15464
rect 1674 14456 1730 14512
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1490 13368 1546 13424
rect 2870 20576 2926 20632
rect 3054 19216 3110 19272
rect 2870 18536 2926 18592
rect 2226 17312 2282 17368
rect 2410 17196 2466 17232
rect 2410 17176 2412 17196
rect 2412 17176 2464 17196
rect 2464 17176 2466 17196
rect 2134 16496 2190 16552
rect 2502 16224 2558 16280
rect 3422 21120 3478 21176
rect 3330 19760 3386 19816
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 4158 19352 4214 19408
rect 3790 18536 3846 18592
rect 3330 18128 3386 18184
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 4158 18944 4214 19000
rect 4158 17856 4214 17912
rect 4434 19896 4490 19952
rect 4434 19624 4490 19680
rect 4158 17584 4214 17640
rect 3238 17448 3294 17504
rect 2686 16360 2742 16416
rect 1858 13796 1914 13832
rect 1858 13776 1860 13796
rect 1860 13776 1912 13796
rect 1912 13776 1914 13796
rect 2042 13776 2098 13832
rect 1490 12824 1546 12880
rect 1490 12416 1546 12472
rect 1398 12144 1454 12200
rect 1490 11328 1546 11384
rect 1490 10784 1546 10840
rect 1950 13368 2006 13424
rect 1858 12008 1914 12064
rect 1858 11192 1914 11248
rect 1674 9988 1730 10024
rect 1674 9968 1676 9988
rect 1676 9968 1728 9988
rect 1728 9968 1730 9988
rect 1582 9696 1638 9752
rect 1306 9016 1362 9072
rect 1306 8200 1362 8256
rect 1306 6976 1362 7032
rect 1490 8608 1546 8664
rect 1582 8472 1638 8528
rect 3146 15952 3202 16008
rect 2686 14184 2742 14240
rect 2134 11600 2190 11656
rect 3238 14900 3240 14920
rect 3240 14900 3292 14920
rect 3292 14900 3294 14920
rect 3238 14864 3294 14900
rect 2962 13504 3018 13560
rect 2778 13232 2834 13288
rect 2686 12144 2742 12200
rect 2410 11600 2466 11656
rect 2042 9560 2098 9616
rect 1950 9444 2006 9480
rect 1950 9424 1952 9444
rect 1952 9424 2004 9444
rect 2004 9424 2006 9444
rect 2594 12008 2650 12064
rect 1766 9016 1822 9072
rect 1490 7420 1492 7440
rect 1492 7420 1544 7440
rect 1544 7420 1546 7440
rect 1490 7384 1546 7420
rect 1674 7248 1730 7304
rect 1858 8880 1914 8936
rect 1582 6840 1638 6896
rect 1398 6568 1454 6624
rect 1306 5888 1362 5944
rect 1490 5480 1546 5536
rect 1306 1944 1362 2000
rect 938 176 994 232
rect 2502 9832 2558 9888
rect 2226 7656 2282 7712
rect 2502 8336 2558 8392
rect 2410 7928 2466 7984
rect 2686 11056 2742 11112
rect 2962 12552 3018 12608
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3974 16768 4030 16824
rect 4802 20168 4858 20224
rect 4986 20032 5042 20088
rect 4710 18300 4712 18320
rect 4712 18300 4764 18320
rect 4764 18300 4766 18320
rect 4710 18264 4766 18300
rect 4618 17992 4674 18048
rect 4618 17040 4674 17096
rect 4526 16904 4582 16960
rect 4250 16496 4306 16552
rect 4158 16224 4214 16280
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3514 13912 3570 13968
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 4066 14220 4068 14240
rect 4068 14220 4120 14240
rect 4120 14220 4122 14240
rect 4066 14184 4122 14220
rect 3882 13368 3938 13424
rect 3054 12416 3110 12472
rect 2778 10376 2834 10432
rect 2686 7792 2742 7848
rect 2594 7520 2650 7576
rect 2226 4800 2282 4856
rect 1950 4140 2006 4176
rect 1950 4120 1952 4140
rect 1952 4120 2004 4140
rect 2004 4120 2006 4140
rect 1858 3576 1914 3632
rect 2870 8744 2926 8800
rect 4342 13388 4398 13424
rect 4342 13368 4344 13388
rect 4344 13368 4396 13388
rect 4396 13368 4398 13388
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3790 11092 3792 11112
rect 3792 11092 3844 11112
rect 3844 11092 3846 11112
rect 3790 11056 3846 11092
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3790 10104 3846 10160
rect 3054 8200 3110 8256
rect 3330 9288 3386 9344
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 4526 13368 4582 13424
rect 3974 10376 4030 10432
rect 3974 9968 4030 10024
rect 2870 5072 2926 5128
rect 3054 5616 3110 5672
rect 3054 4392 3110 4448
rect 2594 3168 2650 3224
rect 2778 2896 2834 2952
rect 2686 2760 2742 2816
rect 3514 8744 3570 8800
rect 4434 12688 4490 12744
rect 4342 10376 4398 10432
rect 4250 10240 4306 10296
rect 4158 9832 4214 9888
rect 4250 9424 4306 9480
rect 4158 9152 4214 9208
rect 4066 9016 4122 9072
rect 3974 8608 4030 8664
rect 3882 8472 3938 8528
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3514 7928 3570 7984
rect 3606 7384 3662 7440
rect 3882 7928 3938 7984
rect 4066 8200 4122 8256
rect 4066 8064 4122 8120
rect 3790 7656 3846 7712
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3514 6860 3570 6896
rect 3514 6840 3516 6860
rect 3516 6840 3568 6860
rect 3568 6840 3570 6860
rect 3698 6840 3754 6896
rect 5170 18264 5226 18320
rect 5078 17720 5134 17776
rect 5262 17992 5318 18048
rect 5446 18536 5502 18592
rect 7746 22752 7802 22808
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6550 20576 6606 20632
rect 6550 20440 6606 20496
rect 6274 20168 6330 20224
rect 6458 20204 6460 20224
rect 6460 20204 6512 20224
rect 6512 20204 6514 20224
rect 6458 20168 6514 20204
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5814 19080 5870 19136
rect 5630 18536 5686 18592
rect 5630 18400 5686 18456
rect 5630 17992 5686 18048
rect 5722 17584 5778 17640
rect 5722 17484 5724 17504
rect 5724 17484 5776 17504
rect 5776 17484 5778 17504
rect 5722 17448 5778 17484
rect 5630 16904 5686 16960
rect 5538 16496 5594 16552
rect 5078 14864 5134 14920
rect 5078 14048 5134 14104
rect 4342 9152 4398 9208
rect 3790 6432 3846 6488
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3606 5788 3608 5808
rect 3608 5788 3660 5808
rect 3660 5788 3662 5808
rect 3606 5752 3662 5788
rect 3790 5752 3846 5808
rect 3790 5208 3846 5264
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3882 4528 3938 4584
rect 3422 3984 3478 4040
rect 3882 4004 3938 4040
rect 3882 3984 3884 4004
rect 3884 3984 3936 4004
rect 3936 3984 3938 4004
rect 3238 856 3294 912
rect 4158 5072 4214 5128
rect 4066 4800 4122 4856
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4526 6840 4582 6896
rect 4434 5072 4490 5128
rect 4342 4548 4398 4584
rect 4342 4528 4344 4548
rect 4344 4528 4396 4548
rect 4396 4528 4398 4548
rect 4342 4256 4398 4312
rect 4250 3576 4306 3632
rect 4158 2760 4214 2816
rect 4250 1808 4306 1864
rect 4710 9288 4766 9344
rect 4710 7792 4766 7848
rect 4618 4392 4674 4448
rect 4526 3712 4582 3768
rect 4894 12144 4950 12200
rect 5078 11500 5080 11520
rect 5080 11500 5132 11520
rect 5132 11500 5134 11520
rect 5078 11464 5134 11500
rect 5630 15408 5686 15464
rect 5538 14728 5594 14784
rect 5538 13776 5594 13832
rect 5446 13504 5502 13560
rect 5354 12552 5410 12608
rect 5354 11736 5410 11792
rect 5170 11192 5226 11248
rect 4986 10784 5042 10840
rect 5262 10260 5318 10296
rect 5262 10240 5264 10260
rect 5264 10240 5316 10260
rect 5316 10240 5318 10260
rect 7746 22072 7802 22128
rect 7470 21936 7526 21992
rect 7470 21664 7526 21720
rect 7194 19760 7250 19816
rect 7102 19624 7158 19680
rect 7102 19488 7158 19544
rect 6918 19216 6974 19272
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6550 17448 6606 17504
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6182 17040 6238 17096
rect 6274 16768 6330 16824
rect 5722 15000 5778 15056
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6734 18536 6790 18592
rect 6734 18400 6790 18456
rect 7010 18400 7066 18456
rect 6734 17992 6790 18048
rect 7470 18400 7526 18456
rect 7286 17856 7342 17912
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 7010 15136 7066 15192
rect 7194 16768 7250 16824
rect 7470 17312 7526 17368
rect 7194 16360 7250 16416
rect 6826 14592 6882 14648
rect 6734 14340 6790 14376
rect 6734 14320 6736 14340
rect 6736 14320 6788 14340
rect 6788 14320 6790 14340
rect 6550 14220 6552 14240
rect 6552 14220 6604 14240
rect 6604 14220 6606 14240
rect 6550 14184 6606 14220
rect 7286 14220 7288 14240
rect 7288 14220 7340 14240
rect 7340 14220 7342 14240
rect 7286 14184 7342 14220
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6826 14048 6882 14104
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5998 12824 6054 12880
rect 5170 9868 5172 9888
rect 5172 9868 5224 9888
rect 5224 9868 5226 9888
rect 5170 9832 5226 9868
rect 4894 9424 4950 9480
rect 5170 9560 5226 9616
rect 5538 9968 5594 10024
rect 5170 8744 5226 8800
rect 5262 8492 5318 8528
rect 5262 8472 5264 8492
rect 5264 8472 5316 8492
rect 5316 8472 5318 8492
rect 4526 2760 4582 2816
rect 5170 6740 5172 6760
rect 5172 6740 5224 6760
rect 5224 6740 5226 6760
rect 5170 6704 5226 6740
rect 4894 3440 4950 3496
rect 4710 2624 4766 2680
rect 5630 9696 5686 9752
rect 5814 11872 5870 11928
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6642 12280 6698 12336
rect 6642 11872 6698 11928
rect 6550 11328 6606 11384
rect 6918 11328 6974 11384
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6550 10376 6606 10432
rect 5906 9968 5962 10024
rect 5630 9016 5686 9072
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6458 9580 6514 9616
rect 6458 9560 6460 9580
rect 6460 9560 6512 9580
rect 6512 9560 6514 9580
rect 6642 10004 6644 10024
rect 6644 10004 6696 10024
rect 6696 10004 6698 10024
rect 6642 9968 6698 10004
rect 6550 9288 6606 9344
rect 5998 9016 6054 9072
rect 5354 7520 5410 7576
rect 5630 7520 5686 7576
rect 6826 10920 6882 10976
rect 7378 12044 7380 12064
rect 7380 12044 7432 12064
rect 7432 12044 7434 12064
rect 7378 12008 7434 12044
rect 7378 11736 7434 11792
rect 7286 11056 7342 11112
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6090 8200 6146 8256
rect 5998 7928 6054 7984
rect 6458 7928 6514 7984
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6734 8608 6790 8664
rect 6550 7112 6606 7168
rect 6458 6976 6514 7032
rect 7010 8608 7066 8664
rect 7286 10512 7342 10568
rect 8114 19896 8170 19952
rect 8114 19660 8116 19680
rect 8116 19660 8168 19680
rect 8168 19660 8170 19680
rect 8114 19624 8170 19660
rect 8390 20304 8446 20360
rect 8114 19080 8170 19136
rect 7746 17740 7802 17776
rect 7746 17720 7748 17740
rect 7748 17720 7800 17740
rect 7800 17720 7802 17740
rect 7746 15816 7802 15872
rect 7654 15680 7710 15736
rect 8114 18400 8170 18456
rect 8114 17720 8170 17776
rect 8574 19896 8630 19952
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 9218 20032 9274 20088
rect 8666 19352 8722 19408
rect 8942 19488 8998 19544
rect 9126 19488 9182 19544
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 9494 18944 9550 19000
rect 8482 18672 8538 18728
rect 8482 18400 8538 18456
rect 8758 18300 8760 18320
rect 8760 18300 8812 18320
rect 8812 18300 8814 18320
rect 8758 18264 8814 18300
rect 9218 18400 9274 18456
rect 9218 18264 9274 18320
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 9402 18128 9458 18184
rect 9586 18128 9642 18184
rect 9126 17856 9182 17912
rect 9218 17196 9274 17232
rect 9218 17176 9220 17196
rect 9220 17176 9272 17196
rect 9272 17176 9274 17196
rect 8298 16904 8354 16960
rect 8850 17060 8906 17096
rect 8850 17040 8852 17060
rect 8852 17040 8904 17060
rect 8904 17040 8906 17060
rect 8022 16224 8078 16280
rect 8482 16224 8538 16280
rect 8022 15136 8078 15192
rect 7286 9832 7342 9888
rect 7378 9152 7434 9208
rect 6826 7420 6828 7440
rect 6828 7420 6880 7440
rect 6880 7420 6882 7440
rect 6826 7384 6882 7420
rect 7470 8608 7526 8664
rect 7378 8200 7434 8256
rect 6734 6976 6790 7032
rect 5722 6568 5778 6624
rect 5814 6452 5870 6488
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 5814 6432 5816 6452
rect 5816 6432 5868 6452
rect 5868 6432 5870 6452
rect 6642 6568 6698 6624
rect 6918 6568 6974 6624
rect 5814 6160 5870 6216
rect 6274 6296 6330 6352
rect 5538 5072 5594 5128
rect 5262 4392 5318 4448
rect 5078 4120 5134 4176
rect 4986 2352 5042 2408
rect 4894 992 4950 1048
rect 5170 3984 5226 4040
rect 5262 3168 5318 3224
rect 5170 1264 5226 1320
rect 5630 4528 5686 4584
rect 5906 5480 5962 5536
rect 5906 5228 5962 5264
rect 5906 5208 5908 5228
rect 5908 5208 5960 5228
rect 5960 5208 5962 5228
rect 6366 6196 6368 6216
rect 6368 6196 6420 6216
rect 6420 6196 6422 6216
rect 6366 6160 6422 6196
rect 6550 6160 6606 6216
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6734 5616 6790 5672
rect 6734 5208 6790 5264
rect 7010 5908 7066 5944
rect 7010 5888 7012 5908
rect 7012 5888 7064 5908
rect 7064 5888 7066 5908
rect 7286 6160 7342 6216
rect 7286 5888 7342 5944
rect 7194 5752 7250 5808
rect 5538 4120 5594 4176
rect 5722 4276 5778 4312
rect 5722 4256 5724 4276
rect 5724 4256 5776 4276
rect 5776 4256 5778 4276
rect 5630 3576 5686 3632
rect 5446 3032 5502 3088
rect 5814 3188 5870 3224
rect 5814 3168 5816 3188
rect 5816 3168 5868 3188
rect 5868 3168 5870 3188
rect 6366 4564 6368 4584
rect 6368 4564 6420 4584
rect 6420 4564 6422 4584
rect 6366 4528 6422 4564
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 5998 4276 6054 4312
rect 5998 4256 6000 4276
rect 6000 4256 6052 4276
rect 6052 4256 6054 4276
rect 7102 5344 7158 5400
rect 7010 4684 7066 4720
rect 7010 4664 7012 4684
rect 7012 4664 7064 4684
rect 7064 4664 7066 4684
rect 7194 4256 7250 4312
rect 6090 3596 6146 3632
rect 6090 3576 6092 3596
rect 6092 3576 6144 3596
rect 6144 3576 6146 3596
rect 5998 3440 6054 3496
rect 5906 2896 5962 2952
rect 6550 3304 6606 3360
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 5814 2624 5870 2680
rect 5722 2216 5778 2272
rect 5630 1536 5686 1592
rect 5078 856 5134 912
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 5998 2100 6054 2136
rect 5998 2080 6000 2100
rect 6000 2080 6052 2100
rect 6052 2080 6054 2100
rect 5998 1808 6054 1864
rect 7010 3712 7066 3768
rect 6734 1672 6790 1728
rect 7470 7520 7526 7576
rect 7470 6604 7472 6624
rect 7472 6604 7524 6624
rect 7524 6604 7526 6624
rect 7470 6568 7526 6604
rect 7470 6160 7526 6216
rect 8022 14592 8078 14648
rect 8022 13232 8078 13288
rect 8574 15852 8576 15872
rect 8576 15852 8628 15872
rect 8628 15852 8630 15872
rect 8574 15816 8630 15852
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8482 15272 8538 15328
rect 8574 14728 8630 14784
rect 8298 12688 8354 12744
rect 8114 12436 8170 12472
rect 8114 12416 8116 12436
rect 8116 12416 8168 12436
rect 8168 12416 8170 12436
rect 8022 11328 8078 11384
rect 7930 10784 7986 10840
rect 7654 8200 7710 8256
rect 7378 4256 7434 4312
rect 7010 2624 7066 2680
rect 7194 2216 7250 2272
rect 6918 1672 6974 1728
rect 7286 1944 7342 2000
rect 7194 1536 7250 1592
rect 8114 8880 8170 8936
rect 8114 8336 8170 8392
rect 8114 7928 8170 7984
rect 8298 12280 8354 12336
rect 8482 14048 8538 14104
rect 8390 12144 8446 12200
rect 9218 14728 9274 14784
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 9126 14592 9182 14648
rect 9862 20576 9918 20632
rect 9862 20304 9918 20360
rect 10138 20032 10194 20088
rect 9954 19352 10010 19408
rect 9862 18964 9918 19000
rect 9862 18944 9864 18964
rect 9864 18944 9916 18964
rect 9916 18944 9918 18964
rect 10322 19352 10378 19408
rect 10138 19216 10194 19272
rect 10414 19216 10470 19272
rect 10322 18944 10378 19000
rect 10138 18672 10194 18728
rect 10966 20168 11022 20224
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11978 20032 12034 20088
rect 10598 19760 10654 19816
rect 10782 19760 10838 19816
rect 11150 19624 11206 19680
rect 10414 17992 10470 18048
rect 10506 17720 10562 17776
rect 9770 17584 9826 17640
rect 9678 16904 9734 16960
rect 9678 15680 9734 15736
rect 9126 13912 9182 13968
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9034 13232 9090 13288
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8390 11756 8446 11792
rect 8390 11736 8392 11756
rect 8392 11736 8444 11756
rect 8444 11736 8446 11756
rect 8390 9696 8446 9752
rect 8390 9152 8446 9208
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8574 10376 8630 10432
rect 9218 11092 9220 11112
rect 9220 11092 9272 11112
rect 9272 11092 9274 11112
rect 9218 11056 9274 11092
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9034 9560 9090 9616
rect 8666 9424 8722 9480
rect 8574 9288 8630 9344
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8390 8880 8446 8936
rect 8574 8880 8630 8936
rect 8574 8200 8630 8256
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8022 6704 8078 6760
rect 8114 6160 8170 6216
rect 8114 5888 8170 5944
rect 8114 5652 8116 5672
rect 8116 5652 8168 5672
rect 8168 5652 8170 5672
rect 8114 5616 8170 5652
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8390 5888 8446 5944
rect 7746 4936 7802 4992
rect 7654 4428 7656 4448
rect 7656 4428 7708 4448
rect 7708 4428 7710 4448
rect 7654 4392 7710 4428
rect 7746 4256 7802 4312
rect 7654 3712 7710 3768
rect 7930 4936 7986 4992
rect 8022 4800 8078 4856
rect 8022 3032 8078 3088
rect 7838 2760 7894 2816
rect 7654 2624 7710 2680
rect 7470 1128 7526 1184
rect 8942 6840 8998 6896
rect 8758 6704 8814 6760
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9862 15272 9918 15328
rect 9678 13640 9734 13696
rect 9678 13504 9734 13560
rect 10506 17040 10562 17096
rect 10046 15000 10102 15056
rect 10690 17992 10746 18048
rect 10690 17584 10746 17640
rect 10690 17312 10746 17368
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 12438 20052 12494 20088
rect 12438 20032 12440 20052
rect 12440 20032 12492 20052
rect 12492 20032 12494 20052
rect 10966 19080 11022 19136
rect 11150 18944 11206 19000
rect 11058 18536 11114 18592
rect 11150 18400 11206 18456
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 10874 17740 10930 17776
rect 10874 17720 10876 17740
rect 10876 17720 10928 17740
rect 10928 17720 10930 17740
rect 11426 17992 11482 18048
rect 11794 17992 11850 18048
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 10782 16516 10838 16552
rect 10782 16496 10784 16516
rect 10784 16496 10836 16516
rect 10836 16496 10838 16516
rect 10138 14456 10194 14512
rect 9862 12688 9918 12744
rect 9678 12416 9734 12472
rect 9678 12280 9734 12336
rect 9678 11872 9734 11928
rect 9586 10240 9642 10296
rect 9494 9832 9550 9888
rect 9586 9696 9642 9752
rect 9494 9152 9550 9208
rect 9402 8744 9458 8800
rect 9310 7928 9366 7984
rect 9310 6976 9366 7032
rect 9586 8336 9642 8392
rect 9678 7656 9734 7712
rect 9310 6840 9366 6896
rect 9310 6604 9312 6624
rect 9312 6604 9364 6624
rect 9364 6604 9366 6624
rect 8850 5652 8852 5672
rect 8852 5652 8904 5672
rect 8904 5652 8906 5672
rect 8850 5616 8906 5652
rect 9034 5616 9090 5672
rect 8390 4936 8446 4992
rect 8298 4800 8354 4856
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8850 4528 8906 4584
rect 7930 1400 7986 1456
rect 8574 3168 8630 3224
rect 8574 2488 8630 2544
rect 8574 1536 8630 1592
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9126 2644 9182 2680
rect 9126 2624 9128 2644
rect 9128 2624 9180 2644
rect 9180 2624 9182 2644
rect 8758 2488 8814 2544
rect 9126 2488 9182 2544
rect 8942 1672 8998 1728
rect 9310 6568 9366 6604
rect 9310 5344 9366 5400
rect 10046 12588 10048 12608
rect 10048 12588 10100 12608
rect 10100 12588 10102 12608
rect 10046 12552 10102 12588
rect 10046 12144 10102 12200
rect 10414 15000 10470 15056
rect 10598 15272 10654 15328
rect 10966 15816 11022 15872
rect 11242 16904 11298 16960
rect 11518 16768 11574 16824
rect 12530 19352 12586 19408
rect 12346 18536 12402 18592
rect 11978 18400 12034 18456
rect 12530 18300 12532 18320
rect 12532 18300 12584 18320
rect 12584 18300 12586 18320
rect 12530 18264 12586 18300
rect 11794 17448 11850 17504
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11702 15544 11758 15600
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11150 15136 11206 15192
rect 10414 13232 10470 13288
rect 10046 11600 10102 11656
rect 9954 10784 10010 10840
rect 10230 11056 10286 11112
rect 10230 10512 10286 10568
rect 10046 10104 10102 10160
rect 9954 8628 10010 8664
rect 9954 8608 9956 8628
rect 9956 8608 10008 8628
rect 10008 8608 10010 8628
rect 9862 6976 9918 7032
rect 9586 6452 9642 6488
rect 9586 6432 9588 6452
rect 9588 6432 9640 6452
rect 9640 6432 9642 6452
rect 9494 4276 9550 4312
rect 9494 4256 9496 4276
rect 9496 4256 9548 4276
rect 9548 4256 9550 4276
rect 10046 7248 10102 7304
rect 11426 15000 11482 15056
rect 11150 14456 11206 14512
rect 11886 15408 11942 15464
rect 12254 17720 12310 17776
rect 12438 17856 12494 17912
rect 11978 14728 12034 14784
rect 12162 16224 12218 16280
rect 12714 18536 12770 18592
rect 10966 13504 11022 13560
rect 10966 12980 11022 13016
rect 10966 12960 10968 12980
rect 10968 12960 11020 12980
rect 11020 12960 11022 12980
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11610 13912 11666 13968
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10966 11192 11022 11248
rect 12070 14184 12126 14240
rect 12162 13640 12218 13696
rect 12346 14048 12402 14104
rect 12346 13776 12402 13832
rect 12162 12960 12218 13016
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11794 10920 11850 10976
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11702 10104 11758 10160
rect 11058 9868 11060 9888
rect 11060 9868 11112 9888
rect 11112 9868 11114 9888
rect 11058 9832 11114 9868
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11334 9560 11390 9616
rect 10414 8780 10416 8800
rect 10416 8780 10468 8800
rect 10468 8780 10470 8800
rect 10414 8744 10470 8780
rect 10322 8472 10378 8528
rect 10322 7928 10378 7984
rect 10322 7656 10378 7712
rect 10322 7520 10378 7576
rect 9862 5616 9918 5672
rect 10322 7248 10378 7304
rect 10322 6840 10378 6896
rect 10138 4936 10194 4992
rect 9494 3848 9550 3904
rect 9494 3304 9550 3360
rect 9678 2896 9734 2952
rect 10230 2896 10286 2952
rect 10414 4800 10470 4856
rect 10690 8472 10746 8528
rect 10874 8628 10930 8664
rect 10874 8608 10876 8628
rect 10876 8608 10928 8628
rect 10928 8608 10930 8628
rect 10598 4800 10654 4856
rect 10414 3576 10470 3632
rect 11610 9288 11666 9344
rect 11702 9152 11758 9208
rect 11334 8880 11390 8936
rect 11702 8880 11758 8936
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11334 7792 11390 7848
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 12070 11328 12126 11384
rect 12254 12144 12310 12200
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 12162 10104 12218 10160
rect 13174 19080 13230 19136
rect 13082 17856 13138 17912
rect 13542 20168 13598 20224
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 12714 14592 12770 14648
rect 12714 14184 12770 14240
rect 12622 12824 12678 12880
rect 12530 12688 12586 12744
rect 12530 12280 12586 12336
rect 12530 12180 12532 12200
rect 12532 12180 12584 12200
rect 12584 12180 12586 12200
rect 12530 12144 12586 12180
rect 12530 12008 12586 12064
rect 12162 9832 12218 9888
rect 12070 6976 12126 7032
rect 11334 5752 11390 5808
rect 11886 6316 11942 6352
rect 11886 6296 11888 6316
rect 11888 6296 11940 6316
rect 11940 6296 11942 6316
rect 12070 6840 12126 6896
rect 12070 6568 12126 6624
rect 12990 15000 13046 15056
rect 12806 12824 12862 12880
rect 12806 11892 12862 11928
rect 12806 11872 12808 11892
rect 12808 11872 12860 11892
rect 12860 11872 12862 11892
rect 12806 11500 12808 11520
rect 12808 11500 12860 11520
rect 12860 11500 12862 11520
rect 12806 11464 12862 11500
rect 12714 11192 12770 11248
rect 12438 8916 12440 8936
rect 12440 8916 12492 8936
rect 12492 8916 12494 8936
rect 12438 8880 12494 8916
rect 12530 8608 12586 8664
rect 12990 13812 12992 13832
rect 12992 13812 13044 13832
rect 13044 13812 13046 13832
rect 12990 13776 13046 13812
rect 13726 18944 13782 19000
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13818 18692 13874 18728
rect 13818 18672 13820 18692
rect 13820 18672 13872 18692
rect 13872 18672 13874 18692
rect 14554 21528 14610 21584
rect 14370 18808 14426 18864
rect 14370 18672 14426 18728
rect 13726 17992 13782 18048
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13634 17720 13690 17776
rect 13818 17756 13820 17776
rect 13820 17756 13872 17776
rect 13872 17756 13874 17776
rect 13818 17720 13874 17756
rect 13542 16904 13598 16960
rect 13266 15680 13322 15736
rect 13174 13368 13230 13424
rect 14278 17448 14334 17504
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 12990 12316 12992 12336
rect 12992 12316 13044 12336
rect 13044 12316 13046 12336
rect 12990 12280 13046 12316
rect 13450 13368 13506 13424
rect 13266 12688 13322 12744
rect 13266 12280 13322 12336
rect 13174 11464 13230 11520
rect 13082 10648 13138 10704
rect 13450 12552 13506 12608
rect 13818 15136 13874 15192
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 14738 19252 14740 19272
rect 14740 19252 14792 19272
rect 14792 19252 14794 19272
rect 14738 19216 14794 19252
rect 14738 19080 14794 19136
rect 14462 14764 14464 14784
rect 14464 14764 14516 14784
rect 14516 14764 14518 14784
rect 14462 14728 14518 14764
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13818 13504 13874 13560
rect 14370 13504 14426 13560
rect 13818 13252 13874 13288
rect 13818 13232 13820 13252
rect 13820 13232 13872 13252
rect 13872 13232 13874 13252
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13450 11636 13452 11656
rect 13452 11636 13504 11656
rect 13504 11636 13506 11656
rect 13450 11600 13506 11636
rect 14094 11600 14150 11656
rect 12990 9696 13046 9752
rect 13818 11464 13874 11520
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13634 10648 13690 10704
rect 13542 10376 13598 10432
rect 13818 10376 13874 10432
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13082 9152 13138 9208
rect 12898 8608 12954 8664
rect 12438 8084 12494 8120
rect 12438 8064 12440 8084
rect 12440 8064 12492 8084
rect 12492 8064 12494 8084
rect 12806 7928 12862 7984
rect 12806 7520 12862 7576
rect 13082 7928 13138 7984
rect 12254 6840 12310 6896
rect 12438 6740 12440 6760
rect 12440 6740 12492 6760
rect 12492 6740 12494 6760
rect 11794 5616 11850 5672
rect 11978 5636 12034 5672
rect 11978 5616 11980 5636
rect 11980 5616 12032 5636
rect 12032 5616 12034 5636
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11794 5344 11850 5400
rect 11610 4800 11666 4856
rect 11334 4528 11390 4584
rect 11150 4392 11206 4448
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11150 4256 11206 4312
rect 10414 1944 10470 2000
rect 10966 3168 11022 3224
rect 11150 3168 11206 3224
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12438 6704 12494 6740
rect 12898 6874 12954 6930
rect 13450 8780 13452 8800
rect 13452 8780 13504 8800
rect 13504 8780 13506 8800
rect 13450 8744 13506 8780
rect 13634 7792 13690 7848
rect 13450 7520 13506 7576
rect 12714 6296 12770 6352
rect 13082 6840 13138 6896
rect 13266 6568 13322 6624
rect 12162 5072 12218 5128
rect 12254 4800 12310 4856
rect 12622 5616 12678 5672
rect 12438 4936 12494 4992
rect 11886 3304 11942 3360
rect 11794 2760 11850 2816
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12346 4392 12402 4448
rect 12530 4528 12586 4584
rect 12254 4020 12256 4040
rect 12256 4020 12308 4040
rect 12308 4020 12310 4040
rect 12254 3984 12310 4020
rect 12162 3576 12218 3632
rect 12070 3168 12126 3224
rect 12438 3304 12494 3360
rect 12898 4820 12954 4856
rect 12898 4800 12900 4820
rect 12900 4800 12952 4820
rect 12952 4800 12954 4820
rect 12714 4528 12770 4584
rect 12622 3576 12678 3632
rect 13174 5888 13230 5944
rect 13174 5616 13230 5672
rect 13082 5208 13138 5264
rect 12990 3712 13046 3768
rect 13082 3576 13138 3632
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14462 12588 14464 12608
rect 14464 12588 14516 12608
rect 14516 12588 14518 12608
rect 14462 12552 14518 12588
rect 14370 12436 14426 12472
rect 14370 12416 14372 12436
rect 14372 12416 14424 12436
rect 14424 12416 14426 12436
rect 14370 9172 14426 9208
rect 14370 9152 14372 9172
rect 14372 9152 14424 9172
rect 14424 9152 14426 9172
rect 14278 9016 14334 9072
rect 15382 20576 15438 20632
rect 15290 20440 15346 20496
rect 15198 19216 15254 19272
rect 15382 19216 15438 19272
rect 15290 18536 15346 18592
rect 15014 14320 15070 14376
rect 14646 9424 14702 9480
rect 14186 8628 14242 8664
rect 14186 8608 14188 8628
rect 14188 8608 14240 8628
rect 14240 8608 14242 8628
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13450 6024 13506 6080
rect 13726 7112 13782 7168
rect 14646 9324 14648 9344
rect 14648 9324 14700 9344
rect 14700 9324 14702 9344
rect 14646 9288 14702 9324
rect 14646 8472 14702 8528
rect 14554 8372 14556 8392
rect 14556 8372 14608 8392
rect 14608 8372 14610 8392
rect 14554 8336 14610 8372
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13726 4256 13782 4312
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 14002 4664 14058 4720
rect 14094 4392 14150 4448
rect 13910 3984 13966 4040
rect 15750 18128 15806 18184
rect 15658 16244 15714 16280
rect 15658 16224 15660 16244
rect 15660 16224 15712 16244
rect 15712 16224 15714 16244
rect 15750 15136 15806 15192
rect 15474 14864 15530 14920
rect 15658 14048 15714 14104
rect 15566 13132 15568 13152
rect 15568 13132 15620 13152
rect 15620 13132 15622 13152
rect 15566 13096 15622 13132
rect 14922 9696 14978 9752
rect 15198 11192 15254 11248
rect 15198 10104 15254 10160
rect 15382 10004 15384 10024
rect 15384 10004 15436 10024
rect 15436 10004 15438 10024
rect 15382 9968 15438 10004
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 17958 22208 18014 22264
rect 17314 20848 17370 20904
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 20534 22616 20590 22672
rect 18878 20304 18934 20360
rect 19706 21800 19762 21856
rect 19430 20440 19486 20496
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 18050 19488 18106 19544
rect 18234 18964 18290 19000
rect 18234 18944 18236 18964
rect 18236 18944 18288 18964
rect 18288 18944 18290 18964
rect 17406 18572 17408 18592
rect 17408 18572 17460 18592
rect 17460 18572 17462 18592
rect 17406 18536 17462 18572
rect 18510 19352 18566 19408
rect 16854 17856 16910 17912
rect 16578 17720 16634 17776
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 15934 12844 15990 12880
rect 15934 12824 15936 12844
rect 15936 12824 15988 12844
rect 15988 12824 15990 12844
rect 15658 11056 15714 11112
rect 15566 10104 15622 10160
rect 15750 10512 15806 10568
rect 15474 9424 15530 9480
rect 14830 9152 14886 9208
rect 14830 7692 14832 7712
rect 14832 7692 14884 7712
rect 14884 7692 14886 7712
rect 14830 7656 14886 7692
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14738 5480 14794 5536
rect 14738 4700 14740 4720
rect 14740 4700 14792 4720
rect 14792 4700 14794 4720
rect 14738 4664 14794 4700
rect 14462 3984 14518 4040
rect 14370 3440 14426 3496
rect 14278 2896 14334 2952
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14646 3848 14702 3904
rect 14646 2624 14702 2680
rect 15382 9152 15438 9208
rect 14922 5888 14978 5944
rect 15382 8608 15438 8664
rect 15658 9716 15714 9752
rect 15658 9696 15660 9716
rect 15660 9696 15712 9716
rect 15712 9696 15714 9716
rect 15566 9288 15622 9344
rect 15198 8200 15254 8256
rect 15934 11192 15990 11248
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16394 15000 16450 15056
rect 16210 12552 16266 12608
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16578 13640 16634 13696
rect 16670 13232 16726 13288
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 17314 18264 17370 18320
rect 17130 15952 17186 16008
rect 17222 14456 17278 14512
rect 17222 14220 17224 14240
rect 17224 14220 17276 14240
rect 17276 14220 17278 14240
rect 17222 14184 17278 14220
rect 17222 14048 17278 14104
rect 17130 13812 17132 13832
rect 17132 13812 17184 13832
rect 17184 13812 17186 13832
rect 17130 13776 17186 13812
rect 17038 13232 17094 13288
rect 16762 12552 16818 12608
rect 16946 12416 17002 12472
rect 15842 7948 15898 7984
rect 15842 7928 15844 7948
rect 15844 7928 15896 7948
rect 15896 7928 15898 7948
rect 15198 7520 15254 7576
rect 15106 6024 15162 6080
rect 14922 5616 14978 5672
rect 14922 3304 14978 3360
rect 15106 3712 15162 3768
rect 15566 7112 15622 7168
rect 15658 6996 15714 7032
rect 16302 12008 16358 12064
rect 16302 11464 16358 11520
rect 16578 12144 16634 12200
rect 16762 12164 16818 12200
rect 16762 12144 16764 12164
rect 16764 12144 16816 12164
rect 16816 12144 16818 12164
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 17038 11872 17094 11928
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16210 9580 16266 9616
rect 16210 9560 16212 9580
rect 16212 9560 16264 9580
rect 16264 9560 16266 9580
rect 16118 8336 16174 8392
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16946 9560 17002 9616
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 15658 6976 15660 6996
rect 15660 6976 15712 6996
rect 15712 6976 15714 6996
rect 15658 6704 15714 6760
rect 15842 6604 15844 6624
rect 15844 6604 15896 6624
rect 15896 6604 15898 6624
rect 15842 6568 15898 6604
rect 15290 5752 15346 5808
rect 15658 5752 15714 5808
rect 15382 4256 15438 4312
rect 16118 6568 16174 6624
rect 16026 6432 16082 6488
rect 15750 5344 15806 5400
rect 15290 4120 15346 4176
rect 15382 3984 15438 4040
rect 15198 3032 15254 3088
rect 15474 3576 15530 3632
rect 15566 2916 15622 2952
rect 15566 2896 15568 2916
rect 15568 2896 15620 2916
rect 15620 2896 15622 2916
rect 15750 3984 15806 4040
rect 15934 3712 15990 3768
rect 15842 3576 15898 3632
rect 14922 1264 14978 1320
rect 17958 17856 18014 17912
rect 17774 17040 17830 17096
rect 17866 16652 17922 16688
rect 17866 16632 17868 16652
rect 17868 16632 17920 16652
rect 17920 16632 17922 16652
rect 17314 13368 17370 13424
rect 17590 13132 17592 13152
rect 17592 13132 17644 13152
rect 17644 13132 17646 13152
rect 17590 13096 17646 13132
rect 17314 12008 17370 12064
rect 17406 10240 17462 10296
rect 18510 18420 18566 18456
rect 18510 18400 18512 18420
rect 18512 18400 18564 18420
rect 18564 18400 18566 18420
rect 18510 18128 18566 18184
rect 18878 19796 18880 19816
rect 18880 19796 18932 19816
rect 18932 19796 18934 19816
rect 18878 19760 18934 19796
rect 18878 19352 18934 19408
rect 18694 18808 18750 18864
rect 19614 20032 19670 20088
rect 19154 19624 19210 19680
rect 19246 19216 19302 19272
rect 19614 19760 19670 19816
rect 19430 19352 19486 19408
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19430 18808 19486 18864
rect 18326 16124 18328 16144
rect 18328 16124 18380 16144
rect 18380 16124 18382 16144
rect 18326 16088 18382 16124
rect 18234 12552 18290 12608
rect 17406 9560 17462 9616
rect 16946 8336 17002 8392
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 17222 7520 17278 7576
rect 16670 7112 16726 7168
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16578 6316 16634 6352
rect 16578 6296 16580 6316
rect 16580 6296 16632 6316
rect 16632 6296 16634 6316
rect 16302 3440 16358 3496
rect 17130 7384 17186 7440
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16210 1944 16266 2000
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17406 6976 17462 7032
rect 17406 4800 17462 4856
rect 17958 8336 18014 8392
rect 17774 6296 17830 6352
rect 17958 6840 18014 6896
rect 18234 9288 18290 9344
rect 18234 7792 18290 7848
rect 17866 5616 17922 5672
rect 18050 5752 18106 5808
rect 18510 15272 18566 15328
rect 18694 14864 18750 14920
rect 18970 18128 19026 18184
rect 18878 16496 18934 16552
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19154 16496 19210 16552
rect 20166 19488 20222 19544
rect 20626 21392 20682 21448
rect 20350 19796 20352 19816
rect 20352 19796 20404 19816
rect 20404 19796 20406 19816
rect 20350 19760 20406 19796
rect 20534 20984 20590 21040
rect 20994 20576 21050 20632
rect 20810 20440 20866 20496
rect 20718 20032 20774 20088
rect 20534 19760 20590 19816
rect 20074 17720 20130 17776
rect 19522 16088 19578 16144
rect 19062 15952 19118 16008
rect 19614 15972 19670 16008
rect 19614 15952 19616 15972
rect 19616 15952 19668 15972
rect 19668 15952 19670 15972
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 18510 13232 18566 13288
rect 18418 12824 18474 12880
rect 18510 8508 18512 8528
rect 18512 8508 18564 8528
rect 18564 8508 18566 8528
rect 18510 8472 18566 8508
rect 18510 7112 18566 7168
rect 18510 6740 18512 6760
rect 18512 6740 18564 6760
rect 18564 6740 18566 6760
rect 18510 6704 18566 6740
rect 18694 13912 18750 13968
rect 19522 14320 19578 14376
rect 19890 16632 19946 16688
rect 20166 16224 20222 16280
rect 20534 17176 20590 17232
rect 20350 15972 20406 16008
rect 20350 15952 20352 15972
rect 20352 15952 20404 15972
rect 20404 15952 20406 15972
rect 20442 15816 20498 15872
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19522 13504 19578 13560
rect 19614 13404 19616 13424
rect 19616 13404 19668 13424
rect 19668 13404 19670 13424
rect 19614 13368 19670 13404
rect 18786 11464 18842 11520
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19614 12164 19670 12200
rect 19614 12144 19616 12164
rect 19616 12144 19668 12164
rect 19668 12144 19670 12164
rect 20074 13812 20076 13832
rect 20076 13812 20128 13832
rect 20128 13812 20130 13832
rect 20074 13776 20130 13812
rect 20074 13132 20076 13152
rect 20076 13132 20128 13152
rect 20128 13132 20130 13152
rect 19430 12008 19486 12064
rect 19798 12008 19854 12064
rect 19338 11892 19394 11928
rect 19338 11872 19340 11892
rect 19340 11872 19392 11892
rect 19392 11872 19394 11892
rect 19706 11872 19762 11928
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 18602 6024 18658 6080
rect 18418 5752 18474 5808
rect 18602 5208 18658 5264
rect 18326 4664 18382 4720
rect 17958 3304 18014 3360
rect 17866 2760 17922 2816
rect 18234 2760 18290 2816
rect 18970 9968 19026 10024
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19430 10004 19432 10024
rect 19432 10004 19484 10024
rect 19484 10004 19486 10024
rect 19430 9968 19486 10004
rect 19614 10512 19670 10568
rect 19154 9560 19210 9616
rect 19062 9424 19118 9480
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19246 9016 19302 9072
rect 18970 8064 19026 8120
rect 18878 7384 18934 7440
rect 18786 7248 18842 7304
rect 20074 13096 20130 13132
rect 20258 12416 20314 12472
rect 19890 11600 19946 11656
rect 19706 10124 19762 10160
rect 19706 10104 19708 10124
rect 19708 10104 19760 10124
rect 19760 10104 19762 10124
rect 19890 9968 19946 10024
rect 19798 9696 19854 9752
rect 19890 9016 19946 9072
rect 19614 8608 19670 8664
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19246 7540 19302 7576
rect 19246 7520 19248 7540
rect 19248 7520 19300 7540
rect 19300 7520 19302 7540
rect 20442 13932 20498 13968
rect 20442 13912 20444 13932
rect 20444 13912 20496 13932
rect 20496 13912 20498 13932
rect 20810 16632 20866 16688
rect 20166 11056 20222 11112
rect 20350 10648 20406 10704
rect 20258 10512 20314 10568
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18970 6296 19026 6352
rect 19430 6160 19486 6216
rect 19522 6024 19578 6080
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19522 5616 19578 5672
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19338 4664 19394 4720
rect 18694 3168 18750 3224
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19706 3712 19762 3768
rect 18418 2488 18474 2544
rect 18970 2760 19026 2816
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19706 3596 19762 3632
rect 19706 3576 19708 3596
rect 19708 3576 19760 3596
rect 19760 3576 19762 3596
rect 19890 4120 19946 4176
rect 19614 3168 19670 3224
rect 19246 1400 19302 1456
rect 18694 856 18750 912
rect 20718 12008 20774 12064
rect 20810 11872 20866 11928
rect 20810 11736 20866 11792
rect 21638 19896 21694 19952
rect 21454 18808 21510 18864
rect 21546 18400 21602 18456
rect 21454 17992 21510 18048
rect 21086 16224 21142 16280
rect 21086 15408 21142 15464
rect 21454 17584 21510 17640
rect 21454 16768 21510 16824
rect 21454 16224 21510 16280
rect 21454 15852 21456 15872
rect 21456 15852 21508 15872
rect 21508 15852 21510 15872
rect 21454 15816 21510 15852
rect 21454 15000 21510 15056
rect 21454 14592 21510 14648
rect 21454 14220 21456 14240
rect 21456 14220 21508 14240
rect 21508 14220 21510 14240
rect 21454 14184 21510 14220
rect 21086 13776 21142 13832
rect 21638 13504 21694 13560
rect 21454 13368 21510 13424
rect 20810 11056 20866 11112
rect 20534 9016 20590 9072
rect 20350 5208 20406 5264
rect 20258 4020 20260 4040
rect 20260 4020 20312 4040
rect 20312 4020 20314 4040
rect 20258 3984 20314 4020
rect 20166 3168 20222 3224
rect 20718 8608 20774 8664
rect 20718 8200 20774 8256
rect 20718 7812 20774 7848
rect 20718 7792 20720 7812
rect 20720 7792 20772 7812
rect 20772 7792 20774 7812
rect 21086 10784 21142 10840
rect 20994 10376 21050 10432
rect 20994 10240 21050 10296
rect 21086 10124 21142 10160
rect 21086 10104 21088 10124
rect 21088 10104 21140 10124
rect 21140 10104 21142 10124
rect 21454 12824 21510 12880
rect 21270 11872 21326 11928
rect 21454 12416 21510 12472
rect 21454 12280 21510 12336
rect 21454 12044 21456 12064
rect 21456 12044 21508 12064
rect 21508 12044 21510 12064
rect 21454 12008 21510 12044
rect 21546 11636 21548 11656
rect 21548 11636 21600 11656
rect 21600 11636 21602 11656
rect 21546 11600 21602 11636
rect 21546 11328 21602 11384
rect 21454 11192 21510 11248
rect 21086 9968 21142 10024
rect 20994 9696 21050 9752
rect 20626 6296 20682 6352
rect 20626 4528 20682 4584
rect 21178 9832 21234 9888
rect 21086 6860 21142 6896
rect 21086 6840 21088 6860
rect 21088 6840 21140 6860
rect 21140 6840 21142 6860
rect 20994 6432 21050 6488
rect 20994 5480 21050 5536
rect 19614 176 19670 232
rect 20718 2624 20774 2680
rect 21454 10376 21510 10432
rect 21270 8608 21326 8664
rect 21362 8084 21418 8120
rect 21362 8064 21364 8084
rect 21364 8064 21416 8084
rect 21416 8064 21418 8084
rect 21638 8200 21694 8256
rect 22282 16496 22338 16552
rect 21822 14320 21878 14376
rect 21822 7792 21878 7848
rect 21454 6432 21510 6488
rect 21454 3440 21510 3496
rect 20718 992 20774 1048
rect 21638 3984 21694 4040
rect 22006 7012 22008 7032
rect 22008 7012 22060 7032
rect 22060 7012 22062 7032
rect 22006 6976 22062 7012
rect 21914 4800 21970 4856
rect 22006 4392 22062 4448
rect 22006 3032 22062 3088
rect 21914 2896 21970 2952
rect 21730 2352 21786 2408
rect 21546 2216 21602 2272
rect 21822 1844 21824 1864
rect 21824 1844 21876 1864
rect 21876 1844 21878 1864
rect 21822 1808 21878 1844
rect 22282 3304 22338 3360
<< metal3 >>
rect 289 22946 355 22949
rect 16982 22946 16988 22948
rect 289 22944 16988 22946
rect 289 22888 294 22944
rect 350 22888 16988 22944
rect 289 22886 16988 22888
rect 289 22883 355 22886
rect 16982 22884 16988 22886
rect 17052 22884 17058 22948
rect 974 22748 980 22812
rect 1044 22810 1050 22812
rect 7741 22810 7807 22813
rect 1044 22808 7807 22810
rect 1044 22752 7746 22808
rect 7802 22752 7807 22808
rect 1044 22750 7807 22752
rect 1044 22748 1050 22750
rect 7741 22747 7807 22750
rect 0 22674 800 22704
rect 2405 22674 2471 22677
rect 0 22672 2471 22674
rect 0 22616 2410 22672
rect 2466 22616 2471 22672
rect 0 22614 2471 22616
rect 0 22584 800 22614
rect 2405 22611 2471 22614
rect 6862 22612 6868 22676
rect 6932 22674 6938 22676
rect 20529 22674 20595 22677
rect 22200 22674 23000 22704
rect 6932 22614 12450 22674
rect 6932 22612 6938 22614
rect 1025 22538 1091 22541
rect 12390 22538 12450 22614
rect 20529 22672 23000 22674
rect 20529 22616 20534 22672
rect 20590 22616 23000 22672
rect 20529 22614 23000 22616
rect 20529 22611 20595 22614
rect 22200 22584 23000 22614
rect 19926 22538 19932 22540
rect 1025 22536 7666 22538
rect 1025 22480 1030 22536
rect 1086 22480 7666 22536
rect 1025 22478 7666 22480
rect 12390 22478 19932 22538
rect 1025 22475 1091 22478
rect 1117 22402 1183 22405
rect 7606 22402 7666 22478
rect 19926 22476 19932 22478
rect 19996 22476 20002 22540
rect 14406 22402 14412 22404
rect 1117 22400 7482 22402
rect 1117 22344 1122 22400
rect 1178 22344 7482 22400
rect 1117 22342 7482 22344
rect 7606 22342 14412 22402
rect 1117 22339 1183 22342
rect 0 22266 800 22296
rect 4153 22266 4219 22269
rect 0 22264 4219 22266
rect 0 22208 4158 22264
rect 4214 22208 4219 22264
rect 0 22206 4219 22208
rect 7422 22266 7482 22342
rect 14406 22340 14412 22342
rect 14476 22340 14482 22404
rect 15326 22266 15332 22268
rect 7422 22206 15332 22266
rect 0 22176 800 22206
rect 4153 22203 4219 22206
rect 15326 22204 15332 22206
rect 15396 22204 15402 22268
rect 17953 22266 18019 22269
rect 22200 22266 23000 22296
rect 17953 22264 23000 22266
rect 17953 22208 17958 22264
rect 18014 22208 23000 22264
rect 17953 22206 23000 22208
rect 17953 22203 18019 22206
rect 22200 22176 23000 22206
rect 974 22068 980 22132
rect 1044 22130 1050 22132
rect 7741 22130 7807 22133
rect 13670 22130 13676 22132
rect 1044 22070 7666 22130
rect 1044 22068 1050 22070
rect 1025 21994 1091 21997
rect 7465 21994 7531 21997
rect 1025 21992 7531 21994
rect 1025 21936 1030 21992
rect 1086 21936 7470 21992
rect 7526 21936 7531 21992
rect 1025 21934 7531 21936
rect 7606 21994 7666 22070
rect 7741 22128 13676 22130
rect 7741 22072 7746 22128
rect 7802 22072 13676 22128
rect 7741 22070 13676 22072
rect 7741 22067 7807 22070
rect 13670 22068 13676 22070
rect 13740 22068 13746 22132
rect 14590 21994 14596 21996
rect 7606 21934 14596 21994
rect 1025 21931 1091 21934
rect 7465 21931 7531 21934
rect 14590 21932 14596 21934
rect 14660 21932 14666 21996
rect 0 21858 800 21888
rect 2221 21858 2287 21861
rect 18086 21858 18092 21860
rect 0 21856 2287 21858
rect 0 21800 2226 21856
rect 2282 21800 2287 21856
rect 0 21798 2287 21800
rect 0 21768 800 21798
rect 2221 21795 2287 21798
rect 2730 21798 18092 21858
rect 2313 21722 2379 21725
rect 2730 21722 2790 21798
rect 18086 21796 18092 21798
rect 18156 21796 18162 21860
rect 19701 21858 19767 21861
rect 22200 21858 23000 21888
rect 19701 21856 23000 21858
rect 19701 21800 19706 21856
rect 19762 21800 23000 21856
rect 19701 21798 23000 21800
rect 19701 21795 19767 21798
rect 22200 21768 23000 21798
rect 2313 21720 2790 21722
rect 2313 21664 2318 21720
rect 2374 21664 2790 21720
rect 2313 21662 2790 21664
rect 7465 21722 7531 21725
rect 15142 21722 15148 21724
rect 7465 21720 15148 21722
rect 7465 21664 7470 21720
rect 7526 21664 15148 21720
rect 7465 21662 15148 21664
rect 2313 21659 2379 21662
rect 7465 21659 7531 21662
rect 15142 21660 15148 21662
rect 15212 21660 15218 21724
rect 1526 21524 1532 21588
rect 1596 21586 1602 21588
rect 14549 21586 14615 21589
rect 1596 21584 14615 21586
rect 1596 21528 14554 21584
rect 14610 21528 14615 21584
rect 1596 21526 14615 21528
rect 1596 21524 1602 21526
rect 14549 21523 14615 21526
rect 0 21450 800 21480
rect 2497 21450 2563 21453
rect 0 21448 2563 21450
rect 0 21392 2502 21448
rect 2558 21392 2563 21448
rect 0 21390 2563 21392
rect 0 21360 800 21390
rect 2497 21387 2563 21390
rect 4654 21388 4660 21452
rect 4724 21450 4730 21452
rect 17902 21450 17908 21452
rect 4724 21390 17908 21450
rect 4724 21388 4730 21390
rect 17902 21388 17908 21390
rect 17972 21388 17978 21452
rect 20621 21450 20687 21453
rect 22200 21450 23000 21480
rect 20621 21448 23000 21450
rect 20621 21392 20626 21448
rect 20682 21392 23000 21448
rect 20621 21390 23000 21392
rect 20621 21387 20687 21390
rect 22200 21360 23000 21390
rect 1158 21252 1164 21316
rect 1228 21314 1234 21316
rect 13486 21314 13492 21316
rect 1228 21254 13492 21314
rect 1228 21252 1234 21254
rect 13486 21252 13492 21254
rect 13556 21252 13562 21316
rect 3417 21178 3483 21181
rect 18454 21178 18460 21180
rect 3417 21176 18460 21178
rect 3417 21120 3422 21176
rect 3478 21120 18460 21176
rect 3417 21118 18460 21120
rect 3417 21115 3483 21118
rect 18454 21116 18460 21118
rect 18524 21116 18530 21180
rect 0 21042 800 21072
rect 1761 21042 1827 21045
rect 17166 21042 17172 21044
rect 0 21040 1827 21042
rect 0 20984 1766 21040
rect 1822 20984 1827 21040
rect 0 20982 1827 20984
rect 0 20952 800 20982
rect 1761 20979 1827 20982
rect 1902 20982 17172 21042
rect 1209 20906 1275 20909
rect 1902 20906 1962 20982
rect 17166 20980 17172 20982
rect 17236 20980 17242 21044
rect 20529 21042 20595 21045
rect 22200 21042 23000 21072
rect 20529 21040 23000 21042
rect 20529 20984 20534 21040
rect 20590 20984 23000 21040
rect 20529 20982 23000 20984
rect 20529 20979 20595 20982
rect 22200 20952 23000 20982
rect 1209 20904 1962 20906
rect 1209 20848 1214 20904
rect 1270 20848 1962 20904
rect 1209 20846 1962 20848
rect 1209 20843 1275 20846
rect 2630 20844 2636 20908
rect 2700 20906 2706 20908
rect 17309 20906 17375 20909
rect 2700 20904 17375 20906
rect 2700 20848 17314 20904
rect 17370 20848 17375 20904
rect 2700 20846 17375 20848
rect 2700 20844 2706 20846
rect 17309 20843 17375 20846
rect 6142 20704 6462 20705
rect 0 20634 800 20664
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 20639 16858 20640
rect 2865 20634 2931 20637
rect 0 20632 2931 20634
rect 0 20576 2870 20632
rect 2926 20576 2931 20632
rect 0 20574 2931 20576
rect 0 20544 800 20574
rect 2865 20571 2931 20574
rect 6545 20634 6611 20637
rect 9857 20634 9923 20637
rect 15377 20634 15443 20637
rect 6545 20632 9923 20634
rect 6545 20576 6550 20632
rect 6606 20576 9862 20632
rect 9918 20576 9923 20632
rect 6545 20574 9923 20576
rect 6545 20571 6611 20574
rect 9857 20571 9923 20574
rect 11838 20632 15443 20634
rect 11838 20576 15382 20632
rect 15438 20576 15443 20632
rect 11838 20574 15443 20576
rect 6545 20498 6611 20501
rect 11838 20498 11898 20574
rect 15377 20571 15443 20574
rect 20989 20634 21055 20637
rect 22200 20634 23000 20664
rect 20989 20632 23000 20634
rect 20989 20576 20994 20632
rect 21050 20576 23000 20632
rect 20989 20574 23000 20576
rect 20989 20571 21055 20574
rect 22200 20544 23000 20574
rect 15285 20498 15351 20501
rect 6545 20496 11898 20498
rect 6545 20440 6550 20496
rect 6606 20440 11898 20496
rect 6545 20438 11898 20440
rect 12390 20496 15351 20498
rect 12390 20440 15290 20496
rect 15346 20440 15351 20496
rect 12390 20438 15351 20440
rect 6545 20435 6611 20438
rect 2037 20362 2103 20365
rect 8385 20362 8451 20365
rect 9857 20362 9923 20365
rect 12390 20362 12450 20438
rect 15285 20435 15351 20438
rect 19425 20498 19491 20501
rect 20805 20498 20871 20501
rect 19425 20496 20871 20498
rect 19425 20440 19430 20496
rect 19486 20440 20810 20496
rect 20866 20440 20871 20496
rect 19425 20438 20871 20440
rect 19425 20435 19491 20438
rect 20805 20435 20871 20438
rect 2037 20360 8451 20362
rect 2037 20304 2042 20360
rect 2098 20304 8390 20360
rect 8446 20304 8451 20360
rect 2037 20302 8451 20304
rect 2037 20299 2103 20302
rect 8385 20299 8451 20302
rect 8526 20302 9322 20362
rect 0 20226 800 20256
rect 1577 20226 1643 20229
rect 4797 20226 4863 20229
rect 6269 20226 6335 20229
rect 0 20224 1643 20226
rect 0 20168 1582 20224
rect 1638 20168 1643 20224
rect 0 20166 1643 20168
rect 0 20136 800 20166
rect 1577 20163 1643 20166
rect 3926 20224 6335 20226
rect 3926 20168 4802 20224
rect 4858 20168 6274 20224
rect 6330 20168 6335 20224
rect 3926 20166 6335 20168
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 3926 19954 3986 20166
rect 4797 20163 4863 20166
rect 6269 20163 6335 20166
rect 6453 20226 6519 20229
rect 6678 20226 6684 20228
rect 6453 20224 6684 20226
rect 6453 20168 6458 20224
rect 6514 20168 6684 20224
rect 6453 20166 6684 20168
rect 6453 20163 6519 20166
rect 6678 20164 6684 20166
rect 6748 20164 6754 20228
rect 7414 20164 7420 20228
rect 7484 20226 7490 20228
rect 8526 20226 8586 20302
rect 7484 20166 8586 20226
rect 9262 20226 9322 20302
rect 9857 20360 12450 20362
rect 9857 20304 9862 20360
rect 9918 20304 12450 20360
rect 9857 20302 12450 20304
rect 18873 20362 18939 20365
rect 18873 20360 19626 20362
rect 18873 20304 18878 20360
rect 18934 20304 19626 20360
rect 18873 20302 19626 20304
rect 9857 20299 9923 20302
rect 18873 20299 18939 20302
rect 10961 20226 11027 20229
rect 13537 20226 13603 20229
rect 9262 20224 13603 20226
rect 9262 20168 10966 20224
rect 11022 20168 13542 20224
rect 13598 20168 13603 20224
rect 9262 20166 13603 20168
rect 19566 20226 19626 20302
rect 22200 20226 23000 20256
rect 19566 20166 23000 20226
rect 7484 20164 7490 20166
rect 10961 20163 11027 20166
rect 13537 20163 13603 20166
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 22200 20136 23000 20166
rect 19137 20095 19457 20096
rect 4981 20090 5047 20093
rect 7782 20090 7788 20092
rect 4981 20088 7788 20090
rect 4981 20032 4986 20088
rect 5042 20032 7788 20088
rect 4981 20030 7788 20032
rect 4981 20027 5047 20030
rect 7782 20028 7788 20030
rect 7852 20028 7858 20092
rect 9213 20090 9279 20093
rect 9622 20090 9628 20092
rect 9213 20088 9628 20090
rect 9213 20032 9218 20088
rect 9274 20032 9628 20088
rect 9213 20030 9628 20032
rect 9213 20027 9279 20030
rect 9622 20028 9628 20030
rect 9692 20028 9698 20092
rect 10133 20090 10199 20093
rect 11973 20090 12039 20093
rect 10133 20088 12039 20090
rect 10133 20032 10138 20088
rect 10194 20032 11978 20088
rect 12034 20032 12039 20088
rect 10133 20030 12039 20032
rect 10133 20027 10199 20030
rect 11973 20027 12039 20030
rect 12198 20028 12204 20092
rect 12268 20090 12274 20092
rect 12433 20090 12499 20093
rect 12268 20088 12499 20090
rect 12268 20032 12438 20088
rect 12494 20032 12499 20088
rect 12268 20030 12499 20032
rect 12268 20028 12274 20030
rect 12433 20027 12499 20030
rect 19609 20090 19675 20093
rect 20713 20090 20779 20093
rect 19609 20088 20779 20090
rect 19609 20032 19614 20088
rect 19670 20032 20718 20088
rect 20774 20032 20779 20088
rect 19609 20030 20779 20032
rect 19609 20027 19675 20030
rect 20713 20027 20779 20030
rect 2730 19894 3986 19954
rect 4429 19954 4495 19957
rect 8109 19954 8175 19957
rect 4429 19952 8175 19954
rect 4429 19896 4434 19952
rect 4490 19896 8114 19952
rect 8170 19896 8175 19952
rect 4429 19894 8175 19896
rect 1485 19818 1551 19821
rect 2730 19818 2790 19894
rect 4429 19891 4495 19894
rect 8109 19891 8175 19894
rect 8569 19954 8635 19957
rect 21633 19954 21699 19957
rect 8569 19952 21699 19954
rect 8569 19896 8574 19952
rect 8630 19896 21638 19952
rect 21694 19896 21699 19952
rect 8569 19894 21699 19896
rect 8569 19891 8635 19894
rect 21633 19891 21699 19894
rect 1485 19816 2790 19818
rect 1485 19760 1490 19816
rect 1546 19760 2790 19816
rect 1485 19758 2790 19760
rect 3325 19820 3391 19821
rect 3325 19816 3372 19820
rect 3436 19818 3442 19820
rect 7189 19818 7255 19821
rect 10593 19818 10659 19821
rect 3325 19760 3330 19816
rect 1485 19755 1551 19758
rect 3325 19756 3372 19760
rect 3436 19758 3482 19818
rect 5950 19816 7255 19818
rect 5950 19760 7194 19816
rect 7250 19760 7255 19816
rect 5950 19758 7255 19760
rect 3436 19756 3442 19758
rect 3325 19755 3391 19756
rect 0 19682 800 19712
rect 1485 19682 1551 19685
rect 0 19680 1551 19682
rect 0 19624 1490 19680
rect 1546 19624 1551 19680
rect 0 19622 1551 19624
rect 0 19592 800 19622
rect 1485 19619 1551 19622
rect 1945 19682 2011 19685
rect 4429 19682 4495 19685
rect 1945 19680 4495 19682
rect 1945 19624 1950 19680
rect 2006 19624 4434 19680
rect 4490 19624 4495 19680
rect 1945 19622 4495 19624
rect 1945 19619 2011 19622
rect 4429 19619 4495 19622
rect 5950 19546 6010 19758
rect 7189 19755 7255 19758
rect 7974 19816 10659 19818
rect 7974 19760 10598 19816
rect 10654 19760 10659 19816
rect 7974 19758 10659 19760
rect 7097 19682 7163 19685
rect 7974 19682 8034 19758
rect 10593 19755 10659 19758
rect 10777 19818 10843 19821
rect 13118 19818 13124 19820
rect 10777 19816 13124 19818
rect 10777 19760 10782 19816
rect 10838 19760 13124 19816
rect 10777 19758 13124 19760
rect 10777 19755 10843 19758
rect 13118 19756 13124 19758
rect 13188 19756 13194 19820
rect 18873 19818 18939 19821
rect 19609 19818 19675 19821
rect 18873 19816 19675 19818
rect 18873 19760 18878 19816
rect 18934 19760 19614 19816
rect 19670 19760 19675 19816
rect 18873 19758 19675 19760
rect 18873 19755 18939 19758
rect 19609 19755 19675 19758
rect 20345 19818 20411 19821
rect 20529 19818 20595 19821
rect 20345 19816 20595 19818
rect 20345 19760 20350 19816
rect 20406 19760 20534 19816
rect 20590 19760 20595 19816
rect 20345 19758 20595 19760
rect 20345 19755 20411 19758
rect 20529 19755 20595 19758
rect 7097 19680 8034 19682
rect 7097 19624 7102 19680
rect 7158 19624 8034 19680
rect 7097 19622 8034 19624
rect 8109 19682 8175 19685
rect 11145 19682 11211 19685
rect 8109 19680 11211 19682
rect 8109 19624 8114 19680
rect 8170 19624 11150 19680
rect 11206 19624 11211 19680
rect 8109 19622 11211 19624
rect 7097 19619 7163 19622
rect 8109 19619 8175 19622
rect 11145 19619 11211 19622
rect 19149 19682 19215 19685
rect 22200 19682 23000 19712
rect 19149 19680 23000 19682
rect 19149 19624 19154 19680
rect 19210 19624 23000 19680
rect 19149 19622 23000 19624
rect 19149 19619 19215 19622
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 22200 19592 23000 19622
rect 16538 19551 16858 19552
rect 2730 19486 6010 19546
rect 7097 19546 7163 19549
rect 8937 19546 9003 19549
rect 7097 19544 9003 19546
rect 7097 19488 7102 19544
rect 7158 19488 8942 19544
rect 8998 19488 9003 19544
rect 7097 19486 9003 19488
rect 1945 19410 2011 19413
rect 2730 19410 2790 19486
rect 7097 19483 7163 19486
rect 8937 19483 9003 19486
rect 9121 19546 9187 19549
rect 18045 19546 18111 19549
rect 20161 19546 20227 19549
rect 9121 19544 10794 19546
rect 9121 19488 9126 19544
rect 9182 19488 10794 19544
rect 9121 19486 10794 19488
rect 9121 19483 9187 19486
rect 1945 19408 2790 19410
rect 1945 19352 1950 19408
rect 2006 19352 2790 19408
rect 1945 19350 2790 19352
rect 4153 19410 4219 19413
rect 7966 19410 7972 19412
rect 4153 19408 7972 19410
rect 4153 19352 4158 19408
rect 4214 19352 7972 19408
rect 4153 19350 7972 19352
rect 1945 19347 2011 19350
rect 4153 19347 4219 19350
rect 7966 19348 7972 19350
rect 8036 19348 8042 19412
rect 8661 19410 8727 19413
rect 9949 19412 10015 19413
rect 10317 19412 10383 19413
rect 9438 19410 9444 19412
rect 8661 19408 9444 19410
rect 8661 19352 8666 19408
rect 8722 19352 9444 19408
rect 8661 19350 9444 19352
rect 8661 19347 8727 19350
rect 9438 19348 9444 19350
rect 9508 19348 9514 19412
rect 9949 19408 9996 19412
rect 10060 19410 10066 19412
rect 9949 19352 9954 19408
rect 9949 19348 9996 19352
rect 10060 19350 10106 19410
rect 10317 19408 10364 19412
rect 10428 19410 10434 19412
rect 10734 19410 10794 19486
rect 18045 19544 20227 19546
rect 18045 19488 18050 19544
rect 18106 19488 20166 19544
rect 20222 19488 20227 19544
rect 18045 19486 20227 19488
rect 18045 19483 18111 19486
rect 20161 19483 20227 19486
rect 12525 19410 12591 19413
rect 10317 19352 10322 19408
rect 10060 19348 10066 19350
rect 10317 19348 10364 19352
rect 10428 19350 10474 19410
rect 10734 19408 12591 19410
rect 10734 19352 12530 19408
rect 12586 19352 12591 19408
rect 10734 19350 12591 19352
rect 10428 19348 10434 19350
rect 9949 19347 10015 19348
rect 10317 19347 10383 19348
rect 12525 19347 12591 19350
rect 18505 19410 18571 19413
rect 18873 19410 18939 19413
rect 18505 19408 18939 19410
rect 18505 19352 18510 19408
rect 18566 19352 18878 19408
rect 18934 19352 18939 19408
rect 18505 19350 18939 19352
rect 18505 19347 18571 19350
rect 18873 19347 18939 19350
rect 19425 19410 19491 19413
rect 19558 19410 19564 19412
rect 19425 19408 19564 19410
rect 19425 19352 19430 19408
rect 19486 19352 19564 19408
rect 19425 19350 19564 19352
rect 19425 19347 19491 19350
rect 19558 19348 19564 19350
rect 19628 19348 19634 19412
rect 0 19274 800 19304
rect 1853 19274 1919 19277
rect 0 19272 1919 19274
rect 0 19216 1858 19272
rect 1914 19216 1919 19272
rect 0 19214 1919 19216
rect 0 19184 800 19214
rect 1853 19211 1919 19214
rect 2313 19274 2379 19277
rect 2630 19274 2636 19276
rect 2313 19272 2636 19274
rect 2313 19216 2318 19272
rect 2374 19216 2636 19272
rect 2313 19214 2636 19216
rect 2313 19211 2379 19214
rect 2630 19212 2636 19214
rect 2700 19212 2706 19276
rect 3049 19274 3115 19277
rect 6913 19274 6979 19277
rect 10133 19274 10199 19277
rect 3049 19272 6979 19274
rect 3049 19216 3054 19272
rect 3110 19216 6918 19272
rect 6974 19216 6979 19272
rect 3049 19214 6979 19216
rect 3049 19211 3115 19214
rect 6913 19211 6979 19214
rect 7054 19272 10199 19274
rect 7054 19216 10138 19272
rect 10194 19216 10199 19272
rect 7054 19214 10199 19216
rect 5809 19138 5875 19141
rect 7054 19138 7114 19214
rect 10133 19211 10199 19214
rect 10409 19274 10475 19277
rect 14733 19274 14799 19277
rect 15193 19276 15259 19277
rect 15377 19276 15443 19277
rect 15142 19274 15148 19276
rect 10409 19272 14799 19274
rect 10409 19216 10414 19272
rect 10470 19216 14738 19272
rect 14794 19216 14799 19272
rect 10409 19214 14799 19216
rect 15102 19214 15148 19274
rect 15212 19272 15259 19276
rect 15254 19216 15259 19272
rect 10409 19211 10475 19214
rect 14733 19211 14799 19214
rect 15142 19212 15148 19214
rect 15212 19212 15259 19216
rect 15326 19212 15332 19276
rect 15396 19274 15443 19276
rect 19241 19274 19307 19277
rect 22200 19274 23000 19304
rect 15396 19272 15488 19274
rect 15438 19216 15488 19272
rect 15396 19214 15488 19216
rect 19241 19272 23000 19274
rect 19241 19216 19246 19272
rect 19302 19216 23000 19272
rect 19241 19214 23000 19216
rect 15396 19212 15443 19214
rect 15193 19211 15259 19212
rect 15377 19211 15443 19212
rect 19241 19211 19307 19214
rect 22200 19184 23000 19214
rect 5809 19136 7114 19138
rect 5809 19080 5814 19136
rect 5870 19080 7114 19136
rect 5809 19078 7114 19080
rect 8109 19136 8175 19141
rect 8109 19080 8114 19136
rect 8170 19080 8175 19136
rect 5809 19075 5875 19078
rect 8109 19075 8175 19080
rect 10961 19138 11027 19141
rect 13169 19138 13235 19141
rect 10961 19136 13235 19138
rect 10961 19080 10966 19136
rect 11022 19080 13174 19136
rect 13230 19080 13235 19136
rect 10961 19078 13235 19080
rect 10961 19075 11027 19078
rect 13169 19075 13235 19078
rect 14590 19076 14596 19140
rect 14660 19138 14666 19140
rect 14733 19138 14799 19141
rect 14660 19136 14799 19138
rect 14660 19080 14738 19136
rect 14794 19080 14799 19136
rect 14660 19078 14799 19080
rect 14660 19076 14666 19078
rect 14733 19075 14799 19078
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 1301 19002 1367 19005
rect 4153 19002 4219 19005
rect 8112 19002 8172 19075
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 1301 19000 1732 19002
rect 1301 18944 1306 19000
rect 1362 18944 1732 19000
rect 1301 18942 1732 18944
rect 1301 18939 1367 18942
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 1672 18866 1732 18942
rect 4153 19000 8172 19002
rect 4153 18944 4158 19000
rect 4214 18944 8172 19000
rect 4153 18942 8172 18944
rect 4153 18939 4219 18942
rect 9254 18940 9260 19004
rect 9324 19002 9330 19004
rect 9489 19002 9555 19005
rect 9324 19000 9555 19002
rect 9324 18944 9494 19000
rect 9550 18944 9555 19000
rect 9324 18942 9555 18944
rect 9324 18940 9330 18942
rect 9489 18939 9555 18942
rect 9857 19002 9923 19005
rect 10317 19002 10383 19005
rect 9857 19000 10383 19002
rect 9857 18944 9862 19000
rect 9918 18944 10322 19000
rect 10378 18944 10383 19000
rect 9857 18942 10383 18944
rect 9857 18939 9923 18942
rect 10317 18939 10383 18942
rect 11145 19002 11211 19005
rect 13721 19002 13787 19005
rect 11145 19000 13787 19002
rect 11145 18944 11150 19000
rect 11206 18944 13726 19000
rect 13782 18944 13787 19000
rect 11145 18942 13787 18944
rect 11145 18939 11211 18942
rect 13721 18939 13787 18942
rect 18086 18940 18092 19004
rect 18156 19002 18162 19004
rect 18229 19002 18295 19005
rect 18156 19000 18295 19002
rect 18156 18944 18234 19000
rect 18290 18944 18295 19000
rect 18156 18942 18295 18944
rect 18156 18940 18162 18942
rect 18229 18939 18295 18942
rect 14365 18866 14431 18869
rect 1672 18806 9460 18866
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 1577 18730 1643 18733
rect 8477 18730 8543 18733
rect 1577 18728 8543 18730
rect 1577 18672 1582 18728
rect 1638 18672 8482 18728
rect 8538 18672 8543 18728
rect 1577 18670 8543 18672
rect 9400 18730 9460 18806
rect 9998 18864 14431 18866
rect 9998 18808 14370 18864
rect 14426 18808 14431 18864
rect 9998 18806 14431 18808
rect 9806 18730 9812 18732
rect 9400 18670 9812 18730
rect 1577 18667 1643 18670
rect 8477 18667 8543 18670
rect 9806 18668 9812 18670
rect 9876 18668 9882 18732
rect 2865 18596 2931 18597
rect 2814 18594 2820 18596
rect 2774 18534 2820 18594
rect 2884 18592 2931 18596
rect 2926 18536 2931 18592
rect 2814 18532 2820 18534
rect 2884 18532 2931 18536
rect 2865 18531 2931 18532
rect 3785 18594 3851 18597
rect 5206 18594 5212 18596
rect 3785 18592 5212 18594
rect 3785 18536 3790 18592
rect 3846 18536 5212 18592
rect 3785 18534 5212 18536
rect 3785 18531 3851 18534
rect 5206 18532 5212 18534
rect 5276 18532 5282 18596
rect 5441 18594 5507 18597
rect 5625 18596 5691 18597
rect 5574 18594 5580 18596
rect 5441 18592 5580 18594
rect 5644 18594 5691 18596
rect 6729 18594 6795 18597
rect 9998 18594 10058 18806
rect 14365 18803 14431 18806
rect 18689 18866 18755 18869
rect 19425 18866 19491 18869
rect 18689 18864 19491 18866
rect 18689 18808 18694 18864
rect 18750 18808 19430 18864
rect 19486 18808 19491 18864
rect 18689 18806 19491 18808
rect 18689 18803 18755 18806
rect 19425 18803 19491 18806
rect 21449 18866 21515 18869
rect 22200 18866 23000 18896
rect 21449 18864 23000 18866
rect 21449 18808 21454 18864
rect 21510 18808 23000 18864
rect 21449 18806 23000 18808
rect 21449 18803 21515 18806
rect 22200 18776 23000 18806
rect 10133 18730 10199 18733
rect 13813 18730 13879 18733
rect 10133 18728 13879 18730
rect 10133 18672 10138 18728
rect 10194 18672 13818 18728
rect 13874 18672 13879 18728
rect 10133 18670 13879 18672
rect 10133 18667 10199 18670
rect 13813 18667 13879 18670
rect 14365 18732 14431 18733
rect 14365 18728 14412 18732
rect 14476 18730 14482 18732
rect 14365 18672 14370 18728
rect 14365 18668 14412 18672
rect 14476 18670 14522 18730
rect 14476 18668 14482 18670
rect 14365 18667 14431 18668
rect 11053 18596 11119 18597
rect 11053 18594 11100 18596
rect 5644 18592 5772 18594
rect 5441 18536 5446 18592
rect 5502 18536 5580 18592
rect 5686 18536 5772 18592
rect 5441 18534 5580 18536
rect 5441 18531 5507 18534
rect 5574 18532 5580 18534
rect 5644 18534 5772 18536
rect 6729 18592 10058 18594
rect 6729 18536 6734 18592
rect 6790 18536 10058 18592
rect 6729 18534 10058 18536
rect 11008 18592 11100 18594
rect 11008 18536 11058 18592
rect 11008 18534 11100 18536
rect 5644 18532 5691 18534
rect 5625 18531 5691 18532
rect 6729 18531 6795 18534
rect 11053 18532 11100 18534
rect 11164 18532 11170 18596
rect 12014 18532 12020 18596
rect 12084 18594 12090 18596
rect 12341 18594 12407 18597
rect 12084 18592 12407 18594
rect 12084 18536 12346 18592
rect 12402 18536 12407 18592
rect 12084 18534 12407 18536
rect 12084 18532 12090 18534
rect 11053 18531 11119 18532
rect 12341 18531 12407 18534
rect 12566 18532 12572 18596
rect 12636 18594 12642 18596
rect 12709 18594 12775 18597
rect 12636 18592 12775 18594
rect 12636 18536 12714 18592
rect 12770 18536 12775 18592
rect 12636 18534 12775 18536
rect 12636 18532 12642 18534
rect 12709 18531 12775 18534
rect 13670 18532 13676 18596
rect 13740 18594 13746 18596
rect 15285 18594 15351 18597
rect 13740 18592 15351 18594
rect 13740 18536 15290 18592
rect 15346 18536 15351 18592
rect 13740 18534 15351 18536
rect 13740 18532 13746 18534
rect 15285 18531 15351 18534
rect 17401 18594 17467 18597
rect 17534 18594 17540 18596
rect 17401 18592 17540 18594
rect 17401 18536 17406 18592
rect 17462 18536 17540 18592
rect 17401 18534 17540 18536
rect 17401 18531 17467 18534
rect 17534 18532 17540 18534
rect 17604 18532 17610 18596
rect 6142 18528 6462 18529
rect 0 18458 800 18488
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 18463 16858 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 2129 18458 2195 18461
rect 5625 18458 5691 18461
rect 2129 18456 5691 18458
rect 2129 18400 2134 18456
rect 2190 18400 5630 18456
rect 5686 18400 5691 18456
rect 2129 18398 5691 18400
rect 2129 18395 2195 18398
rect 5625 18395 5691 18398
rect 6729 18458 6795 18461
rect 6862 18458 6868 18460
rect 6729 18456 6868 18458
rect 6729 18400 6734 18456
rect 6790 18400 6868 18456
rect 6729 18398 6868 18400
rect 6729 18395 6795 18398
rect 6862 18396 6868 18398
rect 6932 18396 6938 18460
rect 7005 18458 7071 18461
rect 7465 18458 7531 18461
rect 7005 18456 7531 18458
rect 7005 18400 7010 18456
rect 7066 18400 7470 18456
rect 7526 18400 7531 18456
rect 7005 18398 7531 18400
rect 7005 18395 7071 18398
rect 7465 18395 7531 18398
rect 7966 18396 7972 18460
rect 8036 18458 8042 18460
rect 8109 18458 8175 18461
rect 8036 18456 8175 18458
rect 8036 18400 8114 18456
rect 8170 18400 8175 18456
rect 8036 18398 8175 18400
rect 8036 18396 8042 18398
rect 8109 18395 8175 18398
rect 8477 18458 8543 18461
rect 9213 18458 9279 18461
rect 11145 18458 11211 18461
rect 8477 18456 9138 18458
rect 8477 18400 8482 18456
rect 8538 18400 9138 18456
rect 8477 18398 9138 18400
rect 8477 18395 8543 18398
rect 4705 18322 4771 18325
rect 5022 18322 5028 18324
rect 4705 18320 5028 18322
rect 4705 18264 4710 18320
rect 4766 18264 5028 18320
rect 4705 18262 5028 18264
rect 4705 18259 4771 18262
rect 5022 18260 5028 18262
rect 5092 18260 5098 18324
rect 5165 18322 5231 18325
rect 8753 18322 8819 18325
rect 5165 18320 8819 18322
rect 5165 18264 5170 18320
rect 5226 18264 8758 18320
rect 8814 18264 8819 18320
rect 5165 18262 8819 18264
rect 9078 18322 9138 18398
rect 9213 18456 11211 18458
rect 9213 18400 9218 18456
rect 9274 18400 11150 18456
rect 11206 18400 11211 18456
rect 9213 18398 11211 18400
rect 9213 18395 9279 18398
rect 11145 18395 11211 18398
rect 11973 18458 12039 18461
rect 18505 18460 18571 18461
rect 11973 18456 12772 18458
rect 11973 18400 11978 18456
rect 12034 18400 12772 18456
rect 11973 18398 12772 18400
rect 11973 18395 12039 18398
rect 9213 18322 9279 18325
rect 12525 18322 12591 18325
rect 9078 18320 12591 18322
rect 9078 18264 9218 18320
rect 9274 18264 12530 18320
rect 12586 18264 12591 18320
rect 9078 18262 12591 18264
rect 12712 18322 12772 18398
rect 18454 18396 18460 18460
rect 18524 18458 18571 18460
rect 21541 18458 21607 18461
rect 22200 18458 23000 18488
rect 18524 18456 18616 18458
rect 18566 18400 18616 18456
rect 18524 18398 18616 18400
rect 21541 18456 23000 18458
rect 21541 18400 21546 18456
rect 21602 18400 23000 18456
rect 21541 18398 23000 18400
rect 18524 18396 18571 18398
rect 18505 18395 18571 18396
rect 21541 18395 21607 18398
rect 22200 18368 23000 18398
rect 17309 18322 17375 18325
rect 12712 18320 17375 18322
rect 12712 18264 17314 18320
rect 17370 18264 17375 18320
rect 12712 18262 17375 18264
rect 5165 18259 5231 18262
rect 8753 18259 8819 18262
rect 9213 18259 9279 18262
rect 12525 18259 12591 18262
rect 17309 18259 17375 18262
rect 3325 18186 3391 18189
rect 3325 18184 9184 18186
rect 3325 18128 3330 18184
rect 3386 18128 9184 18184
rect 3325 18126 9184 18128
rect 3325 18123 3391 18126
rect 0 18050 800 18080
rect 1853 18050 1919 18053
rect 2129 18052 2195 18053
rect 0 18048 1919 18050
rect 0 17992 1858 18048
rect 1914 17992 1919 18048
rect 0 17990 1919 17992
rect 0 17960 800 17990
rect 1853 17987 1919 17990
rect 2078 17988 2084 18052
rect 2148 18050 2195 18052
rect 4613 18050 4679 18053
rect 5257 18050 5323 18053
rect 2148 18048 2240 18050
rect 2190 17992 2240 18048
rect 2148 17990 2240 17992
rect 4613 18048 5323 18050
rect 4613 17992 4618 18048
rect 4674 17992 5262 18048
rect 5318 17992 5323 18048
rect 4613 17990 5323 17992
rect 2148 17988 2195 17990
rect 2129 17987 2195 17988
rect 4613 17987 4679 17990
rect 5257 17987 5323 17990
rect 5625 18050 5691 18053
rect 6729 18050 6795 18053
rect 5625 18048 6795 18050
rect 5625 17992 5630 18048
rect 5686 17992 6734 18048
rect 6790 17992 6795 18048
rect 5625 17990 6795 17992
rect 9124 18050 9184 18126
rect 9254 18124 9260 18188
rect 9324 18186 9330 18188
rect 9397 18186 9463 18189
rect 9324 18184 9463 18186
rect 9324 18128 9402 18184
rect 9458 18128 9463 18184
rect 9324 18126 9463 18128
rect 9324 18124 9330 18126
rect 9397 18123 9463 18126
rect 9581 18188 9647 18189
rect 9581 18184 9628 18188
rect 9692 18186 9698 18188
rect 9581 18128 9586 18184
rect 9581 18124 9628 18128
rect 9692 18126 9738 18186
rect 9692 18124 9698 18126
rect 9806 18124 9812 18188
rect 9876 18186 9882 18188
rect 15745 18186 15811 18189
rect 9876 18184 15811 18186
rect 9876 18128 15750 18184
rect 15806 18128 15811 18184
rect 9876 18126 15811 18128
rect 9876 18124 9882 18126
rect 9581 18123 9647 18124
rect 15745 18123 15811 18126
rect 18505 18186 18571 18189
rect 18965 18186 19031 18189
rect 18505 18184 19031 18186
rect 18505 18128 18510 18184
rect 18566 18128 18970 18184
rect 19026 18128 19031 18184
rect 18505 18126 19031 18128
rect 18505 18123 18571 18126
rect 18965 18123 19031 18126
rect 10409 18050 10475 18053
rect 9124 18048 10475 18050
rect 9124 17992 10414 18048
rect 10470 17992 10475 18048
rect 9124 17990 10475 17992
rect 5625 17987 5691 17990
rect 6729 17987 6795 17990
rect 10409 17987 10475 17990
rect 10685 18050 10751 18053
rect 10910 18050 10916 18052
rect 10685 18048 10916 18050
rect 10685 17992 10690 18048
rect 10746 17992 10916 18048
rect 10685 17990 10916 17992
rect 10685 17987 10751 17990
rect 10910 17988 10916 17990
rect 10980 18050 10986 18052
rect 11421 18050 11487 18053
rect 10980 18048 11487 18050
rect 10980 17992 11426 18048
rect 11482 17992 11487 18048
rect 10980 17990 11487 17992
rect 10980 17988 10986 17990
rect 11421 17987 11487 17990
rect 11789 18050 11855 18053
rect 13721 18050 13787 18053
rect 11789 18048 13787 18050
rect 11789 17992 11794 18048
rect 11850 17992 13726 18048
rect 13782 17992 13787 18048
rect 11789 17990 13787 17992
rect 11789 17987 11855 17990
rect 13721 17987 13787 17990
rect 21449 18050 21515 18053
rect 22200 18050 23000 18080
rect 21449 18048 23000 18050
rect 21449 17992 21454 18048
rect 21510 17992 23000 18048
rect 21449 17990 23000 17992
rect 21449 17987 21515 17990
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 22200 17960 23000 17990
rect 19137 17919 19457 17920
rect 4153 17914 4219 17917
rect 7281 17914 7347 17917
rect 4153 17912 7347 17914
rect 4153 17856 4158 17912
rect 4214 17856 7286 17912
rect 7342 17856 7347 17912
rect 4153 17854 7347 17856
rect 4153 17851 4219 17854
rect 7281 17851 7347 17854
rect 9121 17914 9187 17917
rect 12433 17914 12499 17917
rect 9121 17912 12499 17914
rect 9121 17856 9126 17912
rect 9182 17856 12438 17912
rect 12494 17856 12499 17912
rect 9121 17854 12499 17856
rect 9121 17851 9187 17854
rect 12433 17851 12499 17854
rect 13077 17914 13143 17917
rect 13302 17914 13308 17916
rect 13077 17912 13308 17914
rect 13077 17856 13082 17912
rect 13138 17856 13308 17912
rect 13077 17854 13308 17856
rect 13077 17851 13143 17854
rect 13302 17852 13308 17854
rect 13372 17852 13378 17916
rect 16849 17914 16915 17917
rect 17953 17916 18019 17917
rect 16982 17914 16988 17916
rect 16849 17912 16988 17914
rect 16849 17856 16854 17912
rect 16910 17856 16988 17912
rect 16849 17854 16988 17856
rect 16849 17851 16915 17854
rect 16982 17852 16988 17854
rect 17052 17852 17058 17916
rect 17902 17914 17908 17916
rect 17862 17854 17908 17914
rect 17972 17912 18019 17916
rect 18014 17856 18019 17912
rect 17902 17852 17908 17854
rect 17972 17852 18019 17856
rect 17953 17851 18019 17852
rect 1945 17778 2011 17781
rect 5073 17778 5139 17781
rect 7741 17778 7807 17781
rect 1945 17776 7807 17778
rect 1945 17720 1950 17776
rect 2006 17720 5078 17776
rect 5134 17720 7746 17776
rect 7802 17720 7807 17776
rect 1945 17718 7807 17720
rect 1945 17715 2011 17718
rect 5073 17715 5139 17718
rect 7741 17715 7807 17718
rect 8109 17778 8175 17781
rect 10501 17778 10567 17781
rect 8109 17776 10567 17778
rect 8109 17720 8114 17776
rect 8170 17720 10506 17776
rect 10562 17720 10567 17776
rect 8109 17718 10567 17720
rect 8109 17715 8175 17718
rect 10501 17715 10567 17718
rect 10869 17778 10935 17781
rect 12249 17778 12315 17781
rect 13629 17778 13695 17781
rect 10869 17776 12315 17778
rect 10869 17720 10874 17776
rect 10930 17720 12254 17776
rect 12310 17720 12315 17776
rect 10869 17718 12315 17720
rect 10869 17715 10935 17718
rect 12249 17715 12315 17718
rect 12390 17776 13695 17778
rect 12390 17720 13634 17776
rect 13690 17720 13695 17776
rect 12390 17718 13695 17720
rect 0 17642 800 17672
rect 1485 17642 1551 17645
rect 0 17640 1551 17642
rect 0 17584 1490 17640
rect 1546 17584 1551 17640
rect 0 17582 1551 17584
rect 0 17552 800 17582
rect 1485 17579 1551 17582
rect 3182 17580 3188 17644
rect 3252 17642 3258 17644
rect 4153 17642 4219 17645
rect 5717 17644 5783 17645
rect 5717 17642 5764 17644
rect 3252 17640 4219 17642
rect 3252 17584 4158 17640
rect 4214 17584 4219 17640
rect 3252 17582 4219 17584
rect 5672 17640 5764 17642
rect 5672 17584 5722 17640
rect 5672 17582 5764 17584
rect 3252 17580 3258 17582
rect 4153 17579 4219 17582
rect 5717 17580 5764 17582
rect 5828 17580 5834 17644
rect 9765 17642 9831 17645
rect 10685 17642 10751 17645
rect 12390 17642 12450 17718
rect 13629 17715 13695 17718
rect 13813 17778 13879 17781
rect 14406 17778 14412 17780
rect 13813 17776 14412 17778
rect 13813 17720 13818 17776
rect 13874 17720 14412 17776
rect 13813 17718 14412 17720
rect 13813 17715 13879 17718
rect 14406 17716 14412 17718
rect 14476 17716 14482 17780
rect 16573 17778 16639 17781
rect 19006 17778 19012 17780
rect 16573 17776 19012 17778
rect 16573 17720 16578 17776
rect 16634 17720 19012 17776
rect 16573 17718 19012 17720
rect 16573 17715 16639 17718
rect 19006 17716 19012 17718
rect 19076 17716 19082 17780
rect 19926 17716 19932 17780
rect 19996 17778 20002 17780
rect 20069 17778 20135 17781
rect 19996 17776 20135 17778
rect 19996 17720 20074 17776
rect 20130 17720 20135 17776
rect 19996 17718 20135 17720
rect 19996 17716 20002 17718
rect 20069 17715 20135 17718
rect 5950 17640 10751 17642
rect 5950 17584 9770 17640
rect 9826 17584 10690 17640
rect 10746 17584 10751 17640
rect 5950 17582 10751 17584
rect 5717 17579 5783 17580
rect 3233 17506 3299 17509
rect 5717 17506 5783 17509
rect 3233 17504 5783 17506
rect 3233 17448 3238 17504
rect 3294 17448 5722 17504
rect 5778 17448 5783 17504
rect 3233 17446 5783 17448
rect 3233 17443 3299 17446
rect 5717 17443 5783 17446
rect 2221 17370 2287 17373
rect 5950 17370 6010 17582
rect 9765 17579 9831 17582
rect 10685 17579 10751 17582
rect 10918 17582 12450 17642
rect 21449 17642 21515 17645
rect 22200 17642 23000 17672
rect 21449 17640 23000 17642
rect 21449 17584 21454 17640
rect 21510 17584 23000 17640
rect 21449 17582 23000 17584
rect 6545 17506 6611 17509
rect 10918 17506 10978 17582
rect 21449 17579 21515 17582
rect 22200 17552 23000 17582
rect 6545 17504 10978 17506
rect 6545 17448 6550 17504
rect 6606 17448 10978 17504
rect 6545 17446 10978 17448
rect 11789 17506 11855 17509
rect 14273 17506 14339 17509
rect 11789 17504 14339 17506
rect 11789 17448 11794 17504
rect 11850 17448 14278 17504
rect 14334 17448 14339 17504
rect 11789 17446 14339 17448
rect 6545 17443 6611 17446
rect 11789 17443 11855 17446
rect 14273 17443 14339 17446
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 17375 16858 17376
rect 2221 17368 6010 17370
rect 2221 17312 2226 17368
rect 2282 17312 6010 17368
rect 2221 17310 6010 17312
rect 7465 17370 7531 17373
rect 10685 17370 10751 17373
rect 7465 17368 10751 17370
rect 7465 17312 7470 17368
rect 7526 17312 10690 17368
rect 10746 17312 10751 17368
rect 7465 17310 10751 17312
rect 2221 17307 2287 17310
rect 7465 17307 7531 17310
rect 10685 17307 10751 17310
rect 0 17234 800 17264
rect 1485 17234 1551 17237
rect 0 17232 1551 17234
rect 0 17176 1490 17232
rect 1546 17176 1551 17232
rect 0 17174 1551 17176
rect 0 17144 800 17174
rect 1485 17171 1551 17174
rect 2405 17234 2471 17237
rect 7966 17234 7972 17236
rect 2405 17232 7972 17234
rect 2405 17176 2410 17232
rect 2466 17176 7972 17232
rect 2405 17174 7972 17176
rect 2405 17171 2471 17174
rect 7966 17172 7972 17174
rect 8036 17234 8042 17236
rect 9213 17234 9279 17237
rect 19558 17234 19564 17236
rect 8036 17174 9138 17234
rect 8036 17172 8042 17174
rect 3918 17036 3924 17100
rect 3988 17098 3994 17100
rect 4613 17098 4679 17101
rect 3988 17096 4679 17098
rect 3988 17040 4618 17096
rect 4674 17040 4679 17096
rect 3988 17038 4679 17040
rect 3988 17036 3994 17038
rect 4613 17035 4679 17038
rect 6177 17098 6243 17101
rect 8845 17098 8911 17101
rect 6177 17096 8911 17098
rect 6177 17040 6182 17096
rect 6238 17040 8850 17096
rect 8906 17040 8911 17096
rect 6177 17038 8911 17040
rect 9078 17098 9138 17174
rect 9213 17232 19564 17234
rect 9213 17176 9218 17232
rect 9274 17176 19564 17232
rect 9213 17174 19564 17176
rect 9213 17171 9279 17174
rect 19558 17172 19564 17174
rect 19628 17172 19634 17236
rect 20529 17234 20595 17237
rect 22200 17234 23000 17264
rect 20529 17232 23000 17234
rect 20529 17176 20534 17232
rect 20590 17176 23000 17232
rect 20529 17174 23000 17176
rect 20529 17171 20595 17174
rect 22200 17144 23000 17174
rect 10501 17098 10567 17101
rect 9078 17096 10567 17098
rect 9078 17040 10506 17096
rect 10562 17040 10567 17096
rect 9078 17038 10567 17040
rect 6177 17035 6243 17038
rect 8845 17035 8911 17038
rect 10501 17035 10567 17038
rect 13486 17036 13492 17100
rect 13556 17098 13562 17100
rect 17769 17098 17835 17101
rect 13556 17096 17835 17098
rect 13556 17040 17774 17096
rect 17830 17040 17835 17096
rect 13556 17038 17835 17040
rect 13556 17036 13562 17038
rect 17769 17035 17835 17038
rect 4521 16962 4587 16965
rect 5625 16962 5691 16965
rect 8293 16962 8359 16965
rect 4521 16960 5691 16962
rect 4521 16904 4526 16960
rect 4582 16904 5630 16960
rect 5686 16904 5691 16960
rect 4521 16902 5691 16904
rect 4521 16899 4587 16902
rect 5625 16899 5691 16902
rect 5812 16960 8359 16962
rect 5812 16904 8298 16960
rect 8354 16904 8359 16960
rect 5812 16902 8359 16904
rect 3543 16896 3863 16897
rect 0 16826 800 16856
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 1485 16826 1551 16829
rect 0 16824 1551 16826
rect 0 16768 1490 16824
rect 1546 16768 1551 16824
rect 0 16766 1551 16768
rect 0 16736 800 16766
rect 1485 16763 1551 16766
rect 3969 16826 4035 16829
rect 5812 16826 5872 16902
rect 8293 16899 8359 16902
rect 9673 16962 9739 16965
rect 11237 16962 11303 16965
rect 13537 16962 13603 16965
rect 9673 16960 11303 16962
rect 9673 16904 9678 16960
rect 9734 16904 11242 16960
rect 11298 16904 11303 16960
rect 9673 16902 11303 16904
rect 9673 16899 9739 16902
rect 11237 16899 11303 16902
rect 12390 16960 13603 16962
rect 12390 16904 13542 16960
rect 13598 16904 13603 16960
rect 12390 16902 13603 16904
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 3969 16824 5872 16826
rect 3969 16768 3974 16824
rect 4030 16768 5872 16824
rect 3969 16766 5872 16768
rect 3969 16763 4035 16766
rect 5942 16764 5948 16828
rect 6012 16826 6018 16828
rect 6269 16826 6335 16829
rect 7189 16826 7255 16829
rect 6012 16824 7255 16826
rect 6012 16768 6274 16824
rect 6330 16768 7194 16824
rect 7250 16768 7255 16824
rect 6012 16766 7255 16768
rect 6012 16764 6018 16766
rect 6269 16763 6335 16766
rect 7189 16763 7255 16766
rect 11094 16764 11100 16828
rect 11164 16826 11170 16828
rect 11513 16826 11579 16829
rect 11830 16826 11836 16828
rect 11164 16824 11836 16826
rect 11164 16768 11518 16824
rect 11574 16768 11836 16824
rect 11164 16766 11836 16768
rect 11164 16764 11170 16766
rect 11513 16763 11579 16766
rect 11830 16764 11836 16766
rect 11900 16764 11906 16828
rect 1894 16628 1900 16692
rect 1964 16690 1970 16692
rect 12390 16690 12450 16902
rect 13537 16899 13603 16902
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 21449 16826 21515 16829
rect 22200 16826 23000 16856
rect 21449 16824 23000 16826
rect 21449 16768 21454 16824
rect 21510 16768 23000 16824
rect 21449 16766 23000 16768
rect 21449 16763 21515 16766
rect 22200 16736 23000 16766
rect 1964 16630 12450 16690
rect 1964 16628 1970 16630
rect 12566 16628 12572 16692
rect 12636 16690 12642 16692
rect 17861 16690 17927 16693
rect 12636 16688 17927 16690
rect 12636 16632 17866 16688
rect 17922 16632 17927 16688
rect 12636 16630 17927 16632
rect 12636 16628 12642 16630
rect 17861 16627 17927 16630
rect 19885 16690 19951 16693
rect 20805 16690 20871 16693
rect 19885 16688 20871 16690
rect 19885 16632 19890 16688
rect 19946 16632 20810 16688
rect 20866 16632 20871 16688
rect 19885 16630 20871 16632
rect 19885 16627 19951 16630
rect 20805 16627 20871 16630
rect 2129 16554 2195 16557
rect 4245 16554 4311 16557
rect 2129 16552 4311 16554
rect 2129 16496 2134 16552
rect 2190 16496 4250 16552
rect 4306 16496 4311 16552
rect 2129 16494 4311 16496
rect 2129 16491 2195 16494
rect 4245 16491 4311 16494
rect 5533 16554 5599 16557
rect 10777 16554 10843 16557
rect 18873 16554 18939 16557
rect 5533 16552 10843 16554
rect 5533 16496 5538 16552
rect 5594 16496 10782 16552
rect 10838 16496 10843 16552
rect 5533 16494 10843 16496
rect 5533 16491 5599 16494
rect 10777 16491 10843 16494
rect 10918 16552 18939 16554
rect 10918 16496 18878 16552
rect 18934 16496 18939 16552
rect 10918 16494 18939 16496
rect 2681 16418 2747 16421
rect 7189 16418 7255 16421
rect 10918 16418 10978 16494
rect 18873 16491 18939 16494
rect 19149 16554 19215 16557
rect 22277 16554 22343 16557
rect 19149 16552 22343 16554
rect 19149 16496 19154 16552
rect 19210 16496 22282 16552
rect 22338 16496 22343 16552
rect 19149 16494 22343 16496
rect 19149 16491 19215 16494
rect 22277 16491 22343 16494
rect 2681 16416 5826 16418
rect 2681 16360 2686 16416
rect 2742 16360 5826 16416
rect 2681 16358 5826 16360
rect 2681 16355 2747 16358
rect 0 16282 800 16312
rect 1485 16282 1551 16285
rect 0 16280 1551 16282
rect 0 16224 1490 16280
rect 1546 16224 1551 16280
rect 0 16222 1551 16224
rect 0 16192 800 16222
rect 1485 16219 1551 16222
rect 2497 16282 2563 16285
rect 4153 16282 4219 16285
rect 2497 16280 4219 16282
rect 2497 16224 2502 16280
rect 2558 16224 4158 16280
rect 4214 16224 4219 16280
rect 2497 16222 4219 16224
rect 5766 16282 5826 16358
rect 7189 16416 10978 16418
rect 7189 16360 7194 16416
rect 7250 16360 10978 16416
rect 7189 16358 10978 16360
rect 7189 16355 7255 16358
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 8017 16282 8083 16285
rect 5766 16222 6010 16282
rect 2497 16219 2563 16222
rect 4153 16219 4219 16222
rect 5950 16146 6010 16222
rect 6870 16280 8083 16282
rect 6870 16224 8022 16280
rect 8078 16224 8083 16280
rect 6870 16222 8083 16224
rect 6870 16146 6930 16222
rect 8017 16219 8083 16222
rect 8334 16220 8340 16284
rect 8404 16282 8410 16284
rect 8477 16282 8543 16285
rect 8404 16280 8543 16282
rect 8404 16224 8482 16280
rect 8538 16224 8543 16280
rect 8404 16222 8543 16224
rect 8404 16220 8410 16222
rect 8477 16219 8543 16222
rect 12157 16282 12223 16285
rect 12934 16282 12940 16284
rect 12157 16280 12940 16282
rect 12157 16224 12162 16280
rect 12218 16224 12940 16280
rect 12157 16222 12940 16224
rect 12157 16219 12223 16222
rect 12934 16220 12940 16222
rect 13004 16282 13010 16284
rect 15653 16282 15719 16285
rect 13004 16280 15719 16282
rect 13004 16224 15658 16280
rect 15714 16224 15719 16280
rect 13004 16222 15719 16224
rect 13004 16220 13010 16222
rect 15653 16219 15719 16222
rect 20161 16282 20227 16285
rect 21081 16282 21147 16285
rect 20161 16280 21147 16282
rect 20161 16224 20166 16280
rect 20222 16224 21086 16280
rect 21142 16224 21147 16280
rect 20161 16222 21147 16224
rect 20161 16219 20227 16222
rect 21081 16219 21147 16222
rect 21449 16282 21515 16285
rect 22200 16282 23000 16312
rect 21449 16280 23000 16282
rect 21449 16224 21454 16280
rect 21510 16224 23000 16280
rect 21449 16222 23000 16224
rect 21449 16219 21515 16222
rect 22200 16192 23000 16222
rect 18321 16146 18387 16149
rect 5950 16086 6930 16146
rect 7238 16144 18387 16146
rect 7238 16088 18326 16144
rect 18382 16088 18387 16144
rect 7238 16086 18387 16088
rect 3141 16010 3207 16013
rect 7238 16010 7298 16086
rect 18321 16083 18387 16086
rect 19517 16146 19583 16149
rect 19517 16144 20546 16146
rect 19517 16088 19522 16144
rect 19578 16088 20546 16144
rect 19517 16086 20546 16088
rect 19517 16083 19583 16086
rect 12198 16010 12204 16012
rect 3141 16008 7298 16010
rect 3141 15952 3146 16008
rect 3202 15952 7298 16008
rect 3141 15950 7298 15952
rect 8572 15950 12204 16010
rect 3141 15947 3207 15950
rect 0 15874 800 15904
rect 8572 15877 8632 15950
rect 12198 15948 12204 15950
rect 12268 16010 12274 16012
rect 17125 16010 17191 16013
rect 12268 16008 17191 16010
rect 12268 15952 17130 16008
rect 17186 15952 17191 16008
rect 12268 15950 17191 15952
rect 12268 15948 12274 15950
rect 17125 15947 17191 15950
rect 17902 15948 17908 16012
rect 17972 16010 17978 16012
rect 19057 16010 19123 16013
rect 17972 16008 19123 16010
rect 17972 15952 19062 16008
rect 19118 15952 19123 16008
rect 17972 15950 19123 15952
rect 17972 15948 17978 15950
rect 19057 15947 19123 15950
rect 19609 16010 19675 16013
rect 20345 16010 20411 16013
rect 19609 16008 20411 16010
rect 19609 15952 19614 16008
rect 19670 15952 20350 16008
rect 20406 15952 20411 16008
rect 19609 15950 20411 15952
rect 19609 15947 19675 15950
rect 20345 15947 20411 15950
rect 20486 15877 20546 16086
rect 1485 15874 1551 15877
rect 0 15872 1551 15874
rect 0 15816 1490 15872
rect 1546 15816 1551 15872
rect 0 15814 1551 15816
rect 0 15784 800 15814
rect 1485 15811 1551 15814
rect 7741 15874 7807 15877
rect 8150 15874 8156 15876
rect 7741 15872 8156 15874
rect 7741 15816 7746 15872
rect 7802 15816 8156 15872
rect 7741 15814 8156 15816
rect 7741 15811 7807 15814
rect 8150 15812 8156 15814
rect 8220 15874 8226 15876
rect 8569 15874 8635 15877
rect 8220 15872 8635 15874
rect 8220 15816 8574 15872
rect 8630 15816 8635 15872
rect 8220 15814 8635 15816
rect 8220 15812 8226 15814
rect 8569 15811 8635 15814
rect 10726 15812 10732 15876
rect 10796 15874 10802 15876
rect 10961 15874 11027 15877
rect 10796 15872 11027 15874
rect 10796 15816 10966 15872
rect 11022 15816 11027 15872
rect 10796 15814 11027 15816
rect 10796 15812 10802 15814
rect 10961 15811 11027 15814
rect 20437 15872 20546 15877
rect 20437 15816 20442 15872
rect 20498 15816 20546 15872
rect 20437 15814 20546 15816
rect 21449 15874 21515 15877
rect 22200 15874 23000 15904
rect 21449 15872 23000 15874
rect 21449 15816 21454 15872
rect 21510 15816 23000 15872
rect 21449 15814 23000 15816
rect 20437 15811 20503 15814
rect 21449 15811 21515 15814
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 22200 15784 23000 15814
rect 19137 15743 19457 15744
rect 5206 15676 5212 15740
rect 5276 15738 5282 15740
rect 7649 15738 7715 15741
rect 5276 15736 7715 15738
rect 5276 15680 7654 15736
rect 7710 15680 7715 15736
rect 5276 15678 7715 15680
rect 5276 15676 5282 15678
rect 7649 15675 7715 15678
rect 9673 15738 9739 15741
rect 13261 15738 13327 15741
rect 9673 15736 13327 15738
rect 9673 15680 9678 15736
rect 9734 15680 13266 15736
rect 13322 15680 13327 15736
rect 9673 15678 13327 15680
rect 9673 15675 9739 15678
rect 13261 15675 13327 15678
rect 4102 15540 4108 15604
rect 4172 15602 4178 15604
rect 11697 15602 11763 15605
rect 4172 15600 11763 15602
rect 4172 15544 11702 15600
rect 11758 15544 11763 15600
rect 4172 15542 11763 15544
rect 4172 15540 4178 15542
rect 11697 15539 11763 15542
rect 0 15466 800 15496
rect 1853 15466 1919 15469
rect 0 15464 1919 15466
rect 0 15408 1858 15464
rect 1914 15408 1919 15464
rect 0 15406 1919 15408
rect 0 15376 800 15406
rect 1853 15403 1919 15406
rect 5625 15466 5691 15469
rect 11881 15466 11947 15469
rect 5625 15464 11947 15466
rect 5625 15408 5630 15464
rect 5686 15408 11886 15464
rect 11942 15408 11947 15464
rect 5625 15406 11947 15408
rect 5625 15403 5691 15406
rect 11881 15403 11947 15406
rect 21081 15466 21147 15469
rect 22200 15466 23000 15496
rect 21081 15464 23000 15466
rect 21081 15408 21086 15464
rect 21142 15408 23000 15464
rect 21081 15406 23000 15408
rect 21081 15403 21147 15406
rect 22200 15376 23000 15406
rect 8477 15330 8543 15333
rect 7606 15328 8543 15330
rect 7606 15272 8482 15328
rect 8538 15272 8543 15328
rect 7606 15270 8543 15272
rect 6142 15264 6462 15265
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 7005 15194 7071 15197
rect 7606 15196 7666 15270
rect 8477 15267 8543 15270
rect 9857 15330 9923 15333
rect 10593 15330 10659 15333
rect 9857 15328 10659 15330
rect 9857 15272 9862 15328
rect 9918 15272 10598 15328
rect 10654 15272 10659 15328
rect 9857 15270 10659 15272
rect 9857 15267 9923 15270
rect 10593 15267 10659 15270
rect 18270 15268 18276 15332
rect 18340 15330 18346 15332
rect 18505 15330 18571 15333
rect 18340 15328 18571 15330
rect 18340 15272 18510 15328
rect 18566 15272 18571 15328
rect 18340 15270 18571 15272
rect 18340 15268 18346 15270
rect 18505 15267 18571 15270
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 15199 16858 15200
rect 7598 15194 7604 15196
rect 7005 15192 7604 15194
rect 7005 15136 7010 15192
rect 7066 15136 7604 15192
rect 7005 15134 7604 15136
rect 7005 15131 7071 15134
rect 7598 15132 7604 15134
rect 7668 15132 7674 15196
rect 8017 15194 8083 15197
rect 11145 15194 11211 15197
rect 8017 15192 11211 15194
rect 8017 15136 8022 15192
rect 8078 15136 11150 15192
rect 11206 15136 11211 15192
rect 8017 15134 11211 15136
rect 8017 15131 8083 15134
rect 11145 15131 11211 15134
rect 13302 15132 13308 15196
rect 13372 15194 13378 15196
rect 13813 15194 13879 15197
rect 13372 15192 13879 15194
rect 13372 15136 13818 15192
rect 13874 15136 13879 15192
rect 13372 15134 13879 15136
rect 13372 15132 13378 15134
rect 13813 15131 13879 15134
rect 15326 15132 15332 15196
rect 15396 15194 15402 15196
rect 15745 15194 15811 15197
rect 15396 15192 15811 15194
rect 15396 15136 15750 15192
rect 15806 15136 15811 15192
rect 15396 15134 15811 15136
rect 15396 15132 15402 15134
rect 15745 15131 15811 15134
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 5717 15058 5783 15061
rect 10041 15058 10107 15061
rect 5717 15056 10107 15058
rect 5717 15000 5722 15056
rect 5778 15000 10046 15056
rect 10102 15000 10107 15056
rect 5717 14998 10107 15000
rect 5717 14995 5783 14998
rect 10041 14995 10107 14998
rect 10409 15058 10475 15061
rect 11421 15058 11487 15061
rect 12014 15058 12020 15060
rect 10409 15056 12020 15058
rect 10409 15000 10414 15056
rect 10470 15000 11426 15056
rect 11482 15000 12020 15056
rect 10409 14998 12020 15000
rect 10409 14995 10475 14998
rect 11421 14995 11487 14998
rect 12014 14996 12020 14998
rect 12084 14996 12090 15060
rect 12985 15058 13051 15061
rect 12390 15056 13051 15058
rect 12390 15000 12990 15056
rect 13046 15000 13051 15056
rect 12390 14998 13051 15000
rect 2998 14860 3004 14924
rect 3068 14922 3074 14924
rect 3233 14922 3299 14925
rect 3068 14920 3299 14922
rect 3068 14864 3238 14920
rect 3294 14864 3299 14920
rect 3068 14862 3299 14864
rect 3068 14860 3074 14862
rect 3233 14859 3299 14862
rect 5073 14922 5139 14925
rect 12390 14922 12450 14998
rect 12985 14995 13051 14998
rect 16389 15058 16455 15061
rect 16982 15058 16988 15060
rect 16389 15056 16988 15058
rect 16389 15000 16394 15056
rect 16450 15000 16988 15056
rect 16389 14998 16988 15000
rect 16389 14995 16455 14998
rect 16982 14996 16988 14998
rect 17052 14996 17058 15060
rect 21449 15058 21515 15061
rect 22200 15058 23000 15088
rect 21449 15056 23000 15058
rect 21449 15000 21454 15056
rect 21510 15000 23000 15056
rect 21449 14998 23000 15000
rect 21449 14995 21515 14998
rect 22200 14968 23000 14998
rect 5073 14920 12450 14922
rect 5073 14864 5078 14920
rect 5134 14864 12450 14920
rect 5073 14862 12450 14864
rect 15469 14922 15535 14925
rect 16062 14922 16068 14924
rect 15469 14920 16068 14922
rect 15469 14864 15474 14920
rect 15530 14864 16068 14920
rect 15469 14862 16068 14864
rect 5073 14859 5139 14862
rect 15469 14859 15535 14862
rect 16062 14860 16068 14862
rect 16132 14922 16138 14924
rect 18689 14922 18755 14925
rect 16132 14920 18755 14922
rect 16132 14864 18694 14920
rect 18750 14864 18755 14920
rect 16132 14862 18755 14864
rect 16132 14860 16138 14862
rect 18689 14859 18755 14862
rect 5533 14786 5599 14789
rect 8569 14786 8635 14789
rect 5533 14784 8635 14786
rect 5533 14728 5538 14784
rect 5594 14728 8574 14784
rect 8630 14728 8635 14784
rect 5533 14726 8635 14728
rect 5533 14723 5599 14726
rect 8569 14723 8635 14726
rect 9213 14786 9279 14789
rect 11973 14786 12039 14789
rect 9213 14784 12039 14786
rect 9213 14728 9218 14784
rect 9274 14728 11978 14784
rect 12034 14728 12039 14784
rect 9213 14726 12039 14728
rect 9213 14723 9279 14726
rect 11973 14723 12039 14726
rect 14457 14786 14523 14789
rect 14590 14786 14596 14788
rect 14457 14784 14596 14786
rect 14457 14728 14462 14784
rect 14518 14728 14596 14784
rect 14457 14726 14596 14728
rect 14457 14723 14523 14726
rect 14590 14724 14596 14726
rect 14660 14724 14666 14788
rect 3543 14720 3863 14721
rect 0 14650 800 14680
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 800 14590
rect 1485 14587 1551 14590
rect 6821 14650 6887 14653
rect 8017 14650 8083 14653
rect 6821 14648 8083 14650
rect 6821 14592 6826 14648
rect 6882 14592 8022 14648
rect 8078 14592 8083 14648
rect 6821 14590 8083 14592
rect 6821 14587 6887 14590
rect 8017 14587 8083 14590
rect 9121 14650 9187 14653
rect 12709 14650 12775 14653
rect 9121 14648 12775 14650
rect 9121 14592 9126 14648
rect 9182 14592 12714 14648
rect 12770 14592 12775 14648
rect 9121 14590 12775 14592
rect 9121 14587 9187 14590
rect 12709 14587 12775 14590
rect 21449 14650 21515 14653
rect 22200 14650 23000 14680
rect 21449 14648 23000 14650
rect 21449 14592 21454 14648
rect 21510 14592 23000 14648
rect 21449 14590 23000 14592
rect 21449 14587 21515 14590
rect 22200 14560 23000 14590
rect 1669 14514 1735 14517
rect 10133 14514 10199 14517
rect 1669 14512 10199 14514
rect 1669 14456 1674 14512
rect 1730 14456 10138 14512
rect 10194 14456 10199 14512
rect 1669 14454 10199 14456
rect 1669 14451 1735 14454
rect 10133 14451 10199 14454
rect 11145 14514 11211 14517
rect 17217 14514 17283 14517
rect 11145 14512 17283 14514
rect 11145 14456 11150 14512
rect 11206 14456 17222 14512
rect 17278 14456 17283 14512
rect 11145 14454 17283 14456
rect 11145 14451 11211 14454
rect 17217 14451 17283 14454
rect 6729 14378 6795 14381
rect 15009 14378 15075 14381
rect 6729 14376 15075 14378
rect 6729 14320 6734 14376
rect 6790 14320 15014 14376
rect 15070 14320 15075 14376
rect 6729 14318 15075 14320
rect 6729 14315 6795 14318
rect 15009 14315 15075 14318
rect 19517 14378 19583 14381
rect 21817 14378 21883 14381
rect 19517 14376 21883 14378
rect 19517 14320 19522 14376
rect 19578 14320 21822 14376
rect 21878 14320 21883 14376
rect 19517 14318 21883 14320
rect 19517 14315 19583 14318
rect 21817 14315 21883 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 2681 14242 2747 14245
rect 4061 14242 4127 14245
rect 2681 14240 4127 14242
rect 2681 14184 2686 14240
rect 2742 14184 4066 14240
rect 4122 14184 4127 14240
rect 2681 14182 4127 14184
rect 2681 14179 2747 14182
rect 4061 14179 4127 14182
rect 6545 14242 6611 14245
rect 7281 14242 7347 14245
rect 7414 14242 7420 14244
rect 6545 14240 7420 14242
rect 6545 14184 6550 14240
rect 6606 14184 7286 14240
rect 7342 14184 7420 14240
rect 6545 14182 7420 14184
rect 6545 14179 6611 14182
rect 7281 14179 7347 14182
rect 7414 14180 7420 14182
rect 7484 14180 7490 14244
rect 12065 14242 12131 14245
rect 12566 14242 12572 14244
rect 12065 14240 12572 14242
rect 12065 14184 12070 14240
rect 12126 14184 12572 14240
rect 12065 14182 12572 14184
rect 12065 14179 12131 14182
rect 12566 14180 12572 14182
rect 12636 14180 12642 14244
rect 12709 14242 12775 14245
rect 16246 14242 16252 14244
rect 12709 14240 16252 14242
rect 12709 14184 12714 14240
rect 12770 14184 16252 14240
rect 12709 14182 16252 14184
rect 12709 14179 12775 14182
rect 16246 14180 16252 14182
rect 16316 14180 16322 14244
rect 17217 14242 17283 14245
rect 18454 14242 18460 14244
rect 17217 14240 18460 14242
rect 17217 14184 17222 14240
rect 17278 14184 18460 14240
rect 17217 14182 18460 14184
rect 17217 14179 17283 14182
rect 18454 14180 18460 14182
rect 18524 14180 18530 14244
rect 21449 14242 21515 14245
rect 22200 14242 23000 14272
rect 21449 14240 23000 14242
rect 21449 14184 21454 14240
rect 21510 14184 23000 14240
rect 21449 14182 23000 14184
rect 21449 14179 21515 14182
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 22200 14152 23000 14182
rect 16538 14111 16858 14112
rect 5073 14106 5139 14109
rect 982 14104 5139 14106
rect 841 14072 907 14075
rect 982 14072 5078 14104
rect 841 14070 5078 14072
rect 841 14014 846 14070
rect 902 14048 5078 14070
rect 5134 14048 5139 14104
rect 902 14046 5139 14048
rect 902 14014 1042 14046
rect 5073 14043 5139 14046
rect 6678 14044 6684 14108
rect 6748 14106 6754 14108
rect 6821 14106 6887 14109
rect 6748 14104 6887 14106
rect 6748 14048 6826 14104
rect 6882 14048 6887 14104
rect 6748 14046 6887 14048
rect 6748 14044 6754 14046
rect 6821 14043 6887 14046
rect 7230 14044 7236 14108
rect 7300 14106 7306 14108
rect 8477 14106 8543 14109
rect 7300 14104 8543 14106
rect 7300 14048 8482 14104
rect 8538 14048 8543 14104
rect 7300 14046 8543 14048
rect 7300 14044 7306 14046
rect 8477 14043 8543 14046
rect 12341 14106 12407 14109
rect 15653 14106 15719 14109
rect 17217 14108 17283 14109
rect 17166 14106 17172 14108
rect 12341 14104 15719 14106
rect 12341 14048 12346 14104
rect 12402 14048 15658 14104
rect 15714 14048 15719 14104
rect 12341 14046 15719 14048
rect 17126 14046 17172 14106
rect 17236 14104 17283 14108
rect 17278 14048 17283 14104
rect 12341 14043 12407 14046
rect 15653 14043 15719 14046
rect 17166 14044 17172 14046
rect 17236 14044 17283 14048
rect 17217 14043 17283 14044
rect 841 14012 1042 14014
rect 841 14009 907 14012
rect 3509 13970 3575 13973
rect 7046 13970 7052 13972
rect 2730 13968 7052 13970
rect 2730 13912 3514 13968
rect 3570 13912 7052 13968
rect 2730 13910 7052 13912
rect 0 13834 800 13864
rect 1853 13834 1919 13837
rect 0 13832 1919 13834
rect 0 13776 1858 13832
rect 1914 13776 1919 13832
rect 0 13774 1919 13776
rect 0 13744 800 13774
rect 1853 13771 1919 13774
rect 2037 13834 2103 13837
rect 2730 13834 2790 13910
rect 3509 13907 3575 13910
rect 7046 13908 7052 13910
rect 7116 13970 7122 13972
rect 9121 13970 9187 13973
rect 7116 13968 9187 13970
rect 7116 13912 9126 13968
rect 9182 13912 9187 13968
rect 7116 13910 9187 13912
rect 7116 13908 7122 13910
rect 9121 13907 9187 13910
rect 11605 13970 11671 13973
rect 18689 13970 18755 13973
rect 20437 13970 20503 13973
rect 11605 13968 15946 13970
rect 11605 13912 11610 13968
rect 11666 13912 15946 13968
rect 11605 13910 15946 13912
rect 11605 13907 11671 13910
rect 2037 13832 2790 13834
rect 2037 13776 2042 13832
rect 2098 13776 2790 13832
rect 2037 13774 2790 13776
rect 5533 13834 5599 13837
rect 7414 13834 7420 13836
rect 5533 13832 7420 13834
rect 5533 13776 5538 13832
rect 5594 13776 7420 13832
rect 5533 13774 7420 13776
rect 2037 13771 2103 13774
rect 5533 13771 5599 13774
rect 7414 13772 7420 13774
rect 7484 13772 7490 13836
rect 9806 13834 9812 13836
rect 7606 13774 9812 13834
rect 4838 13636 4844 13700
rect 4908 13698 4914 13700
rect 5942 13698 5948 13700
rect 4908 13638 5948 13698
rect 4908 13636 4914 13638
rect 5942 13636 5948 13638
rect 6012 13636 6018 13700
rect 7606 13698 7666 13774
rect 9806 13772 9812 13774
rect 9876 13834 9882 13836
rect 12341 13834 12407 13837
rect 9876 13832 12407 13834
rect 9876 13776 12346 13832
rect 12402 13776 12407 13832
rect 9876 13774 12407 13776
rect 9876 13772 9882 13774
rect 12341 13771 12407 13774
rect 12750 13772 12756 13836
rect 12820 13834 12826 13836
rect 12985 13834 13051 13837
rect 12820 13832 13051 13834
rect 12820 13776 12990 13832
rect 13046 13776 13051 13832
rect 12820 13774 13051 13776
rect 15886 13834 15946 13910
rect 18689 13968 20503 13970
rect 18689 13912 18694 13968
rect 18750 13912 20442 13968
rect 20498 13912 20503 13968
rect 18689 13910 20503 13912
rect 18689 13907 18755 13910
rect 20437 13907 20503 13910
rect 17125 13836 17191 13837
rect 15886 13774 17050 13834
rect 12820 13772 12826 13774
rect 12985 13771 13051 13774
rect 7238 13638 7666 13698
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 2957 13562 3023 13565
rect 2730 13560 3023 13562
rect 2730 13504 2962 13560
rect 3018 13504 3023 13560
rect 2730 13502 3023 13504
rect 0 13426 800 13456
rect 1485 13426 1551 13429
rect 0 13424 1551 13426
rect 0 13368 1490 13424
rect 1546 13368 1551 13424
rect 0 13366 1551 13368
rect 0 13336 800 13366
rect 1485 13363 1551 13366
rect 1945 13426 2011 13429
rect 2730 13426 2790 13502
rect 2957 13499 3023 13502
rect 5441 13562 5507 13565
rect 7238 13562 7298 13638
rect 9438 13636 9444 13700
rect 9508 13698 9514 13700
rect 9673 13698 9739 13701
rect 9508 13696 9739 13698
rect 9508 13640 9678 13696
rect 9734 13640 9739 13696
rect 9508 13638 9739 13640
rect 9508 13636 9514 13638
rect 9673 13635 9739 13638
rect 10910 13636 10916 13700
rect 10980 13698 10986 13700
rect 12157 13698 12223 13701
rect 10980 13696 12223 13698
rect 10980 13640 12162 13696
rect 12218 13640 12223 13696
rect 10980 13638 12223 13640
rect 10980 13636 10986 13638
rect 12157 13635 12223 13638
rect 15326 13636 15332 13700
rect 15396 13698 15402 13700
rect 16573 13698 16639 13701
rect 15396 13696 16639 13698
rect 15396 13640 16578 13696
rect 16634 13640 16639 13696
rect 15396 13638 16639 13640
rect 16990 13698 17050 13774
rect 17125 13832 17172 13836
rect 17236 13834 17242 13836
rect 20069 13834 20135 13837
rect 17125 13776 17130 13832
rect 17125 13772 17172 13776
rect 17236 13774 17282 13834
rect 17358 13832 20135 13834
rect 17358 13776 20074 13832
rect 20130 13776 20135 13832
rect 17358 13774 20135 13776
rect 17236 13772 17242 13774
rect 17125 13771 17191 13772
rect 17358 13698 17418 13774
rect 20069 13771 20135 13774
rect 21081 13834 21147 13837
rect 22200 13834 23000 13864
rect 21081 13832 23000 13834
rect 21081 13776 21086 13832
rect 21142 13776 23000 13832
rect 21081 13774 23000 13776
rect 21081 13771 21147 13774
rect 22200 13744 23000 13774
rect 16990 13638 17418 13698
rect 15396 13636 15402 13638
rect 16573 13635 16639 13638
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 5441 13560 7298 13562
rect 5441 13504 5446 13560
rect 5502 13504 7298 13560
rect 5441 13502 7298 13504
rect 5441 13499 5507 13502
rect 9254 13500 9260 13564
rect 9324 13562 9330 13564
rect 9673 13562 9739 13565
rect 9324 13560 9739 13562
rect 9324 13504 9678 13560
rect 9734 13504 9739 13560
rect 9324 13502 9739 13504
rect 9324 13500 9330 13502
rect 9673 13499 9739 13502
rect 10961 13562 11027 13565
rect 12198 13562 12204 13564
rect 10961 13560 12204 13562
rect 10961 13504 10966 13560
rect 11022 13504 12204 13560
rect 10961 13502 12204 13504
rect 10961 13499 11027 13502
rect 12198 13500 12204 13502
rect 12268 13500 12274 13564
rect 13486 13500 13492 13564
rect 13556 13562 13562 13564
rect 13813 13562 13879 13565
rect 13556 13560 13879 13562
rect 13556 13504 13818 13560
rect 13874 13504 13879 13560
rect 13556 13502 13879 13504
rect 13556 13500 13562 13502
rect 13813 13499 13879 13502
rect 14365 13562 14431 13565
rect 19517 13564 19583 13565
rect 14365 13560 17556 13562
rect 14365 13504 14370 13560
rect 14426 13504 17556 13560
rect 14365 13502 17556 13504
rect 14365 13499 14431 13502
rect 1945 13424 2790 13426
rect 1945 13368 1950 13424
rect 2006 13368 2790 13424
rect 1945 13366 2790 13368
rect 3877 13426 3943 13429
rect 4337 13426 4403 13429
rect 3877 13424 4403 13426
rect 3877 13368 3882 13424
rect 3938 13368 4342 13424
rect 4398 13368 4403 13424
rect 3877 13366 4403 13368
rect 1945 13363 2011 13366
rect 3877 13363 3943 13366
rect 4337 13363 4403 13366
rect 4521 13426 4587 13429
rect 13169 13426 13235 13429
rect 4521 13424 13235 13426
rect 4521 13368 4526 13424
rect 4582 13368 13174 13424
rect 13230 13368 13235 13424
rect 4521 13366 13235 13368
rect 4521 13363 4587 13366
rect 13169 13363 13235 13366
rect 13445 13426 13511 13429
rect 17309 13426 17375 13429
rect 13445 13424 17375 13426
rect 13445 13368 13450 13424
rect 13506 13368 17314 13424
rect 17370 13368 17375 13424
rect 13445 13366 17375 13368
rect 17496 13426 17556 13502
rect 19517 13560 19564 13564
rect 19628 13562 19634 13564
rect 21633 13562 21699 13565
rect 19628 13560 21699 13562
rect 19517 13504 19522 13560
rect 19628 13504 21638 13560
rect 21694 13504 21699 13560
rect 19517 13500 19564 13504
rect 19628 13502 21699 13504
rect 19628 13500 19634 13502
rect 19517 13499 19583 13500
rect 21633 13499 21699 13502
rect 19609 13426 19675 13429
rect 17496 13424 19675 13426
rect 17496 13368 19614 13424
rect 19670 13368 19675 13424
rect 17496 13366 19675 13368
rect 13445 13363 13511 13366
rect 17309 13363 17375 13366
rect 19609 13363 19675 13366
rect 21449 13426 21515 13429
rect 22200 13426 23000 13456
rect 21449 13424 23000 13426
rect 21449 13368 21454 13424
rect 21510 13368 23000 13424
rect 21449 13366 23000 13368
rect 21449 13363 21515 13366
rect 22200 13336 23000 13366
rect 2773 13290 2839 13293
rect 8017 13290 8083 13293
rect 9029 13290 9095 13293
rect 2773 13288 9095 13290
rect 2773 13232 2778 13288
rect 2834 13232 8022 13288
rect 8078 13232 9034 13288
rect 9090 13232 9095 13288
rect 2773 13230 9095 13232
rect 2773 13227 2839 13230
rect 8017 13227 8083 13230
rect 9029 13227 9095 13230
rect 9622 13228 9628 13292
rect 9692 13290 9698 13292
rect 10409 13290 10475 13293
rect 9692 13288 10475 13290
rect 9692 13232 10414 13288
rect 10470 13232 10475 13288
rect 9692 13230 10475 13232
rect 9692 13228 9698 13230
rect 10409 13227 10475 13230
rect 11102 13230 12450 13290
rect 790 13092 796 13156
rect 860 13154 866 13156
rect 860 13094 1042 13154
rect 860 13092 866 13094
rect 982 13018 1042 13094
rect 3366 13092 3372 13156
rect 3436 13154 3442 13156
rect 3436 13094 4170 13154
rect 3436 13092 3442 13094
rect 4110 13018 4170 13094
rect 6678 13092 6684 13156
rect 6748 13154 6754 13156
rect 11102 13154 11162 13230
rect 6748 13094 11162 13154
rect 12390 13154 12450 13230
rect 13670 13228 13676 13292
rect 13740 13290 13746 13292
rect 13813 13290 13879 13293
rect 13740 13288 13879 13290
rect 13740 13232 13818 13288
rect 13874 13232 13879 13288
rect 13740 13230 13879 13232
rect 13740 13228 13746 13230
rect 13813 13227 13879 13230
rect 14774 13228 14780 13292
rect 14844 13290 14850 13292
rect 16665 13290 16731 13293
rect 14844 13288 16731 13290
rect 14844 13232 16670 13288
rect 16726 13232 16731 13288
rect 14844 13230 16731 13232
rect 14844 13228 14850 13230
rect 16665 13227 16731 13230
rect 17033 13290 17099 13293
rect 18505 13290 18571 13293
rect 17033 13288 18571 13290
rect 17033 13232 17038 13288
rect 17094 13232 18510 13288
rect 18566 13232 18571 13288
rect 17033 13230 18571 13232
rect 17033 13227 17099 13230
rect 18505 13227 18571 13230
rect 15561 13154 15627 13157
rect 12390 13152 15627 13154
rect 12390 13096 15566 13152
rect 15622 13096 15627 13152
rect 12390 13094 15627 13096
rect 6748 13092 6754 13094
rect 15561 13091 15627 13094
rect 17585 13154 17651 13157
rect 18086 13154 18092 13156
rect 17585 13152 18092 13154
rect 17585 13096 17590 13152
rect 17646 13096 18092 13152
rect 17585 13094 18092 13096
rect 17585 13091 17651 13094
rect 18086 13092 18092 13094
rect 18156 13092 18162 13156
rect 20069 13154 20135 13157
rect 21398 13154 21404 13156
rect 20069 13152 21404 13154
rect 20069 13096 20074 13152
rect 20130 13096 21404 13152
rect 20069 13094 21404 13096
rect 20069 13091 20135 13094
rect 21398 13092 21404 13094
rect 21468 13092 21474 13156
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 5390 13018 5396 13020
rect 982 12958 1778 13018
rect 4110 12958 5396 13018
rect 0 12882 800 12912
rect 1485 12882 1551 12885
rect 0 12880 1551 12882
rect 0 12824 1490 12880
rect 1546 12824 1551 12880
rect 0 12822 1551 12824
rect 1718 12882 1778 12958
rect 5390 12956 5396 12958
rect 5460 12956 5466 13020
rect 10961 13018 11027 13021
rect 6548 13016 11027 13018
rect 6548 12960 10966 13016
rect 11022 12960 11027 13016
rect 6548 12958 11027 12960
rect 5993 12882 6059 12885
rect 6548 12882 6608 12958
rect 10961 12955 11027 12958
rect 12157 13018 12223 13021
rect 12157 13016 16452 13018
rect 12157 12960 12162 13016
rect 12218 12960 16452 13016
rect 12157 12958 16452 12960
rect 12157 12955 12223 12958
rect 1718 12822 2790 12882
rect 0 12792 800 12822
rect 1485 12819 1551 12822
rect 2730 12746 2790 12822
rect 5993 12880 6608 12882
rect 5993 12824 5998 12880
rect 6054 12824 6608 12880
rect 5993 12822 6608 12824
rect 5993 12819 6059 12822
rect 8518 12820 8524 12884
rect 8588 12882 8594 12884
rect 12617 12882 12683 12885
rect 12801 12882 12867 12885
rect 15694 12882 15700 12884
rect 8588 12880 12683 12882
rect 8588 12824 12622 12880
rect 12678 12824 12683 12880
rect 8588 12822 12683 12824
rect 8588 12820 8594 12822
rect 12617 12819 12683 12822
rect 12758 12880 15700 12882
rect 12758 12824 12806 12880
rect 12862 12824 15700 12880
rect 12758 12822 15700 12824
rect 12758 12819 12867 12822
rect 15694 12820 15700 12822
rect 15764 12820 15770 12884
rect 15929 12882 15995 12885
rect 16062 12882 16068 12884
rect 15929 12880 16068 12882
rect 15929 12824 15934 12880
rect 15990 12824 16068 12880
rect 15929 12822 16068 12824
rect 15929 12819 15995 12822
rect 16062 12820 16068 12822
rect 16132 12820 16138 12884
rect 16392 12882 16452 12958
rect 18413 12882 18479 12885
rect 16392 12880 18479 12882
rect 16392 12824 18418 12880
rect 18474 12824 18479 12880
rect 16392 12822 18479 12824
rect 18413 12819 18479 12822
rect 21449 12882 21515 12885
rect 22200 12882 23000 12912
rect 21449 12880 23000 12882
rect 21449 12824 21454 12880
rect 21510 12824 23000 12880
rect 21449 12822 23000 12824
rect 21449 12819 21515 12822
rect 4286 12746 4292 12748
rect 2730 12686 4292 12746
rect 4286 12684 4292 12686
rect 4356 12684 4362 12748
rect 4429 12746 4495 12749
rect 8293 12746 8359 12749
rect 9857 12746 9923 12749
rect 12382 12746 12388 12748
rect 4429 12744 8359 12746
rect 4429 12688 4434 12744
rect 4490 12688 8298 12744
rect 8354 12688 8359 12744
rect 4429 12686 8359 12688
rect 4429 12683 4495 12686
rect 8293 12683 8359 12686
rect 8480 12744 12388 12746
rect 8480 12688 9862 12744
rect 9918 12688 12388 12744
rect 8480 12686 12388 12688
rect 2814 12548 2820 12612
rect 2884 12610 2890 12612
rect 2957 12610 3023 12613
rect 2884 12608 3023 12610
rect 2884 12552 2962 12608
rect 3018 12552 3023 12608
rect 2884 12550 3023 12552
rect 2884 12548 2890 12550
rect 2957 12547 3023 12550
rect 5349 12610 5415 12613
rect 8480 12610 8540 12686
rect 9857 12683 9923 12686
rect 12382 12684 12388 12686
rect 12452 12684 12458 12748
rect 12525 12746 12591 12749
rect 12758 12746 12818 12819
rect 22200 12792 23000 12822
rect 12525 12744 12818 12746
rect 12525 12688 12530 12744
rect 12586 12688 12818 12744
rect 12525 12686 12818 12688
rect 13261 12746 13327 12749
rect 17902 12746 17908 12748
rect 13261 12744 17908 12746
rect 13261 12688 13266 12744
rect 13322 12688 17908 12744
rect 13261 12686 17908 12688
rect 12525 12683 12591 12686
rect 13261 12683 13327 12686
rect 17902 12684 17908 12686
rect 17972 12684 17978 12748
rect 5349 12608 8540 12610
rect 5349 12552 5354 12608
rect 5410 12552 8540 12608
rect 5349 12550 8540 12552
rect 10041 12610 10107 12613
rect 10174 12610 10180 12612
rect 10041 12608 10180 12610
rect 10041 12552 10046 12608
rect 10102 12552 10180 12608
rect 10041 12550 10180 12552
rect 5349 12547 5415 12550
rect 10041 12547 10107 12550
rect 10174 12548 10180 12550
rect 10244 12548 10250 12612
rect 11094 12548 11100 12612
rect 11164 12610 11170 12612
rect 13445 12610 13511 12613
rect 11164 12608 13511 12610
rect 11164 12552 13450 12608
rect 13506 12552 13511 12608
rect 11164 12550 13511 12552
rect 11164 12548 11170 12550
rect 13445 12547 13511 12550
rect 14457 12610 14523 12613
rect 15142 12610 15148 12612
rect 14457 12608 15148 12610
rect 14457 12552 14462 12608
rect 14518 12552 15148 12608
rect 14457 12550 15148 12552
rect 14457 12547 14523 12550
rect 15142 12548 15148 12550
rect 15212 12548 15218 12612
rect 15326 12548 15332 12612
rect 15396 12548 15402 12612
rect 15878 12548 15884 12612
rect 15948 12610 15954 12612
rect 16205 12610 16271 12613
rect 15948 12608 16271 12610
rect 15948 12552 16210 12608
rect 16266 12552 16271 12608
rect 15948 12550 16271 12552
rect 15948 12548 15954 12550
rect 3543 12544 3863 12545
rect 0 12474 800 12504
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 1485 12474 1551 12477
rect 0 12472 1551 12474
rect 0 12416 1490 12472
rect 1546 12416 1551 12472
rect 0 12414 1551 12416
rect 0 12384 800 12414
rect 1485 12411 1551 12414
rect 2814 12412 2820 12476
rect 2884 12474 2890 12476
rect 3049 12474 3115 12477
rect 8109 12474 8175 12477
rect 2884 12472 3115 12474
rect 2884 12416 3054 12472
rect 3110 12416 3115 12472
rect 2884 12414 3115 12416
rect 2884 12412 2890 12414
rect 3049 12411 3115 12414
rect 6502 12472 8175 12474
rect 6502 12416 8114 12472
rect 8170 12416 8175 12472
rect 6502 12414 8175 12416
rect 2998 12276 3004 12340
rect 3068 12338 3074 12340
rect 6502 12338 6562 12414
rect 8109 12411 8175 12414
rect 9673 12474 9739 12477
rect 14365 12474 14431 12477
rect 15334 12474 15394 12548
rect 16205 12547 16271 12550
rect 16757 12610 16823 12613
rect 17350 12610 17356 12612
rect 16757 12608 17356 12610
rect 16757 12552 16762 12608
rect 16818 12552 17356 12608
rect 16757 12550 17356 12552
rect 16757 12547 16823 12550
rect 17350 12548 17356 12550
rect 17420 12610 17426 12612
rect 18229 12610 18295 12613
rect 17420 12608 18295 12610
rect 17420 12552 18234 12608
rect 18290 12552 18295 12608
rect 17420 12550 18295 12552
rect 17420 12548 17426 12550
rect 18229 12547 18295 12550
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 12479 19457 12480
rect 9673 12472 12772 12474
rect 9673 12416 9678 12472
rect 9734 12416 12772 12472
rect 9673 12414 12772 12416
rect 9673 12411 9739 12414
rect 3068 12278 6562 12338
rect 6637 12338 6703 12341
rect 8293 12338 8359 12341
rect 6637 12336 8359 12338
rect 6637 12280 6642 12336
rect 6698 12280 8298 12336
rect 8354 12280 8359 12336
rect 6637 12278 8359 12280
rect 3068 12276 3074 12278
rect 6637 12275 6703 12278
rect 8293 12275 8359 12278
rect 9673 12338 9739 12341
rect 12525 12338 12591 12341
rect 9673 12336 12591 12338
rect 9673 12280 9678 12336
rect 9734 12280 12530 12336
rect 12586 12280 12591 12336
rect 9673 12278 12591 12280
rect 9673 12275 9739 12278
rect 12525 12275 12591 12278
rect 1393 12202 1459 12205
rect 2681 12202 2747 12205
rect 4889 12202 4955 12205
rect 8385 12202 8451 12205
rect 10041 12204 10107 12205
rect 1393 12200 8451 12202
rect 1393 12144 1398 12200
rect 1454 12144 2686 12200
rect 2742 12144 4894 12200
rect 4950 12144 8390 12200
rect 8446 12144 8451 12200
rect 1393 12142 8451 12144
rect 1393 12139 1459 12142
rect 2681 12139 2747 12142
rect 4889 12139 4955 12142
rect 8385 12139 8451 12142
rect 9990 12140 9996 12204
rect 10060 12202 10107 12204
rect 12249 12202 12315 12205
rect 12525 12202 12591 12205
rect 10060 12200 10152 12202
rect 10102 12144 10152 12200
rect 10060 12142 10152 12144
rect 12249 12200 12591 12202
rect 12249 12144 12254 12200
rect 12310 12144 12530 12200
rect 12586 12144 12591 12200
rect 12249 12142 12591 12144
rect 12712 12202 12772 12414
rect 14365 12472 15394 12474
rect 14365 12416 14370 12472
rect 14426 12416 15394 12472
rect 14365 12414 15394 12416
rect 14365 12411 14431 12414
rect 15694 12412 15700 12476
rect 15764 12474 15770 12476
rect 16941 12474 17007 12477
rect 15764 12472 17007 12474
rect 15764 12416 16946 12472
rect 17002 12416 17007 12472
rect 15764 12414 17007 12416
rect 15764 12412 15770 12414
rect 16941 12411 17007 12414
rect 20253 12474 20319 12477
rect 20478 12474 20484 12476
rect 20253 12472 20484 12474
rect 20253 12416 20258 12472
rect 20314 12416 20484 12472
rect 20253 12414 20484 12416
rect 20253 12411 20319 12414
rect 20478 12412 20484 12414
rect 20548 12412 20554 12476
rect 21449 12474 21515 12477
rect 22200 12474 23000 12504
rect 21449 12472 23000 12474
rect 21449 12416 21454 12472
rect 21510 12416 23000 12472
rect 21449 12414 23000 12416
rect 21449 12411 21515 12414
rect 22200 12384 23000 12414
rect 12985 12340 13051 12341
rect 12934 12276 12940 12340
rect 13004 12338 13051 12340
rect 13261 12338 13327 12341
rect 21449 12338 21515 12341
rect 13004 12336 13096 12338
rect 13046 12280 13096 12336
rect 13004 12278 13096 12280
rect 13261 12336 21515 12338
rect 13261 12280 13266 12336
rect 13322 12280 21454 12336
rect 21510 12280 21515 12336
rect 13261 12278 21515 12280
rect 13004 12276 13051 12278
rect 12985 12275 13051 12276
rect 13261 12275 13327 12278
rect 21449 12275 21515 12278
rect 16573 12202 16639 12205
rect 12712 12200 16639 12202
rect 12712 12144 16578 12200
rect 16634 12144 16639 12200
rect 12712 12142 16639 12144
rect 10060 12140 10107 12142
rect 10041 12139 10107 12140
rect 12249 12139 12315 12142
rect 12525 12139 12591 12142
rect 16573 12139 16639 12142
rect 16757 12202 16823 12205
rect 17718 12202 17724 12204
rect 16757 12200 17724 12202
rect 16757 12144 16762 12200
rect 16818 12144 17724 12200
rect 16757 12142 17724 12144
rect 16757 12139 16823 12142
rect 17718 12140 17724 12142
rect 17788 12140 17794 12204
rect 19609 12202 19675 12205
rect 21214 12202 21220 12204
rect 19609 12200 21220 12202
rect 19609 12144 19614 12200
rect 19670 12144 21220 12200
rect 19609 12142 21220 12144
rect 19609 12139 19675 12142
rect 21214 12140 21220 12142
rect 21284 12140 21290 12204
rect 0 12066 800 12096
rect 1853 12066 1919 12069
rect 0 12064 1919 12066
rect 0 12008 1858 12064
rect 1914 12008 1919 12064
rect 0 12006 1919 12008
rect 0 11976 800 12006
rect 1853 12003 1919 12006
rect 2589 12066 2655 12069
rect 2814 12066 2820 12068
rect 2589 12064 2820 12066
rect 2589 12008 2594 12064
rect 2650 12008 2820 12064
rect 2589 12006 2820 12008
rect 2589 12003 2655 12006
rect 2814 12004 2820 12006
rect 2884 12004 2890 12068
rect 7373 12066 7439 12069
rect 10910 12066 10916 12068
rect 7373 12064 10916 12066
rect 7373 12008 7378 12064
rect 7434 12008 10916 12064
rect 7373 12006 10916 12008
rect 7373 12003 7439 12006
rect 10910 12004 10916 12006
rect 10980 12004 10986 12068
rect 12525 12066 12591 12069
rect 16297 12068 16363 12069
rect 15694 12066 15700 12068
rect 12525 12064 15700 12066
rect 12525 12008 12530 12064
rect 12586 12008 15700 12064
rect 12525 12006 15700 12008
rect 12525 12003 12591 12006
rect 15694 12004 15700 12006
rect 15764 12004 15770 12068
rect 16246 12004 16252 12068
rect 16316 12066 16363 12068
rect 17309 12066 17375 12069
rect 19425 12066 19491 12069
rect 16316 12064 16408 12066
rect 16358 12008 16408 12064
rect 16316 12006 16408 12008
rect 17309 12064 19491 12066
rect 17309 12008 17314 12064
rect 17370 12008 19430 12064
rect 19486 12008 19491 12064
rect 17309 12006 19491 12008
rect 16316 12004 16363 12006
rect 16297 12003 16363 12004
rect 17309 12003 17375 12006
rect 19425 12003 19491 12006
rect 19793 12066 19859 12069
rect 20713 12066 20779 12069
rect 19793 12064 20779 12066
rect 19793 12008 19798 12064
rect 19854 12008 20718 12064
rect 20774 12008 20779 12064
rect 19793 12006 20779 12008
rect 19793 12003 19859 12006
rect 20713 12003 20779 12006
rect 21449 12066 21515 12069
rect 22200 12066 23000 12096
rect 21449 12064 23000 12066
rect 21449 12008 21454 12064
rect 21510 12008 23000 12064
rect 21449 12006 23000 12008
rect 21449 12003 21515 12006
rect 6142 12000 6462 12001
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 22200 11976 23000 12006
rect 16538 11935 16858 11936
rect 5206 11868 5212 11932
rect 5276 11930 5282 11932
rect 5809 11930 5875 11933
rect 6637 11932 6703 11933
rect 6637 11930 6684 11932
rect 5276 11928 5875 11930
rect 5276 11872 5814 11928
rect 5870 11872 5875 11928
rect 5276 11870 5875 11872
rect 6592 11928 6684 11930
rect 6592 11872 6642 11928
rect 6592 11870 6684 11872
rect 5276 11868 5282 11870
rect 5809 11867 5875 11870
rect 6637 11868 6684 11870
rect 6748 11868 6754 11932
rect 7414 11868 7420 11932
rect 7484 11930 7490 11932
rect 9673 11930 9739 11933
rect 7484 11928 9739 11930
rect 7484 11872 9678 11928
rect 9734 11872 9739 11928
rect 7484 11870 9739 11872
rect 7484 11868 7490 11870
rect 6637 11867 6703 11868
rect 9673 11867 9739 11870
rect 12801 11930 12867 11933
rect 17033 11930 17099 11933
rect 18638 11930 18644 11932
rect 12801 11928 16268 11930
rect 12801 11872 12806 11928
rect 12862 11872 16268 11928
rect 12801 11870 16268 11872
rect 12801 11867 12867 11870
rect 5349 11794 5415 11797
rect 7373 11794 7439 11797
rect 5349 11792 7439 11794
rect 5349 11736 5354 11792
rect 5410 11736 7378 11792
rect 7434 11736 7439 11792
rect 5349 11734 7439 11736
rect 5349 11731 5415 11734
rect 7373 11731 7439 11734
rect 8385 11794 8451 11797
rect 16208 11794 16268 11870
rect 17033 11928 18644 11930
rect 17033 11872 17038 11928
rect 17094 11872 18644 11928
rect 17033 11870 18644 11872
rect 17033 11867 17099 11870
rect 18638 11868 18644 11870
rect 18708 11868 18714 11932
rect 19333 11930 19399 11933
rect 19701 11932 19767 11933
rect 19701 11930 19748 11932
rect 19333 11928 19748 11930
rect 19333 11872 19338 11928
rect 19394 11872 19706 11928
rect 19333 11870 19748 11872
rect 19333 11867 19399 11870
rect 19701 11868 19748 11870
rect 19812 11868 19818 11932
rect 20805 11930 20871 11933
rect 21265 11930 21331 11933
rect 20805 11928 21331 11930
rect 20805 11872 20810 11928
rect 20866 11872 21270 11928
rect 21326 11872 21331 11928
rect 20805 11870 21331 11872
rect 19701 11867 19767 11868
rect 20805 11867 20871 11870
rect 21265 11867 21331 11870
rect 20805 11794 20871 11797
rect 8385 11792 16130 11794
rect 8385 11736 8390 11792
rect 8446 11736 16130 11792
rect 8385 11734 16130 11736
rect 16208 11792 20871 11794
rect 16208 11736 20810 11792
rect 20866 11736 20871 11792
rect 16208 11734 20871 11736
rect 8385 11731 8451 11734
rect 0 11658 800 11688
rect 2129 11658 2195 11661
rect 0 11656 2195 11658
rect 0 11600 2134 11656
rect 2190 11600 2195 11656
rect 0 11598 2195 11600
rect 0 11568 800 11598
rect 2129 11595 2195 11598
rect 2405 11658 2471 11661
rect 5942 11658 5948 11660
rect 2405 11656 5948 11658
rect 2405 11600 2410 11656
rect 2466 11600 5948 11656
rect 2405 11598 5948 11600
rect 2405 11595 2471 11598
rect 5942 11596 5948 11598
rect 6012 11658 6018 11660
rect 10041 11658 10107 11661
rect 12014 11658 12020 11660
rect 6012 11598 9920 11658
rect 6012 11596 6018 11598
rect 5073 11522 5139 11525
rect 7414 11522 7420 11524
rect 5073 11520 7420 11522
rect 5073 11464 5078 11520
rect 5134 11464 7420 11520
rect 5073 11462 7420 11464
rect 5073 11459 5139 11462
rect 7414 11460 7420 11462
rect 7484 11460 7490 11524
rect 9860 11522 9920 11598
rect 10041 11656 12020 11658
rect 10041 11600 10046 11656
rect 10102 11600 12020 11656
rect 10041 11598 12020 11600
rect 10041 11595 10107 11598
rect 12014 11596 12020 11598
rect 12084 11658 12090 11660
rect 13118 11658 13124 11660
rect 12084 11598 13124 11658
rect 12084 11596 12090 11598
rect 13118 11596 13124 11598
rect 13188 11658 13194 11660
rect 13445 11658 13511 11661
rect 13188 11656 13511 11658
rect 13188 11600 13450 11656
rect 13506 11600 13511 11656
rect 13188 11598 13511 11600
rect 13188 11596 13194 11598
rect 13445 11595 13511 11598
rect 13670 11596 13676 11660
rect 13740 11658 13746 11660
rect 14089 11658 14155 11661
rect 13740 11656 14155 11658
rect 13740 11600 14094 11656
rect 14150 11600 14155 11656
rect 13740 11598 14155 11600
rect 16070 11658 16130 11734
rect 20805 11731 20871 11734
rect 19885 11660 19951 11661
rect 17718 11658 17724 11660
rect 16070 11598 17724 11658
rect 13740 11596 13746 11598
rect 14089 11595 14155 11598
rect 17718 11596 17724 11598
rect 17788 11596 17794 11660
rect 19885 11658 19932 11660
rect 19840 11656 19932 11658
rect 19840 11600 19890 11656
rect 19840 11598 19932 11600
rect 19885 11596 19932 11598
rect 19996 11596 20002 11660
rect 21541 11658 21607 11661
rect 22200 11658 23000 11688
rect 21541 11656 23000 11658
rect 21541 11600 21546 11656
rect 21602 11600 23000 11656
rect 21541 11598 23000 11600
rect 19885 11595 19951 11596
rect 21541 11595 21607 11598
rect 22200 11568 23000 11598
rect 12566 11522 12572 11524
rect 9860 11462 12572 11522
rect 12566 11460 12572 11462
rect 12636 11522 12642 11524
rect 12801 11522 12867 11525
rect 12636 11520 12867 11522
rect 12636 11464 12806 11520
rect 12862 11464 12867 11520
rect 12636 11462 12867 11464
rect 12636 11460 12642 11462
rect 12801 11459 12867 11462
rect 13169 11522 13235 11525
rect 13813 11522 13879 11525
rect 13169 11520 13879 11522
rect 13169 11464 13174 11520
rect 13230 11464 13818 11520
rect 13874 11464 13879 11520
rect 13169 11462 13879 11464
rect 13169 11459 13235 11462
rect 13813 11459 13879 11462
rect 16297 11522 16363 11525
rect 18781 11522 18847 11525
rect 16297 11520 18847 11522
rect 16297 11464 16302 11520
rect 16358 11464 18786 11520
rect 18842 11464 18847 11520
rect 16297 11462 18847 11464
rect 16297 11459 16363 11462
rect 18781 11459 18847 11462
rect 3543 11456 3863 11457
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 1485 11386 1551 11389
rect 6545 11386 6611 11389
rect 1485 11384 2100 11386
rect 1485 11328 1490 11384
rect 1546 11328 2100 11384
rect 1485 11326 2100 11328
rect 1485 11323 1551 11326
rect 0 11250 800 11280
rect 1853 11250 1919 11253
rect 0 11248 1919 11250
rect 0 11192 1858 11248
rect 1914 11192 1919 11248
rect 0 11190 1919 11192
rect 2040 11250 2100 11326
rect 3926 11384 6611 11386
rect 3926 11328 6550 11384
rect 6606 11328 6611 11384
rect 3926 11326 6611 11328
rect 3926 11250 3986 11326
rect 6545 11323 6611 11326
rect 6678 11324 6684 11388
rect 6748 11386 6754 11388
rect 6913 11386 6979 11389
rect 8017 11388 8083 11389
rect 6748 11384 6979 11386
rect 6748 11328 6918 11384
rect 6974 11328 6979 11384
rect 6748 11326 6979 11328
rect 6748 11324 6754 11326
rect 6913 11323 6979 11326
rect 7966 11324 7972 11388
rect 8036 11386 8083 11388
rect 8036 11384 8128 11386
rect 8078 11328 8128 11384
rect 8036 11326 8128 11328
rect 8036 11324 8083 11326
rect 9254 11324 9260 11388
rect 9324 11386 9330 11388
rect 9806 11386 9812 11388
rect 9324 11326 9812 11386
rect 9324 11324 9330 11326
rect 9806 11324 9812 11326
rect 9876 11324 9882 11388
rect 11830 11324 11836 11388
rect 11900 11386 11906 11388
rect 12065 11386 12131 11389
rect 11900 11384 12131 11386
rect 11900 11328 12070 11384
rect 12126 11328 12131 11384
rect 11900 11326 12131 11328
rect 11900 11324 11906 11326
rect 8017 11323 8083 11324
rect 12065 11323 12131 11326
rect 14958 11324 14964 11388
rect 15028 11386 15034 11388
rect 18270 11386 18276 11388
rect 15028 11326 18276 11386
rect 15028 11324 15034 11326
rect 18270 11324 18276 11326
rect 18340 11324 18346 11388
rect 21541 11386 21607 11389
rect 19566 11384 21607 11386
rect 19566 11328 21546 11384
rect 21602 11328 21607 11384
rect 19566 11326 21607 11328
rect 2040 11190 3986 11250
rect 5165 11250 5231 11253
rect 10174 11250 10180 11252
rect 5165 11248 10180 11250
rect 5165 11192 5170 11248
rect 5226 11192 10180 11248
rect 5165 11190 10180 11192
rect 0 11160 800 11190
rect 1853 11187 1919 11190
rect 5165 11187 5231 11190
rect 10174 11188 10180 11190
rect 10244 11188 10250 11252
rect 10961 11250 11027 11253
rect 12566 11250 12572 11252
rect 10961 11248 12572 11250
rect 10961 11192 10966 11248
rect 11022 11192 12572 11248
rect 10961 11190 12572 11192
rect 10961 11187 11027 11190
rect 12566 11188 12572 11190
rect 12636 11250 12642 11252
rect 12709 11250 12775 11253
rect 12636 11248 12775 11250
rect 12636 11192 12714 11248
rect 12770 11192 12775 11248
rect 12636 11190 12775 11192
rect 12636 11188 12642 11190
rect 12709 11187 12775 11190
rect 13118 11188 13124 11252
rect 13188 11250 13194 11252
rect 15193 11250 15259 11253
rect 13188 11248 15259 11250
rect 13188 11192 15198 11248
rect 15254 11192 15259 11248
rect 13188 11190 15259 11192
rect 13188 11188 13194 11190
rect 15193 11187 15259 11190
rect 15929 11250 15995 11253
rect 19566 11250 19626 11326
rect 21541 11323 21607 11326
rect 15929 11248 19626 11250
rect 15929 11192 15934 11248
rect 15990 11192 19626 11248
rect 15929 11190 19626 11192
rect 21449 11250 21515 11253
rect 22200 11250 23000 11280
rect 21449 11248 23000 11250
rect 21449 11192 21454 11248
rect 21510 11192 23000 11248
rect 21449 11190 23000 11192
rect 15929 11187 15995 11190
rect 21449 11187 21515 11190
rect 22200 11160 23000 11190
rect 2681 11114 2747 11117
rect 2814 11114 2820 11116
rect 2681 11112 2820 11114
rect 2681 11056 2686 11112
rect 2742 11056 2820 11112
rect 2681 11054 2820 11056
rect 2681 11051 2747 11054
rect 2814 11052 2820 11054
rect 2884 11052 2890 11116
rect 3366 11052 3372 11116
rect 3436 11114 3442 11116
rect 3785 11114 3851 11117
rect 7281 11114 7347 11117
rect 9213 11116 9279 11117
rect 3436 11112 7347 11114
rect 3436 11056 3790 11112
rect 3846 11056 7286 11112
rect 7342 11056 7347 11112
rect 3436 11054 7347 11056
rect 3436 11052 3442 11054
rect 3785 11051 3851 11054
rect 7281 11051 7347 11054
rect 7414 11052 7420 11116
rect 7484 11114 7490 11116
rect 8518 11114 8524 11116
rect 7484 11054 8524 11114
rect 7484 11052 7490 11054
rect 8518 11052 8524 11054
rect 8588 11052 8594 11116
rect 9213 11114 9260 11116
rect 9168 11112 9260 11114
rect 9168 11056 9218 11112
rect 9168 11054 9260 11056
rect 9213 11052 9260 11054
rect 9324 11052 9330 11116
rect 10225 11114 10291 11117
rect 10358 11114 10364 11116
rect 10225 11112 10364 11114
rect 10225 11056 10230 11112
rect 10286 11056 10364 11112
rect 10225 11054 10364 11056
rect 9213 11051 9279 11052
rect 10225 11051 10291 11054
rect 10358 11052 10364 11054
rect 10428 11052 10434 11116
rect 15653 11114 15719 11117
rect 18086 11114 18092 11116
rect 10550 11112 15719 11114
rect 10550 11056 15658 11112
rect 15714 11056 15719 11112
rect 10550 11054 15719 11056
rect 1025 10978 1091 10981
rect 1710 10978 1716 10980
rect 1025 10976 1716 10978
rect 1025 10920 1030 10976
rect 1086 10920 1716 10976
rect 1025 10918 1716 10920
rect 1025 10915 1091 10918
rect 1710 10916 1716 10918
rect 1780 10916 1786 10980
rect 6821 10978 6887 10981
rect 10550 10978 10610 11054
rect 15653 11051 15719 11054
rect 15886 11054 18092 11114
rect 6821 10976 10610 10978
rect 6821 10920 6826 10976
rect 6882 10920 10610 10976
rect 6821 10918 10610 10920
rect 11789 10978 11855 10981
rect 15886 10978 15946 11054
rect 18086 11052 18092 11054
rect 18156 11052 18162 11116
rect 19558 11052 19564 11116
rect 19628 11114 19634 11116
rect 20161 11114 20227 11117
rect 19628 11112 20227 11114
rect 19628 11056 20166 11112
rect 20222 11056 20227 11112
rect 19628 11054 20227 11056
rect 19628 11052 19634 11054
rect 20161 11051 20227 11054
rect 20805 11114 20871 11117
rect 21950 11114 21956 11116
rect 20805 11112 21956 11114
rect 20805 11056 20810 11112
rect 20866 11056 21956 11112
rect 20805 11054 21956 11056
rect 20805 11051 20871 11054
rect 21950 11052 21956 11054
rect 22020 11052 22026 11116
rect 11789 10976 15946 10978
rect 11789 10920 11794 10976
rect 11850 10920 15946 10976
rect 11789 10918 15946 10920
rect 6821 10915 6887 10918
rect 11789 10915 11855 10918
rect 6142 10912 6462 10913
rect 0 10842 800 10872
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 1485 10842 1551 10845
rect 4981 10842 5047 10845
rect 5942 10842 5948 10844
rect 0 10840 2790 10842
rect 0 10784 1490 10840
rect 1546 10784 2790 10840
rect 0 10782 2790 10784
rect 0 10752 800 10782
rect 1485 10779 1551 10782
rect 2730 10706 2790 10782
rect 4981 10840 5948 10842
rect 4981 10784 4986 10840
rect 5042 10784 5948 10840
rect 4981 10782 5948 10784
rect 4981 10779 5047 10782
rect 5942 10780 5948 10782
rect 6012 10780 6018 10844
rect 7925 10842 7991 10845
rect 9949 10842 10015 10845
rect 7925 10840 10015 10842
rect 7925 10784 7930 10840
rect 7986 10784 9954 10840
rect 10010 10784 10015 10840
rect 7925 10782 10015 10784
rect 7925 10779 7991 10782
rect 9949 10779 10015 10782
rect 12198 10780 12204 10844
rect 12268 10842 12274 10844
rect 21081 10842 21147 10845
rect 22200 10842 23000 10872
rect 12268 10782 16314 10842
rect 12268 10780 12274 10782
rect 13077 10706 13143 10709
rect 2730 10704 13143 10706
rect 2730 10648 13082 10704
rect 13138 10648 13143 10704
rect 2730 10646 13143 10648
rect 13077 10643 13143 10646
rect 13629 10706 13695 10709
rect 16254 10706 16314 10782
rect 21081 10840 23000 10842
rect 21081 10784 21086 10840
rect 21142 10784 23000 10840
rect 21081 10782 23000 10784
rect 21081 10779 21147 10782
rect 22200 10752 23000 10782
rect 20345 10706 20411 10709
rect 13629 10704 15946 10706
rect 13629 10648 13634 10704
rect 13690 10648 15946 10704
rect 13629 10646 15946 10648
rect 16254 10704 20411 10706
rect 16254 10648 20350 10704
rect 20406 10648 20411 10704
rect 16254 10646 20411 10648
rect 13629 10643 13695 10646
rect 7281 10570 7347 10573
rect 3374 10568 7347 10570
rect 3374 10512 7286 10568
rect 7342 10512 7347 10568
rect 3374 10510 7347 10512
rect 0 10434 800 10464
rect 2773 10434 2839 10437
rect 0 10432 2839 10434
rect 0 10376 2778 10432
rect 2834 10376 2839 10432
rect 0 10374 2839 10376
rect 0 10344 800 10374
rect 2773 10371 2839 10374
rect 1669 10026 1735 10029
rect 3374 10026 3434 10510
rect 7281 10507 7347 10510
rect 7782 10508 7788 10572
rect 7852 10570 7858 10572
rect 10225 10570 10291 10573
rect 12198 10570 12204 10572
rect 7852 10510 10104 10570
rect 7852 10508 7858 10510
rect 3969 10434 4035 10437
rect 4337 10434 4403 10437
rect 6545 10434 6611 10437
rect 6678 10434 6684 10436
rect 3969 10432 5964 10434
rect 3969 10376 3974 10432
rect 4030 10376 4342 10432
rect 4398 10376 5964 10432
rect 3969 10374 5964 10376
rect 3969 10371 4035 10374
rect 4337 10371 4403 10374
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 4245 10298 4311 10301
rect 5257 10298 5323 10301
rect 4245 10296 5323 10298
rect 4245 10240 4250 10296
rect 4306 10240 5262 10296
rect 5318 10240 5323 10296
rect 4245 10238 5323 10240
rect 4245 10235 4311 10238
rect 5257 10235 5323 10238
rect 5390 10236 5396 10300
rect 5460 10298 5466 10300
rect 5758 10298 5764 10300
rect 5460 10238 5764 10298
rect 5460 10236 5466 10238
rect 5758 10236 5764 10238
rect 5828 10236 5834 10300
rect 5904 10298 5964 10374
rect 6545 10432 6684 10434
rect 6545 10376 6550 10432
rect 6606 10376 6684 10432
rect 6545 10374 6684 10376
rect 6545 10371 6611 10374
rect 6678 10372 6684 10374
rect 6748 10372 6754 10436
rect 7598 10372 7604 10436
rect 7668 10434 7674 10436
rect 8569 10434 8635 10437
rect 7668 10432 8635 10434
rect 7668 10376 8574 10432
rect 8630 10376 8635 10432
rect 7668 10374 8635 10376
rect 10044 10434 10104 10510
rect 10225 10568 12204 10570
rect 10225 10512 10230 10568
rect 10286 10512 12204 10568
rect 10225 10510 12204 10512
rect 10225 10507 10291 10510
rect 12198 10508 12204 10510
rect 12268 10508 12274 10572
rect 15745 10570 15811 10573
rect 13356 10568 15811 10570
rect 13356 10512 15750 10568
rect 15806 10512 15811 10568
rect 13356 10510 15811 10512
rect 15886 10570 15946 10646
rect 20345 10643 20411 10646
rect 19609 10570 19675 10573
rect 15886 10568 19675 10570
rect 15886 10512 19614 10568
rect 19670 10512 19675 10568
rect 15886 10510 19675 10512
rect 13356 10434 13416 10510
rect 15745 10507 15811 10510
rect 19609 10507 19675 10510
rect 20253 10570 20319 10573
rect 20478 10570 20484 10572
rect 20253 10568 20484 10570
rect 20253 10512 20258 10568
rect 20314 10512 20484 10568
rect 20253 10510 20484 10512
rect 20253 10507 20319 10510
rect 20478 10508 20484 10510
rect 20548 10508 20554 10572
rect 10044 10374 13416 10434
rect 13537 10434 13603 10437
rect 13813 10434 13879 10437
rect 13537 10432 13879 10434
rect 13537 10376 13542 10432
rect 13598 10376 13818 10432
rect 13874 10376 13879 10432
rect 13537 10374 13879 10376
rect 7668 10372 7674 10374
rect 8569 10371 8635 10374
rect 13537 10371 13603 10374
rect 13813 10371 13879 10374
rect 15510 10372 15516 10436
rect 15580 10434 15586 10436
rect 17350 10434 17356 10436
rect 15580 10374 17356 10434
rect 15580 10372 15586 10374
rect 17350 10372 17356 10374
rect 17420 10372 17426 10436
rect 20989 10434 21055 10437
rect 21449 10434 21515 10437
rect 22200 10434 23000 10464
rect 20989 10432 23000 10434
rect 20989 10376 20994 10432
rect 21050 10376 21454 10432
rect 21510 10376 23000 10432
rect 20989 10374 23000 10376
rect 20989 10371 21055 10374
rect 21449 10371 21515 10374
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 22200 10344 23000 10374
rect 19137 10303 19457 10304
rect 6540 10298 6546 10300
rect 5904 10238 6546 10298
rect 6540 10236 6546 10238
rect 6610 10236 6616 10300
rect 9581 10298 9647 10301
rect 9581 10296 13876 10298
rect 9581 10240 9586 10296
rect 9642 10240 13876 10296
rect 9581 10238 13876 10240
rect 9581 10235 9647 10238
rect 3785 10162 3851 10165
rect 10041 10162 10107 10165
rect 3785 10160 10107 10162
rect 3785 10104 3790 10160
rect 3846 10104 10046 10160
rect 10102 10104 10107 10160
rect 3785 10102 10107 10104
rect 3785 10099 3851 10102
rect 10041 10099 10107 10102
rect 11697 10162 11763 10165
rect 12157 10164 12223 10165
rect 12157 10162 12204 10164
rect 11697 10160 12204 10162
rect 11697 10104 11702 10160
rect 11758 10104 12162 10160
rect 11697 10102 12204 10104
rect 11697 10099 11763 10102
rect 12157 10100 12204 10102
rect 12268 10100 12274 10164
rect 13816 10162 13876 10238
rect 15694 10236 15700 10300
rect 15764 10298 15770 10300
rect 17401 10298 17467 10301
rect 15764 10296 17467 10298
rect 15764 10240 17406 10296
rect 17462 10240 17467 10296
rect 15764 10238 17467 10240
rect 15764 10236 15770 10238
rect 17401 10235 17467 10238
rect 20846 10236 20852 10300
rect 20916 10298 20922 10300
rect 20989 10298 21055 10301
rect 20916 10296 21055 10298
rect 20916 10240 20994 10296
rect 21050 10240 21055 10296
rect 20916 10238 21055 10240
rect 20916 10236 20922 10238
rect 20989 10235 21055 10238
rect 15193 10162 15259 10165
rect 13816 10160 15259 10162
rect 13816 10104 15198 10160
rect 15254 10104 15259 10160
rect 13816 10102 15259 10104
rect 12157 10099 12223 10100
rect 15193 10099 15259 10102
rect 15561 10162 15627 10165
rect 16062 10162 16068 10164
rect 15561 10160 16068 10162
rect 15561 10104 15566 10160
rect 15622 10104 16068 10160
rect 15561 10102 16068 10104
rect 15561 10099 15627 10102
rect 16062 10100 16068 10102
rect 16132 10100 16138 10164
rect 19701 10162 19767 10165
rect 21081 10162 21147 10165
rect 19701 10160 21147 10162
rect 19701 10104 19706 10160
rect 19762 10104 21086 10160
rect 21142 10104 21147 10160
rect 19701 10102 21147 10104
rect 19701 10099 19767 10102
rect 21081 10099 21147 10102
rect 1669 10024 3434 10026
rect 1669 9968 1674 10024
rect 1730 9968 3434 10024
rect 1669 9966 3434 9968
rect 3969 10026 4035 10029
rect 5533 10026 5599 10029
rect 5901 10026 5967 10029
rect 6637 10026 6703 10029
rect 15377 10026 15443 10029
rect 17534 10026 17540 10028
rect 3969 10024 5599 10026
rect 3969 9968 3974 10024
rect 4030 9968 5538 10024
rect 5594 9968 5599 10024
rect 3969 9966 5599 9968
rect 1669 9963 1735 9966
rect 3969 9963 4035 9966
rect 5533 9963 5599 9966
rect 5766 10024 15443 10026
rect 5766 9968 5906 10024
rect 5962 9968 6642 10024
rect 6698 9968 15382 10024
rect 15438 9968 15443 10024
rect 5766 9966 15443 9968
rect 0 9890 800 9920
rect 2497 9890 2563 9893
rect 2998 9890 3004 9892
rect 0 9830 1640 9890
rect 0 9800 800 9830
rect 1580 9757 1640 9830
rect 2497 9888 3004 9890
rect 2497 9832 2502 9888
rect 2558 9832 3004 9888
rect 2497 9830 3004 9832
rect 2497 9827 2563 9830
rect 2998 9828 3004 9830
rect 3068 9828 3074 9892
rect 4153 9890 4219 9893
rect 4286 9890 4292 9892
rect 4153 9888 4292 9890
rect 4153 9832 4158 9888
rect 4214 9832 4292 9888
rect 4153 9830 4292 9832
rect 4153 9827 4219 9830
rect 4286 9828 4292 9830
rect 4356 9828 4362 9892
rect 5165 9890 5231 9893
rect 5766 9890 5826 9966
rect 5901 9963 5967 9966
rect 6637 9963 6703 9966
rect 15377 9963 15443 9966
rect 15518 9966 17540 10026
rect 5165 9888 5826 9890
rect 5165 9832 5170 9888
rect 5226 9832 5826 9888
rect 5165 9830 5826 9832
rect 7281 9890 7347 9893
rect 9489 9890 9555 9893
rect 11053 9890 11119 9893
rect 7281 9888 11119 9890
rect 7281 9832 7286 9888
rect 7342 9832 9494 9888
rect 9550 9832 11058 9888
rect 11114 9832 11119 9888
rect 7281 9830 11119 9832
rect 5165 9827 5231 9830
rect 7281 9827 7347 9830
rect 9489 9827 9555 9830
rect 11053 9827 11119 9830
rect 12157 9890 12223 9893
rect 12382 9890 12388 9892
rect 12157 9888 12388 9890
rect 12157 9832 12162 9888
rect 12218 9832 12388 9888
rect 12157 9830 12388 9832
rect 12157 9827 12223 9830
rect 12382 9828 12388 9830
rect 12452 9890 12458 9892
rect 15518 9890 15578 9966
rect 17534 9964 17540 9966
rect 17604 10026 17610 10028
rect 18965 10026 19031 10029
rect 17604 10024 19031 10026
rect 17604 9968 18970 10024
rect 19026 9968 19031 10024
rect 17604 9966 19031 9968
rect 17604 9964 17610 9966
rect 18965 9963 19031 9966
rect 19425 10026 19491 10029
rect 19885 10026 19951 10029
rect 21081 10026 21147 10029
rect 19425 10024 21147 10026
rect 19425 9968 19430 10024
rect 19486 9968 19890 10024
rect 19946 9968 21086 10024
rect 21142 9968 21147 10024
rect 19425 9966 21147 9968
rect 19425 9963 19491 9966
rect 19885 9963 19951 9966
rect 21081 9963 21147 9966
rect 12452 9830 15578 9890
rect 12452 9828 12458 9830
rect 18822 9828 18828 9892
rect 18892 9890 18898 9892
rect 20110 9890 20116 9892
rect 18892 9830 20116 9890
rect 18892 9828 18898 9830
rect 20110 9828 20116 9830
rect 20180 9828 20186 9892
rect 21173 9890 21239 9893
rect 22200 9890 23000 9920
rect 21173 9888 23000 9890
rect 21173 9832 21178 9888
rect 21234 9832 23000 9888
rect 21173 9830 23000 9832
rect 21173 9827 21239 9830
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 22200 9800 23000 9830
rect 16538 9759 16858 9760
rect 1577 9754 1643 9757
rect 4102 9754 4108 9756
rect 1577 9752 4108 9754
rect 1577 9696 1582 9752
rect 1638 9696 4108 9752
rect 1577 9694 4108 9696
rect 1577 9691 1643 9694
rect 4102 9692 4108 9694
rect 4172 9692 4178 9756
rect 4470 9692 4476 9756
rect 4540 9754 4546 9756
rect 5206 9754 5212 9756
rect 4540 9694 5212 9754
rect 4540 9692 4546 9694
rect 5206 9692 5212 9694
rect 5276 9754 5282 9756
rect 5625 9754 5691 9757
rect 5758 9754 5764 9756
rect 5276 9694 5458 9754
rect 5276 9692 5282 9694
rect 2037 9618 2103 9621
rect 5165 9618 5231 9621
rect 2037 9616 5231 9618
rect 2037 9560 2042 9616
rect 2098 9560 5170 9616
rect 5226 9560 5231 9616
rect 2037 9558 5231 9560
rect 5398 9618 5458 9694
rect 5625 9752 5764 9754
rect 5625 9696 5630 9752
rect 5686 9696 5764 9752
rect 5625 9694 5764 9696
rect 5625 9691 5691 9694
rect 5758 9692 5764 9694
rect 5828 9692 5834 9756
rect 7046 9692 7052 9756
rect 7116 9754 7122 9756
rect 7598 9754 7604 9756
rect 7116 9694 7604 9754
rect 7116 9692 7122 9694
rect 7598 9692 7604 9694
rect 7668 9692 7674 9756
rect 7966 9692 7972 9756
rect 8036 9754 8042 9756
rect 8385 9754 8451 9757
rect 9581 9756 9647 9757
rect 8036 9752 8451 9754
rect 8036 9696 8390 9752
rect 8446 9696 8451 9752
rect 8036 9694 8451 9696
rect 8036 9692 8042 9694
rect 8385 9691 8451 9694
rect 8518 9692 8524 9756
rect 8588 9754 8594 9756
rect 9438 9754 9444 9756
rect 8588 9694 9444 9754
rect 8588 9692 8594 9694
rect 9438 9692 9444 9694
rect 9508 9692 9514 9756
rect 9581 9752 9628 9756
rect 9692 9754 9698 9756
rect 12985 9754 13051 9757
rect 14917 9754 14983 9757
rect 9581 9696 9586 9752
rect 9581 9692 9628 9696
rect 9692 9694 9738 9754
rect 12985 9752 14983 9754
rect 12985 9696 12990 9752
rect 13046 9696 14922 9752
rect 14978 9696 14983 9752
rect 12985 9694 14983 9696
rect 9692 9692 9698 9694
rect 9581 9691 9647 9692
rect 12985 9691 13051 9694
rect 14917 9691 14983 9694
rect 15653 9754 15719 9757
rect 16062 9754 16068 9756
rect 15653 9752 16068 9754
rect 15653 9696 15658 9752
rect 15714 9696 16068 9752
rect 15653 9694 16068 9696
rect 15653 9691 15719 9694
rect 16062 9692 16068 9694
rect 16132 9692 16138 9756
rect 19793 9754 19859 9757
rect 20989 9754 21055 9757
rect 19793 9752 21055 9754
rect 19793 9696 19798 9752
rect 19854 9696 20994 9752
rect 21050 9696 21055 9752
rect 19793 9694 21055 9696
rect 19793 9691 19859 9694
rect 20989 9691 21055 9694
rect 6453 9618 6519 9621
rect 5398 9616 6519 9618
rect 5398 9560 6458 9616
rect 6514 9560 6519 9616
rect 5398 9558 6519 9560
rect 2037 9555 2103 9558
rect 5165 9555 5231 9558
rect 6453 9555 6519 9558
rect 6862 9556 6868 9620
rect 6932 9618 6938 9620
rect 9029 9618 9095 9621
rect 10542 9618 10548 9620
rect 6932 9558 8954 9618
rect 6932 9556 6938 9558
rect 0 9482 800 9512
rect 1025 9482 1091 9485
rect 0 9480 1091 9482
rect 0 9424 1030 9480
rect 1086 9424 1091 9480
rect 0 9422 1091 9424
rect 0 9392 800 9422
rect 1025 9419 1091 9422
rect 1945 9482 2011 9485
rect 2078 9482 2084 9484
rect 1945 9480 2084 9482
rect 1945 9424 1950 9480
rect 2006 9424 2084 9480
rect 1945 9422 2084 9424
rect 1945 9419 2011 9422
rect 2078 9420 2084 9422
rect 2148 9420 2154 9484
rect 4102 9420 4108 9484
rect 4172 9482 4178 9484
rect 4245 9482 4311 9485
rect 4172 9480 4311 9482
rect 4172 9424 4250 9480
rect 4306 9424 4311 9480
rect 4172 9422 4311 9424
rect 4172 9420 4178 9422
rect 4245 9419 4311 9422
rect 4889 9482 4955 9485
rect 5206 9482 5212 9484
rect 4889 9480 5212 9482
rect 4889 9424 4894 9480
rect 4950 9424 5212 9480
rect 4889 9422 5212 9424
rect 4889 9419 4955 9422
rect 5206 9420 5212 9422
rect 5276 9420 5282 9484
rect 7046 9420 7052 9484
rect 7116 9482 7122 9484
rect 8150 9482 8156 9484
rect 7116 9422 8156 9482
rect 7116 9420 7122 9422
rect 8150 9420 8156 9422
rect 8220 9482 8226 9484
rect 8661 9482 8727 9485
rect 8220 9480 8727 9482
rect 8220 9424 8666 9480
rect 8722 9424 8727 9480
rect 8220 9422 8727 9424
rect 8894 9482 8954 9558
rect 9029 9616 10548 9618
rect 9029 9560 9034 9616
rect 9090 9560 10548 9616
rect 9029 9558 10548 9560
rect 9029 9555 9095 9558
rect 10542 9556 10548 9558
rect 10612 9556 10618 9620
rect 11329 9618 11395 9621
rect 16205 9618 16271 9621
rect 11329 9616 16271 9618
rect 11329 9560 11334 9616
rect 11390 9560 16210 9616
rect 16266 9560 16271 9616
rect 11329 9558 16271 9560
rect 11329 9555 11395 9558
rect 16205 9555 16271 9558
rect 16941 9618 17007 9621
rect 17401 9618 17467 9621
rect 16941 9616 17467 9618
rect 16941 9560 16946 9616
rect 17002 9560 17406 9616
rect 17462 9560 17467 9616
rect 16941 9558 17467 9560
rect 16941 9555 17007 9558
rect 17401 9555 17467 9558
rect 19006 9556 19012 9620
rect 19076 9618 19082 9620
rect 19149 9618 19215 9621
rect 19076 9616 19215 9618
rect 19076 9560 19154 9616
rect 19210 9560 19215 9616
rect 19076 9558 19215 9560
rect 19076 9556 19082 9558
rect 19149 9555 19215 9558
rect 14641 9482 14707 9485
rect 8894 9480 14707 9482
rect 8894 9424 14646 9480
rect 14702 9424 14707 9480
rect 8894 9422 14707 9424
rect 8220 9420 8226 9422
rect 8661 9419 8727 9422
rect 14641 9419 14707 9422
rect 15469 9482 15535 9485
rect 19057 9482 19123 9485
rect 22200 9482 23000 9512
rect 15469 9480 18292 9482
rect 15469 9424 15474 9480
rect 15530 9424 18292 9480
rect 15469 9422 18292 9424
rect 15469 9419 15535 9422
rect 18232 9349 18292 9422
rect 19057 9480 23000 9482
rect 19057 9424 19062 9480
rect 19118 9424 23000 9480
rect 19057 9422 23000 9424
rect 19057 9419 19123 9422
rect 22200 9392 23000 9422
rect 2078 9284 2084 9348
rect 2148 9346 2154 9348
rect 3325 9346 3391 9349
rect 2148 9344 3391 9346
rect 2148 9288 3330 9344
rect 3386 9288 3391 9344
rect 2148 9286 3391 9288
rect 2148 9284 2154 9286
rect 3325 9283 3391 9286
rect 4705 9344 4771 9349
rect 4705 9288 4710 9344
rect 4766 9288 4771 9344
rect 4705 9283 4771 9288
rect 6545 9346 6611 9349
rect 8569 9346 8635 9349
rect 6545 9344 8635 9346
rect 6545 9288 6550 9344
rect 6606 9288 8574 9344
rect 8630 9288 8635 9344
rect 6545 9286 8635 9288
rect 6545 9283 6611 9286
rect 8569 9283 8635 9286
rect 11605 9346 11671 9349
rect 14641 9346 14707 9349
rect 15561 9346 15627 9349
rect 11605 9344 11898 9346
rect 11605 9288 11610 9344
rect 11666 9288 11898 9344
rect 11605 9286 11898 9288
rect 11605 9283 11671 9286
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 4153 9210 4219 9213
rect 4337 9210 4403 9213
rect 4153 9208 4403 9210
rect 4153 9152 4158 9208
rect 4214 9152 4342 9208
rect 4398 9152 4403 9208
rect 4153 9150 4403 9152
rect 4708 9210 4768 9283
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 7373 9210 7439 9213
rect 4708 9208 7439 9210
rect 4708 9152 7378 9208
rect 7434 9152 7439 9208
rect 4708 9150 7439 9152
rect 4153 9147 4219 9150
rect 4337 9147 4403 9150
rect 7373 9147 7439 9150
rect 8150 9148 8156 9212
rect 8220 9210 8226 9212
rect 8385 9210 8451 9213
rect 8220 9208 8451 9210
rect 8220 9152 8390 9208
rect 8446 9152 8451 9208
rect 8220 9150 8451 9152
rect 8220 9148 8226 9150
rect 8385 9147 8451 9150
rect 9489 9210 9555 9213
rect 11697 9210 11763 9213
rect 9489 9208 11763 9210
rect 9489 9152 9494 9208
rect 9550 9152 11702 9208
rect 11758 9152 11763 9208
rect 9489 9150 11763 9152
rect 11838 9210 11898 9286
rect 14641 9344 15627 9346
rect 14641 9288 14646 9344
rect 14702 9288 15566 9344
rect 15622 9288 15627 9344
rect 14641 9286 15627 9288
rect 14641 9283 14707 9286
rect 15561 9283 15627 9286
rect 18229 9344 18295 9349
rect 18229 9288 18234 9344
rect 18290 9288 18295 9344
rect 18229 9283 18295 9288
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 9215 19457 9216
rect 12382 9210 12388 9212
rect 11838 9150 12388 9210
rect 9489 9147 9555 9150
rect 11697 9147 11763 9150
rect 12382 9148 12388 9150
rect 12452 9148 12458 9212
rect 13077 9210 13143 9213
rect 13302 9210 13308 9212
rect 13077 9208 13308 9210
rect 13077 9152 13082 9208
rect 13138 9152 13308 9208
rect 13077 9150 13308 9152
rect 13077 9147 13143 9150
rect 13302 9148 13308 9150
rect 13372 9148 13378 9212
rect 14365 9210 14431 9213
rect 14365 9208 14474 9210
rect 14365 9152 14370 9208
rect 14426 9152 14474 9208
rect 14365 9147 14474 9152
rect 14590 9148 14596 9212
rect 14660 9210 14666 9212
rect 14825 9210 14891 9213
rect 14660 9208 14891 9210
rect 14660 9152 14830 9208
rect 14886 9152 14891 9208
rect 14660 9150 14891 9152
rect 14660 9148 14666 9150
rect 14825 9147 14891 9150
rect 15377 9210 15443 9213
rect 18454 9210 18460 9212
rect 15377 9208 18460 9210
rect 15377 9152 15382 9208
rect 15438 9152 18460 9208
rect 15377 9150 18460 9152
rect 15377 9147 15443 9150
rect 18454 9148 18460 9150
rect 18524 9148 18530 9212
rect 0 9074 800 9104
rect 1301 9074 1367 9077
rect 0 9072 1367 9074
rect 0 9016 1306 9072
rect 1362 9016 1367 9072
rect 0 9014 1367 9016
rect 0 8984 800 9014
rect 1301 9011 1367 9014
rect 1761 9074 1827 9077
rect 4061 9074 4127 9077
rect 5625 9074 5691 9077
rect 1761 9072 5691 9074
rect 1761 9016 1766 9072
rect 1822 9016 4066 9072
rect 4122 9016 5630 9072
rect 5686 9016 5691 9072
rect 1761 9014 5691 9016
rect 1761 9011 1827 9014
rect 4061 9011 4127 9014
rect 5625 9011 5691 9014
rect 5993 9074 6059 9077
rect 14273 9074 14339 9077
rect 5993 9072 14339 9074
rect 5993 9016 5998 9072
rect 6054 9016 14278 9072
rect 14334 9016 14339 9072
rect 5993 9014 14339 9016
rect 14414 9074 14474 9147
rect 19241 9074 19307 9077
rect 14414 9072 19307 9074
rect 14414 9016 19246 9072
rect 19302 9016 19307 9072
rect 14414 9014 19307 9016
rect 5993 9011 6059 9014
rect 14273 9011 14339 9014
rect 19241 9011 19307 9014
rect 19885 9074 19951 9077
rect 20529 9074 20595 9077
rect 22200 9074 23000 9104
rect 19885 9072 23000 9074
rect 19885 9016 19890 9072
rect 19946 9016 20534 9072
rect 20590 9016 23000 9072
rect 19885 9014 23000 9016
rect 19885 9011 19951 9014
rect 20529 9011 20595 9014
rect 22200 8984 23000 9014
rect 1853 8938 1919 8941
rect 1853 8936 6930 8938
rect 1853 8880 1858 8936
rect 1914 8880 6930 8936
rect 1853 8878 6930 8880
rect 1853 8875 1919 8878
rect 2865 8804 2931 8805
rect 2814 8740 2820 8804
rect 2884 8802 2931 8804
rect 3509 8802 3575 8805
rect 5165 8802 5231 8805
rect 2884 8800 2976 8802
rect 2926 8744 2976 8800
rect 2884 8742 2976 8744
rect 3509 8800 5231 8802
rect 3509 8744 3514 8800
rect 3570 8744 5170 8800
rect 5226 8744 5231 8800
rect 3509 8742 5231 8744
rect 6870 8802 6930 8878
rect 7782 8876 7788 8940
rect 7852 8938 7858 8940
rect 8109 8938 8175 8941
rect 8385 8938 8451 8941
rect 7852 8936 8451 8938
rect 7852 8880 8114 8936
rect 8170 8880 8390 8936
rect 8446 8880 8451 8936
rect 7852 8878 8451 8880
rect 7852 8876 7858 8878
rect 8109 8875 8175 8878
rect 8385 8875 8451 8878
rect 8569 8938 8635 8941
rect 11329 8938 11395 8941
rect 8569 8936 11395 8938
rect 8569 8880 8574 8936
rect 8630 8880 11334 8936
rect 11390 8880 11395 8936
rect 8569 8878 11395 8880
rect 8569 8875 8635 8878
rect 11329 8875 11395 8878
rect 11697 8938 11763 8941
rect 12433 8938 12499 8941
rect 18822 8938 18828 8940
rect 11697 8936 11898 8938
rect 11697 8880 11702 8936
rect 11758 8880 11898 8936
rect 11697 8878 11898 8880
rect 11697 8875 11763 8878
rect 9397 8802 9463 8805
rect 10409 8802 10475 8805
rect 6870 8800 10475 8802
rect 6870 8744 9402 8800
rect 9458 8744 10414 8800
rect 10470 8744 10475 8800
rect 6870 8742 10475 8744
rect 11838 8802 11898 8878
rect 12433 8936 18828 8938
rect 12433 8880 12438 8936
rect 12494 8880 18828 8936
rect 12433 8878 18828 8880
rect 12433 8875 12499 8878
rect 18822 8876 18828 8878
rect 18892 8876 18898 8940
rect 13445 8802 13511 8805
rect 15142 8802 15148 8804
rect 11838 8800 15148 8802
rect 11838 8744 13450 8800
rect 13506 8744 15148 8800
rect 11838 8742 15148 8744
rect 2884 8740 2931 8742
rect 2865 8739 2931 8740
rect 3509 8739 3575 8742
rect 5165 8739 5231 8742
rect 9397 8739 9463 8742
rect 10409 8739 10475 8742
rect 13445 8739 13511 8742
rect 15142 8740 15148 8742
rect 15212 8740 15218 8804
rect 6142 8736 6462 8737
rect 0 8666 800 8696
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 1485 8666 1551 8669
rect 3969 8666 4035 8669
rect 0 8664 4035 8666
rect 0 8608 1490 8664
rect 1546 8608 3974 8664
rect 4030 8608 4035 8664
rect 0 8606 4035 8608
rect 0 8576 800 8606
rect 1485 8603 1551 8606
rect 3969 8603 4035 8606
rect 6729 8666 6795 8669
rect 7005 8666 7071 8669
rect 6729 8664 7071 8666
rect 6729 8608 6734 8664
rect 6790 8608 7010 8664
rect 7066 8608 7071 8664
rect 6729 8606 7071 8608
rect 6729 8603 6795 8606
rect 7005 8603 7071 8606
rect 7465 8666 7531 8669
rect 9254 8666 9260 8668
rect 7465 8664 9260 8666
rect 7465 8608 7470 8664
rect 7526 8608 9260 8664
rect 7465 8606 9260 8608
rect 7465 8603 7531 8606
rect 9254 8604 9260 8606
rect 9324 8604 9330 8668
rect 9438 8604 9444 8668
rect 9508 8666 9514 8668
rect 9949 8666 10015 8669
rect 10869 8668 10935 8669
rect 10869 8666 10916 8668
rect 9508 8664 10015 8666
rect 9508 8608 9954 8664
rect 10010 8608 10015 8664
rect 9508 8606 10015 8608
rect 10824 8664 10916 8666
rect 10824 8608 10874 8664
rect 10824 8606 10916 8608
rect 9508 8604 9514 8606
rect 9949 8603 10015 8606
rect 10869 8604 10916 8606
rect 10980 8604 10986 8668
rect 12382 8604 12388 8668
rect 12452 8666 12458 8668
rect 12525 8666 12591 8669
rect 12452 8664 12591 8666
rect 12452 8608 12530 8664
rect 12586 8608 12591 8664
rect 12452 8606 12591 8608
rect 12452 8604 12458 8606
rect 10869 8603 10935 8604
rect 5260 8533 5458 8564
rect 1577 8530 1643 8533
rect 3877 8530 3943 8533
rect 5257 8532 5458 8533
rect 4838 8530 4844 8532
rect 1577 8528 4844 8530
rect 1577 8472 1582 8528
rect 1638 8472 3882 8528
rect 3938 8472 4844 8528
rect 1577 8470 4844 8472
rect 1577 8467 1643 8470
rect 3877 8467 3943 8470
rect 4838 8468 4844 8470
rect 4908 8468 4914 8532
rect 5206 8530 5212 8532
rect 5130 8470 5212 8530
rect 5276 8530 5458 8532
rect 10317 8532 10383 8533
rect 10317 8530 10364 8532
rect 5276 8528 10364 8530
rect 5318 8504 10322 8528
rect 5318 8472 5323 8504
rect 5206 8468 5212 8470
rect 5276 8468 5323 8472
rect 5398 8472 10322 8504
rect 5398 8470 10364 8472
rect 5257 8467 5323 8468
rect 10317 8468 10364 8470
rect 10428 8468 10434 8532
rect 10542 8468 10548 8532
rect 10612 8530 10618 8532
rect 10685 8530 10751 8533
rect 12390 8530 12450 8604
rect 12525 8603 12591 8606
rect 12893 8668 12959 8669
rect 12893 8664 12940 8668
rect 13004 8666 13010 8668
rect 14181 8666 14247 8669
rect 15377 8666 15443 8669
rect 12893 8608 12898 8664
rect 12893 8604 12940 8608
rect 13004 8606 13050 8666
rect 14181 8664 15443 8666
rect 14181 8608 14186 8664
rect 14242 8608 15382 8664
rect 15438 8608 15443 8664
rect 14181 8606 15443 8608
rect 13004 8604 13010 8606
rect 12893 8603 12959 8604
rect 14181 8603 14247 8606
rect 15377 8603 15443 8606
rect 19006 8604 19012 8668
rect 19076 8666 19082 8668
rect 19609 8666 19675 8669
rect 19076 8664 19675 8666
rect 19076 8608 19614 8664
rect 19670 8608 19675 8664
rect 19076 8606 19675 8608
rect 19076 8604 19082 8606
rect 19609 8603 19675 8606
rect 20713 8666 20779 8669
rect 21265 8666 21331 8669
rect 22200 8666 23000 8696
rect 20713 8664 23000 8666
rect 20713 8608 20718 8664
rect 20774 8608 21270 8664
rect 21326 8608 23000 8664
rect 20713 8606 23000 8608
rect 20713 8603 20779 8606
rect 21265 8603 21331 8606
rect 22200 8576 23000 8606
rect 14641 8530 14707 8533
rect 10612 8528 12450 8530
rect 10612 8472 10690 8528
rect 10746 8472 12450 8528
rect 10612 8470 12450 8472
rect 14368 8528 14707 8530
rect 14368 8472 14646 8528
rect 14702 8472 14707 8528
rect 14368 8470 14707 8472
rect 10612 8468 10618 8470
rect 10317 8467 10383 8468
rect 10685 8467 10751 8470
rect 2497 8394 2563 8397
rect 4654 8394 4660 8396
rect 2497 8392 4660 8394
rect 2497 8336 2502 8392
rect 2558 8336 4660 8392
rect 2497 8334 4660 8336
rect 2497 8331 2563 8334
rect 4654 8332 4660 8334
rect 4724 8332 4730 8396
rect 5206 8332 5212 8396
rect 5276 8394 5282 8396
rect 7414 8394 7420 8396
rect 5276 8334 7420 8394
rect 5276 8332 5282 8334
rect 7414 8332 7420 8334
rect 7484 8332 7490 8396
rect 8109 8394 8175 8397
rect 9581 8394 9647 8397
rect 14368 8394 14428 8470
rect 14641 8467 14707 8470
rect 16246 8468 16252 8532
rect 16316 8530 16322 8532
rect 18505 8530 18571 8533
rect 16316 8528 18571 8530
rect 16316 8472 18510 8528
rect 18566 8472 18571 8528
rect 16316 8470 18571 8472
rect 16316 8468 16322 8470
rect 18505 8467 18571 8470
rect 14549 8396 14615 8397
rect 14549 8394 14596 8396
rect 8109 8392 9184 8394
rect 8109 8336 8114 8392
rect 8170 8336 9184 8392
rect 8109 8334 9184 8336
rect 8109 8331 8175 8334
rect 0 8258 800 8288
rect 974 8258 980 8260
rect 0 8198 980 8258
rect 0 8168 800 8198
rect 974 8196 980 8198
rect 1044 8196 1050 8260
rect 1301 8258 1367 8261
rect 3049 8258 3115 8261
rect 1301 8256 3115 8258
rect 1301 8200 1306 8256
rect 1362 8200 3054 8256
rect 3110 8200 3115 8256
rect 1301 8198 3115 8200
rect 1301 8195 1367 8198
rect 3049 8195 3115 8198
rect 4061 8258 4127 8261
rect 6085 8258 6151 8261
rect 7373 8258 7439 8261
rect 4061 8256 7439 8258
rect 4061 8200 4066 8256
rect 4122 8200 6090 8256
rect 6146 8200 7378 8256
rect 7434 8200 7439 8256
rect 4061 8198 7439 8200
rect 4061 8195 4127 8198
rect 6085 8195 6151 8198
rect 7373 8195 7439 8198
rect 7649 8256 7715 8261
rect 7649 8200 7654 8256
rect 7710 8200 7715 8256
rect 7649 8195 7715 8200
rect 7966 8196 7972 8260
rect 8036 8258 8042 8260
rect 8036 8198 8264 8258
rect 8036 8196 8042 8198
rect 3543 8192 3863 8193
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 4061 8122 4127 8125
rect 7652 8122 7712 8195
rect 7966 8122 7972 8124
rect 4061 8120 7972 8122
rect 4061 8064 4066 8120
rect 4122 8064 7972 8120
rect 4061 8062 7972 8064
rect 4061 8059 4127 8062
rect 7966 8060 7972 8062
rect 8036 8060 8042 8124
rect 8204 8122 8264 8198
rect 8334 8196 8340 8260
rect 8404 8258 8410 8260
rect 8569 8258 8635 8261
rect 8404 8256 8635 8258
rect 8404 8200 8574 8256
rect 8630 8200 8635 8256
rect 8404 8198 8635 8200
rect 9124 8258 9184 8334
rect 9581 8392 14428 8394
rect 9581 8336 9586 8392
rect 9642 8336 14428 8392
rect 9581 8334 14428 8336
rect 14504 8392 14596 8394
rect 14504 8336 14554 8392
rect 14504 8334 14596 8336
rect 9581 8331 9647 8334
rect 14549 8332 14596 8334
rect 14660 8332 14666 8396
rect 16113 8394 16179 8397
rect 16941 8394 17007 8397
rect 17953 8394 18019 8397
rect 16113 8392 18019 8394
rect 16113 8336 16118 8392
rect 16174 8336 16946 8392
rect 17002 8336 17958 8392
rect 18014 8336 18019 8392
rect 16113 8334 18019 8336
rect 14549 8331 14615 8332
rect 16113 8331 16179 8334
rect 16941 8331 17007 8334
rect 17953 8331 18019 8334
rect 19014 8334 19626 8394
rect 15193 8258 15259 8261
rect 19014 8258 19074 8334
rect 9124 8198 13554 8258
rect 8404 8196 8410 8198
rect 8569 8195 8635 8198
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 8334 8122 8340 8124
rect 8204 8062 8340 8122
rect 8334 8060 8340 8062
rect 8404 8060 8410 8124
rect 12433 8122 12499 8125
rect 13118 8122 13124 8124
rect 9124 8120 12499 8122
rect 9124 8064 12438 8120
rect 12494 8064 12499 8120
rect 9124 8062 12499 8064
rect 2405 7986 2471 7989
rect 3509 7986 3575 7989
rect 3877 7986 3943 7989
rect 5993 7986 6059 7989
rect 2405 7984 3250 7986
rect 2405 7928 2410 7984
rect 2466 7928 3250 7984
rect 2405 7926 3250 7928
rect 2405 7923 2471 7926
rect 0 7850 800 7880
rect 1025 7850 1091 7853
rect 2681 7852 2747 7853
rect 0 7848 1091 7850
rect 0 7792 1030 7848
rect 1086 7792 1091 7848
rect 0 7790 1091 7792
rect 0 7760 800 7790
rect 1025 7787 1091 7790
rect 2630 7788 2636 7852
rect 2700 7850 2747 7852
rect 3190 7850 3250 7926
rect 3509 7984 6059 7986
rect 3509 7928 3514 7984
rect 3570 7928 3882 7984
rect 3938 7928 5998 7984
rect 6054 7928 6059 7984
rect 3509 7926 6059 7928
rect 3509 7923 3575 7926
rect 3877 7923 3943 7926
rect 5993 7923 6059 7926
rect 6453 7986 6519 7989
rect 8109 7986 8175 7989
rect 6453 7984 8175 7986
rect 6453 7928 6458 7984
rect 6514 7928 8114 7984
rect 8170 7928 8175 7984
rect 6453 7926 8175 7928
rect 6453 7923 6519 7926
rect 8109 7923 8175 7926
rect 4705 7850 4771 7853
rect 9124 7850 9184 8062
rect 12433 8059 12499 8062
rect 12804 8062 13124 8122
rect 12804 7989 12864 8062
rect 13118 8060 13124 8062
rect 13188 8060 13194 8124
rect 9305 7986 9371 7989
rect 10317 7986 10383 7989
rect 11830 7986 11836 7988
rect 9305 7984 10383 7986
rect 9305 7928 9310 7984
rect 9366 7928 10322 7984
rect 10378 7928 10383 7984
rect 9305 7926 10383 7928
rect 9305 7923 9371 7926
rect 10317 7923 10383 7926
rect 11056 7926 11836 7986
rect 2700 7848 2792 7850
rect 2742 7792 2792 7848
rect 2700 7790 2792 7792
rect 3190 7848 4771 7850
rect 3190 7792 4710 7848
rect 4766 7792 4771 7848
rect 3190 7790 4771 7792
rect 2700 7788 2747 7790
rect 2681 7787 2747 7788
rect 4705 7787 4771 7790
rect 4846 7790 9184 7850
rect 1025 7716 1091 7717
rect 974 7652 980 7716
rect 1044 7714 1091 7716
rect 2221 7714 2287 7717
rect 3785 7714 3851 7717
rect 4846 7714 4906 7790
rect 9254 7788 9260 7852
rect 9324 7850 9330 7852
rect 10542 7850 10548 7852
rect 9324 7790 10548 7850
rect 9324 7788 9330 7790
rect 10542 7788 10548 7790
rect 10612 7788 10618 7852
rect 9673 7714 9739 7717
rect 1044 7712 1136 7714
rect 1086 7656 1136 7712
rect 1044 7654 1136 7656
rect 2221 7712 2882 7714
rect 2221 7656 2226 7712
rect 2282 7656 2882 7712
rect 2221 7654 2882 7656
rect 1044 7652 1091 7654
rect 1025 7651 1091 7652
rect 2221 7651 2287 7654
rect 2589 7580 2655 7581
rect 2589 7576 2636 7580
rect 2700 7578 2706 7580
rect 2822 7578 2882 7654
rect 3785 7712 4906 7714
rect 3785 7656 3790 7712
rect 3846 7656 4906 7712
rect 3785 7654 4906 7656
rect 6548 7712 9739 7714
rect 6548 7656 9678 7712
rect 9734 7656 9739 7712
rect 6548 7654 9739 7656
rect 3785 7651 3851 7654
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 5349 7578 5415 7581
rect 2589 7520 2594 7576
rect 2589 7516 2636 7520
rect 2700 7518 2746 7578
rect 2822 7576 5415 7578
rect 2822 7520 5354 7576
rect 5410 7520 5415 7576
rect 2822 7518 5415 7520
rect 2700 7516 2706 7518
rect 2589 7515 2655 7516
rect 5349 7515 5415 7518
rect 5625 7578 5691 7581
rect 5758 7578 5764 7580
rect 5625 7576 5764 7578
rect 5625 7520 5630 7576
rect 5686 7520 5764 7576
rect 5625 7518 5764 7520
rect 5625 7515 5691 7518
rect 5758 7516 5764 7518
rect 5828 7516 5834 7580
rect 0 7442 800 7472
rect 1485 7444 1551 7445
rect 1485 7442 1532 7444
rect 0 7440 1532 7442
rect 0 7384 1490 7440
rect 0 7382 1532 7384
rect 0 7352 800 7382
rect 1485 7380 1532 7382
rect 1596 7380 1602 7444
rect 3601 7442 3667 7445
rect 6548 7442 6608 7654
rect 9673 7651 9739 7654
rect 10174 7652 10180 7716
rect 10244 7714 10250 7716
rect 10317 7714 10383 7717
rect 10244 7712 10383 7714
rect 10244 7656 10322 7712
rect 10378 7656 10383 7712
rect 10244 7654 10383 7656
rect 10244 7652 10250 7654
rect 10317 7651 10383 7654
rect 10726 7652 10732 7716
rect 10796 7714 10802 7716
rect 11056 7714 11116 7926
rect 11830 7924 11836 7926
rect 11900 7924 11906 7988
rect 12801 7984 12867 7989
rect 12801 7928 12806 7984
rect 12862 7928 12867 7984
rect 12801 7923 12867 7928
rect 13077 7986 13143 7989
rect 13494 7988 13554 8198
rect 15193 8256 19074 8258
rect 15193 8200 15198 8256
rect 15254 8200 19074 8256
rect 15193 8198 19074 8200
rect 15193 8195 15259 8198
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 16982 8122 16988 8124
rect 15150 8062 16988 8122
rect 13077 7984 13186 7986
rect 13077 7928 13082 7984
rect 13138 7928 13186 7984
rect 13077 7923 13186 7928
rect 13486 7924 13492 7988
rect 13556 7986 13562 7988
rect 15150 7986 15210 8062
rect 16982 8060 16988 8062
rect 17052 8060 17058 8124
rect 18454 8060 18460 8124
rect 18524 8122 18530 8124
rect 18965 8122 19031 8125
rect 18524 8120 19031 8122
rect 18524 8064 18970 8120
rect 19026 8064 19031 8120
rect 18524 8062 19031 8064
rect 19566 8122 19626 8334
rect 20713 8258 20779 8261
rect 21633 8258 21699 8261
rect 22200 8258 23000 8288
rect 20713 8256 23000 8258
rect 20713 8200 20718 8256
rect 20774 8200 21638 8256
rect 21694 8200 23000 8256
rect 20713 8198 23000 8200
rect 20713 8195 20779 8198
rect 21633 8195 21699 8198
rect 22200 8168 23000 8198
rect 21357 8122 21423 8125
rect 19566 8120 21423 8122
rect 19566 8064 21362 8120
rect 21418 8064 21423 8120
rect 19566 8062 21423 8064
rect 18524 8060 18530 8062
rect 18965 8059 19031 8062
rect 21357 8059 21423 8062
rect 13556 7926 15210 7986
rect 15837 7986 15903 7989
rect 18270 7986 18276 7988
rect 15837 7984 18276 7986
rect 15837 7928 15842 7984
rect 15898 7928 18276 7984
rect 15837 7926 18276 7928
rect 13556 7924 13562 7926
rect 15837 7923 15903 7926
rect 18270 7924 18276 7926
rect 18340 7986 18346 7988
rect 21214 7986 21220 7988
rect 18340 7926 21220 7986
rect 18340 7924 18346 7926
rect 21214 7924 21220 7926
rect 21284 7924 21290 7988
rect 11329 7850 11395 7853
rect 13126 7852 13186 7923
rect 11329 7848 13048 7850
rect 11329 7792 11334 7848
rect 11390 7792 13048 7848
rect 11329 7790 13048 7792
rect 11329 7787 11395 7790
rect 10796 7654 11116 7714
rect 12988 7714 13048 7790
rect 13118 7788 13124 7852
rect 13188 7850 13194 7852
rect 13629 7850 13695 7853
rect 16982 7850 16988 7852
rect 13188 7848 13695 7850
rect 13188 7792 13634 7848
rect 13690 7792 13695 7848
rect 13188 7790 13695 7792
rect 13188 7788 13194 7790
rect 13629 7787 13695 7790
rect 13816 7790 16988 7850
rect 13816 7714 13876 7790
rect 16982 7788 16988 7790
rect 17052 7788 17058 7852
rect 18229 7850 18295 7853
rect 20713 7850 20779 7853
rect 18229 7848 20779 7850
rect 18229 7792 18234 7848
rect 18290 7792 20718 7848
rect 20774 7792 20779 7848
rect 18229 7790 20779 7792
rect 18229 7787 18295 7790
rect 20713 7787 20779 7790
rect 21817 7850 21883 7853
rect 22200 7850 23000 7880
rect 21817 7848 23000 7850
rect 21817 7792 21822 7848
rect 21878 7792 23000 7848
rect 21817 7790 23000 7792
rect 21817 7787 21883 7790
rect 22200 7760 23000 7790
rect 14825 7716 14891 7717
rect 14774 7714 14780 7716
rect 12988 7654 13876 7714
rect 14734 7654 14780 7714
rect 14844 7712 14891 7716
rect 14886 7656 14891 7712
rect 10796 7652 10802 7654
rect 14774 7652 14780 7654
rect 14844 7652 14891 7656
rect 14825 7651 14891 7652
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 7465 7578 7531 7581
rect 10317 7578 10383 7581
rect 7465 7576 10383 7578
rect 7465 7520 7470 7576
rect 7526 7520 10322 7576
rect 10378 7520 10383 7576
rect 7465 7518 10383 7520
rect 7465 7515 7531 7518
rect 10317 7515 10383 7518
rect 12801 7578 12867 7581
rect 13302 7578 13308 7580
rect 12801 7576 13308 7578
rect 12801 7520 12806 7576
rect 12862 7520 13308 7576
rect 12801 7518 13308 7520
rect 12801 7515 12867 7518
rect 13302 7516 13308 7518
rect 13372 7516 13378 7580
rect 13445 7578 13511 7581
rect 15193 7578 15259 7581
rect 13445 7576 15259 7578
rect 13445 7520 13450 7576
rect 13506 7520 15198 7576
rect 15254 7520 15259 7576
rect 13445 7518 15259 7520
rect 13445 7515 13511 7518
rect 15193 7515 15259 7518
rect 17217 7578 17283 7581
rect 18822 7578 18828 7580
rect 17217 7576 18828 7578
rect 17217 7520 17222 7576
rect 17278 7520 18828 7576
rect 17217 7518 18828 7520
rect 17217 7515 17283 7518
rect 18822 7516 18828 7518
rect 18892 7578 18898 7580
rect 19241 7578 19307 7581
rect 18892 7576 19307 7578
rect 18892 7520 19246 7576
rect 19302 7520 19307 7576
rect 18892 7518 19307 7520
rect 18892 7516 18898 7518
rect 19241 7515 19307 7518
rect 3601 7440 6608 7442
rect 3601 7384 3606 7440
rect 3662 7384 6608 7440
rect 3601 7382 6608 7384
rect 6821 7442 6887 7445
rect 12014 7442 12020 7444
rect 6821 7440 12020 7442
rect 6821 7384 6826 7440
rect 6882 7384 12020 7440
rect 6821 7382 12020 7384
rect 1485 7379 1551 7380
rect 3601 7379 3667 7382
rect 6821 7379 6887 7382
rect 12014 7380 12020 7382
rect 12084 7442 12090 7444
rect 17125 7442 17191 7445
rect 12084 7440 17191 7442
rect 12084 7384 17130 7440
rect 17186 7384 17191 7440
rect 12084 7382 17191 7384
rect 12084 7380 12090 7382
rect 17125 7379 17191 7382
rect 18873 7442 18939 7445
rect 22200 7442 23000 7472
rect 18873 7440 23000 7442
rect 18873 7384 18878 7440
rect 18934 7384 23000 7440
rect 18873 7382 23000 7384
rect 18873 7379 18939 7382
rect 22200 7352 23000 7382
rect 1669 7306 1735 7309
rect 10041 7306 10107 7309
rect 1669 7304 10107 7306
rect 1669 7248 1674 7304
rect 1730 7248 10046 7304
rect 10102 7248 10107 7304
rect 1669 7246 10107 7248
rect 1669 7243 1735 7246
rect 10041 7243 10107 7246
rect 10317 7306 10383 7309
rect 18781 7306 18847 7309
rect 10317 7304 18847 7306
rect 10317 7248 10322 7304
rect 10378 7248 18786 7304
rect 18842 7248 18847 7304
rect 10317 7246 18847 7248
rect 10317 7243 10383 7246
rect 18781 7243 18847 7246
rect 5758 7108 5764 7172
rect 5828 7170 5834 7172
rect 6545 7170 6611 7173
rect 13721 7170 13787 7173
rect 5828 7168 6611 7170
rect 5828 7112 6550 7168
rect 6606 7112 6611 7168
rect 5828 7110 6611 7112
rect 5828 7108 5834 7110
rect 6545 7107 6611 7110
rect 10964 7168 13787 7170
rect 10964 7112 13726 7168
rect 13782 7112 13787 7168
rect 10964 7110 13787 7112
rect 3543 7104 3863 7105
rect 0 7034 800 7064
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 1301 7034 1367 7037
rect 0 7032 1367 7034
rect 0 6976 1306 7032
rect 1362 6976 1367 7032
rect 0 6974 1367 6976
rect 0 6944 800 6974
rect 1301 6971 1367 6974
rect 4838 6972 4844 7036
rect 4908 7034 4914 7036
rect 6453 7034 6519 7037
rect 4908 7032 6519 7034
rect 4908 6976 6458 7032
rect 6514 6976 6519 7032
rect 4908 6974 6519 6976
rect 4908 6972 4914 6974
rect 6453 6971 6519 6974
rect 6729 7034 6795 7037
rect 9305 7036 9371 7037
rect 9857 7036 9923 7037
rect 7414 7034 7420 7036
rect 6729 7032 7420 7034
rect 6729 6976 6734 7032
rect 6790 6976 7420 7032
rect 6729 6974 7420 6976
rect 6729 6971 6795 6974
rect 7414 6972 7420 6974
rect 7484 6972 7490 7036
rect 7598 6972 7604 7036
rect 7668 7034 7674 7036
rect 8150 7034 8156 7036
rect 7668 6974 8156 7034
rect 7668 6972 7674 6974
rect 8150 6972 8156 6974
rect 8220 6972 8226 7036
rect 9254 7034 9260 7036
rect 9214 6974 9260 7034
rect 9324 7032 9371 7036
rect 9806 7034 9812 7036
rect 9366 6976 9371 7032
rect 9254 6972 9260 6974
rect 9324 6972 9371 6976
rect 9730 6974 9812 7034
rect 9876 7034 9923 7036
rect 10964 7034 11024 7110
rect 13721 7107 13787 7110
rect 15561 7170 15627 7173
rect 16062 7170 16068 7172
rect 15561 7168 16068 7170
rect 15561 7112 15566 7168
rect 15622 7112 16068 7168
rect 15561 7110 16068 7112
rect 15561 7107 15627 7110
rect 16062 7108 16068 7110
rect 16132 7170 16138 7172
rect 16665 7170 16731 7173
rect 16132 7168 16731 7170
rect 16132 7112 16670 7168
rect 16726 7112 16731 7168
rect 16132 7110 16731 7112
rect 16132 7108 16138 7110
rect 16665 7107 16731 7110
rect 17718 7108 17724 7172
rect 17788 7170 17794 7172
rect 18505 7170 18571 7173
rect 17788 7168 18571 7170
rect 17788 7112 18510 7168
rect 18566 7112 18571 7168
rect 17788 7110 18571 7112
rect 17788 7108 17794 7110
rect 18505 7107 18571 7110
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 9876 7032 11024 7034
rect 9918 6976 11024 7032
rect 9806 6972 9812 6974
rect 9876 6974 11024 6976
rect 9876 6972 9923 6974
rect 11094 6972 11100 7036
rect 11164 7034 11170 7036
rect 12065 7034 12131 7037
rect 11164 7032 12131 7034
rect 11164 6976 12070 7032
rect 12126 6976 12131 7032
rect 11164 6974 12131 6976
rect 11164 6972 11170 6974
rect 9305 6971 9371 6972
rect 9857 6971 9923 6972
rect 12065 6971 12131 6974
rect 12382 6972 12388 7036
rect 12452 7034 12458 7036
rect 15653 7034 15719 7037
rect 17401 7034 17467 7037
rect 12452 6974 12772 7034
rect 12452 6972 12458 6974
rect 12712 6932 12772 6974
rect 15653 7032 17467 7034
rect 15653 6976 15658 7032
rect 15714 6976 17406 7032
rect 17462 6976 17467 7032
rect 15653 6974 17467 6976
rect 15653 6971 15719 6974
rect 17401 6971 17467 6974
rect 22001 7034 22067 7037
rect 22200 7034 23000 7064
rect 22001 7032 23000 7034
rect 22001 6976 22006 7032
rect 22062 6976 23000 7032
rect 22001 6974 23000 6976
rect 22001 6971 22067 6974
rect 22200 6944 23000 6974
rect 12893 6932 12959 6935
rect 12712 6930 12959 6932
rect 1577 6898 1643 6901
rect 3509 6898 3575 6901
rect 1577 6896 3575 6898
rect 1577 6840 1582 6896
rect 1638 6840 3514 6896
rect 3570 6840 3575 6896
rect 1577 6838 3575 6840
rect 1577 6835 1643 6838
rect 3509 6835 3575 6838
rect 3693 6898 3759 6901
rect 4521 6898 4587 6901
rect 8937 6898 9003 6901
rect 3693 6896 9003 6898
rect 3693 6840 3698 6896
rect 3754 6840 4526 6896
rect 4582 6840 8942 6896
rect 8998 6840 9003 6896
rect 3693 6838 9003 6840
rect 3693 6835 3759 6838
rect 4521 6835 4587 6838
rect 8937 6835 9003 6838
rect 9305 6898 9371 6901
rect 9438 6898 9444 6900
rect 9305 6896 9444 6898
rect 9305 6840 9310 6896
rect 9366 6840 9444 6896
rect 9305 6838 9444 6840
rect 9305 6835 9371 6838
rect 9438 6836 9444 6838
rect 9508 6836 9514 6900
rect 9990 6836 9996 6900
rect 10060 6898 10066 6900
rect 10317 6898 10383 6901
rect 10060 6896 10383 6898
rect 10060 6840 10322 6896
rect 10378 6840 10383 6896
rect 10060 6838 10383 6840
rect 10060 6836 10066 6838
rect 10317 6835 10383 6838
rect 12065 6898 12131 6901
rect 12249 6898 12315 6901
rect 12065 6896 12315 6898
rect 12065 6840 12070 6896
rect 12126 6840 12254 6896
rect 12310 6840 12315 6896
rect 12712 6874 12898 6930
rect 12954 6874 12959 6930
rect 12712 6872 12959 6874
rect 12893 6869 12959 6872
rect 13077 6898 13143 6901
rect 17953 6898 18019 6901
rect 21081 6898 21147 6901
rect 13077 6896 18019 6898
rect 12065 6838 12315 6840
rect 12065 6835 12131 6838
rect 12249 6835 12315 6838
rect 13077 6840 13082 6896
rect 13138 6840 17958 6896
rect 18014 6840 18019 6896
rect 13077 6838 18019 6840
rect 13077 6835 13143 6838
rect 17953 6835 18019 6838
rect 18094 6896 21147 6898
rect 18094 6840 21086 6896
rect 21142 6840 21147 6896
rect 18094 6838 21147 6840
rect 289 6762 355 6765
rect 5165 6764 5231 6765
rect 4102 6762 4108 6764
rect 289 6760 4108 6762
rect 289 6704 294 6760
rect 350 6704 4108 6760
rect 289 6702 4108 6704
rect 289 6699 355 6702
rect 4102 6700 4108 6702
rect 4172 6700 4178 6764
rect 5165 6762 5212 6764
rect 5120 6760 5212 6762
rect 5120 6704 5170 6760
rect 5120 6702 5212 6704
rect 5165 6700 5212 6702
rect 5276 6700 5282 6764
rect 8017 6762 8083 6765
rect 5490 6760 8083 6762
rect 5490 6704 8022 6760
rect 8078 6704 8083 6760
rect 5490 6702 8083 6704
rect 5165 6699 5231 6700
rect 1393 6626 1459 6629
rect 5490 6626 5550 6702
rect 8017 6699 8083 6702
rect 8753 6762 8819 6765
rect 12433 6764 12499 6765
rect 12382 6762 12388 6764
rect 8753 6760 11898 6762
rect 8753 6704 8758 6760
rect 8814 6704 11898 6760
rect 8753 6702 11898 6704
rect 12342 6702 12388 6762
rect 12452 6760 12499 6764
rect 12494 6704 12499 6760
rect 8753 6699 8819 6702
rect 1393 6624 5550 6626
rect 1393 6568 1398 6624
rect 1454 6568 5550 6624
rect 1393 6566 5550 6568
rect 5717 6626 5783 6629
rect 6637 6626 6703 6629
rect 6913 6626 6979 6629
rect 5717 6624 6056 6626
rect 5717 6568 5722 6624
rect 5778 6568 6056 6624
rect 5717 6566 6056 6568
rect 1393 6563 1459 6566
rect 5717 6563 5783 6566
rect 0 6490 800 6520
rect 3785 6490 3851 6493
rect 0 6488 3851 6490
rect 0 6432 3790 6488
rect 3846 6432 3851 6488
rect 0 6430 3851 6432
rect 0 6400 800 6430
rect 3785 6427 3851 6430
rect 5574 6428 5580 6492
rect 5644 6490 5650 6492
rect 5809 6490 5875 6493
rect 5644 6488 5875 6490
rect 5644 6432 5814 6488
rect 5870 6432 5875 6488
rect 5644 6430 5875 6432
rect 5644 6428 5650 6430
rect 5809 6427 5875 6430
rect 5022 6156 5028 6220
rect 5092 6218 5098 6220
rect 5809 6218 5875 6221
rect 5092 6216 5875 6218
rect 5092 6160 5814 6216
rect 5870 6160 5875 6216
rect 5092 6158 5875 6160
rect 5996 6218 6056 6566
rect 6637 6624 6979 6626
rect 6637 6568 6642 6624
rect 6698 6568 6918 6624
rect 6974 6568 6979 6624
rect 6637 6566 6979 6568
rect 6637 6563 6703 6566
rect 6913 6563 6979 6566
rect 7046 6564 7052 6628
rect 7116 6626 7122 6628
rect 7465 6626 7531 6629
rect 7116 6624 7531 6626
rect 7116 6568 7470 6624
rect 7526 6568 7531 6624
rect 7116 6566 7531 6568
rect 7116 6564 7122 6566
rect 7465 6563 7531 6566
rect 9305 6626 9371 6629
rect 9622 6626 9628 6628
rect 9305 6624 9628 6626
rect 9305 6568 9310 6624
rect 9366 6568 9628 6624
rect 9305 6566 9628 6568
rect 9305 6563 9371 6566
rect 9622 6564 9628 6566
rect 9692 6564 9698 6628
rect 11838 6626 11898 6702
rect 12382 6700 12388 6702
rect 12452 6700 12499 6704
rect 15142 6700 15148 6764
rect 15212 6762 15218 6764
rect 15653 6762 15719 6765
rect 18094 6762 18154 6838
rect 21081 6835 21147 6838
rect 15212 6760 15719 6762
rect 15212 6704 15658 6760
rect 15714 6704 15719 6760
rect 15212 6702 15719 6704
rect 15212 6700 15218 6702
rect 12433 6699 12499 6700
rect 15653 6699 15719 6702
rect 16254 6702 18154 6762
rect 18505 6762 18571 6765
rect 18638 6762 18644 6764
rect 18505 6760 18644 6762
rect 18505 6704 18510 6760
rect 18566 6704 18644 6760
rect 18505 6702 18644 6704
rect 12065 6626 12131 6629
rect 11838 6624 12131 6626
rect 11838 6568 12070 6624
rect 12126 6568 12131 6624
rect 11838 6566 12131 6568
rect 12065 6563 12131 6566
rect 13261 6626 13327 6629
rect 15326 6626 15332 6628
rect 13261 6624 15332 6626
rect 13261 6568 13266 6624
rect 13322 6568 15332 6624
rect 13261 6566 15332 6568
rect 13261 6563 13327 6566
rect 15326 6564 15332 6566
rect 15396 6564 15402 6628
rect 15837 6626 15903 6629
rect 16113 6626 16179 6629
rect 15837 6624 16179 6626
rect 15837 6568 15842 6624
rect 15898 6568 16118 6624
rect 16174 6568 16179 6624
rect 15837 6566 16179 6568
rect 15837 6563 15903 6566
rect 16113 6563 16179 6566
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 6678 6428 6684 6492
rect 6748 6490 6754 6492
rect 9254 6490 9260 6492
rect 6748 6430 9260 6490
rect 6748 6428 6754 6430
rect 9254 6428 9260 6430
rect 9324 6428 9330 6492
rect 9581 6490 9647 6493
rect 9990 6490 9996 6492
rect 9581 6488 9996 6490
rect 9581 6432 9586 6488
rect 9642 6432 9996 6488
rect 9581 6430 9996 6432
rect 9581 6427 9647 6430
rect 9990 6428 9996 6430
rect 10060 6428 10066 6492
rect 11830 6428 11836 6492
rect 11900 6490 11906 6492
rect 16021 6490 16087 6493
rect 11900 6488 16087 6490
rect 11900 6432 16026 6488
rect 16082 6432 16087 6488
rect 11900 6430 16087 6432
rect 11900 6428 11906 6430
rect 16021 6427 16087 6430
rect 6269 6354 6335 6357
rect 11881 6354 11947 6357
rect 12709 6354 12775 6357
rect 16254 6354 16314 6702
rect 18505 6699 18571 6702
rect 18638 6700 18644 6702
rect 18708 6700 18714 6764
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 6495 16858 6496
rect 18830 6430 20546 6490
rect 6269 6352 16314 6354
rect 6269 6296 6274 6352
rect 6330 6296 11886 6352
rect 11942 6296 12714 6352
rect 12770 6296 16314 6352
rect 6269 6294 16314 6296
rect 16573 6354 16639 6357
rect 17769 6354 17835 6357
rect 16573 6352 17835 6354
rect 16573 6296 16578 6352
rect 16634 6296 17774 6352
rect 17830 6296 17835 6352
rect 16573 6294 17835 6296
rect 6269 6291 6335 6294
rect 11881 6291 11947 6294
rect 12709 6291 12775 6294
rect 16573 6291 16639 6294
rect 17769 6291 17835 6294
rect 6361 6218 6427 6221
rect 5996 6216 6427 6218
rect 5996 6160 6366 6216
rect 6422 6160 6427 6216
rect 5996 6158 6427 6160
rect 5092 6156 5098 6158
rect 5809 6155 5875 6158
rect 6361 6155 6427 6158
rect 6545 6218 6611 6221
rect 7281 6218 7347 6221
rect 6545 6216 7347 6218
rect 6545 6160 6550 6216
rect 6606 6160 7286 6216
rect 7342 6160 7347 6216
rect 6545 6158 7347 6160
rect 6545 6155 6611 6158
rect 7281 6155 7347 6158
rect 7465 6218 7531 6221
rect 7782 6218 7788 6220
rect 7465 6216 7788 6218
rect 7465 6160 7470 6216
rect 7526 6160 7788 6216
rect 7465 6158 7788 6160
rect 7465 6155 7531 6158
rect 7782 6156 7788 6158
rect 7852 6156 7858 6220
rect 8109 6218 8175 6221
rect 18830 6218 18890 6430
rect 18965 6354 19031 6357
rect 19558 6354 19564 6356
rect 18965 6352 19564 6354
rect 18965 6296 18970 6352
rect 19026 6296 19564 6352
rect 18965 6294 19564 6296
rect 18965 6291 19031 6294
rect 19558 6292 19564 6294
rect 19628 6292 19634 6356
rect 20486 6354 20546 6430
rect 20662 6428 20668 6492
rect 20732 6490 20738 6492
rect 20989 6490 21055 6493
rect 20732 6488 21055 6490
rect 20732 6432 20994 6488
rect 21050 6432 21055 6488
rect 20732 6430 21055 6432
rect 20732 6428 20738 6430
rect 20989 6427 21055 6430
rect 21449 6490 21515 6493
rect 22200 6490 23000 6520
rect 21449 6488 23000 6490
rect 21449 6432 21454 6488
rect 21510 6432 23000 6488
rect 21449 6430 23000 6432
rect 21449 6427 21515 6430
rect 22200 6400 23000 6430
rect 20621 6354 20687 6357
rect 21398 6354 21404 6356
rect 20486 6352 21404 6354
rect 20486 6296 20626 6352
rect 20682 6296 21404 6352
rect 20486 6294 21404 6296
rect 20621 6291 20687 6294
rect 21398 6292 21404 6294
rect 21468 6292 21474 6356
rect 8109 6216 18890 6218
rect 8109 6160 8114 6216
rect 8170 6160 18890 6216
rect 8109 6158 18890 6160
rect 19425 6218 19491 6221
rect 19558 6218 19564 6220
rect 19425 6216 19564 6218
rect 19425 6160 19430 6216
rect 19486 6160 19564 6216
rect 19425 6158 19564 6160
rect 8109 6155 8175 6158
rect 19425 6155 19491 6158
rect 19558 6156 19564 6158
rect 19628 6156 19634 6220
rect 0 6082 800 6112
rect 933 6082 999 6085
rect 8518 6082 8524 6084
rect 0 6080 999 6082
rect 0 6024 938 6080
rect 994 6024 999 6080
rect 0 6022 999 6024
rect 0 5992 800 6022
rect 933 6019 999 6022
rect 3926 6022 8524 6082
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 1301 5946 1367 5949
rect 1894 5946 1900 5948
rect 1301 5944 1900 5946
rect 1301 5888 1306 5944
rect 1362 5888 1900 5944
rect 1301 5886 1900 5888
rect 1301 5883 1367 5886
rect 1894 5884 1900 5886
rect 1964 5884 1970 5948
rect 3182 5748 3188 5812
rect 3252 5810 3258 5812
rect 3601 5810 3667 5813
rect 3252 5808 3667 5810
rect 3252 5752 3606 5808
rect 3662 5752 3667 5808
rect 3252 5750 3667 5752
rect 3252 5748 3258 5750
rect 3601 5747 3667 5750
rect 3785 5810 3851 5813
rect 3926 5810 3986 6022
rect 8518 6020 8524 6022
rect 8588 6020 8594 6084
rect 9622 6020 9628 6084
rect 9692 6082 9698 6084
rect 13445 6082 13511 6085
rect 15101 6084 15167 6085
rect 15101 6082 15148 6084
rect 9692 6080 13511 6082
rect 9692 6024 13450 6080
rect 13506 6024 13511 6080
rect 9692 6022 13511 6024
rect 15056 6080 15148 6082
rect 15056 6024 15106 6080
rect 15056 6022 15148 6024
rect 9692 6020 9698 6022
rect 13445 6019 13511 6022
rect 15101 6020 15148 6022
rect 15212 6020 15218 6084
rect 18086 6020 18092 6084
rect 18156 6082 18162 6084
rect 18597 6082 18663 6085
rect 18156 6080 18663 6082
rect 18156 6024 18602 6080
rect 18658 6024 18663 6080
rect 18156 6022 18663 6024
rect 18156 6020 18162 6022
rect 15101 6019 15167 6020
rect 18597 6019 18663 6022
rect 19517 6082 19583 6085
rect 19926 6082 19932 6084
rect 19517 6080 19932 6082
rect 19517 6024 19522 6080
rect 19578 6024 19932 6080
rect 19517 6022 19932 6024
rect 19517 6019 19583 6022
rect 19926 6020 19932 6022
rect 19996 6082 20002 6084
rect 22200 6082 23000 6112
rect 19996 6022 23000 6082
rect 19996 6020 20002 6022
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 22200 5992 23000 6022
rect 19137 5951 19457 5952
rect 7005 5946 7071 5949
rect 7281 5948 7347 5949
rect 8109 5948 8175 5949
rect 3785 5808 3986 5810
rect 3785 5752 3790 5808
rect 3846 5752 3986 5808
rect 3785 5750 3986 5752
rect 4110 5944 7071 5946
rect 4110 5888 7010 5944
rect 7066 5888 7071 5944
rect 4110 5886 7071 5888
rect 3785 5747 3851 5750
rect 0 5674 800 5704
rect 2446 5674 2452 5676
rect 0 5614 2452 5674
rect 0 5584 800 5614
rect 1534 5541 1594 5614
rect 2446 5612 2452 5614
rect 2516 5612 2522 5676
rect 3049 5674 3115 5677
rect 4110 5674 4170 5886
rect 7005 5883 7071 5886
rect 7230 5884 7236 5948
rect 7300 5946 7347 5948
rect 7782 5946 7788 5948
rect 7300 5944 7788 5946
rect 7342 5888 7788 5944
rect 7300 5886 7788 5888
rect 7300 5884 7347 5886
rect 7782 5884 7788 5886
rect 7852 5884 7858 5948
rect 8109 5944 8156 5948
rect 8220 5946 8226 5948
rect 8385 5946 8451 5949
rect 8518 5946 8524 5948
rect 8109 5888 8114 5944
rect 8109 5884 8156 5888
rect 8220 5886 8266 5946
rect 8385 5944 8524 5946
rect 8385 5888 8390 5944
rect 8446 5888 8524 5944
rect 8385 5886 8524 5888
rect 8220 5884 8226 5886
rect 7281 5883 7347 5884
rect 8109 5883 8175 5884
rect 8385 5883 8451 5886
rect 8518 5884 8524 5886
rect 8588 5884 8594 5948
rect 13169 5946 13235 5949
rect 9630 5944 13235 5946
rect 9630 5888 13174 5944
rect 13230 5888 13235 5944
rect 9630 5886 13235 5888
rect 5206 5748 5212 5812
rect 5276 5810 5282 5812
rect 7189 5810 7255 5813
rect 9630 5810 9690 5886
rect 13169 5883 13235 5886
rect 14917 5946 14983 5949
rect 18638 5946 18644 5948
rect 14917 5944 18644 5946
rect 14917 5888 14922 5944
rect 14978 5888 18644 5944
rect 14917 5886 18644 5888
rect 14917 5883 14983 5886
rect 18638 5884 18644 5886
rect 18708 5884 18714 5948
rect 5276 5808 7255 5810
rect 5276 5752 7194 5808
rect 7250 5752 7255 5808
rect 5276 5750 7255 5752
rect 5276 5748 5282 5750
rect 7189 5747 7255 5750
rect 7468 5750 9690 5810
rect 11329 5810 11395 5813
rect 15285 5810 15351 5813
rect 11329 5808 15351 5810
rect 11329 5752 11334 5808
rect 11390 5752 15290 5808
rect 15346 5752 15351 5808
rect 11329 5750 15351 5752
rect 3049 5672 4170 5674
rect 3049 5616 3054 5672
rect 3110 5616 4170 5672
rect 3049 5614 4170 5616
rect 3049 5611 3115 5614
rect 4654 5612 4660 5676
rect 4724 5674 4730 5676
rect 6729 5674 6795 5677
rect 7468 5674 7528 5750
rect 11329 5747 11395 5750
rect 15285 5747 15351 5750
rect 15653 5810 15719 5813
rect 18045 5810 18111 5813
rect 15653 5808 18111 5810
rect 15653 5752 15658 5808
rect 15714 5752 18050 5808
rect 18106 5752 18111 5808
rect 15653 5750 18111 5752
rect 15653 5747 15719 5750
rect 18045 5747 18111 5750
rect 18413 5810 18479 5813
rect 18413 5808 20362 5810
rect 18413 5752 18418 5808
rect 18474 5752 20362 5808
rect 18413 5750 20362 5752
rect 18413 5747 18479 5750
rect 4724 5614 6608 5674
rect 4724 5612 4730 5614
rect 1485 5536 1594 5541
rect 1485 5480 1490 5536
rect 1546 5480 1594 5536
rect 1485 5478 1594 5480
rect 1485 5475 1551 5478
rect 5758 5476 5764 5540
rect 5828 5538 5834 5540
rect 5901 5538 5967 5541
rect 5828 5536 5967 5538
rect 5828 5480 5906 5536
rect 5962 5480 5967 5536
rect 5828 5478 5967 5480
rect 6548 5538 6608 5614
rect 6729 5672 7528 5674
rect 6729 5616 6734 5672
rect 6790 5616 7528 5672
rect 6729 5614 7528 5616
rect 6729 5611 6795 5614
rect 7966 5612 7972 5676
rect 8036 5674 8042 5676
rect 8109 5674 8175 5677
rect 8036 5672 8175 5674
rect 8036 5616 8114 5672
rect 8170 5616 8175 5672
rect 8036 5614 8175 5616
rect 8036 5612 8042 5614
rect 8109 5611 8175 5614
rect 8334 5612 8340 5676
rect 8404 5674 8410 5676
rect 8845 5674 8911 5677
rect 9029 5674 9095 5677
rect 9438 5674 9444 5676
rect 8404 5672 8954 5674
rect 8404 5616 8850 5672
rect 8906 5616 8954 5672
rect 8404 5614 8954 5616
rect 8404 5612 8410 5614
rect 8845 5611 8954 5614
rect 9029 5672 9444 5674
rect 9029 5616 9034 5672
rect 9090 5616 9444 5672
rect 9029 5614 9444 5616
rect 9029 5611 9095 5614
rect 9438 5612 9444 5614
rect 9508 5612 9514 5676
rect 9857 5674 9923 5677
rect 9630 5672 9923 5674
rect 9630 5616 9862 5672
rect 9918 5616 9923 5672
rect 9630 5614 9923 5616
rect 8894 5538 8954 5611
rect 6548 5478 8954 5538
rect 5828 5476 5834 5478
rect 5901 5475 5967 5478
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 7097 5402 7163 5405
rect 9305 5402 9371 5405
rect 9630 5402 9690 5614
rect 9857 5611 9923 5614
rect 11789 5672 11855 5677
rect 11789 5616 11794 5672
rect 11850 5616 11855 5672
rect 11789 5611 11855 5616
rect 11973 5674 12039 5677
rect 12617 5676 12683 5677
rect 12566 5674 12572 5676
rect 11973 5672 12572 5674
rect 12636 5672 12683 5676
rect 11973 5616 11978 5672
rect 12034 5616 12572 5672
rect 12678 5616 12683 5672
rect 11973 5614 12572 5616
rect 11973 5611 12039 5614
rect 12566 5612 12572 5614
rect 12636 5612 12683 5616
rect 12617 5611 12683 5612
rect 13169 5674 13235 5677
rect 14917 5674 14983 5677
rect 13169 5672 14983 5674
rect 13169 5616 13174 5672
rect 13230 5616 14922 5672
rect 14978 5616 14983 5672
rect 13169 5614 14983 5616
rect 13169 5611 13235 5614
rect 14917 5611 14983 5614
rect 17861 5674 17927 5677
rect 19517 5674 19583 5677
rect 17861 5672 19583 5674
rect 17861 5616 17866 5672
rect 17922 5616 19522 5672
rect 19578 5616 19583 5672
rect 17861 5614 19583 5616
rect 20302 5674 20362 5750
rect 22200 5674 23000 5704
rect 20302 5614 23000 5674
rect 17861 5611 17927 5614
rect 19517 5611 19583 5614
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 11792 5405 11852 5611
rect 22200 5584 23000 5614
rect 14733 5538 14799 5541
rect 15142 5538 15148 5540
rect 14733 5536 15148 5538
rect 14733 5480 14738 5536
rect 14794 5480 15148 5536
rect 14733 5478 15148 5480
rect 14733 5475 14799 5478
rect 15142 5476 15148 5478
rect 15212 5476 15218 5540
rect 16982 5476 16988 5540
rect 17052 5538 17058 5540
rect 20989 5538 21055 5541
rect 17052 5536 21055 5538
rect 17052 5480 20994 5536
rect 21050 5480 21055 5536
rect 17052 5478 21055 5480
rect 17052 5476 17058 5478
rect 20989 5475 21055 5478
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 7097 5400 9690 5402
rect 7097 5344 7102 5400
rect 7158 5344 9310 5400
rect 9366 5344 9690 5400
rect 7097 5342 9690 5344
rect 11789 5400 11855 5405
rect 11789 5344 11794 5400
rect 11850 5344 11855 5400
rect 7097 5339 7163 5342
rect 9305 5339 9371 5342
rect 11789 5339 11855 5344
rect 13302 5340 13308 5404
rect 13372 5402 13378 5404
rect 15745 5402 15811 5405
rect 13372 5400 15811 5402
rect 13372 5344 15750 5400
rect 15806 5344 15811 5400
rect 13372 5342 15811 5344
rect 13372 5340 13378 5342
rect 15745 5339 15811 5342
rect 0 5266 800 5296
rect 3785 5266 3851 5269
rect 0 5264 3851 5266
rect 0 5208 3790 5264
rect 3846 5208 3851 5264
rect 0 5206 3851 5208
rect 0 5176 800 5206
rect 3785 5203 3851 5206
rect 5390 5204 5396 5268
rect 5460 5266 5466 5268
rect 5901 5266 5967 5269
rect 5460 5264 5967 5266
rect 5460 5208 5906 5264
rect 5962 5208 5967 5264
rect 5460 5206 5967 5208
rect 5460 5204 5466 5206
rect 5901 5203 5967 5206
rect 6729 5266 6795 5269
rect 10726 5266 10732 5268
rect 6729 5264 10732 5266
rect 6729 5208 6734 5264
rect 6790 5208 10732 5264
rect 6729 5206 10732 5208
rect 6729 5203 6795 5206
rect 10726 5204 10732 5206
rect 10796 5266 10802 5268
rect 10918 5266 11484 5300
rect 13077 5266 13143 5269
rect 10796 5264 13143 5266
rect 10796 5240 13082 5264
rect 10796 5206 10978 5240
rect 11424 5208 13082 5240
rect 13138 5208 13143 5264
rect 11424 5206 13143 5208
rect 10796 5204 10802 5206
rect 13077 5203 13143 5206
rect 18597 5266 18663 5269
rect 20345 5266 20411 5269
rect 22200 5266 23000 5296
rect 18597 5264 23000 5266
rect 18597 5208 18602 5264
rect 18658 5208 20350 5264
rect 20406 5208 23000 5264
rect 18597 5206 23000 5208
rect 18597 5203 18663 5206
rect 20345 5203 20411 5206
rect 22200 5176 23000 5206
rect 2865 5130 2931 5133
rect 4153 5130 4219 5133
rect 4429 5130 4495 5133
rect 2865 5128 3986 5130
rect 2865 5072 2870 5128
rect 2926 5072 3986 5128
rect 2865 5070 3986 5072
rect 2865 5067 2931 5070
rect 3926 4994 3986 5070
rect 4153 5128 4495 5130
rect 4153 5072 4158 5128
rect 4214 5072 4434 5128
rect 4490 5072 4495 5128
rect 4153 5070 4495 5072
rect 4153 5067 4219 5070
rect 4429 5067 4495 5070
rect 5533 5130 5599 5133
rect 12157 5130 12223 5133
rect 5533 5128 12223 5130
rect 5533 5072 5538 5128
rect 5594 5072 12162 5128
rect 12218 5072 12223 5128
rect 5533 5070 12223 5072
rect 5533 5067 5599 5070
rect 12157 5067 12223 5070
rect 12566 5068 12572 5132
rect 12636 5130 12642 5132
rect 12636 5070 15210 5130
rect 12636 5068 12642 5070
rect 7741 4994 7807 4997
rect 7925 4996 7991 4997
rect 7925 4994 7972 4996
rect 3926 4992 7807 4994
rect 3926 4936 7746 4992
rect 7802 4936 7807 4992
rect 3926 4934 7807 4936
rect 7880 4992 7972 4994
rect 7880 4936 7930 4992
rect 7880 4934 7972 4936
rect 7741 4931 7807 4934
rect 7925 4932 7972 4934
rect 8036 4932 8042 4996
rect 8385 4994 8451 4997
rect 8518 4994 8524 4996
rect 8385 4992 8524 4994
rect 8385 4936 8390 4992
rect 8446 4936 8524 4992
rect 8385 4934 8524 4936
rect 7925 4931 7991 4932
rect 8385 4931 8451 4934
rect 8518 4932 8524 4934
rect 8588 4932 8594 4996
rect 10133 4994 10199 4997
rect 12433 4994 12499 4997
rect 10133 4992 12499 4994
rect 10133 4936 10138 4992
rect 10194 4936 12438 4992
rect 12494 4936 12499 4992
rect 10133 4934 12499 4936
rect 10133 4931 10199 4934
rect 12433 4931 12499 4934
rect 3543 4928 3863 4929
rect 0 4858 800 4888
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 974 4858 980 4860
rect 0 4798 980 4858
rect 0 4768 800 4798
rect 974 4796 980 4798
rect 1044 4858 1050 4860
rect 2221 4858 2287 4861
rect 1044 4856 2287 4858
rect 1044 4800 2226 4856
rect 2282 4800 2287 4856
rect 1044 4798 2287 4800
rect 1044 4796 1050 4798
rect 2221 4795 2287 4798
rect 4061 4858 4127 4861
rect 8017 4858 8083 4861
rect 4061 4856 8083 4858
rect 4061 4800 4066 4856
rect 4122 4800 8022 4856
rect 8078 4800 8083 4856
rect 4061 4798 8083 4800
rect 4061 4795 4127 4798
rect 8017 4795 8083 4798
rect 8293 4860 8359 4861
rect 10409 4860 10475 4861
rect 8293 4856 8340 4860
rect 8404 4858 8410 4860
rect 8293 4800 8298 4856
rect 8293 4796 8340 4800
rect 8404 4798 8450 4858
rect 8404 4796 8410 4798
rect 10358 4796 10364 4860
rect 10428 4858 10475 4860
rect 10593 4858 10659 4861
rect 11605 4858 11671 4861
rect 12249 4858 12315 4861
rect 10428 4856 10520 4858
rect 10470 4800 10520 4856
rect 10428 4798 10520 4800
rect 10593 4856 11671 4858
rect 10593 4800 10598 4856
rect 10654 4800 11610 4856
rect 11666 4800 11671 4856
rect 10593 4798 11671 4800
rect 10428 4796 10475 4798
rect 8293 4795 8359 4796
rect 10409 4795 10475 4796
rect 10593 4795 10659 4798
rect 11605 4795 11671 4798
rect 11884 4856 12315 4858
rect 11884 4800 12254 4856
rect 12310 4800 12315 4856
rect 11884 4798 12315 4800
rect 7005 4722 7071 4725
rect 11884 4722 11944 4798
rect 12249 4795 12315 4798
rect 12893 4858 12959 4861
rect 15150 4858 15210 5070
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 17401 4858 17467 4861
rect 21909 4858 21975 4861
rect 22200 4858 23000 4888
rect 12893 4856 13738 4858
rect 12893 4800 12898 4856
rect 12954 4800 13738 4856
rect 12893 4798 13738 4800
rect 15150 4856 18890 4858
rect 15150 4800 17406 4856
rect 17462 4800 18890 4856
rect 15150 4798 18890 4800
rect 12893 4795 12959 4798
rect 4110 4720 11944 4722
rect 4110 4664 7010 4720
rect 7066 4664 11944 4720
rect 4110 4662 11944 4664
rect 1117 4586 1183 4589
rect 3877 4586 3943 4589
rect 1117 4584 3943 4586
rect 1117 4528 1122 4584
rect 1178 4528 3882 4584
rect 3938 4528 3943 4584
rect 1117 4526 3943 4528
rect 1117 4523 1183 4526
rect 3877 4523 3943 4526
rect 0 4450 800 4480
rect 1158 4450 1164 4452
rect 0 4390 1164 4450
rect 0 4360 800 4390
rect 1158 4388 1164 4390
rect 1228 4450 1234 4452
rect 3049 4450 3115 4453
rect 1228 4448 3115 4450
rect 1228 4392 3054 4448
rect 3110 4392 3115 4448
rect 1228 4390 3115 4392
rect 1228 4388 1234 4390
rect 3049 4387 3115 4390
rect 4110 4314 4170 4662
rect 7005 4659 7071 4662
rect 12014 4660 12020 4724
rect 12084 4722 12090 4724
rect 13302 4722 13308 4724
rect 12084 4662 13308 4722
rect 12084 4660 12090 4662
rect 13302 4660 13308 4662
rect 13372 4660 13378 4724
rect 13678 4722 13738 4798
rect 17401 4795 17467 4798
rect 13997 4722 14063 4725
rect 13678 4720 14063 4722
rect 13678 4664 14002 4720
rect 14058 4664 14063 4720
rect 13678 4662 14063 4664
rect 13997 4659 14063 4662
rect 14733 4722 14799 4725
rect 18321 4722 18387 4725
rect 18638 4722 18644 4724
rect 14733 4720 15210 4722
rect 14733 4664 14738 4720
rect 14794 4664 15210 4720
rect 14733 4662 15210 4664
rect 14733 4659 14799 4662
rect 4337 4588 4403 4589
rect 4286 4524 4292 4588
rect 4356 4586 4403 4588
rect 5625 4586 5691 4589
rect 6361 4586 6427 4589
rect 8845 4586 8911 4589
rect 4356 4584 4448 4586
rect 4398 4528 4448 4584
rect 4356 4526 4448 4528
rect 5260 4584 8911 4586
rect 5260 4528 5630 4584
rect 5686 4528 6366 4584
rect 6422 4528 8850 4584
rect 8906 4528 8911 4584
rect 5260 4526 8911 4528
rect 4356 4524 4403 4526
rect 4337 4523 4403 4524
rect 5260 4453 5320 4526
rect 5625 4523 5691 4526
rect 6361 4523 6427 4526
rect 8845 4523 8911 4526
rect 11329 4586 11395 4589
rect 12525 4588 12591 4589
rect 12525 4586 12572 4588
rect 11329 4584 11852 4586
rect 11329 4528 11334 4584
rect 11390 4528 11852 4584
rect 11329 4526 11852 4528
rect 12480 4584 12572 4586
rect 12480 4528 12530 4584
rect 12480 4526 12572 4528
rect 11329 4523 11395 4526
rect 4470 4388 4476 4452
rect 4540 4450 4546 4452
rect 4613 4450 4679 4453
rect 4540 4448 4679 4450
rect 4540 4392 4618 4448
rect 4674 4392 4679 4448
rect 4540 4390 4679 4392
rect 4540 4388 4546 4390
rect 4613 4387 4679 4390
rect 5257 4448 5323 4453
rect 5257 4392 5262 4448
rect 5318 4392 5323 4448
rect 5257 4387 5323 4392
rect 7649 4450 7715 4453
rect 11145 4450 11211 4453
rect 7649 4448 11211 4450
rect 7649 4392 7654 4448
rect 7710 4392 11150 4448
rect 11206 4392 11211 4448
rect 7649 4390 11211 4392
rect 7649 4387 7715 4390
rect 11145 4387 11211 4390
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 2730 4254 4170 4314
rect 4337 4314 4403 4317
rect 5390 4314 5396 4316
rect 4337 4312 5396 4314
rect 4337 4256 4342 4312
rect 4398 4256 5396 4312
rect 4337 4254 5396 4256
rect 1945 4178 2011 4181
rect 2730 4178 2790 4254
rect 4337 4251 4403 4254
rect 5390 4252 5396 4254
rect 5460 4252 5466 4316
rect 5717 4314 5783 4317
rect 5993 4314 6059 4317
rect 5717 4312 6059 4314
rect 5717 4256 5722 4312
rect 5778 4256 5998 4312
rect 6054 4256 6059 4312
rect 5717 4254 6059 4256
rect 5717 4251 5783 4254
rect 5993 4251 6059 4254
rect 6862 4252 6868 4316
rect 6932 4314 6938 4316
rect 7189 4314 7255 4317
rect 6932 4312 7255 4314
rect 6932 4256 7194 4312
rect 7250 4256 7255 4312
rect 6932 4254 7255 4256
rect 6932 4252 6938 4254
rect 7189 4251 7255 4254
rect 7373 4314 7439 4317
rect 7598 4314 7604 4316
rect 7373 4312 7604 4314
rect 7373 4256 7378 4312
rect 7434 4256 7604 4312
rect 7373 4254 7604 4256
rect 7373 4251 7439 4254
rect 7598 4252 7604 4254
rect 7668 4252 7674 4316
rect 7741 4314 7807 4317
rect 9489 4314 9555 4317
rect 11145 4314 11211 4317
rect 7741 4312 11211 4314
rect 7741 4256 7746 4312
rect 7802 4256 9494 4312
rect 9550 4256 11150 4312
rect 11206 4256 11211 4312
rect 7741 4254 11211 4256
rect 11792 4314 11852 4526
rect 12525 4524 12572 4526
rect 12636 4524 12642 4588
rect 12709 4586 12775 4589
rect 14958 4586 14964 4588
rect 12709 4584 14964 4586
rect 12709 4528 12714 4584
rect 12770 4528 14964 4584
rect 12709 4526 14964 4528
rect 12525 4523 12591 4524
rect 12709 4523 12775 4526
rect 14958 4524 14964 4526
rect 15028 4524 15034 4588
rect 15150 4586 15210 4662
rect 18321 4720 18644 4722
rect 18321 4664 18326 4720
rect 18382 4664 18644 4720
rect 18321 4662 18644 4664
rect 18321 4659 18387 4662
rect 18638 4660 18644 4662
rect 18708 4660 18714 4724
rect 18830 4722 18890 4798
rect 21909 4856 23000 4858
rect 21909 4800 21914 4856
rect 21970 4800 23000 4856
rect 21909 4798 23000 4800
rect 21909 4795 21975 4798
rect 22200 4768 23000 4798
rect 19333 4722 19399 4725
rect 18830 4720 19399 4722
rect 18830 4664 19338 4720
rect 19394 4664 19399 4720
rect 18830 4662 19399 4664
rect 19333 4659 19399 4662
rect 20621 4586 20687 4589
rect 15150 4584 20687 4586
rect 15150 4528 20626 4584
rect 20682 4528 20687 4584
rect 15150 4526 20687 4528
rect 20621 4523 20687 4526
rect 12341 4450 12407 4453
rect 14089 4450 14155 4453
rect 12341 4448 14155 4450
rect 12341 4392 12346 4448
rect 12402 4392 14094 4448
rect 14150 4392 14155 4448
rect 12341 4390 14155 4392
rect 12341 4387 12407 4390
rect 14089 4387 14155 4390
rect 22001 4450 22067 4453
rect 22200 4450 23000 4480
rect 22001 4448 23000 4450
rect 22001 4392 22006 4448
rect 22062 4392 23000 4448
rect 22001 4390 23000 4392
rect 22001 4387 22067 4390
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 22200 4360 23000 4390
rect 16538 4319 16858 4320
rect 13721 4314 13787 4317
rect 15377 4314 15443 4317
rect 11792 4312 13787 4314
rect 11792 4256 13726 4312
rect 13782 4256 13787 4312
rect 11792 4254 13787 4256
rect 7741 4251 7807 4254
rect 9489 4251 9555 4254
rect 11145 4251 11211 4254
rect 13721 4251 13787 4254
rect 15150 4312 15443 4314
rect 15150 4256 15382 4312
rect 15438 4256 15443 4312
rect 15150 4254 15443 4256
rect 5073 4178 5139 4181
rect 1945 4176 2790 4178
rect 1945 4120 1950 4176
rect 2006 4120 2790 4176
rect 1945 4118 2790 4120
rect 3558 4176 5139 4178
rect 3558 4120 5078 4176
rect 5134 4120 5139 4176
rect 3558 4118 5139 4120
rect 1945 4115 2011 4118
rect 0 4042 800 4072
rect 933 4042 999 4045
rect 0 4040 999 4042
rect 0 3984 938 4040
rect 994 3984 999 4040
rect 0 3982 999 3984
rect 0 3952 800 3982
rect 933 3979 999 3982
rect 3417 4042 3483 4045
rect 3558 4042 3618 4118
rect 5073 4115 5139 4118
rect 5533 4178 5599 4181
rect 15150 4178 15210 4254
rect 15377 4251 15443 4254
rect 5533 4176 15210 4178
rect 5533 4120 5538 4176
rect 5594 4120 15210 4176
rect 5533 4118 15210 4120
rect 15285 4180 15351 4181
rect 15285 4176 15332 4180
rect 15396 4178 15402 4180
rect 19885 4178 19951 4181
rect 15396 4176 19951 4178
rect 15285 4120 15290 4176
rect 15396 4120 19890 4176
rect 19946 4120 19951 4176
rect 5533 4115 5599 4118
rect 15285 4116 15332 4120
rect 15396 4118 19951 4120
rect 15396 4116 15402 4118
rect 15285 4115 15351 4116
rect 19885 4115 19951 4118
rect 3877 4044 3943 4045
rect 3877 4042 3924 4044
rect 3417 4040 3618 4042
rect 3417 3984 3422 4040
rect 3478 3984 3618 4040
rect 3417 3982 3618 3984
rect 3832 4040 3924 4042
rect 3832 3984 3882 4040
rect 3832 3982 3924 3984
rect 3417 3979 3483 3982
rect 3877 3980 3924 3982
rect 3988 3980 3994 4044
rect 5165 4042 5231 4045
rect 12249 4042 12315 4045
rect 13905 4042 13971 4045
rect 5165 4040 12315 4042
rect 5165 3984 5170 4040
rect 5226 3984 12254 4040
rect 12310 3984 12315 4040
rect 5165 3982 12315 3984
rect 3877 3979 3943 3980
rect 5165 3979 5231 3982
rect 12249 3979 12315 3982
rect 12390 4040 13971 4042
rect 12390 3984 13910 4040
rect 13966 3984 13971 4040
rect 12390 3982 13971 3984
rect 8518 3906 8524 3908
rect 3926 3846 8524 3906
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 0 3634 800 3664
rect 1853 3634 1919 3637
rect 3926 3634 3986 3846
rect 8518 3844 8524 3846
rect 8588 3844 8594 3908
rect 9489 3906 9555 3909
rect 12390 3906 12450 3982
rect 13905 3979 13971 3982
rect 14457 4040 14523 4045
rect 14457 3984 14462 4040
rect 14518 3984 14523 4040
rect 14457 3979 14523 3984
rect 15377 4042 15443 4045
rect 15510 4042 15516 4044
rect 15377 4040 15516 4042
rect 15377 3984 15382 4040
rect 15438 3984 15516 4040
rect 15377 3982 15516 3984
rect 15377 3979 15443 3982
rect 15510 3980 15516 3982
rect 15580 3980 15586 4044
rect 15745 4042 15811 4045
rect 15878 4042 15884 4044
rect 15745 4040 15884 4042
rect 15745 3984 15750 4040
rect 15806 3984 15884 4040
rect 15745 3982 15884 3984
rect 15745 3979 15811 3982
rect 15878 3980 15884 3982
rect 15948 3980 15954 4044
rect 20253 4042 20319 4045
rect 16070 4040 20319 4042
rect 16070 3984 20258 4040
rect 20314 3984 20319 4040
rect 16070 3982 20319 3984
rect 9489 3904 12450 3906
rect 9489 3848 9494 3904
rect 9550 3848 12450 3904
rect 9489 3846 12450 3848
rect 9489 3843 9555 3846
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 4521 3770 4587 3773
rect 6862 3770 6868 3772
rect 4521 3768 6868 3770
rect 4521 3712 4526 3768
rect 4582 3712 6868 3768
rect 4521 3710 6868 3712
rect 4521 3707 4587 3710
rect 6862 3708 6868 3710
rect 6932 3708 6938 3772
rect 7005 3770 7071 3773
rect 7414 3770 7420 3772
rect 7005 3768 7420 3770
rect 7005 3712 7010 3768
rect 7066 3712 7420 3768
rect 7005 3710 7420 3712
rect 7005 3707 7071 3710
rect 7414 3708 7420 3710
rect 7484 3708 7490 3772
rect 7649 3770 7715 3773
rect 8150 3770 8156 3772
rect 7649 3768 8156 3770
rect 7649 3712 7654 3768
rect 7710 3712 8156 3768
rect 7649 3710 8156 3712
rect 7649 3707 7715 3710
rect 8150 3708 8156 3710
rect 8220 3708 8226 3772
rect 12985 3770 13051 3773
rect 9124 3768 13051 3770
rect 9124 3712 12990 3768
rect 13046 3712 13051 3768
rect 9124 3710 13051 3712
rect 14460 3770 14520 3979
rect 14641 3906 14707 3909
rect 16070 3906 16130 3982
rect 20253 3979 20319 3982
rect 21633 4042 21699 4045
rect 22200 4042 23000 4072
rect 21633 4040 23000 4042
rect 21633 3984 21638 4040
rect 21694 3984 23000 4040
rect 21633 3982 23000 3984
rect 21633 3979 21699 3982
rect 22200 3952 23000 3982
rect 14641 3904 16130 3906
rect 14641 3848 14646 3904
rect 14702 3848 16130 3904
rect 14641 3846 16130 3848
rect 14641 3843 14707 3846
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 15101 3770 15167 3773
rect 14460 3768 15167 3770
rect 14460 3712 15106 3768
rect 15162 3712 15167 3768
rect 14460 3710 15167 3712
rect 0 3574 1778 3634
rect 0 3544 800 3574
rect 1718 3498 1778 3574
rect 1853 3632 3986 3634
rect 1853 3576 1858 3632
rect 1914 3576 3986 3632
rect 1853 3574 3986 3576
rect 4245 3634 4311 3637
rect 5625 3634 5691 3637
rect 4245 3632 5691 3634
rect 4245 3576 4250 3632
rect 4306 3576 5630 3632
rect 5686 3576 5691 3632
rect 4245 3574 5691 3576
rect 1853 3571 1919 3574
rect 4245 3571 4311 3574
rect 5625 3571 5691 3574
rect 6085 3634 6151 3637
rect 9124 3634 9184 3710
rect 12985 3707 13051 3710
rect 15101 3707 15167 3710
rect 15929 3770 15995 3773
rect 17902 3770 17908 3772
rect 15929 3768 17908 3770
rect 15929 3712 15934 3768
rect 15990 3712 17908 3768
rect 15929 3710 17908 3712
rect 15929 3707 15995 3710
rect 17902 3708 17908 3710
rect 17972 3708 17978 3772
rect 19701 3770 19767 3773
rect 19701 3768 19994 3770
rect 19701 3712 19706 3768
rect 19762 3712 19994 3768
rect 19701 3710 19994 3712
rect 19701 3707 19767 3710
rect 6085 3632 9184 3634
rect 6085 3576 6090 3632
rect 6146 3576 9184 3632
rect 6085 3574 9184 3576
rect 10409 3634 10475 3637
rect 10542 3634 10548 3636
rect 10409 3632 10548 3634
rect 10409 3576 10414 3632
rect 10470 3576 10548 3632
rect 10409 3574 10548 3576
rect 6085 3571 6151 3574
rect 10409 3571 10475 3574
rect 10542 3572 10548 3574
rect 10612 3572 10618 3636
rect 10726 3572 10732 3636
rect 10796 3634 10802 3636
rect 12014 3634 12020 3636
rect 10796 3574 12020 3634
rect 10796 3572 10802 3574
rect 12014 3572 12020 3574
rect 12084 3572 12090 3636
rect 12157 3634 12223 3637
rect 12617 3634 12683 3637
rect 12157 3632 12683 3634
rect 12157 3576 12162 3632
rect 12218 3576 12622 3632
rect 12678 3576 12683 3632
rect 12157 3574 12683 3576
rect 12157 3571 12223 3574
rect 12617 3571 12683 3574
rect 13077 3634 13143 3637
rect 15469 3634 15535 3637
rect 13077 3632 15535 3634
rect 13077 3576 13082 3632
rect 13138 3576 15474 3632
rect 15530 3576 15535 3632
rect 13077 3574 15535 3576
rect 13077 3571 13143 3574
rect 15469 3571 15535 3574
rect 15837 3634 15903 3637
rect 19701 3634 19767 3637
rect 15837 3632 19767 3634
rect 15837 3576 15842 3632
rect 15898 3576 19706 3632
rect 19762 3576 19767 3632
rect 15837 3574 19767 3576
rect 19934 3634 19994 3710
rect 22200 3634 23000 3664
rect 19934 3574 23000 3634
rect 15837 3571 15903 3574
rect 19701 3571 19767 3574
rect 22200 3544 23000 3574
rect 4889 3498 4955 3501
rect 1718 3496 4955 3498
rect 1718 3440 4894 3496
rect 4950 3440 4955 3496
rect 1718 3438 4955 3440
rect 4889 3435 4955 3438
rect 5993 3498 6059 3501
rect 14365 3498 14431 3501
rect 5993 3496 14431 3498
rect 5993 3440 5998 3496
rect 6054 3440 14370 3496
rect 14426 3440 14431 3496
rect 5993 3438 14431 3440
rect 5993 3435 6059 3438
rect 14365 3435 14431 3438
rect 16297 3498 16363 3501
rect 21449 3498 21515 3501
rect 16297 3496 21515 3498
rect 16297 3440 16302 3496
rect 16358 3440 21454 3496
rect 21510 3440 21515 3496
rect 16297 3438 21515 3440
rect 16297 3435 16363 3438
rect 21449 3435 21515 3438
rect 6545 3362 6611 3365
rect 9489 3362 9555 3365
rect 6545 3360 9555 3362
rect 6545 3304 6550 3360
rect 6606 3304 9494 3360
rect 9550 3304 9555 3360
rect 6545 3302 9555 3304
rect 6545 3299 6611 3302
rect 9489 3299 9555 3302
rect 11881 3362 11947 3365
rect 12198 3362 12204 3364
rect 11881 3360 12204 3362
rect 11881 3304 11886 3360
rect 11942 3304 12204 3360
rect 11881 3302 12204 3304
rect 11881 3299 11947 3302
rect 12198 3300 12204 3302
rect 12268 3300 12274 3364
rect 12433 3362 12499 3365
rect 13486 3362 13492 3364
rect 12433 3360 13492 3362
rect 12433 3304 12438 3360
rect 12494 3304 13492 3360
rect 12433 3302 13492 3304
rect 12433 3299 12499 3302
rect 13486 3300 13492 3302
rect 13556 3300 13562 3364
rect 14917 3362 14983 3365
rect 15142 3362 15148 3364
rect 14917 3360 15148 3362
rect 14917 3304 14922 3360
rect 14978 3304 15148 3360
rect 14917 3302 15148 3304
rect 14917 3299 14983 3302
rect 15142 3300 15148 3302
rect 15212 3300 15218 3364
rect 17953 3362 18019 3365
rect 19006 3362 19012 3364
rect 17953 3360 19012 3362
rect 17953 3304 17958 3360
rect 18014 3304 19012 3360
rect 17953 3302 19012 3304
rect 17953 3299 18019 3302
rect 19006 3300 19012 3302
rect 19076 3300 19082 3364
rect 21950 3300 21956 3364
rect 22020 3362 22026 3364
rect 22277 3362 22343 3365
rect 22020 3360 22343 3362
rect 22020 3304 22282 3360
rect 22338 3304 22343 3360
rect 22020 3302 22343 3304
rect 22020 3300 22026 3302
rect 22277 3299 22343 3302
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 3231 16858 3232
rect 2589 3228 2655 3229
rect 2589 3226 2636 3228
rect 2544 3224 2636 3226
rect 2700 3226 2706 3228
rect 5257 3226 5323 3229
rect 2700 3224 5323 3226
rect 2544 3168 2594 3224
rect 2700 3168 5262 3224
rect 5318 3168 5323 3224
rect 2544 3166 2636 3168
rect 2589 3164 2636 3166
rect 2700 3166 5323 3168
rect 2700 3164 2706 3166
rect 2589 3163 2655 3164
rect 5257 3163 5323 3166
rect 5574 3164 5580 3228
rect 5644 3226 5650 3228
rect 5809 3226 5875 3229
rect 5644 3224 5875 3226
rect 5644 3168 5814 3224
rect 5870 3168 5875 3224
rect 5644 3166 5875 3168
rect 5644 3164 5650 3166
rect 5809 3163 5875 3166
rect 8569 3226 8635 3229
rect 10961 3226 11027 3229
rect 11145 3228 11211 3229
rect 8569 3224 11027 3226
rect 8569 3168 8574 3224
rect 8630 3168 10966 3224
rect 11022 3168 11027 3224
rect 8569 3166 11027 3168
rect 8569 3163 8635 3166
rect 10961 3163 11027 3166
rect 11094 3164 11100 3228
rect 11164 3226 11211 3228
rect 12065 3226 12131 3229
rect 12382 3226 12388 3228
rect 11164 3224 11256 3226
rect 11206 3168 11256 3224
rect 11164 3166 11256 3168
rect 12065 3224 12388 3226
rect 12065 3168 12070 3224
rect 12126 3168 12388 3224
rect 12065 3166 12388 3168
rect 11164 3164 11211 3166
rect 11145 3163 11211 3164
rect 12065 3163 12131 3166
rect 12382 3164 12388 3166
rect 12452 3164 12458 3228
rect 18689 3226 18755 3229
rect 19609 3226 19675 3229
rect 18689 3224 19675 3226
rect 18689 3168 18694 3224
rect 18750 3168 19614 3224
rect 19670 3168 19675 3224
rect 18689 3166 19675 3168
rect 18689 3163 18755 3166
rect 19609 3163 19675 3166
rect 20161 3226 20227 3229
rect 20161 3224 22202 3226
rect 20161 3168 20166 3224
rect 20222 3168 22202 3224
rect 20161 3166 22202 3168
rect 20161 3163 20227 3166
rect 22142 3120 22202 3166
rect 0 3090 800 3120
rect 5206 3090 5212 3092
rect 0 3030 5212 3090
rect 0 3000 800 3030
rect 5206 3028 5212 3030
rect 5276 3028 5282 3092
rect 5441 3090 5507 3093
rect 7414 3090 7420 3092
rect 5441 3088 7420 3090
rect 5441 3032 5446 3088
rect 5502 3032 7420 3088
rect 5441 3030 7420 3032
rect 5441 3027 5507 3030
rect 7414 3028 7420 3030
rect 7484 3028 7490 3092
rect 8017 3090 8083 3093
rect 12566 3090 12572 3092
rect 8017 3088 12572 3090
rect 8017 3032 8022 3088
rect 8078 3032 12572 3088
rect 8017 3030 12572 3032
rect 8017 3027 8083 3030
rect 12566 3028 12572 3030
rect 12636 3028 12642 3092
rect 15193 3090 15259 3093
rect 22001 3090 22067 3093
rect 15193 3088 22067 3090
rect 15193 3032 15198 3088
rect 15254 3032 22006 3088
rect 22062 3032 22067 3088
rect 15193 3030 22067 3032
rect 22142 3030 23000 3120
rect 15193 3027 15259 3030
rect 22001 3027 22067 3030
rect 22200 3000 23000 3030
rect 1342 2892 1348 2956
rect 1412 2954 1418 2956
rect 2773 2954 2839 2957
rect 5901 2954 5967 2957
rect 1412 2952 2839 2954
rect 1412 2896 2778 2952
rect 2834 2896 2839 2952
rect 1412 2894 2839 2896
rect 1412 2892 1418 2894
rect 2773 2891 2839 2894
rect 3420 2952 5967 2954
rect 3420 2896 5906 2952
rect 5962 2896 5967 2952
rect 3420 2894 5967 2896
rect 1710 2756 1716 2820
rect 1780 2818 1786 2820
rect 2681 2818 2747 2821
rect 1780 2816 2747 2818
rect 1780 2760 2686 2816
rect 2742 2760 2747 2816
rect 1780 2758 2747 2760
rect 1780 2756 1786 2758
rect 2681 2755 2747 2758
rect 0 2682 800 2712
rect 3420 2682 3480 2894
rect 5901 2891 5967 2894
rect 9673 2954 9739 2957
rect 10225 2954 10291 2957
rect 14273 2954 14339 2957
rect 9673 2952 14339 2954
rect 9673 2896 9678 2952
rect 9734 2896 10230 2952
rect 10286 2896 14278 2952
rect 14334 2896 14339 2952
rect 9673 2894 14339 2896
rect 9673 2891 9739 2894
rect 10225 2891 10291 2894
rect 14273 2891 14339 2894
rect 15561 2954 15627 2957
rect 21909 2954 21975 2957
rect 15561 2952 21975 2954
rect 15561 2896 15566 2952
rect 15622 2896 21914 2952
rect 21970 2896 21975 2952
rect 15561 2894 21975 2896
rect 15561 2891 15627 2894
rect 21909 2891 21975 2894
rect 4153 2818 4219 2821
rect 4521 2818 4587 2821
rect 4153 2816 4587 2818
rect 4153 2760 4158 2816
rect 4214 2760 4526 2816
rect 4582 2760 4587 2816
rect 4153 2758 4587 2760
rect 4153 2755 4219 2758
rect 4521 2755 4587 2758
rect 7046 2756 7052 2820
rect 7116 2818 7122 2820
rect 7833 2818 7899 2821
rect 7116 2816 7899 2818
rect 7116 2760 7838 2816
rect 7894 2760 7899 2816
rect 7116 2758 7899 2760
rect 7116 2756 7122 2758
rect 7833 2755 7899 2758
rect 9254 2756 9260 2820
rect 9324 2818 9330 2820
rect 11789 2818 11855 2821
rect 9324 2816 11855 2818
rect 9324 2760 11794 2816
rect 11850 2760 11855 2816
rect 9324 2758 11855 2760
rect 9324 2756 9330 2758
rect 11789 2755 11855 2758
rect 17861 2818 17927 2821
rect 18229 2818 18295 2821
rect 18965 2818 19031 2821
rect 17861 2816 19031 2818
rect 17861 2760 17866 2816
rect 17922 2760 18234 2816
rect 18290 2760 18970 2816
rect 19026 2760 19031 2816
rect 17861 2758 19031 2760
rect 17861 2755 17927 2758
rect 18229 2755 18295 2758
rect 18965 2755 19031 2758
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 0 2622 3480 2682
rect 4705 2682 4771 2685
rect 5809 2682 5875 2685
rect 5942 2682 5948 2684
rect 4705 2680 4906 2682
rect 4705 2624 4710 2680
rect 4766 2624 4906 2680
rect 4705 2622 4906 2624
rect 0 2592 800 2622
rect 4705 2619 4771 2622
rect 4846 2546 4906 2622
rect 5809 2680 5948 2682
rect 5809 2624 5814 2680
rect 5870 2624 5948 2680
rect 5809 2622 5948 2624
rect 5809 2619 5875 2622
rect 5942 2620 5948 2622
rect 6012 2620 6018 2684
rect 7005 2682 7071 2685
rect 7649 2684 7715 2685
rect 7230 2682 7236 2684
rect 7005 2680 7236 2682
rect 7005 2624 7010 2680
rect 7066 2624 7236 2680
rect 7005 2622 7236 2624
rect 7005 2619 7071 2622
rect 7230 2620 7236 2622
rect 7300 2620 7306 2684
rect 7598 2620 7604 2684
rect 7668 2682 7715 2684
rect 9121 2682 9187 2685
rect 14641 2684 14707 2685
rect 11830 2682 11836 2684
rect 7668 2680 7760 2682
rect 7710 2624 7760 2680
rect 7668 2622 7760 2624
rect 9121 2680 11836 2682
rect 9121 2624 9126 2680
rect 9182 2624 11836 2680
rect 9121 2622 11836 2624
rect 7668 2620 7715 2622
rect 7649 2619 7715 2620
rect 9121 2619 9187 2622
rect 11830 2620 11836 2622
rect 11900 2620 11906 2684
rect 14590 2682 14596 2684
rect 14550 2622 14596 2682
rect 14660 2680 14707 2684
rect 14702 2624 14707 2680
rect 14590 2620 14596 2622
rect 14660 2620 14707 2624
rect 14641 2619 14707 2620
rect 20713 2682 20779 2685
rect 22200 2682 23000 2712
rect 20713 2680 23000 2682
rect 20713 2624 20718 2680
rect 20774 2624 23000 2680
rect 20713 2622 23000 2624
rect 20713 2619 20779 2622
rect 22200 2592 23000 2622
rect 8569 2546 8635 2549
rect 4846 2544 8635 2546
rect 4846 2488 8574 2544
rect 8630 2488 8635 2544
rect 4846 2486 8635 2488
rect 8569 2483 8635 2486
rect 8753 2546 8819 2549
rect 9121 2546 9187 2549
rect 12750 2546 12756 2548
rect 8753 2544 12756 2546
rect 8753 2488 8758 2544
rect 8814 2488 9126 2544
rect 9182 2488 12756 2544
rect 8753 2486 12756 2488
rect 8753 2483 8819 2486
rect 9121 2483 9187 2486
rect 12750 2484 12756 2486
rect 12820 2484 12826 2548
rect 18270 2484 18276 2548
rect 18340 2546 18346 2548
rect 18413 2546 18479 2549
rect 18340 2544 18479 2546
rect 18340 2488 18418 2544
rect 18474 2488 18479 2544
rect 18340 2486 18479 2488
rect 18340 2484 18346 2486
rect 18413 2483 18479 2486
rect 4981 2410 5047 2413
rect 10726 2410 10732 2412
rect 4981 2408 10732 2410
rect 4981 2352 4986 2408
rect 5042 2352 10732 2408
rect 4981 2350 10732 2352
rect 4981 2347 5047 2350
rect 10726 2348 10732 2350
rect 10796 2348 10802 2412
rect 21725 2410 21791 2413
rect 10872 2408 21791 2410
rect 10872 2352 21730 2408
rect 21786 2352 21791 2408
rect 10872 2350 21791 2352
rect 0 2274 800 2304
rect 5717 2276 5783 2277
rect 4654 2274 4660 2276
rect 0 2214 4660 2274
rect 0 2184 800 2214
rect 4654 2212 4660 2214
rect 4724 2212 4730 2276
rect 5717 2272 5764 2276
rect 5828 2274 5834 2276
rect 7189 2274 7255 2277
rect 10872 2274 10932 2350
rect 21725 2347 21791 2350
rect 5717 2216 5722 2272
rect 5717 2212 5764 2216
rect 5828 2214 5874 2274
rect 7189 2272 10932 2274
rect 7189 2216 7194 2272
rect 7250 2216 10932 2272
rect 7189 2214 10932 2216
rect 21541 2274 21607 2277
rect 22200 2274 23000 2304
rect 21541 2272 23000 2274
rect 21541 2216 21546 2272
rect 21602 2216 23000 2272
rect 21541 2214 23000 2216
rect 5828 2212 5834 2214
rect 5717 2211 5783 2212
rect 7189 2211 7255 2214
rect 21541 2211 21607 2214
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 22200 2184 23000 2214
rect 16538 2143 16858 2144
rect 4838 2076 4844 2140
rect 4908 2138 4914 2140
rect 5993 2138 6059 2141
rect 4908 2136 6059 2138
rect 4908 2080 5998 2136
rect 6054 2080 6059 2136
rect 4908 2078 6059 2080
rect 4908 2076 4914 2078
rect 5993 2075 6059 2078
rect 1301 2002 1367 2005
rect 7281 2002 7347 2005
rect 1301 2000 7347 2002
rect 1301 1944 1306 2000
rect 1362 1944 7286 2000
rect 7342 1944 7347 2000
rect 1301 1942 7347 1944
rect 1301 1939 1367 1942
rect 7281 1939 7347 1942
rect 10409 2002 10475 2005
rect 16205 2002 16271 2005
rect 19558 2002 19564 2004
rect 10409 2000 19564 2002
rect 10409 1944 10414 2000
rect 10470 1944 16210 2000
rect 16266 1944 19564 2000
rect 10409 1942 19564 1944
rect 10409 1939 10475 1942
rect 16205 1939 16271 1942
rect 19558 1940 19564 1942
rect 19628 1940 19634 2004
rect 0 1866 800 1896
rect 4245 1866 4311 1869
rect 5993 1866 6059 1869
rect 10910 1866 10916 1868
rect 0 1806 3940 1866
rect 0 1776 800 1806
rect 3880 1730 3940 1806
rect 4245 1864 10916 1866
rect 4245 1808 4250 1864
rect 4306 1808 5998 1864
rect 6054 1808 10916 1864
rect 4245 1806 10916 1808
rect 4245 1803 4311 1806
rect 5993 1803 6059 1806
rect 10910 1804 10916 1806
rect 10980 1804 10986 1868
rect 21817 1866 21883 1869
rect 22200 1866 23000 1896
rect 21817 1864 23000 1866
rect 21817 1808 21822 1864
rect 21878 1808 23000 1864
rect 21817 1806 23000 1808
rect 21817 1803 21883 1806
rect 22200 1776 23000 1806
rect 6729 1730 6795 1733
rect 3880 1728 6795 1730
rect 3880 1672 6734 1728
rect 6790 1672 6795 1728
rect 3880 1670 6795 1672
rect 6729 1667 6795 1670
rect 6913 1730 6979 1733
rect 8937 1730 9003 1733
rect 14406 1730 14412 1732
rect 6913 1728 14412 1730
rect 6913 1672 6918 1728
rect 6974 1672 8942 1728
rect 8998 1672 14412 1728
rect 6913 1670 14412 1672
rect 6913 1667 6979 1670
rect 8937 1667 9003 1670
rect 14406 1668 14412 1670
rect 14476 1668 14482 1732
rect 5625 1594 5691 1597
rect 7189 1594 7255 1597
rect 5625 1592 7255 1594
rect 5625 1536 5630 1592
rect 5686 1536 7194 1592
rect 7250 1536 7255 1592
rect 5625 1534 7255 1536
rect 5625 1531 5691 1534
rect 7189 1531 7255 1534
rect 7782 1532 7788 1596
rect 7852 1594 7858 1596
rect 8569 1594 8635 1597
rect 15326 1594 15332 1596
rect 7852 1592 15332 1594
rect 7852 1536 8574 1592
rect 8630 1536 15332 1592
rect 7852 1534 15332 1536
rect 7852 1532 7858 1534
rect 8569 1531 8635 1534
rect 15326 1532 15332 1534
rect 15396 1532 15402 1596
rect 0 1458 800 1488
rect 2078 1458 2084 1460
rect 0 1398 2084 1458
rect 0 1368 800 1398
rect 2078 1396 2084 1398
rect 2148 1396 2154 1460
rect 7925 1458 7991 1461
rect 17718 1458 17724 1460
rect 7925 1456 17724 1458
rect 7925 1400 7930 1456
rect 7986 1400 17724 1456
rect 7925 1398 17724 1400
rect 7925 1395 7991 1398
rect 17718 1396 17724 1398
rect 17788 1396 17794 1460
rect 19241 1458 19307 1461
rect 22200 1458 23000 1488
rect 19241 1456 23000 1458
rect 19241 1400 19246 1456
rect 19302 1400 23000 1456
rect 19241 1398 23000 1400
rect 19241 1395 19307 1398
rect 22200 1368 23000 1398
rect 5165 1322 5231 1325
rect 14917 1322 14983 1325
rect 5165 1320 14983 1322
rect 5165 1264 5170 1320
rect 5226 1264 14922 1320
rect 14978 1264 14983 1320
rect 5165 1262 14983 1264
rect 5165 1259 5231 1262
rect 14917 1259 14983 1262
rect 7465 1186 7531 1189
rect 15142 1186 15148 1188
rect 7465 1184 15148 1186
rect 7465 1128 7470 1184
rect 7526 1128 15148 1184
rect 7465 1126 15148 1128
rect 7465 1123 7531 1126
rect 15142 1124 15148 1126
rect 15212 1124 15218 1188
rect 0 1050 800 1080
rect 3366 1050 3372 1052
rect 0 990 3372 1050
rect 0 960 800 990
rect 3366 988 3372 990
rect 3436 988 3442 1052
rect 4889 1050 4955 1053
rect 13670 1050 13676 1052
rect 4889 1048 13676 1050
rect 4889 992 4894 1048
rect 4950 992 13676 1048
rect 4889 990 13676 992
rect 4889 987 4955 990
rect 13670 988 13676 990
rect 13740 988 13746 1052
rect 20713 1050 20779 1053
rect 22200 1050 23000 1080
rect 20713 1048 23000 1050
rect 20713 992 20718 1048
rect 20774 992 23000 1048
rect 20713 990 23000 992
rect 20713 987 20779 990
rect 22200 960 23000 990
rect 3233 914 3299 917
rect 2454 912 3299 914
rect 2454 856 3238 912
rect 3294 856 3299 912
rect 2454 854 3299 856
rect 0 642 800 672
rect 2454 642 2514 854
rect 3233 851 3299 854
rect 5073 914 5139 917
rect 18454 914 18460 916
rect 5073 912 18460 914
rect 5073 856 5078 912
rect 5134 856 18460 912
rect 5073 854 18460 856
rect 5073 851 5139 854
rect 18454 852 18460 854
rect 18524 852 18530 916
rect 18689 912 18755 917
rect 18689 856 18694 912
rect 18750 856 18755 912
rect 18689 851 18755 856
rect 0 582 2514 642
rect 18692 642 18752 851
rect 22200 642 23000 672
rect 18692 582 23000 642
rect 0 552 800 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 933 234 999 237
rect 0 232 999 234
rect 0 176 938 232
rect 994 176 999 232
rect 0 174 999 176
rect 0 144 800 174
rect 933 171 999 174
rect 19609 234 19675 237
rect 22200 234 23000 264
rect 19609 232 23000 234
rect 19609 176 19614 232
rect 19670 176 23000 232
rect 19609 174 23000 176
rect 19609 171 19675 174
rect 22200 144 23000 174
<< via3 >>
rect 16988 22884 17052 22948
rect 980 22748 1044 22812
rect 6868 22612 6932 22676
rect 19932 22476 19996 22540
rect 14412 22340 14476 22404
rect 15332 22204 15396 22268
rect 980 22068 1044 22132
rect 13676 22068 13740 22132
rect 14596 21932 14660 21996
rect 18092 21796 18156 21860
rect 15148 21660 15212 21724
rect 1532 21524 1596 21588
rect 4660 21388 4724 21452
rect 17908 21388 17972 21452
rect 1164 21252 1228 21316
rect 13492 21252 13556 21316
rect 18460 21116 18524 21180
rect 17172 20980 17236 21044
rect 2636 20844 2700 20908
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 6684 20164 6748 20228
rect 7420 20164 7484 20228
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 7788 20028 7852 20092
rect 9628 20028 9692 20092
rect 12204 20028 12268 20092
rect 3372 19816 3436 19820
rect 3372 19760 3386 19816
rect 3386 19760 3436 19816
rect 3372 19756 3436 19760
rect 13124 19756 13188 19820
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 7972 19348 8036 19412
rect 9444 19348 9508 19412
rect 9996 19408 10060 19412
rect 9996 19352 10010 19408
rect 10010 19352 10060 19408
rect 9996 19348 10060 19352
rect 10364 19408 10428 19412
rect 10364 19352 10378 19408
rect 10378 19352 10428 19408
rect 10364 19348 10428 19352
rect 19564 19348 19628 19412
rect 2636 19212 2700 19276
rect 15148 19272 15212 19276
rect 15148 19216 15198 19272
rect 15198 19216 15212 19272
rect 15148 19212 15212 19216
rect 15332 19272 15396 19276
rect 15332 19216 15382 19272
rect 15382 19216 15396 19272
rect 15332 19212 15396 19216
rect 14596 19076 14660 19140
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 9260 18940 9324 19004
rect 18092 18940 18156 19004
rect 9812 18668 9876 18732
rect 2820 18592 2884 18596
rect 2820 18536 2870 18592
rect 2870 18536 2884 18592
rect 2820 18532 2884 18536
rect 5212 18532 5276 18596
rect 5580 18592 5644 18596
rect 14412 18728 14476 18732
rect 14412 18672 14426 18728
rect 14426 18672 14476 18728
rect 14412 18668 14476 18672
rect 5580 18536 5630 18592
rect 5630 18536 5644 18592
rect 5580 18532 5644 18536
rect 11100 18592 11164 18596
rect 11100 18536 11114 18592
rect 11114 18536 11164 18592
rect 11100 18532 11164 18536
rect 12020 18532 12084 18596
rect 12572 18532 12636 18596
rect 13676 18532 13740 18596
rect 17540 18532 17604 18596
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 6868 18396 6932 18460
rect 7972 18396 8036 18460
rect 5028 18260 5092 18324
rect 18460 18456 18524 18460
rect 18460 18400 18510 18456
rect 18510 18400 18524 18456
rect 18460 18396 18524 18400
rect 2084 18048 2148 18052
rect 2084 17992 2134 18048
rect 2134 17992 2148 18048
rect 2084 17988 2148 17992
rect 9260 18124 9324 18188
rect 9628 18184 9692 18188
rect 9628 18128 9642 18184
rect 9642 18128 9692 18184
rect 9628 18124 9692 18128
rect 9812 18124 9876 18188
rect 10916 17988 10980 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 13308 17852 13372 17916
rect 16988 17852 17052 17916
rect 17908 17912 17972 17916
rect 17908 17856 17958 17912
rect 17958 17856 17972 17912
rect 17908 17852 17972 17856
rect 3188 17580 3252 17644
rect 5764 17640 5828 17644
rect 5764 17584 5778 17640
rect 5778 17584 5828 17640
rect 5764 17580 5828 17584
rect 14412 17716 14476 17780
rect 19012 17716 19076 17780
rect 19932 17716 19996 17780
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 7972 17172 8036 17236
rect 3924 17036 3988 17100
rect 19564 17172 19628 17236
rect 13492 17036 13556 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 5948 16764 6012 16828
rect 11100 16764 11164 16828
rect 11836 16764 11900 16828
rect 1900 16628 1964 16692
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 12572 16628 12636 16692
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 8340 16220 8404 16284
rect 12940 16220 13004 16284
rect 12204 15948 12268 16012
rect 17908 15948 17972 16012
rect 8156 15812 8220 15876
rect 10732 15812 10796 15876
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 5212 15676 5276 15740
rect 4108 15540 4172 15604
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 18276 15268 18340 15332
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 7604 15132 7668 15196
rect 13308 15132 13372 15196
rect 15332 15132 15396 15196
rect 12020 14996 12084 15060
rect 3004 14860 3068 14924
rect 16988 14996 17052 15060
rect 16068 14860 16132 14924
rect 14596 14724 14660 14788
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 7420 14180 7484 14244
rect 12572 14180 12636 14244
rect 16252 14180 16316 14244
rect 18460 14180 18524 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 6684 14044 6748 14108
rect 7236 14044 7300 14108
rect 17172 14104 17236 14108
rect 17172 14048 17222 14104
rect 17222 14048 17236 14104
rect 17172 14044 17236 14048
rect 7052 13908 7116 13972
rect 7420 13772 7484 13836
rect 4844 13636 4908 13700
rect 5948 13636 6012 13700
rect 9812 13772 9876 13836
rect 12756 13772 12820 13836
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 9444 13636 9508 13700
rect 10916 13636 10980 13700
rect 15332 13636 15396 13700
rect 17172 13832 17236 13836
rect 17172 13776 17186 13832
rect 17186 13776 17236 13832
rect 17172 13772 17236 13776
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 9260 13500 9324 13564
rect 12204 13500 12268 13564
rect 13492 13500 13556 13564
rect 19564 13560 19628 13564
rect 19564 13504 19578 13560
rect 19578 13504 19628 13560
rect 19564 13500 19628 13504
rect 9628 13228 9692 13292
rect 796 13092 860 13156
rect 3372 13092 3436 13156
rect 6684 13092 6748 13156
rect 13676 13228 13740 13292
rect 14780 13228 14844 13292
rect 18092 13092 18156 13156
rect 21404 13092 21468 13156
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 5396 12956 5460 13020
rect 8524 12820 8588 12884
rect 15700 12820 15764 12884
rect 16068 12820 16132 12884
rect 4292 12684 4356 12748
rect 2820 12548 2884 12612
rect 12388 12684 12452 12748
rect 17908 12684 17972 12748
rect 10180 12548 10244 12612
rect 11100 12548 11164 12612
rect 15148 12548 15212 12612
rect 15332 12548 15396 12612
rect 15884 12548 15948 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 2820 12412 2884 12476
rect 3004 12276 3068 12340
rect 17356 12548 17420 12612
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 9996 12200 10060 12204
rect 9996 12144 10046 12200
rect 10046 12144 10060 12200
rect 9996 12140 10060 12144
rect 15700 12412 15764 12476
rect 20484 12412 20548 12476
rect 12940 12336 13004 12340
rect 12940 12280 12990 12336
rect 12990 12280 13004 12336
rect 12940 12276 13004 12280
rect 17724 12140 17788 12204
rect 21220 12140 21284 12204
rect 2820 12004 2884 12068
rect 10916 12004 10980 12068
rect 15700 12004 15764 12068
rect 16252 12064 16316 12068
rect 16252 12008 16302 12064
rect 16302 12008 16316 12064
rect 16252 12004 16316 12008
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 5212 11868 5276 11932
rect 6684 11928 6748 11932
rect 6684 11872 6698 11928
rect 6698 11872 6748 11928
rect 6684 11868 6748 11872
rect 7420 11868 7484 11932
rect 18644 11868 18708 11932
rect 19748 11928 19812 11932
rect 19748 11872 19762 11928
rect 19762 11872 19812 11928
rect 19748 11868 19812 11872
rect 5948 11596 6012 11660
rect 7420 11460 7484 11524
rect 12020 11596 12084 11660
rect 13124 11596 13188 11660
rect 13676 11596 13740 11660
rect 17724 11596 17788 11660
rect 19932 11656 19996 11660
rect 19932 11600 19946 11656
rect 19946 11600 19996 11656
rect 19932 11596 19996 11600
rect 12572 11460 12636 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6684 11324 6748 11388
rect 7972 11384 8036 11388
rect 7972 11328 8022 11384
rect 8022 11328 8036 11384
rect 7972 11324 8036 11328
rect 9260 11324 9324 11388
rect 9812 11324 9876 11388
rect 11836 11324 11900 11388
rect 14964 11324 15028 11388
rect 18276 11324 18340 11388
rect 10180 11188 10244 11252
rect 12572 11188 12636 11252
rect 13124 11188 13188 11252
rect 2820 11052 2884 11116
rect 3372 11052 3436 11116
rect 7420 11052 7484 11116
rect 8524 11052 8588 11116
rect 9260 11112 9324 11116
rect 9260 11056 9274 11112
rect 9274 11056 9324 11112
rect 9260 11052 9324 11056
rect 10364 11052 10428 11116
rect 1716 10916 1780 10980
rect 18092 11052 18156 11116
rect 19564 11052 19628 11116
rect 21956 11052 22020 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 5948 10780 6012 10844
rect 12204 10780 12268 10844
rect 7788 10508 7852 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 5396 10236 5460 10300
rect 5764 10236 5828 10300
rect 6684 10372 6748 10436
rect 7604 10372 7668 10436
rect 12204 10508 12268 10572
rect 20484 10508 20548 10572
rect 15516 10372 15580 10436
rect 17356 10372 17420 10436
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6546 10236 6610 10300
rect 12204 10160 12268 10164
rect 12204 10104 12218 10160
rect 12218 10104 12268 10160
rect 12204 10100 12268 10104
rect 15700 10236 15764 10300
rect 20852 10236 20916 10300
rect 16068 10100 16132 10164
rect 3004 9828 3068 9892
rect 4292 9828 4356 9892
rect 12388 9828 12452 9892
rect 17540 9964 17604 10028
rect 18828 9828 18892 9892
rect 20116 9828 20180 9892
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 4108 9692 4172 9756
rect 4476 9692 4540 9756
rect 5212 9692 5276 9756
rect 5764 9692 5828 9756
rect 7052 9692 7116 9756
rect 7604 9692 7668 9756
rect 7972 9692 8036 9756
rect 8524 9692 8588 9756
rect 9444 9692 9508 9756
rect 9628 9752 9692 9756
rect 9628 9696 9642 9752
rect 9642 9696 9692 9752
rect 9628 9692 9692 9696
rect 16068 9692 16132 9756
rect 6868 9556 6932 9620
rect 2084 9420 2148 9484
rect 4108 9420 4172 9484
rect 5212 9420 5276 9484
rect 7052 9420 7116 9484
rect 8156 9420 8220 9484
rect 10548 9556 10612 9620
rect 19012 9556 19076 9620
rect 2084 9284 2148 9348
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 8156 9148 8220 9212
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 12388 9148 12452 9212
rect 13308 9148 13372 9212
rect 14596 9148 14660 9212
rect 18460 9148 18524 9212
rect 2820 8800 2884 8804
rect 2820 8744 2870 8800
rect 2870 8744 2884 8800
rect 2820 8740 2884 8744
rect 7788 8876 7852 8940
rect 18828 8876 18892 8940
rect 15148 8740 15212 8804
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 9260 8604 9324 8668
rect 9444 8604 9508 8668
rect 10916 8664 10980 8668
rect 10916 8608 10930 8664
rect 10930 8608 10980 8664
rect 10916 8604 10980 8608
rect 12388 8604 12452 8668
rect 4844 8468 4908 8532
rect 5212 8528 5276 8532
rect 10364 8528 10428 8532
rect 5212 8472 5262 8528
rect 5262 8472 5276 8528
rect 5212 8468 5276 8472
rect 10364 8472 10378 8528
rect 10378 8472 10428 8528
rect 10364 8468 10428 8472
rect 10548 8468 10612 8532
rect 12940 8664 13004 8668
rect 12940 8608 12954 8664
rect 12954 8608 13004 8664
rect 12940 8604 13004 8608
rect 19012 8604 19076 8668
rect 4660 8332 4724 8396
rect 5212 8332 5276 8396
rect 7420 8332 7484 8396
rect 16252 8468 16316 8532
rect 980 8196 1044 8260
rect 7972 8196 8036 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 7972 8060 8036 8124
rect 8340 8196 8404 8260
rect 14596 8392 14660 8396
rect 14596 8336 14610 8392
rect 14610 8336 14660 8392
rect 14596 8332 14660 8336
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 8340 8060 8404 8124
rect 2636 7848 2700 7852
rect 13124 8060 13188 8124
rect 2636 7792 2686 7848
rect 2686 7792 2700 7848
rect 2636 7788 2700 7792
rect 980 7712 1044 7716
rect 9260 7788 9324 7852
rect 10548 7788 10612 7852
rect 980 7656 1030 7712
rect 1030 7656 1044 7712
rect 980 7652 1044 7656
rect 2636 7576 2700 7580
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 2636 7520 2650 7576
rect 2650 7520 2700 7576
rect 2636 7516 2700 7520
rect 5764 7516 5828 7580
rect 1532 7440 1596 7444
rect 1532 7384 1546 7440
rect 1546 7384 1596 7440
rect 1532 7380 1596 7384
rect 10180 7652 10244 7716
rect 10732 7652 10796 7716
rect 11836 7924 11900 7988
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 13492 7924 13556 7988
rect 16988 8060 17052 8124
rect 18460 8060 18524 8124
rect 18276 7924 18340 7988
rect 21220 7924 21284 7988
rect 13124 7788 13188 7852
rect 16988 7788 17052 7852
rect 14780 7712 14844 7716
rect 14780 7656 14830 7712
rect 14830 7656 14844 7712
rect 14780 7652 14844 7656
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 13308 7516 13372 7580
rect 18828 7516 18892 7580
rect 12020 7380 12084 7444
rect 5764 7108 5828 7172
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 4844 6972 4908 7036
rect 7420 6972 7484 7036
rect 7604 6972 7668 7036
rect 8156 6972 8220 7036
rect 9260 7032 9324 7036
rect 9260 6976 9310 7032
rect 9310 6976 9324 7032
rect 9260 6972 9324 6976
rect 9812 7032 9876 7036
rect 16068 7108 16132 7172
rect 17724 7108 17788 7172
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 9812 6976 9862 7032
rect 9862 6976 9876 7032
rect 9812 6972 9876 6976
rect 11100 6972 11164 7036
rect 12388 6972 12452 7036
rect 9444 6836 9508 6900
rect 9996 6836 10060 6900
rect 4108 6700 4172 6764
rect 5212 6760 5276 6764
rect 5212 6704 5226 6760
rect 5226 6704 5276 6760
rect 5212 6700 5276 6704
rect 12388 6760 12452 6764
rect 12388 6704 12438 6760
rect 12438 6704 12452 6760
rect 5580 6428 5644 6492
rect 5028 6156 5092 6220
rect 7052 6564 7116 6628
rect 9628 6564 9692 6628
rect 12388 6700 12452 6704
rect 15148 6700 15212 6764
rect 15332 6564 15396 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 6684 6428 6748 6492
rect 9260 6428 9324 6492
rect 9996 6428 10060 6492
rect 11836 6428 11900 6492
rect 18644 6700 18708 6764
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 7788 6156 7852 6220
rect 19564 6292 19628 6356
rect 20668 6428 20732 6492
rect 21404 6292 21468 6356
rect 19564 6156 19628 6220
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 1900 5884 1964 5948
rect 3188 5748 3252 5812
rect 8524 6020 8588 6084
rect 9628 6020 9692 6084
rect 15148 6080 15212 6084
rect 15148 6024 15162 6080
rect 15162 6024 15212 6080
rect 15148 6020 15212 6024
rect 18092 6020 18156 6084
rect 19932 6020 19996 6084
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 2452 5612 2516 5676
rect 7236 5944 7300 5948
rect 7236 5888 7286 5944
rect 7286 5888 7300 5944
rect 7236 5884 7300 5888
rect 7788 5884 7852 5948
rect 8156 5944 8220 5948
rect 8156 5888 8170 5944
rect 8170 5888 8220 5944
rect 8156 5884 8220 5888
rect 8524 5884 8588 5948
rect 5212 5748 5276 5812
rect 18644 5884 18708 5948
rect 4660 5612 4724 5676
rect 5764 5476 5828 5540
rect 7972 5612 8036 5676
rect 8340 5612 8404 5676
rect 9444 5612 9508 5676
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 12572 5672 12636 5676
rect 12572 5616 12622 5672
rect 12622 5616 12636 5672
rect 12572 5612 12636 5616
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 15148 5476 15212 5540
rect 16988 5476 17052 5540
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 13308 5340 13372 5404
rect 5396 5204 5460 5268
rect 10732 5204 10796 5268
rect 12572 5068 12636 5132
rect 7972 4992 8036 4996
rect 7972 4936 7986 4992
rect 7986 4936 8036 4992
rect 7972 4932 8036 4936
rect 8524 4932 8588 4996
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 980 4796 1044 4860
rect 8340 4856 8404 4860
rect 8340 4800 8354 4856
rect 8354 4800 8404 4856
rect 8340 4796 8404 4800
rect 10364 4856 10428 4860
rect 10364 4800 10414 4856
rect 10414 4800 10428 4856
rect 10364 4796 10428 4800
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 1164 4388 1228 4452
rect 12020 4660 12084 4724
rect 13308 4660 13372 4724
rect 4292 4584 4356 4588
rect 4292 4528 4342 4584
rect 4342 4528 4356 4584
rect 4292 4524 4356 4528
rect 12572 4584 12636 4588
rect 12572 4528 12586 4584
rect 12586 4528 12636 4584
rect 4476 4388 4540 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 5396 4252 5460 4316
rect 6868 4252 6932 4316
rect 7604 4252 7668 4316
rect 12572 4524 12636 4528
rect 14964 4524 15028 4588
rect 18644 4660 18708 4724
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 15332 4176 15396 4180
rect 15332 4120 15346 4176
rect 15346 4120 15396 4176
rect 15332 4116 15396 4120
rect 3924 4040 3988 4044
rect 3924 3984 3938 4040
rect 3938 3984 3988 4040
rect 3924 3980 3988 3984
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8524 3844 8588 3908
rect 15516 3980 15580 4044
rect 15884 3980 15948 4044
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 6868 3708 6932 3772
rect 7420 3708 7484 3772
rect 8156 3708 8220 3772
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 17908 3708 17972 3772
rect 10548 3572 10612 3636
rect 10732 3572 10796 3636
rect 12020 3572 12084 3636
rect 12204 3300 12268 3364
rect 13492 3300 13556 3364
rect 15148 3300 15212 3364
rect 19012 3300 19076 3364
rect 21956 3300 22020 3364
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 2636 3224 2700 3228
rect 2636 3168 2650 3224
rect 2650 3168 2700 3224
rect 2636 3164 2700 3168
rect 5580 3164 5644 3228
rect 11100 3224 11164 3228
rect 11100 3168 11150 3224
rect 11150 3168 11164 3224
rect 11100 3164 11164 3168
rect 12388 3164 12452 3228
rect 5212 3028 5276 3092
rect 7420 3028 7484 3092
rect 12572 3028 12636 3092
rect 1348 2892 1412 2956
rect 1716 2756 1780 2820
rect 7052 2756 7116 2820
rect 9260 2756 9324 2820
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 5948 2620 6012 2684
rect 7236 2620 7300 2684
rect 7604 2680 7668 2684
rect 7604 2624 7654 2680
rect 7654 2624 7668 2680
rect 7604 2620 7668 2624
rect 11836 2620 11900 2684
rect 14596 2680 14660 2684
rect 14596 2624 14646 2680
rect 14646 2624 14660 2680
rect 14596 2620 14660 2624
rect 12756 2484 12820 2548
rect 18276 2484 18340 2548
rect 10732 2348 10796 2412
rect 4660 2212 4724 2276
rect 5764 2272 5828 2276
rect 5764 2216 5778 2272
rect 5778 2216 5828 2272
rect 5764 2212 5828 2216
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 4844 2076 4908 2140
rect 19564 1940 19628 2004
rect 10916 1804 10980 1868
rect 14412 1668 14476 1732
rect 7788 1532 7852 1596
rect 15332 1532 15396 1596
rect 2084 1396 2148 1460
rect 17724 1396 17788 1460
rect 15148 1124 15212 1188
rect 3372 988 3436 1052
rect 13676 988 13740 1052
rect 18460 852 18524 916
<< metal4 >>
rect 16987 22948 17053 22949
rect 16987 22884 16988 22948
rect 17052 22884 17053 22948
rect 16987 22883 17053 22884
rect 979 22812 1045 22813
rect 979 22810 980 22812
rect 62 22750 980 22810
rect 62 6930 122 22750
rect 979 22748 980 22750
rect 1044 22748 1045 22812
rect 979 22747 1045 22748
rect 6867 22676 6933 22677
rect 6867 22612 6868 22676
rect 6932 22612 6933 22676
rect 6867 22611 6933 22612
rect 979 22132 1045 22133
rect 979 22068 980 22132
rect 1044 22068 1045 22132
rect 979 22067 1045 22068
rect 795 13156 861 13157
rect 795 13092 796 13156
rect 860 13092 861 13156
rect 795 13091 861 13092
rect 798 8394 858 13091
rect 982 11930 1042 22067
rect 1531 21588 1597 21589
rect 1531 21524 1532 21588
rect 1596 21524 1597 21588
rect 1531 21523 1597 21524
rect 1163 21316 1229 21317
rect 1163 21252 1164 21316
rect 1228 21252 1229 21316
rect 1163 21251 1229 21252
rect 1166 16590 1226 21251
rect 1166 16530 1410 16590
rect 982 11870 1226 11930
rect 798 8334 1042 8394
rect 982 8261 1042 8334
rect 979 8260 1045 8261
rect 979 8196 980 8260
rect 1044 8196 1045 8260
rect 979 8195 1045 8196
rect 982 7717 1042 8195
rect 979 7716 1045 7717
rect 979 7652 980 7716
rect 1044 7652 1045 7716
rect 979 7651 1045 7652
rect 62 6870 1042 6930
rect 982 4861 1042 6870
rect 979 4860 1045 4861
rect 979 4796 980 4860
rect 1044 4796 1045 4860
rect 979 4795 1045 4796
rect 1166 4453 1226 11870
rect 1163 4452 1229 4453
rect 1163 4388 1164 4452
rect 1228 4388 1229 4452
rect 1163 4387 1229 4388
rect 1350 2957 1410 16530
rect 1534 7445 1594 21523
rect 4659 21452 4725 21453
rect 4659 21388 4660 21452
rect 4724 21388 4725 21452
rect 4659 21387 4725 21388
rect 2635 20908 2701 20909
rect 2635 20844 2636 20908
rect 2700 20844 2701 20908
rect 2635 20843 2701 20844
rect 2638 19277 2698 20843
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3371 19820 3437 19821
rect 3371 19756 3372 19820
rect 3436 19756 3437 19820
rect 3371 19755 3437 19756
rect 2635 19276 2701 19277
rect 2635 19212 2636 19276
rect 2700 19212 2701 19276
rect 2635 19211 2701 19212
rect 2819 18596 2885 18597
rect 2819 18532 2820 18596
rect 2884 18532 2885 18596
rect 2819 18531 2885 18532
rect 2083 18052 2149 18053
rect 2083 17988 2084 18052
rect 2148 17988 2149 18052
rect 2083 17987 2149 17988
rect 1899 16692 1965 16693
rect 1899 16628 1900 16692
rect 1964 16628 1965 16692
rect 1899 16627 1965 16628
rect 1715 10980 1781 10981
rect 1715 10916 1716 10980
rect 1780 10916 1781 10980
rect 1715 10915 1781 10916
rect 1531 7444 1597 7445
rect 1531 7380 1532 7444
rect 1596 7380 1597 7444
rect 1531 7379 1597 7380
rect 1347 2956 1413 2957
rect 1347 2892 1348 2956
rect 1412 2892 1413 2956
rect 1347 2891 1413 2892
rect 1718 2821 1778 10915
rect 1902 5949 1962 16627
rect 2086 9485 2146 17987
rect 2083 9484 2149 9485
rect 2083 9420 2084 9484
rect 2148 9420 2149 9484
rect 2083 9419 2149 9420
rect 2083 9348 2149 9349
rect 2083 9284 2084 9348
rect 2148 9284 2149 9348
rect 2083 9283 2149 9284
rect 1899 5948 1965 5949
rect 1899 5884 1900 5948
rect 1964 5884 1965 5948
rect 1899 5883 1965 5884
rect 1715 2820 1781 2821
rect 1715 2756 1716 2820
rect 1780 2756 1781 2820
rect 1715 2755 1781 2756
rect 2086 1461 2146 9283
rect 2454 8394 2514 13822
rect 2822 12613 2882 18531
rect 3187 17644 3253 17645
rect 3187 17580 3188 17644
rect 3252 17580 3253 17644
rect 3187 17579 3253 17580
rect 3003 14924 3069 14925
rect 3003 14860 3004 14924
rect 3068 14860 3069 14924
rect 3003 14859 3069 14860
rect 2819 12612 2885 12613
rect 2819 12548 2820 12612
rect 2884 12548 2885 12612
rect 2819 12547 2885 12548
rect 2819 12476 2885 12477
rect 2819 12412 2820 12476
rect 2884 12412 2885 12476
rect 2819 12411 2885 12412
rect 2822 12069 2882 12411
rect 3006 12341 3066 14859
rect 3003 12340 3069 12341
rect 3003 12276 3004 12340
rect 3068 12276 3069 12340
rect 3003 12275 3069 12276
rect 2819 12068 2885 12069
rect 2819 12004 2820 12068
rect 2884 12004 2885 12068
rect 2819 12003 2885 12004
rect 2819 11116 2885 11117
rect 2819 11052 2820 11116
rect 2884 11052 2885 11116
rect 2819 11051 2885 11052
rect 2822 8805 2882 11051
rect 3006 9893 3066 12275
rect 3003 9892 3069 9893
rect 3003 9828 3004 9892
rect 3068 9828 3069 9892
rect 3003 9827 3069 9828
rect 2819 8804 2885 8805
rect 2819 8740 2820 8804
rect 2884 8740 2885 8804
rect 2819 8739 2885 8740
rect 2270 8334 2514 8394
rect 2270 6930 2330 8334
rect 2635 7580 2701 7581
rect 2635 7516 2636 7580
rect 2700 7516 2701 7580
rect 2635 7515 2701 7516
rect 2270 6870 2514 6930
rect 2454 5677 2514 6870
rect 2451 5676 2517 5677
rect 2451 5612 2452 5676
rect 2516 5612 2517 5676
rect 2451 5611 2517 5612
rect 2638 3229 2698 7515
rect 3190 5813 3250 17579
rect 3374 13157 3434 19755
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3923 17100 3989 17101
rect 3923 17036 3924 17100
rect 3988 17036 3989 17100
rect 3923 17035 3989 17036
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3371 13156 3437 13157
rect 3371 13092 3372 13156
rect 3436 13092 3437 13156
rect 3371 13091 3437 13092
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3371 11116 3437 11117
rect 3371 11052 3372 11116
rect 3436 11052 3437 11116
rect 3371 11051 3437 11052
rect 3187 5812 3253 5813
rect 3187 5748 3188 5812
rect 3252 5748 3253 5812
rect 3187 5747 3253 5748
rect 2635 3228 2701 3229
rect 2635 3164 2636 3228
rect 2700 3164 2701 3228
rect 2635 3163 2701 3164
rect 2083 1460 2149 1461
rect 2083 1396 2084 1460
rect 2148 1396 2149 1460
rect 2083 1395 2149 1396
rect 3374 1053 3434 11051
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3926 4045 3986 17035
rect 4107 15604 4173 15605
rect 4107 15540 4108 15604
rect 4172 15540 4173 15604
rect 4107 15539 4173 15540
rect 4110 9757 4170 15539
rect 4294 12749 4354 15862
rect 4291 12748 4357 12749
rect 4291 12684 4292 12748
rect 4356 12684 4357 12748
rect 4291 12683 4357 12684
rect 4291 9892 4357 9893
rect 4291 9828 4292 9892
rect 4356 9828 4357 9892
rect 4291 9827 4357 9828
rect 4107 9756 4173 9757
rect 4107 9692 4108 9756
rect 4172 9692 4173 9756
rect 4107 9691 4173 9692
rect 4107 9484 4173 9485
rect 4107 9420 4108 9484
rect 4172 9420 4173 9484
rect 4107 9419 4173 9420
rect 4110 6765 4170 9419
rect 4107 6764 4173 6765
rect 4107 6700 4108 6764
rect 4172 6700 4173 6764
rect 4107 6699 4173 6700
rect 4294 4589 4354 9827
rect 4475 9756 4541 9757
rect 4475 9692 4476 9756
rect 4540 9692 4541 9756
rect 4475 9691 4541 9692
rect 4291 4588 4357 4589
rect 4291 4524 4292 4588
rect 4356 4524 4357 4588
rect 4291 4523 4357 4524
rect 4478 4453 4538 9691
rect 4662 8397 4722 21387
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6683 20228 6749 20229
rect 6683 20164 6684 20228
rect 6748 20164 6749 20228
rect 6683 20163 6749 20164
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 5211 18596 5277 18597
rect 5211 18532 5212 18596
rect 5276 18532 5277 18596
rect 5211 18531 5277 18532
rect 5579 18532 5580 18582
rect 5644 18532 5645 18582
rect 5579 18531 5645 18532
rect 5027 18324 5093 18325
rect 5027 18260 5028 18324
rect 5092 18260 5093 18324
rect 5027 18259 5093 18260
rect 4843 13700 4909 13701
rect 4843 13636 4844 13700
rect 4908 13636 4909 13700
rect 4843 13635 4909 13636
rect 4846 8533 4906 13635
rect 4843 8532 4909 8533
rect 4843 8468 4844 8532
rect 4908 8468 4909 8532
rect 4843 8467 4909 8468
rect 4659 8396 4725 8397
rect 4659 8332 4660 8396
rect 4724 8332 4725 8396
rect 4659 8331 4725 8332
rect 4843 7036 4909 7037
rect 4843 6972 4844 7036
rect 4908 6972 4909 7036
rect 4843 6971 4909 6972
rect 4659 5676 4725 5677
rect 4659 5612 4660 5676
rect 4724 5612 4725 5676
rect 4659 5611 4725 5612
rect 4475 4452 4541 4453
rect 4475 4388 4476 4452
rect 4540 4388 4541 4452
rect 4475 4387 4541 4388
rect 3923 4044 3989 4045
rect 3923 3980 3924 4044
rect 3988 3980 3989 4044
rect 3923 3979 3989 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 4662 2277 4722 5611
rect 4659 2276 4725 2277
rect 4659 2212 4660 2276
rect 4724 2212 4725 2276
rect 4659 2211 4725 2212
rect 4846 2141 4906 6971
rect 5030 6221 5090 18259
rect 5214 15741 5274 18531
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5763 17644 5829 17645
rect 5763 17580 5764 17644
rect 5828 17580 5829 17644
rect 5763 17579 5829 17580
rect 5211 15740 5277 15741
rect 5211 15676 5212 15740
rect 5276 15676 5277 15740
rect 5211 15675 5277 15676
rect 5766 13562 5826 17579
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 5947 16828 6013 16829
rect 5947 16764 5948 16828
rect 6012 16764 6013 16828
rect 5947 16763 6013 16764
rect 5950 13701 6010 16763
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 5947 13700 6013 13701
rect 5947 13636 5948 13700
rect 6012 13636 6013 13700
rect 5947 13635 6013 13636
rect 5766 13502 6010 13562
rect 5395 13020 5461 13021
rect 5395 12956 5396 13020
rect 5460 12956 5461 13020
rect 5395 12955 5461 12956
rect 5211 11932 5277 11933
rect 5211 11868 5212 11932
rect 5276 11868 5277 11932
rect 5211 11867 5277 11868
rect 5214 9757 5274 11867
rect 5398 10434 5458 12955
rect 5582 11930 5642 13142
rect 5582 11870 5826 11930
rect 5398 10374 5642 10434
rect 5395 10300 5461 10301
rect 5395 10236 5396 10300
rect 5460 10236 5461 10300
rect 5395 10235 5461 10236
rect 5211 9756 5277 9757
rect 5211 9692 5212 9756
rect 5276 9692 5277 9756
rect 5211 9691 5277 9692
rect 5211 9484 5277 9485
rect 5211 9420 5212 9484
rect 5276 9420 5277 9484
rect 5211 9419 5277 9420
rect 5214 8533 5274 9419
rect 5211 8532 5277 8533
rect 5211 8468 5212 8532
rect 5276 8468 5277 8532
rect 5211 8467 5277 8468
rect 5211 8396 5277 8397
rect 5211 8332 5212 8396
rect 5276 8332 5277 8396
rect 5211 8331 5277 8332
rect 5214 6765 5274 8331
rect 5211 6764 5277 6765
rect 5211 6700 5212 6764
rect 5276 6700 5277 6764
rect 5211 6699 5277 6700
rect 5027 6220 5093 6221
rect 5027 6156 5028 6220
rect 5092 6156 5093 6220
rect 5027 6155 5093 6156
rect 5211 5812 5277 5813
rect 5211 5748 5212 5812
rect 5276 5748 5277 5812
rect 5211 5747 5277 5748
rect 5214 3093 5274 5747
rect 5398 5269 5458 10235
rect 5582 6493 5642 10374
rect 5766 10301 5826 11870
rect 5950 11661 6010 13502
rect 6142 13088 6462 14112
rect 6686 14109 6746 20163
rect 6870 18461 6930 22611
rect 14411 22404 14477 22405
rect 14411 22340 14412 22404
rect 14476 22340 14477 22404
rect 14411 22339 14477 22340
rect 13675 22132 13741 22133
rect 13675 22068 13676 22132
rect 13740 22068 13741 22132
rect 13675 22067 13741 22068
rect 13491 21316 13557 21317
rect 13491 21252 13492 21316
rect 13556 21252 13557 21316
rect 13491 21251 13557 21252
rect 7419 20228 7485 20229
rect 7419 20164 7420 20228
rect 7484 20164 7485 20228
rect 7419 20163 7485 20164
rect 6867 18460 6933 18461
rect 6867 18396 6868 18460
rect 6932 18396 6933 18460
rect 6867 18395 6933 18396
rect 7422 14245 7482 20163
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 7787 20092 7853 20093
rect 7787 20028 7788 20092
rect 7852 20028 7853 20092
rect 7787 20027 7853 20028
rect 7603 15196 7669 15197
rect 7603 15132 7604 15196
rect 7668 15132 7669 15196
rect 7603 15131 7669 15132
rect 7419 14244 7485 14245
rect 7419 14180 7420 14244
rect 7484 14180 7485 14244
rect 7419 14179 7485 14180
rect 6683 14108 6749 14109
rect 6683 14044 6684 14108
rect 6748 14044 6749 14108
rect 6683 14043 6749 14044
rect 7235 14108 7301 14109
rect 7235 14044 7236 14108
rect 7300 14044 7301 14108
rect 7235 14043 7301 14044
rect 6686 13157 6746 14043
rect 7051 13972 7117 13973
rect 7051 13908 7052 13972
rect 7116 13908 7117 13972
rect 7051 13907 7117 13908
rect 6683 13156 6749 13157
rect 6683 13092 6684 13156
rect 6748 13092 6749 13156
rect 6683 13091 6749 13092
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 5947 11660 6013 11661
rect 5947 11596 5948 11660
rect 6012 11596 6013 11660
rect 5947 11595 6013 11596
rect 6142 10912 6462 11936
rect 6683 11388 6749 11389
rect 6683 11386 6684 11388
rect 6640 11324 6684 11386
rect 6748 11324 6749 11388
rect 6640 11323 6749 11324
rect 6640 10978 6700 11323
rect 6640 10918 6746 10978
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 5947 10844 6013 10845
rect 5947 10780 5948 10844
rect 6012 10780 6013 10844
rect 5947 10779 6013 10780
rect 5763 10300 5829 10301
rect 5763 10236 5764 10300
rect 5828 10236 5829 10300
rect 5763 10235 5829 10236
rect 5763 9756 5829 9757
rect 5763 9692 5764 9756
rect 5828 9692 5829 9756
rect 5763 9691 5829 9692
rect 5766 7581 5826 9691
rect 5763 7580 5829 7581
rect 5763 7516 5764 7580
rect 5828 7516 5829 7580
rect 5763 7515 5829 7516
rect 5763 7172 5829 7173
rect 5763 7108 5764 7172
rect 5828 7108 5829 7172
rect 5763 7107 5829 7108
rect 5579 6492 5645 6493
rect 5579 6428 5580 6492
rect 5644 6428 5645 6492
rect 5579 6427 5645 6428
rect 5766 6218 5826 7107
rect 5582 6158 5826 6218
rect 5395 5268 5461 5269
rect 5395 5204 5396 5268
rect 5460 5204 5461 5268
rect 5395 5203 5461 5204
rect 5398 4317 5458 5203
rect 5395 4316 5461 4317
rect 5395 4252 5396 4316
rect 5460 4252 5461 4316
rect 5395 4251 5461 4252
rect 5582 3229 5642 6158
rect 5763 5540 5829 5541
rect 5763 5476 5764 5540
rect 5828 5476 5829 5540
rect 5763 5475 5829 5476
rect 5579 3228 5645 3229
rect 5579 3164 5580 3228
rect 5644 3164 5645 3228
rect 5579 3163 5645 3164
rect 5211 3092 5277 3093
rect 5211 3028 5212 3092
rect 5276 3028 5277 3092
rect 5211 3027 5277 3028
rect 5766 2277 5826 5475
rect 5950 2685 6010 10779
rect 6142 9824 6462 10848
rect 6686 10437 6746 10918
rect 6683 10436 6749 10437
rect 6683 10372 6684 10436
rect 6748 10372 6749 10436
rect 6683 10371 6749 10372
rect 6545 10300 6611 10301
rect 6545 10236 6546 10300
rect 6610 10298 6611 10300
rect 6610 10238 6746 10298
rect 6610 10236 6611 10238
rect 6545 10235 6611 10236
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6686 6493 6746 10238
rect 7054 9757 7114 13907
rect 7051 9756 7117 9757
rect 7051 9692 7052 9756
rect 7116 9692 7117 9756
rect 7051 9691 7117 9692
rect 6867 9620 6933 9621
rect 6867 9556 6868 9620
rect 6932 9556 6933 9620
rect 6867 9555 6933 9556
rect 6683 6492 6749 6493
rect 6683 6428 6684 6492
rect 6748 6428 6749 6492
rect 6683 6427 6749 6428
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6870 4317 6930 9555
rect 7051 9484 7117 9485
rect 7051 9420 7052 9484
rect 7116 9420 7117 9484
rect 7051 9419 7117 9420
rect 7054 6629 7114 9419
rect 7051 6628 7117 6629
rect 7051 6564 7052 6628
rect 7116 6564 7117 6628
rect 7051 6563 7117 6564
rect 6867 4316 6933 4317
rect 6867 4252 6868 4316
rect 6932 4252 6933 4316
rect 6867 4251 6933 4252
rect 6867 3772 6933 3773
rect 6867 3708 6868 3772
rect 6932 3770 6933 3772
rect 7054 3770 7114 6563
rect 7238 5949 7298 14043
rect 7419 13836 7485 13837
rect 7419 13772 7420 13836
rect 7484 13772 7485 13836
rect 7419 13771 7485 13772
rect 7422 11933 7482 13771
rect 7419 11932 7485 11933
rect 7419 11868 7420 11932
rect 7484 11868 7485 11932
rect 7419 11867 7485 11868
rect 7422 11525 7482 11867
rect 7419 11524 7485 11525
rect 7419 11460 7420 11524
rect 7484 11460 7485 11524
rect 7419 11459 7485 11460
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 7422 8397 7482 11051
rect 7606 10437 7666 15131
rect 7790 10573 7850 20027
rect 7971 19412 8037 19413
rect 7971 19348 7972 19412
rect 8036 19348 8037 19412
rect 7971 19347 8037 19348
rect 7974 18461 8034 19347
rect 8741 19072 9061 20096
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 9627 20092 9693 20093
rect 9627 20028 9628 20092
rect 9692 20028 9693 20092
rect 9627 20027 9693 20028
rect 9443 19412 9509 19413
rect 9443 19348 9444 19412
rect 9508 19348 9509 19412
rect 9443 19347 9509 19348
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 7971 18460 8037 18461
rect 7971 18396 7972 18460
rect 8036 18396 8037 18460
rect 7971 18395 8037 18396
rect 8741 17984 9061 19008
rect 9259 19004 9325 19005
rect 9259 18940 9260 19004
rect 9324 18940 9325 19004
rect 9259 18939 9325 18940
rect 9262 18189 9322 18939
rect 9259 18188 9325 18189
rect 9259 18124 9260 18188
rect 9324 18124 9325 18188
rect 9259 18123 9325 18124
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 7971 17236 8037 17237
rect 7971 17172 7972 17236
rect 8036 17172 8037 17236
rect 7971 17171 8037 17172
rect 7974 11389 8034 17171
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8339 16284 8405 16285
rect 8339 16220 8340 16284
rect 8404 16220 8405 16284
rect 8339 16219 8405 16220
rect 8155 15876 8221 15877
rect 8155 15812 8156 15876
rect 8220 15812 8221 15876
rect 8155 15811 8221 15812
rect 7971 11388 8037 11389
rect 7971 11324 7972 11388
rect 8036 11324 8037 11388
rect 7971 11323 8037 11324
rect 7787 10572 7853 10573
rect 7787 10508 7788 10572
rect 7852 10508 7853 10572
rect 7787 10507 7853 10508
rect 7603 10436 7669 10437
rect 7603 10372 7604 10436
rect 7668 10372 7669 10436
rect 7603 10371 7669 10372
rect 7603 9756 7669 9757
rect 7603 9692 7604 9756
rect 7668 9692 7669 9756
rect 7603 9691 7669 9692
rect 7419 8396 7485 8397
rect 7419 8332 7420 8396
rect 7484 8332 7485 8396
rect 7419 8331 7485 8332
rect 7606 7170 7666 9691
rect 7790 8941 7850 10507
rect 7971 9756 8037 9757
rect 7971 9692 7972 9756
rect 8036 9692 8037 9756
rect 7971 9691 8037 9692
rect 7787 8940 7853 8941
rect 7787 8876 7788 8940
rect 7852 8876 7853 8940
rect 7787 8875 7853 8876
rect 7974 8261 8034 9691
rect 8158 9485 8218 15811
rect 8155 9484 8221 9485
rect 8155 9420 8156 9484
rect 8220 9420 8221 9484
rect 8155 9419 8221 9420
rect 8155 9212 8221 9213
rect 8155 9148 8156 9212
rect 8220 9148 8221 9212
rect 8155 9147 8221 9148
rect 7971 8260 8037 8261
rect 7971 8196 7972 8260
rect 8036 8196 8037 8260
rect 7971 8195 8037 8196
rect 7971 8124 8037 8125
rect 7971 8060 7972 8124
rect 8036 8060 8037 8124
rect 7971 8059 8037 8060
rect 7606 7110 7850 7170
rect 7419 7036 7485 7037
rect 7419 6972 7420 7036
rect 7484 6972 7485 7036
rect 7419 6971 7485 6972
rect 7603 7036 7669 7037
rect 7603 6972 7604 7036
rect 7668 6972 7669 7036
rect 7603 6971 7669 6972
rect 7235 5948 7301 5949
rect 7235 5884 7236 5948
rect 7300 5884 7301 5948
rect 7235 5883 7301 5884
rect 7422 5810 7482 6971
rect 6932 3710 7114 3770
rect 6932 3708 6933 3710
rect 6867 3707 6933 3708
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5947 2684 6013 2685
rect 5947 2620 5948 2684
rect 6012 2620 6013 2684
rect 5947 2619 6013 2620
rect 5763 2276 5829 2277
rect 5763 2212 5764 2276
rect 5828 2212 5829 2276
rect 5763 2211 5829 2212
rect 6142 2208 6462 3232
rect 7054 2821 7114 3710
rect 7238 5750 7482 5810
rect 7051 2820 7117 2821
rect 7051 2756 7052 2820
rect 7116 2756 7117 2820
rect 7051 2755 7117 2756
rect 7238 2685 7298 5750
rect 7606 4450 7666 6971
rect 7790 6221 7850 7110
rect 7787 6220 7853 6221
rect 7787 6156 7788 6220
rect 7852 6156 7853 6220
rect 7787 6155 7853 6156
rect 7787 5948 7853 5949
rect 7787 5884 7788 5948
rect 7852 5884 7853 5948
rect 7787 5883 7853 5884
rect 7422 4390 7666 4450
rect 7422 3773 7482 4390
rect 7603 4316 7669 4317
rect 7603 4252 7604 4316
rect 7668 4252 7669 4316
rect 7603 4251 7669 4252
rect 7419 3772 7485 3773
rect 7419 3708 7420 3772
rect 7484 3708 7485 3772
rect 7419 3707 7485 3708
rect 7419 3092 7485 3093
rect 7419 3028 7420 3092
rect 7484 3028 7485 3092
rect 7419 3027 7485 3028
rect 7235 2684 7301 2685
rect 7235 2620 7236 2684
rect 7300 2620 7301 2684
rect 7235 2619 7301 2620
rect 7422 2546 7482 3027
rect 7606 2685 7666 4251
rect 7603 2684 7669 2685
rect 7603 2620 7604 2684
rect 7668 2620 7669 2684
rect 7603 2619 7669 2620
rect 7790 2546 7850 5883
rect 7974 5677 8034 8059
rect 8158 7037 8218 9147
rect 8342 8261 8402 16219
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 9446 13834 9506 19347
rect 9630 18189 9690 20027
rect 11340 19616 11660 20640
rect 12203 20092 12269 20093
rect 12203 20028 12204 20092
rect 12268 20028 12269 20092
rect 12203 20027 12269 20028
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 9995 19412 10061 19413
rect 9995 19348 9996 19412
rect 10060 19348 10061 19412
rect 9995 19347 10061 19348
rect 10363 19412 10429 19413
rect 10363 19348 10364 19412
rect 10428 19348 10429 19412
rect 10363 19347 10429 19348
rect 9811 18732 9877 18733
rect 9811 18668 9812 18732
rect 9876 18668 9877 18732
rect 9811 18667 9877 18668
rect 9814 18189 9874 18667
rect 9627 18188 9693 18189
rect 9627 18124 9628 18188
rect 9692 18124 9693 18188
rect 9627 18123 9693 18124
rect 9811 18188 9877 18189
rect 9811 18124 9812 18188
rect 9876 18124 9877 18188
rect 9811 18123 9877 18124
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8523 12884 8589 12885
rect 8523 12820 8524 12884
rect 8588 12820 8589 12884
rect 8523 12819 8589 12820
rect 8526 11117 8586 12819
rect 8741 12544 9061 13568
rect 9262 13774 9506 13834
rect 9811 13836 9877 13837
rect 9262 13565 9322 13774
rect 9811 13772 9812 13836
rect 9876 13772 9877 13836
rect 9811 13771 9877 13772
rect 9443 13700 9509 13701
rect 9443 13636 9444 13700
rect 9508 13636 9509 13700
rect 9443 13635 9509 13636
rect 9259 13564 9325 13565
rect 9259 13500 9260 13564
rect 9324 13500 9325 13564
rect 9259 13499 9325 13500
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8523 11116 8589 11117
rect 8523 11052 8524 11116
rect 8588 11052 8589 11116
rect 8523 11051 8589 11052
rect 8741 10368 9061 11392
rect 9259 11388 9325 11389
rect 9259 11324 9260 11388
rect 9324 11324 9325 11388
rect 9259 11323 9325 11324
rect 9262 11117 9322 11323
rect 9259 11116 9325 11117
rect 9259 11052 9260 11116
rect 9324 11052 9325 11116
rect 9259 11051 9325 11052
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8523 9756 8589 9757
rect 8523 9692 8524 9756
rect 8588 9692 8589 9756
rect 8523 9691 8589 9692
rect 8339 8260 8405 8261
rect 8339 8196 8340 8260
rect 8404 8196 8405 8260
rect 8339 8195 8405 8196
rect 8339 8124 8405 8125
rect 8339 8060 8340 8124
rect 8404 8060 8405 8124
rect 8339 8059 8405 8060
rect 8155 7036 8221 7037
rect 8155 6972 8156 7036
rect 8220 6972 8221 7036
rect 8155 6971 8221 6972
rect 8155 5948 8221 5949
rect 8155 5884 8156 5948
rect 8220 5884 8221 5948
rect 8155 5883 8221 5884
rect 7971 5676 8037 5677
rect 7971 5612 7972 5676
rect 8036 5612 8037 5676
rect 7971 5611 8037 5612
rect 8158 5130 8218 5883
rect 8342 5677 8402 8059
rect 8526 6085 8586 9691
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 9262 8669 9322 11051
rect 9446 9757 9506 13635
rect 9627 13292 9693 13293
rect 9627 13228 9628 13292
rect 9692 13228 9693 13292
rect 9627 13227 9693 13228
rect 9630 11250 9690 13227
rect 9814 11389 9874 13771
rect 9998 12205 10058 19347
rect 10179 12612 10245 12613
rect 10179 12548 10180 12612
rect 10244 12548 10245 12612
rect 10179 12547 10245 12548
rect 9995 12204 10061 12205
rect 9995 12140 9996 12204
rect 10060 12140 10061 12204
rect 9995 12139 10061 12140
rect 10182 11930 10242 12547
rect 9998 11870 10242 11930
rect 9811 11388 9877 11389
rect 9811 11324 9812 11388
rect 9876 11324 9877 11388
rect 9811 11323 9877 11324
rect 9630 11190 9874 11250
rect 9443 9756 9509 9757
rect 9443 9692 9444 9756
rect 9508 9692 9509 9756
rect 9443 9691 9509 9692
rect 9627 9756 9693 9757
rect 9627 9692 9628 9756
rect 9692 9692 9693 9756
rect 9627 9691 9693 9692
rect 9259 8668 9325 8669
rect 9259 8604 9260 8668
rect 9324 8604 9325 8668
rect 9259 8603 9325 8604
rect 9443 8668 9509 8669
rect 9443 8604 9444 8668
rect 9508 8604 9509 8668
rect 9443 8603 9509 8604
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 9262 7853 9322 8603
rect 9259 7852 9325 7853
rect 9259 7788 9260 7852
rect 9324 7788 9325 7852
rect 9259 7787 9325 7788
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8523 6084 8589 6085
rect 8523 6020 8524 6084
rect 8588 6020 8589 6084
rect 8523 6019 8589 6020
rect 8741 6016 9061 7040
rect 9259 7036 9325 7037
rect 9259 6972 9260 7036
rect 9324 6972 9325 7036
rect 9259 6971 9325 6972
rect 9262 6626 9322 6971
rect 9446 6901 9506 8603
rect 9443 6900 9509 6901
rect 9443 6836 9444 6900
rect 9508 6836 9509 6900
rect 9443 6835 9509 6836
rect 9630 6629 9690 9691
rect 9814 7037 9874 11190
rect 9811 7036 9877 7037
rect 9811 6972 9812 7036
rect 9876 6972 9877 7036
rect 9811 6971 9877 6972
rect 9998 6901 10058 11870
rect 10179 11252 10245 11253
rect 10179 11188 10180 11252
rect 10244 11188 10245 11252
rect 10179 11187 10245 11188
rect 10182 7717 10242 11187
rect 10366 11117 10426 19347
rect 11099 18596 11165 18597
rect 11099 18532 11100 18596
rect 11164 18532 11165 18596
rect 11099 18531 11165 18532
rect 10915 18052 10981 18053
rect 10915 17988 10916 18052
rect 10980 17988 10981 18052
rect 10915 17987 10981 17988
rect 10731 15876 10797 15877
rect 10731 15812 10732 15876
rect 10796 15812 10797 15876
rect 10731 15811 10797 15812
rect 10363 11116 10429 11117
rect 10363 11052 10364 11116
rect 10428 11052 10429 11116
rect 10363 11051 10429 11052
rect 10734 10658 10794 15811
rect 10918 13701 10978 17987
rect 11102 16829 11162 18531
rect 11340 18528 11660 19552
rect 12019 18596 12085 18597
rect 12019 18532 12020 18596
rect 12084 18532 12085 18596
rect 12019 18531 12085 18532
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11099 16828 11165 16829
rect 11099 16764 11100 16828
rect 11164 16764 11165 16828
rect 11099 16763 11165 16764
rect 11340 16352 11660 17376
rect 11835 16828 11901 16829
rect 11835 16764 11836 16828
rect 11900 16764 11901 16828
rect 11835 16763 11901 16764
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 10915 13700 10981 13701
rect 10915 13636 10916 13700
rect 10980 13636 10981 13700
rect 10915 13635 10981 13636
rect 10918 12069 10978 13635
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11099 12612 11165 12613
rect 11099 12548 11100 12612
rect 11164 12548 11165 12612
rect 11099 12547 11165 12548
rect 10915 12068 10981 12069
rect 10915 12004 10916 12068
rect 10980 12004 10981 12068
rect 10915 12003 10981 12004
rect 10547 9620 10613 9621
rect 10547 9556 10548 9620
rect 10612 9556 10613 9620
rect 10547 9555 10613 9556
rect 10550 8533 10610 9555
rect 10734 9074 10794 10422
rect 10734 9014 10932 9074
rect 10872 8669 10932 9014
rect 10872 8668 10981 8669
rect 10872 8606 10916 8668
rect 10915 8604 10916 8606
rect 10980 8604 10981 8668
rect 10915 8603 10981 8604
rect 10363 8532 10429 8533
rect 10363 8468 10364 8532
rect 10428 8468 10429 8532
rect 10363 8467 10429 8468
rect 10547 8532 10613 8533
rect 10547 8468 10548 8532
rect 10612 8468 10613 8532
rect 10547 8467 10613 8468
rect 10179 7716 10245 7717
rect 10179 7652 10180 7716
rect 10244 7652 10245 7716
rect 10179 7651 10245 7652
rect 9995 6900 10061 6901
rect 9995 6836 9996 6900
rect 10060 6836 10061 6900
rect 9995 6835 10061 6836
rect 10182 6762 10242 7651
rect 9998 6702 10242 6762
rect 9627 6628 9693 6629
rect 9262 6566 9506 6626
rect 9259 6492 9325 6493
rect 9259 6428 9260 6492
rect 9324 6428 9325 6492
rect 9259 6427 9325 6428
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8523 5948 8589 5949
rect 8523 5884 8524 5948
rect 8588 5884 8589 5948
rect 8523 5883 8589 5884
rect 8339 5676 8405 5677
rect 8339 5612 8340 5676
rect 8404 5612 8405 5676
rect 8339 5611 8405 5612
rect 7974 5070 8218 5130
rect 7974 4997 8034 5070
rect 8526 4997 8586 5883
rect 7971 4996 8037 4997
rect 7971 4932 7972 4996
rect 8036 4932 8037 4996
rect 7971 4931 8037 4932
rect 8523 4996 8589 4997
rect 8523 4932 8524 4996
rect 8588 4932 8589 4996
rect 8523 4931 8589 4932
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8339 4860 8405 4861
rect 8339 4796 8340 4860
rect 8404 4796 8405 4860
rect 8339 4795 8405 4796
rect 8342 4450 8402 4795
rect 8342 4390 8586 4450
rect 8526 3909 8586 4390
rect 8523 3908 8589 3909
rect 8523 3844 8524 3908
rect 8588 3844 8589 3908
rect 8523 3843 8589 3844
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7422 2486 7850 2546
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 4843 2140 4909 2141
rect 4843 2076 4844 2140
rect 4908 2076 4909 2140
rect 6142 2128 6462 2144
rect 4843 2075 4909 2076
rect 7790 1597 7850 2486
rect 8741 2752 9061 3776
rect 9262 2821 9322 6427
rect 9446 5677 9506 6566
rect 9627 6564 9628 6628
rect 9692 6564 9693 6628
rect 9998 6578 10058 6702
rect 9627 6563 9693 6564
rect 9630 6085 9690 6563
rect 9627 6084 9693 6085
rect 9627 6020 9628 6084
rect 9692 6020 9693 6084
rect 9627 6019 9693 6020
rect 9443 5676 9509 5677
rect 9443 5612 9444 5676
rect 9508 5612 9509 5676
rect 9443 5611 9509 5612
rect 10366 4861 10426 8467
rect 10547 7852 10613 7853
rect 10547 7788 10548 7852
rect 10612 7788 10613 7852
rect 10547 7787 10613 7788
rect 10363 4860 10429 4861
rect 10363 4796 10364 4860
rect 10428 4796 10429 4860
rect 10363 4795 10429 4796
rect 10550 3637 10610 7787
rect 10731 7716 10797 7717
rect 10731 7652 10732 7716
rect 10796 7652 10797 7716
rect 10731 7651 10797 7652
rect 10734 5269 10794 7651
rect 11102 7578 11162 12547
rect 10918 7518 11162 7578
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11838 11389 11898 16763
rect 12022 15061 12082 18531
rect 12206 16013 12266 20027
rect 13123 19820 13189 19821
rect 13123 19756 13124 19820
rect 13188 19756 13189 19820
rect 13123 19755 13189 19756
rect 12571 18532 12572 18582
rect 12636 18532 12637 18582
rect 12571 18531 12637 18532
rect 12571 16692 12637 16693
rect 12571 16628 12572 16692
rect 12636 16628 12637 16692
rect 12571 16627 12637 16628
rect 12203 16012 12269 16013
rect 12203 15948 12204 16012
rect 12268 15948 12269 16012
rect 12203 15947 12269 15948
rect 12019 15060 12085 15061
rect 12019 14996 12020 15060
rect 12084 14996 12085 15060
rect 12019 14995 12085 14996
rect 12574 14738 12634 16627
rect 12939 16284 13005 16285
rect 12939 16220 12940 16284
rect 13004 16220 13005 16284
rect 12939 16219 13005 16220
rect 12571 14244 12637 14245
rect 12571 14180 12572 14244
rect 12636 14180 12637 14244
rect 12571 14179 12637 14180
rect 12203 13564 12269 13565
rect 12203 13500 12204 13564
rect 12268 13500 12269 13564
rect 12203 13499 12269 13500
rect 12019 11660 12085 11661
rect 12019 11596 12020 11660
rect 12084 11596 12085 11660
rect 12019 11595 12085 11596
rect 11835 11388 11901 11389
rect 11835 11324 11836 11388
rect 11900 11324 11901 11388
rect 11835 11323 11901 11324
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11838 7989 11898 11323
rect 11835 7988 11901 7989
rect 11835 7924 11836 7988
rect 11900 7924 11901 7988
rect 11835 7923 11901 7924
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 10731 5268 10797 5269
rect 10731 5204 10732 5268
rect 10796 5204 10797 5268
rect 10731 5203 10797 5204
rect 10547 3636 10613 3637
rect 10547 3572 10548 3636
rect 10612 3572 10613 3636
rect 10547 3571 10613 3572
rect 10731 3636 10797 3637
rect 10731 3572 10732 3636
rect 10796 3572 10797 3636
rect 10731 3571 10797 3572
rect 9259 2820 9325 2821
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 10734 2413 10794 3571
rect 10731 2412 10797 2413
rect 10731 2348 10732 2412
rect 10796 2348 10797 2412
rect 10731 2347 10797 2348
rect 10918 1869 10978 7518
rect 11099 7036 11165 7037
rect 11099 6972 11100 7036
rect 11164 6972 11165 7036
rect 11099 6971 11165 6972
rect 11102 3229 11162 6971
rect 11340 6560 11660 7584
rect 12022 7445 12082 11595
rect 12206 10845 12266 13499
rect 12387 12748 12453 12749
rect 12387 12684 12388 12748
rect 12452 12684 12453 12748
rect 12387 12683 12453 12684
rect 12203 10844 12269 10845
rect 12203 10780 12204 10844
rect 12268 10780 12269 10844
rect 12203 10779 12269 10780
rect 12206 10573 12266 10779
rect 12203 10572 12269 10573
rect 12203 10508 12204 10572
rect 12268 10508 12269 10572
rect 12203 10507 12269 10508
rect 12203 10164 12269 10165
rect 12203 10100 12204 10164
rect 12268 10100 12269 10164
rect 12203 10099 12269 10100
rect 12019 7444 12085 7445
rect 12019 7380 12020 7444
rect 12084 7380 12085 7444
rect 12019 7379 12085 7380
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11835 6492 11901 6493
rect 11835 6428 11836 6492
rect 11900 6428 11901 6492
rect 11835 6427 11901 6428
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11099 3228 11165 3229
rect 11099 3164 11100 3228
rect 11164 3164 11165 3228
rect 11099 3163 11165 3164
rect 11340 2208 11660 3232
rect 11838 2685 11898 6427
rect 12019 4724 12085 4725
rect 12019 4660 12020 4724
rect 12084 4660 12085 4724
rect 12019 4659 12085 4660
rect 12022 3637 12082 4659
rect 12019 3636 12085 3637
rect 12019 3572 12020 3636
rect 12084 3572 12085 3636
rect 12019 3571 12085 3572
rect 12206 3365 12266 10099
rect 12390 9893 12450 12683
rect 12574 11525 12634 14179
rect 12755 13836 12821 13837
rect 12755 13772 12756 13836
rect 12820 13772 12821 13836
rect 12755 13771 12821 13772
rect 12571 11524 12637 11525
rect 12571 11460 12572 11524
rect 12636 11460 12637 11524
rect 12571 11459 12637 11460
rect 12571 11252 12637 11253
rect 12571 11188 12572 11252
rect 12636 11188 12637 11252
rect 12571 11187 12637 11188
rect 12387 9892 12453 9893
rect 12387 9828 12388 9892
rect 12452 9828 12453 9892
rect 12387 9827 12453 9828
rect 12387 9212 12453 9213
rect 12387 9148 12388 9212
rect 12452 9210 12453 9212
rect 12574 9210 12634 11187
rect 12452 9150 12634 9210
rect 12452 9148 12453 9150
rect 12387 9147 12453 9148
rect 12387 8668 12453 8669
rect 12387 8604 12388 8668
rect 12452 8604 12453 8668
rect 12387 8603 12453 8604
rect 12390 7037 12450 8603
rect 12387 7036 12453 7037
rect 12387 6972 12388 7036
rect 12452 6972 12453 7036
rect 12387 6971 12453 6972
rect 12387 6764 12453 6765
rect 12387 6700 12388 6764
rect 12452 6700 12453 6764
rect 12387 6699 12453 6700
rect 12203 3364 12269 3365
rect 12203 3300 12204 3364
rect 12268 3300 12269 3364
rect 12203 3299 12269 3300
rect 12390 3229 12450 6699
rect 12574 5677 12634 9150
rect 12571 5676 12637 5677
rect 12571 5612 12572 5676
rect 12636 5612 12637 5676
rect 12571 5611 12637 5612
rect 12571 5132 12637 5133
rect 12571 5068 12572 5132
rect 12636 5068 12637 5132
rect 12571 5067 12637 5068
rect 12574 4589 12634 5067
rect 12571 4588 12637 4589
rect 12571 4524 12572 4588
rect 12636 4524 12637 4588
rect 12571 4523 12637 4524
rect 12387 3228 12453 3229
rect 12387 3164 12388 3228
rect 12452 3164 12453 3228
rect 12387 3163 12453 3164
rect 12574 3093 12634 4523
rect 12571 3092 12637 3093
rect 12571 3028 12572 3092
rect 12636 3028 12637 3092
rect 12571 3027 12637 3028
rect 11835 2684 11901 2685
rect 11835 2620 11836 2684
rect 11900 2620 11901 2684
rect 11835 2619 11901 2620
rect 12758 2549 12818 13771
rect 12942 12341 13002 16219
rect 12939 12340 13005 12341
rect 12939 12276 12940 12340
rect 13004 12276 13005 12340
rect 12939 12275 13005 12276
rect 12942 8669 13002 12275
rect 13126 11661 13186 19755
rect 13307 17916 13373 17917
rect 13307 17852 13308 17916
rect 13372 17852 13373 17916
rect 13307 17851 13373 17852
rect 13310 16010 13370 17851
rect 13494 17101 13554 21251
rect 13678 18597 13738 22067
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13675 18596 13741 18597
rect 13675 18532 13676 18596
rect 13740 18532 13741 18596
rect 13675 18531 13741 18532
rect 13939 17984 14259 19008
rect 14414 18733 14474 22339
rect 15331 22268 15397 22269
rect 15331 22204 15332 22268
rect 15396 22204 15397 22268
rect 15331 22203 15397 22204
rect 14595 21996 14661 21997
rect 14595 21932 14596 21996
rect 14660 21932 14661 21996
rect 14595 21931 14661 21932
rect 14598 19141 14658 21931
rect 15147 21724 15213 21725
rect 15147 21660 15148 21724
rect 15212 21660 15213 21724
rect 15147 21659 15213 21660
rect 15150 19277 15210 21659
rect 15334 19277 15394 22203
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 15147 19276 15213 19277
rect 15147 19212 15148 19276
rect 15212 19212 15213 19276
rect 15147 19211 15213 19212
rect 15331 19276 15397 19277
rect 15331 19212 15332 19276
rect 15396 19212 15397 19276
rect 15331 19211 15397 19212
rect 14595 19140 14661 19141
rect 14595 19076 14596 19140
rect 14660 19076 14661 19140
rect 14595 19075 14661 19076
rect 14411 18732 14477 18733
rect 14411 18668 14412 18732
rect 14476 18668 14477 18732
rect 14411 18667 14477 18668
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13491 17100 13557 17101
rect 13491 17036 13492 17100
rect 13556 17036 13557 17100
rect 13491 17035 13557 17036
rect 13939 16896 14259 17920
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 14411 17780 14477 17781
rect 14411 17716 14412 17780
rect 14476 17716 14477 17780
rect 14411 17715 14477 17716
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13310 15950 13554 16010
rect 13307 15196 13373 15197
rect 13307 15132 13308 15196
rect 13372 15132 13373 15196
rect 13307 15131 13373 15132
rect 13123 11660 13189 11661
rect 13123 11596 13124 11660
rect 13188 11596 13189 11660
rect 13123 11595 13189 11596
rect 13123 11252 13189 11253
rect 13123 11188 13124 11252
rect 13188 11188 13189 11252
rect 13123 11187 13189 11188
rect 12939 8668 13005 8669
rect 12939 8604 12940 8668
rect 13004 8604 13005 8668
rect 12939 8603 13005 8604
rect 13126 8125 13186 11187
rect 13310 9213 13370 15131
rect 13494 13565 13554 15950
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13491 13564 13557 13565
rect 13491 13500 13492 13564
rect 13556 13500 13557 13564
rect 13491 13499 13557 13500
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13675 11660 13741 11661
rect 13675 11596 13676 11660
rect 13740 11596 13741 11660
rect 13675 11595 13741 11596
rect 13307 9212 13373 9213
rect 13307 9148 13308 9212
rect 13372 9148 13373 9212
rect 13307 9147 13373 9148
rect 13123 8124 13189 8125
rect 13123 8060 13124 8124
rect 13188 8060 13189 8124
rect 13123 8059 13189 8060
rect 13491 7988 13557 7989
rect 13491 7924 13492 7988
rect 13556 7924 13557 7988
rect 13491 7923 13557 7924
rect 13307 7580 13373 7581
rect 13307 7516 13308 7580
rect 13372 7516 13373 7580
rect 13307 7515 13373 7516
rect 13310 5405 13370 7515
rect 13307 5404 13373 5405
rect 13307 5340 13308 5404
rect 13372 5340 13373 5404
rect 13307 5339 13373 5340
rect 13310 4725 13370 5339
rect 13307 4724 13373 4725
rect 13307 4660 13308 4724
rect 13372 4660 13373 4724
rect 13307 4659 13373 4660
rect 13494 3365 13554 7923
rect 13491 3364 13557 3365
rect 13491 3300 13492 3364
rect 13556 3300 13557 3364
rect 13491 3299 13557 3300
rect 12755 2548 12821 2549
rect 12755 2484 12756 2548
rect 12820 2484 12821 2548
rect 12755 2483 12821 2484
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 10915 1868 10981 1869
rect 10915 1804 10916 1868
rect 10980 1804 10981 1868
rect 10915 1803 10981 1804
rect 7787 1596 7853 1597
rect 7787 1532 7788 1596
rect 7852 1532 7853 1596
rect 7787 1531 7853 1532
rect 13678 1053 13738 11595
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 14414 1733 14474 17715
rect 16538 17440 16858 18464
rect 16990 17917 17050 22883
rect 19931 22540 19997 22541
rect 19931 22476 19932 22540
rect 19996 22476 19997 22540
rect 19931 22475 19997 22476
rect 18091 21860 18157 21861
rect 18091 21796 18092 21860
rect 18156 21796 18157 21860
rect 18091 21795 18157 21796
rect 17907 21452 17973 21453
rect 17907 21388 17908 21452
rect 17972 21388 17973 21452
rect 17907 21387 17973 21388
rect 17171 21044 17237 21045
rect 17171 20980 17172 21044
rect 17236 20980 17237 21044
rect 17171 20979 17237 20980
rect 16987 17916 17053 17917
rect 16987 17852 16988 17916
rect 17052 17852 17053 17916
rect 16987 17851 17053 17852
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 15331 15196 15397 15197
rect 15331 15132 15332 15196
rect 15396 15132 15397 15196
rect 15331 15131 15397 15132
rect 14595 14788 14661 14789
rect 14595 14724 14596 14788
rect 14660 14724 14661 14788
rect 14595 14723 14661 14724
rect 14598 9213 14658 14723
rect 15334 13701 15394 15131
rect 16067 14924 16133 14925
rect 16067 14860 16068 14924
rect 16132 14860 16133 14924
rect 16067 14859 16133 14860
rect 15331 13700 15397 13701
rect 15331 13636 15332 13700
rect 15396 13636 15397 13700
rect 15331 13635 15397 13636
rect 14779 13292 14845 13293
rect 14779 13228 14780 13292
rect 14844 13228 14845 13292
rect 14779 13227 14845 13228
rect 14595 9212 14661 9213
rect 14595 9148 14596 9212
rect 14660 9148 14661 9212
rect 14595 9147 14661 9148
rect 14595 8396 14661 8397
rect 14595 8332 14596 8396
rect 14660 8332 14661 8396
rect 14595 8331 14661 8332
rect 14598 2685 14658 8331
rect 14782 7717 14842 13227
rect 15334 12613 15394 13635
rect 16070 12885 16130 14859
rect 16251 14244 16317 14245
rect 16251 14180 16252 14244
rect 16316 14180 16317 14244
rect 16251 14179 16317 14180
rect 15699 12884 15765 12885
rect 15699 12820 15700 12884
rect 15764 12820 15765 12884
rect 15699 12819 15765 12820
rect 16067 12884 16133 12885
rect 16067 12820 16068 12884
rect 16132 12820 16133 12884
rect 16067 12819 16133 12820
rect 15147 12612 15213 12613
rect 15147 12548 15148 12612
rect 15212 12548 15213 12612
rect 15147 12547 15213 12548
rect 15331 12612 15397 12613
rect 15331 12548 15332 12612
rect 15396 12548 15397 12612
rect 15331 12547 15397 12548
rect 15150 11658 15210 12547
rect 15702 12477 15762 12819
rect 15883 12612 15949 12613
rect 15883 12548 15884 12612
rect 15948 12548 15949 12612
rect 15883 12547 15949 12548
rect 15699 12476 15765 12477
rect 15699 12412 15700 12476
rect 15764 12412 15765 12476
rect 15699 12411 15765 12412
rect 15699 12068 15765 12069
rect 15699 12004 15700 12068
rect 15764 12004 15765 12068
rect 15699 12003 15765 12004
rect 15150 11598 15394 11658
rect 14963 11388 15029 11389
rect 14963 11324 14964 11388
rect 15028 11324 15029 11388
rect 14963 11323 15029 11324
rect 14779 7716 14845 7717
rect 14779 7652 14780 7716
rect 14844 7652 14845 7716
rect 14779 7651 14845 7652
rect 14966 4589 15026 11323
rect 15147 8804 15213 8805
rect 15147 8740 15148 8804
rect 15212 8740 15213 8804
rect 15147 8739 15213 8740
rect 15150 6765 15210 8739
rect 15147 6764 15213 6765
rect 15147 6700 15148 6764
rect 15212 6700 15213 6764
rect 15147 6699 15213 6700
rect 15334 6629 15394 11598
rect 15515 10436 15581 10437
rect 15515 10372 15516 10436
rect 15580 10372 15581 10436
rect 15515 10371 15581 10372
rect 15331 6628 15397 6629
rect 15331 6564 15332 6628
rect 15396 6564 15397 6628
rect 15331 6563 15397 6564
rect 15147 6084 15213 6085
rect 15147 6020 15148 6084
rect 15212 6020 15213 6084
rect 15147 6019 15213 6020
rect 15150 5541 15210 6019
rect 15147 5540 15213 5541
rect 15147 5476 15148 5540
rect 15212 5476 15213 5540
rect 15147 5475 15213 5476
rect 14963 4588 15029 4589
rect 14963 4524 14964 4588
rect 15028 4524 15029 4588
rect 14963 4523 15029 4524
rect 15331 4180 15397 4181
rect 15331 4116 15332 4180
rect 15396 4116 15397 4180
rect 15331 4115 15397 4116
rect 15147 3364 15213 3365
rect 15147 3300 15148 3364
rect 15212 3300 15213 3364
rect 15147 3299 15213 3300
rect 14595 2684 14661 2685
rect 14595 2620 14596 2684
rect 14660 2620 14661 2684
rect 14595 2619 14661 2620
rect 14411 1732 14477 1733
rect 14411 1668 14412 1732
rect 14476 1668 14477 1732
rect 14411 1667 14477 1668
rect 15150 1189 15210 3299
rect 15334 1597 15394 4115
rect 15518 4045 15578 10371
rect 15702 10301 15762 12003
rect 15699 10300 15765 10301
rect 15699 10236 15700 10300
rect 15764 10236 15765 10300
rect 15699 10235 15765 10236
rect 15886 4045 15946 12547
rect 16070 10165 16130 12819
rect 16254 12069 16314 14179
rect 16538 14176 16858 15200
rect 16987 15060 17053 15061
rect 16987 14996 16988 15060
rect 17052 14996 17053 15060
rect 16987 14995 17053 14996
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16251 12068 16317 12069
rect 16251 12004 16252 12068
rect 16316 12004 16317 12068
rect 16251 12003 16317 12004
rect 16067 10164 16133 10165
rect 16067 10100 16068 10164
rect 16132 10100 16133 10164
rect 16067 10099 16133 10100
rect 16067 9756 16133 9757
rect 16067 9692 16068 9756
rect 16132 9692 16133 9756
rect 16067 9691 16133 9692
rect 16070 7173 16130 9691
rect 16254 8533 16314 12003
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16251 8532 16317 8533
rect 16251 8468 16252 8532
rect 16316 8468 16317 8532
rect 16251 8467 16317 8468
rect 16538 7648 16858 8672
rect 16990 8125 17050 14995
rect 17174 14109 17234 20979
rect 17539 18596 17605 18597
rect 17539 18532 17540 18596
rect 17604 18532 17605 18596
rect 17539 18531 17605 18532
rect 17171 14108 17237 14109
rect 17171 14044 17172 14108
rect 17236 14044 17237 14108
rect 17171 14043 17237 14044
rect 17171 13836 17237 13837
rect 17171 13772 17172 13836
rect 17236 13772 17237 13836
rect 17171 13771 17237 13772
rect 16987 8124 17053 8125
rect 16987 8060 16988 8124
rect 17052 8060 17053 8124
rect 16987 8059 17053 8060
rect 16987 7852 17053 7853
rect 16987 7788 16988 7852
rect 17052 7788 17053 7852
rect 16987 7787 17053 7788
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16067 7172 16133 7173
rect 16067 7108 16068 7172
rect 16132 7108 16133 7172
rect 16067 7107 16133 7108
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16990 5541 17050 7787
rect 16987 5540 17053 5541
rect 16987 5476 16988 5540
rect 17052 5476 17053 5540
rect 16987 5475 17053 5476
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 15515 4044 15581 4045
rect 15515 3980 15516 4044
rect 15580 3980 15581 4044
rect 15515 3979 15581 3980
rect 15883 4044 15949 4045
rect 15883 3980 15884 4044
rect 15948 3980 15949 4044
rect 15883 3979 15949 3980
rect 16538 3296 16858 4320
rect 17174 3858 17234 13771
rect 17355 12612 17421 12613
rect 17355 12548 17356 12612
rect 17420 12548 17421 12612
rect 17355 12547 17421 12548
rect 17358 10437 17418 12547
rect 17355 10436 17421 10437
rect 17355 10372 17356 10436
rect 17420 10372 17421 10436
rect 17355 10371 17421 10372
rect 17542 10029 17602 18531
rect 17910 17917 17970 21387
rect 18094 19005 18154 21795
rect 18459 21180 18525 21181
rect 18459 21116 18460 21180
rect 18524 21116 18525 21180
rect 18459 21115 18525 21116
rect 18091 19004 18157 19005
rect 18091 18940 18092 19004
rect 18156 18940 18157 19004
rect 18091 18939 18157 18940
rect 18462 18461 18522 21115
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19563 19412 19629 19413
rect 19563 19348 19564 19412
rect 19628 19348 19629 19412
rect 19563 19347 19629 19348
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 18459 18460 18525 18461
rect 18459 18396 18460 18460
rect 18524 18396 18525 18460
rect 18459 18395 18525 18396
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 17907 17916 17973 17917
rect 17907 17852 17908 17916
rect 17972 17852 17973 17916
rect 17907 17851 17973 17852
rect 19011 17780 19077 17781
rect 19011 17716 19012 17780
rect 19076 17716 19077 17780
rect 19011 17715 19077 17716
rect 18275 15332 18341 15333
rect 18275 15268 18276 15332
rect 18340 15268 18341 15332
rect 18275 15267 18341 15268
rect 18091 13156 18157 13157
rect 18091 13092 18092 13156
rect 18156 13092 18157 13156
rect 18091 13091 18157 13092
rect 17907 12748 17973 12749
rect 17907 12684 17908 12748
rect 17972 12684 17973 12748
rect 17907 12683 17973 12684
rect 17723 12204 17789 12205
rect 17723 12140 17724 12204
rect 17788 12140 17789 12204
rect 17723 12139 17789 12140
rect 17726 11661 17786 12139
rect 17723 11660 17789 11661
rect 17723 11596 17724 11660
rect 17788 11596 17789 11660
rect 17723 11595 17789 11596
rect 17539 10028 17605 10029
rect 17539 9964 17540 10028
rect 17604 9964 17605 10028
rect 17539 9963 17605 9964
rect 17726 7173 17786 11595
rect 17723 7172 17789 7173
rect 17723 7108 17724 7172
rect 17788 7108 17789 7172
rect 17723 7107 17789 7108
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 15331 1596 15397 1597
rect 15331 1532 15332 1596
rect 15396 1532 15397 1596
rect 15331 1531 15397 1532
rect 17726 1461 17786 7107
rect 17910 3773 17970 12683
rect 18094 11117 18154 13091
rect 18278 11389 18338 15267
rect 18459 14244 18525 14245
rect 18459 14180 18460 14244
rect 18524 14180 18525 14244
rect 18459 14179 18525 14180
rect 18275 11388 18341 11389
rect 18275 11324 18276 11388
rect 18340 11324 18341 11388
rect 18275 11323 18341 11324
rect 18091 11116 18157 11117
rect 18091 11052 18092 11116
rect 18156 11052 18157 11116
rect 18091 11051 18157 11052
rect 18094 6085 18154 11051
rect 18462 9213 18522 14179
rect 18643 11932 18709 11933
rect 18643 11868 18644 11932
rect 18708 11868 18709 11932
rect 18643 11867 18709 11868
rect 18459 9212 18525 9213
rect 18459 9148 18460 9212
rect 18524 9148 18525 9212
rect 18459 9147 18525 9148
rect 18462 8125 18522 9147
rect 18459 8124 18525 8125
rect 18459 8060 18460 8124
rect 18524 8060 18525 8124
rect 18459 8059 18525 8060
rect 18275 7988 18341 7989
rect 18275 7924 18276 7988
rect 18340 7924 18341 7988
rect 18275 7923 18341 7924
rect 18091 6084 18157 6085
rect 18091 6020 18092 6084
rect 18156 6020 18157 6084
rect 18091 6019 18157 6020
rect 17907 3772 17973 3773
rect 17907 3708 17908 3772
rect 17972 3708 17973 3772
rect 17907 3707 17973 3708
rect 18278 2549 18338 7923
rect 18275 2548 18341 2549
rect 18275 2484 18276 2548
rect 18340 2484 18341 2548
rect 18275 2483 18341 2484
rect 17723 1460 17789 1461
rect 17723 1396 17724 1460
rect 17788 1396 17789 1460
rect 17723 1395 17789 1396
rect 15147 1188 15213 1189
rect 15147 1124 15148 1188
rect 15212 1124 15213 1188
rect 15147 1123 15213 1124
rect 3371 1052 3437 1053
rect 3371 988 3372 1052
rect 3436 988 3437 1052
rect 3371 987 3437 988
rect 13675 1052 13741 1053
rect 13675 988 13676 1052
rect 13740 988 13741 1052
rect 13675 987 13741 988
rect 18462 917 18522 8059
rect 18646 6765 18706 11867
rect 18827 9892 18893 9893
rect 18827 9828 18828 9892
rect 18892 9828 18893 9892
rect 18827 9827 18893 9828
rect 18830 8941 18890 9827
rect 19014 9621 19074 17715
rect 19137 16896 19457 17920
rect 19566 17237 19626 19347
rect 19934 17781 19994 22475
rect 19931 17780 19997 17781
rect 19931 17716 19932 17780
rect 19996 17716 19997 17780
rect 19931 17715 19997 17716
rect 19563 17236 19629 17237
rect 19563 17172 19564 17236
rect 19628 17172 19629 17236
rect 19563 17171 19629 17172
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19563 13564 19629 13565
rect 19563 13500 19564 13564
rect 19628 13500 19629 13564
rect 19563 13499 19629 13500
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19566 12450 19626 13499
rect 21403 13156 21469 13157
rect 21403 13092 21404 13156
rect 21468 13092 21469 13156
rect 21403 13091 21469 13092
rect 20483 12476 20549 12477
rect 19566 12390 20178 12450
rect 20483 12412 20484 12476
rect 20548 12412 20549 12476
rect 20483 12411 20549 12412
rect 19931 11660 19997 11661
rect 19931 11596 19932 11660
rect 19996 11596 19997 11660
rect 19931 11595 19997 11596
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19563 11116 19629 11117
rect 19563 11052 19564 11116
rect 19628 11052 19629 11116
rect 19563 11051 19629 11052
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19011 9620 19077 9621
rect 19011 9556 19012 9620
rect 19076 9556 19077 9620
rect 19011 9555 19077 9556
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 18827 8940 18893 8941
rect 18827 8876 18828 8940
rect 18892 8876 18893 8940
rect 18827 8875 18893 8876
rect 18830 7581 18890 8875
rect 19011 8668 19077 8669
rect 19011 8604 19012 8668
rect 19076 8604 19077 8668
rect 19011 8603 19077 8604
rect 18827 7580 18893 7581
rect 18827 7516 18828 7580
rect 18892 7516 18893 7580
rect 18827 7515 18893 7516
rect 18643 6764 18709 6765
rect 18643 6700 18644 6764
rect 18708 6700 18709 6764
rect 18643 6699 18709 6700
rect 18646 5949 18706 6699
rect 18643 5948 18709 5949
rect 18643 5884 18644 5948
rect 18708 5884 18709 5948
rect 18643 5883 18709 5884
rect 18646 4725 18706 5883
rect 18643 4724 18709 4725
rect 18643 4660 18644 4724
rect 18708 4660 18709 4724
rect 18643 4659 18709 4660
rect 19014 3365 19074 8603
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19566 6357 19626 11051
rect 19563 6356 19629 6357
rect 19563 6292 19564 6356
rect 19628 6292 19629 6356
rect 19563 6291 19629 6292
rect 19563 6220 19629 6221
rect 19563 6156 19564 6220
rect 19628 6156 19629 6220
rect 19563 6155 19629 6156
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19011 3364 19077 3365
rect 19011 3300 19012 3364
rect 19076 3300 19077 3364
rect 19011 3299 19077 3300
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 19566 2005 19626 6155
rect 19934 6085 19994 11595
rect 20118 9893 20178 12390
rect 20486 10573 20546 12411
rect 21219 12204 21285 12205
rect 21219 12140 21220 12204
rect 21284 12140 21285 12204
rect 21219 12139 21285 12140
rect 20483 10572 20549 10573
rect 20483 10508 20484 10572
rect 20548 10508 20549 10572
rect 20483 10507 20549 10508
rect 20854 10301 20914 10422
rect 20851 10300 20917 10301
rect 20851 10236 20852 10300
rect 20916 10236 20917 10300
rect 20851 10235 20917 10236
rect 20115 9892 20181 9893
rect 20115 9828 20116 9892
rect 20180 9828 20181 9892
rect 20115 9827 20181 9828
rect 21222 7989 21282 12139
rect 21219 7988 21285 7989
rect 21219 7924 21220 7988
rect 21284 7924 21285 7988
rect 21219 7923 21285 7924
rect 21406 6357 21466 13091
rect 21955 11116 22021 11117
rect 21955 11052 21956 11116
rect 22020 11052 22021 11116
rect 21955 11051 22021 11052
rect 21403 6356 21469 6357
rect 21403 6292 21404 6356
rect 21468 6292 21469 6356
rect 21403 6291 21469 6292
rect 19931 6084 19997 6085
rect 19931 6020 19932 6084
rect 19996 6020 19997 6084
rect 19931 6019 19997 6020
rect 21958 3365 22018 11051
rect 21955 3364 22021 3365
rect 21955 3300 21956 3364
rect 22020 3300 22021 3364
rect 21955 3299 22021 3300
rect 19563 2004 19629 2005
rect 19563 1940 19564 2004
rect 19628 1940 19629 2004
rect 19563 1939 19629 1940
rect 18459 916 18525 917
rect 18459 852 18460 916
rect 18524 852 18525 916
rect 18459 851 18525 852
<< via4 >>
rect 2366 13822 2602 14058
rect 2550 7852 2786 7938
rect 2550 7788 2636 7852
rect 2636 7788 2700 7852
rect 2700 7788 2786 7852
rect 2550 7702 2786 7788
rect 4206 15862 4442 16098
rect 5494 18596 5730 18818
rect 5494 18582 5580 18596
rect 5580 18582 5644 18596
rect 5644 18582 5730 18596
rect 5494 13142 5730 13378
rect 6598 11932 6834 12018
rect 6598 11868 6684 11932
rect 6684 11868 6748 11932
rect 6748 11868 6834 11932
rect 6598 11782 6834 11868
rect 10646 10422 10882 10658
rect 8070 3772 8306 3858
rect 8070 3708 8156 3772
rect 8156 3708 8220 3772
rect 8220 3708 8306 3772
rect 8070 3622 8306 3708
rect 9910 6492 10146 6578
rect 9910 6428 9996 6492
rect 9996 6428 10060 6492
rect 10060 6428 10146 6492
rect 9910 6342 10146 6428
rect 12486 18596 12722 18818
rect 12486 18582 12572 18596
rect 12572 18582 12636 18596
rect 12636 18582 12722 18596
rect 12486 14502 12722 14738
rect 13590 13292 13826 13378
rect 13590 13228 13676 13292
rect 13676 13228 13740 13292
rect 13740 13228 13826 13292
rect 13590 13142 13826 13228
rect 13038 7852 13274 7938
rect 13038 7788 13124 7852
rect 13124 7788 13188 7852
rect 13188 7788 13274 7852
rect 13038 7702 13274 7788
rect 17822 16012 18058 16098
rect 17822 15948 17908 16012
rect 17908 15948 17972 16012
rect 17972 15948 18058 16012
rect 17822 15862 18058 15948
rect 17086 3622 17322 3858
rect 19662 11932 19898 12018
rect 19662 11868 19748 11932
rect 19748 11868 19812 11932
rect 19812 11868 19898 11932
rect 19662 11782 19898 11868
rect 20766 10422 21002 10658
rect 20582 6492 20818 6578
rect 20582 6428 20668 6492
rect 20668 6428 20732 6492
rect 20732 6428 20818 6492
rect 20582 6342 20818 6428
<< metal5 >>
rect 5452 18818 12764 18860
rect 5452 18582 5494 18818
rect 5730 18582 12486 18818
rect 12722 18582 12764 18818
rect 5452 18540 12764 18582
rect 4164 16098 18100 16140
rect 4164 15862 4206 16098
rect 4442 15862 17822 16098
rect 18058 15862 18100 16098
rect 4164 15820 18100 15862
rect 12260 14738 12764 14780
rect 12260 14502 12486 14738
rect 12722 14502 12764 14738
rect 12260 14460 12764 14502
rect 12260 14100 12580 14460
rect 2324 14058 12580 14100
rect 2324 13822 2366 14058
rect 2602 13822 12580 14058
rect 2324 13780 12580 13822
rect 5452 13378 13868 13420
rect 5452 13142 5494 13378
rect 5730 13142 13590 13378
rect 13826 13142 13868 13378
rect 5452 13100 13868 13142
rect 6556 12018 19940 12060
rect 6556 11782 6598 12018
rect 6834 11782 19662 12018
rect 19898 11782 19940 12018
rect 6556 11740 19940 11782
rect 10604 10658 21044 10700
rect 10604 10422 10646 10658
rect 10882 10422 20766 10658
rect 21002 10422 21044 10658
rect 10604 10380 21044 10422
rect 2508 7938 13316 7980
rect 2508 7702 2550 7938
rect 2786 7702 13038 7938
rect 13274 7702 13316 7938
rect 2508 7660 13316 7702
rect 9868 6578 20860 6620
rect 9868 6342 9910 6578
rect 10146 6342 20582 6578
rect 20818 6342 20860 6578
rect 9868 6300 20860 6342
rect 8028 3858 17364 3900
rect 8028 3622 8070 3858
rect 8306 3622 17086 3858
rect 17322 3622 17364 3858
rect 8028 3580 17364 3622
use sky130_fd_sc_hd__diode_2  ANTENNA__059__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A
timestamp 1649977179
transform 1 0 5612 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform -1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A
timestamp 1649977179
transform -1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 1932 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform 1 0 15180 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1649977179
transform -1 0 2668 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform 1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform -1 0 13432 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__A
timestamp 1649977179
transform -1 0 21252 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__A
timestamp 1649977179
transform 1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform 1 0 20424 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 21252 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__A
timestamp 1649977179
transform -1 0 21252 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 19780 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform -1 0 21252 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__A
timestamp 1649977179
transform -1 0 20516 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform 1 0 19872 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__A
timestamp 1649977179
transform 1 0 18768 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 19320 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 20332 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A
timestamp 1649977179
transform -1 0 20700 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1649977179
transform 1 0 16284 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A
timestamp 1649977179
transform -1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform 1 0 18768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform 1 0 15548 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform 1 0 16468 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1649977179
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A
timestamp 1649977179
transform 1 0 13432 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__A
timestamp 1649977179
transform -1 0 12604 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__A
timestamp 1649977179
transform 1 0 13248 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A
timestamp 1649977179
transform -1 0 13984 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A
timestamp 1649977179
transform -1 0 14996 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A
timestamp 1649977179
transform -1 0 14444 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A
timestamp 1649977179
transform -1 0 15640 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A
timestamp 1649977179
transform 1 0 14996 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A
timestamp 1649977179
transform 1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1649977179
transform 1 0 16284 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A
timestamp 1649977179
transform 1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A
timestamp 1649977179
transform -1 0 19964 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__A
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_2_N_in_A
timestamp 1649977179
transform -1 0 21252 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 19964 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 18124 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 18676 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 11684 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 10120 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 15640 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 17940 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 14536 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 19136 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 13708 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 11868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 8740 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 10120 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 16928 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 14904 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 15456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13708 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 17756 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 14720 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 15088 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14720 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 13064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 20700 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 20884 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 19964 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 20608 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 21068 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 20792 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 21252 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 21252 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 20332 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 20148 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 20332 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 20516 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 19136 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 20148 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 13984 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 13892 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 10764 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 10580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 12144 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 4508 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 14720 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 15272 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 18492 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 16284 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 17572 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 17388 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 13708 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 14904 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 14720 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 14168 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 3956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 14352 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 11408 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 13800 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 14260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 10120 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 14904 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 15548 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 12880 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 13984 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 14536 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 17664 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1649977179
transform -1 0 17296 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1649977179
transform -1 0 18400 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1649977179
transform -1 0 10212 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1649977179
transform -1 0 8372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1649977179
transform -1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1649977179
transform -1 0 9292 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1649977179
transform -1 0 9200 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1649977179
transform -1 0 8740 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1649977179
transform -1 0 19688 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1649977179
transform -1 0 18216 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1649977179
transform -1 0 19780 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1649977179
transform -1 0 15916 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1649977179
transform -1 0 19228 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1649977179
transform -1 0 19596 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1649977179
transform -1 0 20148 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1649977179
transform -1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1649977179
transform -1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1649977179
transform -1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1649977179
transform -1 0 5428 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1649977179
transform 1 0 9292 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1649977179
transform -1 0 15916 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1649977179
transform -1 0 12696 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1649977179
transform -1 0 11960 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1649977179
transform -1 0 6532 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1649977179
transform -1 0 5428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14904 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 10580 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 13064 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 14076 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13432 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12052 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13524 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 8280 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 6992 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 3772 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 12972 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_4__A0
timestamp 1649977179
transform -1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_5__A1
timestamp 1649977179
transform -1 0 14352 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 9752 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_6__A1
timestamp 1649977179
transform -1 0 8556 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9844 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 10120 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9936 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 11960 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11592 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_33.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11500 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13340 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 16468 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 17020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 13800 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13708 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8464 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A0
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 9108 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8372 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 6532 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 3220 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l2_in_5__A0
timestamp 1649977179
transform -1 0 11868 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 6624 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6440 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5060 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 5244 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 9752 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 9844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7176 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 8372 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 8832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 3680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 13248 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13064 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18400 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 13248 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform -1 0 19780 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 15364 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16652 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17296 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 19412 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 19596 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 19780 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 19412 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A0
timestamp 1649977179
transform -1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 16836 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l2_in_7__A1
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16100 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15732 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17480 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 19412 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 19780 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16836 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 19780 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 19044 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 20148 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 14168 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 16192 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 21252 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 8740 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 6164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 8464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 5980 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 6440 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 9200 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 9384 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A0
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 7912 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A0
timestamp 1649977179
transform -1 0 4232 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 8740 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12144 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_3__A0
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A0
timestamp 1649977179
transform 1 0 5152 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_4__A1
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A0
timestamp 1649977179
transform -1 0 3588 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_5__A1
timestamp 1649977179
transform 1 0 5428 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A0
timestamp 1649977179
transform 1 0 3956 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l2_in_6__A1
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9016 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 11684 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12328 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11408 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 10580 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11592 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13800 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14168 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 13984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11960 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16284 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13984 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_32.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 14352 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output211_A
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output221_A
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67
timestamp 1649977179
transform 1 0 7268 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_151
timestamp 1649977179
transform 1 0 14996 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_23
timestamp 1649977179
transform 1 0 3220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_74
timestamp 1649977179
transform 1 0 7912 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_218
timestamp 1649977179
transform 1 0 21160 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_87
timestamp 1649977179
transform 1 0 9108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_212
timestamp 1649977179
transform 1 0 20608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_150
timestamp 1649977179
transform 1 0 14904 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_85
timestamp 1649977179
transform 1 0 8924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_212
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_104
timestamp 1649977179
transform 1 0 10672 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_222
timestamp 1649977179
transform 1 0 21528 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_99
timestamp 1649977179
transform 1 0 10212 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_153
timestamp 1649977179
transform 1 0 15180 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_172
timestamp 1649977179
transform 1 0 16928 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_161
timestamp 1649977179
transform 1 0 15916 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1649977179
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_98
timestamp 1649977179
transform 1 0 10120 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_102
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_158
timestamp 1649977179
transform 1 0 15640 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_125
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_176
timestamp 1649977179
transform 1 0 17296 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_206
timestamp 1649977179
transform 1 0 20056 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_150
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_196
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_89
timestamp 1649977179
transform 1 0 9292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_186
timestamp 1649977179
transform 1 0 18216 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_222
timestamp 1649977179
transform 1 0 21528 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_36
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_222
timestamp 1649977179
transform 1 0 21528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_7
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_35
timestamp 1649977179
transform 1 0 4324 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_137
timestamp 1649977179
transform 1 0 13708 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_52
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_72
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_91
timestamp 1649977179
transform 1 0 9476 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1649977179
transform 1 0 4048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_60
timestamp 1649977179
transform 1 0 6624 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_89
timestamp 1649977179
transform 1 0 9292 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_128
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 1649977179
transform 1 0 15272 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_205
timestamp 1649977179
transform 1 0 19964 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_17
timestamp 1649977179
transform 1 0 2668 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_41
timestamp 1649977179
transform 1 0 4876 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_46
timestamp 1649977179
transform 1 0 5336 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_126
timestamp 1649977179
transform 1 0 12696 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_163
timestamp 1649977179
transform 1 0 16100 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_42
timestamp 1649977179
transform 1 0 4968 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_126
timestamp 1649977179
transform 1 0 12696 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_145
timestamp 1649977179
transform 1 0 14444 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_148
timestamp 1649977179
transform 1 0 14720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_46
timestamp 1649977179
transform 1 0 5336 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_80
timestamp 1649977179
transform 1 0 8464 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_100
timestamp 1649977179
transform 1 0 10304 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_150
timestamp 1649977179
transform 1 0 14904 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_178
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_33
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_37
timestamp 1649977179
transform 1 0 4508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_17
timestamp 1649977179
transform 1 0 2668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_53
timestamp 1649977179
transform 1 0 5980 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_82
timestamp 1649977179
transform 1 0 8648 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_177
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_209
timestamp 1649977179
transform 1 0 20332 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_17
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_46
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_106
timestamp 1649977179
transform 1 0 10856 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_131
timestamp 1649977179
transform 1 0 13156 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_218
timestamp 1649977179
transform 1 0 21160 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_17
timestamp 1649977179
transform 1 0 2668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_30
timestamp 1649977179
transform 1 0 3864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp 1649977179
transform 1 0 19872 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_11
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1649977179
transform 1 0 9476 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_112
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_182
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_208
timestamp 1649977179
transform 1 0 20240 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_119
timestamp 1649977179
transform 1 0 12052 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_191 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18676 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_74
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_90
timestamp 1649977179
transform 1 0 9384 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_137
timestamp 1649977179
transform 1 0 13708 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_197 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_203
timestamp 1649977179
transform 1 0 19780 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_206
timestamp 1649977179
transform 1 0 20056 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_89
timestamp 1649977179
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_147
timestamp 1649977179
transform 1 0 14628 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_178 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_190
timestamp 1649977179
transform 1 0 18584 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_62
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_122
timestamp 1649977179
transform 1 0 12328 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_166
timestamp 1649977179
transform 1 0 16376 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_172
timestamp 1649977179
transform 1 0 16928 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_184
timestamp 1649977179
transform 1 0 18032 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_40
timestamp 1649977179
transform 1 0 4784 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_134
timestamp 1649977179
transform 1 0 13432 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_158
timestamp 1649977179
transform 1 0 15640 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_180
timestamp 1649977179
transform 1 0 17664 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_188
timestamp 1649977179
transform 1 0 18400 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1649977179
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1649977179
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_151
timestamp 1649977179
transform 1 0 14996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_163
timestamp 1649977179
transform 1 0 16100 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_169
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_173
timestamp 1649977179
transform 1 0 17020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_200
timestamp 1649977179
transform 1 0 19504 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_150
timestamp 1649977179
transform 1 0 14904 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_180
timestamp 1649977179
transform 1 0 17664 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_46
timestamp 1649977179
transform 1 0 5336 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_103
timestamp 1649977179
transform 1 0 10580 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_128
timestamp 1649977179
transform 1 0 12880 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_148
timestamp 1649977179
transform 1 0 14720 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1649977179
transform 1 0 15088 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_158
timestamp 1649977179
transform 1 0 15640 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_162
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_166
timestamp 1649977179
transform 1 0 16376 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_46
timestamp 1649977179
transform 1 0 5336 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  Test_en_N_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1649977179
transform 1 0 4416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform 1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform 1 0 3404 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 2392 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform -1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 1840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 2116 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 2392 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 3312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 4048 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 2116 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 5612 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform -1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 20700 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 21068 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 21068 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 20792 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 21068 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 20884 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 20792 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 20516 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 21068 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 21068 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform 1 0 20516 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 20792 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 20056 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 17664 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 19504 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform 1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform 1 0 14168 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 15272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 16560 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 15548 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 13984 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 9384 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 8832 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1649977179
transform -1 0 11776 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 11224 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 10948 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 12880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1649977179
transform -1 0 13248 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform -1 0 13800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1649977179
transform -1 0 13524 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 14444 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1649977179
transform -1 0 14720 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform -1 0 15088 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1649977179
transform -1 0 14812 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform -1 0 15456 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1649977179
transform -1 0 16744 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1649977179
transform -1 0 16652 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform -1 0 17664 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform -1 0 17020 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_E_FTB01
timestamp 1649977179
transform -1 0 17940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_1_W_FTB01
timestamp 1649977179
transform 1 0 18216 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_E_FTB01
timestamp 1649977179
transform -1 0 18860 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_N_FTB01
timestamp 1649977179
transform -1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_S_FTB01
timestamp 1649977179
transform 1 0 20424 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_2_W_FTB01
timestamp 1649977179
transform 1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_E_FTB01
timestamp 1649977179
transform -1 0 19136 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_N_FTB01
timestamp 1649977179
transform -1 0 18584 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_S_FTB01
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clk_3_W_FTB01
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_2_N_in .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21620 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_2_N_in
timestamp 1649977179
transform 1 0 19780 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_2_N_in
timestamp 1649977179
transform -1 0 19136 0 -1 20672
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 18860 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 4416 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1649977179
transform -1 0 3220 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 5428 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 5704 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input14 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input15
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 2300 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform -1 0 2300 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input23
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 3496 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 21620 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform 1 0 20700 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 20700 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 19228 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 20976 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 21620 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform -1 0 21620 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 20700 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 21620 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 20700 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 18768 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 20424 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 19136 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform 1 0 20700 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 21620 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 19136 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 6256 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform -1 0 9292 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 6256 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input54
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1649977179
transform -1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input56
timestamp 1649977179
transform -1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 11408 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input58
timestamp 1649977179
transform 1 0 11224 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 14996 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform -1 0 6164 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input64
timestamp 1649977179
transform -1 0 7268 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input65
timestamp 1649977179
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input68
timestamp 1649977179
transform -1 0 8280 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input69
timestamp 1649977179
transform -1 0 6808 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input70
timestamp 1649977179
transform 1 0 6532 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform -1 0 3680 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input72
timestamp 1649977179
transform -1 0 9292 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform -1 0 6624 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1649977179
transform -1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1649977179
transform 1 0 8096 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1649977179
transform -1 0 8832 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1649977179
transform -1 0 9936 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input78
timestamp 1649977179
transform -1 0 9844 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1649977179
transform -1 0 10212 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input80
timestamp 1649977179
transform -1 0 10580 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1649977179
transform 1 0 10488 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1649977179
transform -1 0 3680 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1649977179
transform -1 0 5336 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1649977179
transform -1 0 5244 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1649977179
transform 1 0 2392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 4048 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input89
timestamp 1649977179
transform 1 0 4048 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input90
timestamp 1649977179
transform -1 0 6808 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1649977179
transform -1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1649977179
transform -1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1649977179
transform -1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1649977179
transform 1 0 4048 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1649977179
transform -1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1649977179
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input98
timestamp 1649977179
transform 1 0 7268 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input99
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1649977179
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1649977179
transform 1 0 7176 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input102
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input103
timestamp 1649977179
transform 1 0 19504 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input104
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1649977179
transform 1 0 17664 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1649977179
transform -1 0 15548 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input108
timestamp 1649977179
transform -1 0 14444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1649977179
transform -1 0 20700 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input110
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input113
timestamp 1649977179
transform -1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input114
timestamp 1649977179
transform -1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input115
timestamp 1649977179
transform -1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input116
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1649977179
transform 1 0 9200 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input118
timestamp 1649977179
transform 1 0 9476 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input119
timestamp 1649977179
transform -1 0 6256 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input120
timestamp 1649977179
transform -1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 12972 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10948 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11592 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14076 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11960 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11408 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9200 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6440 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9108 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9108 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10120 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11592 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12696 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15272 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13984 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9016 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7820 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1840 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3312 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3220 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3772 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform -1 0 3036 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3680 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 3036 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7820 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 7084 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8464 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5796 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4324 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5704 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5704 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14444 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 15640 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16560 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17664 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19504 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 19228 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 20976 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17664 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17848 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17480 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18124 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17020 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14996 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 17020 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4784 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 6900 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 7912 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8280 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 7176 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 6900 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5336 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5428 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 3312 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_4_
timestamp 1649977179
transform 1 0 2668 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4140 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9476 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11224 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11776 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13800 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14260 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13800 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform -1 0 11592 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_4_
timestamp 1649977179
transform 1 0 13248 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12052 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13708 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_3__294 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13248 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11592 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 13064 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11408 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11408 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14076 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12420 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform -1 0 12144 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_4_
timestamp 1649977179
transform -1 0 12604 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13248 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13156 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l2_in_3__297
timestamp 1649977179
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14168 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13340 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 14168 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 10028 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9200 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 7176 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_6_
timestamp 1649977179
transform -1 0 8556 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_7__299
timestamp 1649977179
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_7_
timestamp 1649977179
transform -1 0 8556 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_2_
timestamp 1649977179
transform -1 0 6256 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_3_
timestamp 1649977179
transform 1 0 7820 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l4_in_1_
timestamp 1649977179
transform -1 0 7728 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l5_in_0_
timestamp 1649977179
transform -1 0 9108 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8004 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9016 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10396 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_3__300
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9844 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11132 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11224 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11776 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform -1 0 11408 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_2_
timestamp 1649977179
transform -1 0 10948 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12604 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_2_
timestamp 1649977179
transform -1 0 11408 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l2_in_3__295
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11960 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12696 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14628 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_3__296
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_3_
timestamp 1649977179
transform -1 0 13800 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12972 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13800 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16192 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10764 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 10120 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_33.mux_l1_in_3__298
timestamp 1649977179
transform 1 0 10212 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l1_in_3_
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11132 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10212 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11316 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16468 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5980 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6072 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_3_
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_4_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10948 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4784 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12328 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform -1 0 8832 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__301
timestamp 1649977179
transform -1 0 4232 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 4600 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 7176 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_4_
timestamp 1649977179
transform 1 0 2760 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 1932 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__304
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform -1 0 2208 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4508 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 4232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4232 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_4_
timestamp 1649977179
transform 1 0 2668 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_5_
timestamp 1649977179
transform 1 0 2852 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_6_
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_7__278
timestamp 1649977179
transform -1 0 4140 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_7_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_2_
timestamp 1649977179
transform 1 0 2116 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_3_
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_1_
timestamp 1649977179
transform 1 0 1840 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l5_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7268 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4508 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__279
timestamp 1649977179
transform 1 0 4232 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4508 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4048 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8004 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8004 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_3_
timestamp 1649977179
transform -1 0 5796 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_3__302
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6808 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5796 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7820 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6992 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7360 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_2_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l2_in_3__303
timestamp 1649977179
transform 1 0 6716 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5520 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5428 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5336 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l1_in_3__277
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_3_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3128 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3956 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15180 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16836 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_3_
timestamp 1649977179
transform -1 0 16100 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_4_
timestamp 1649977179
transform -1 0 15732 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16836 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 16560 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 17664 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__280
timestamp 1649977179
transform -1 0 17296 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 17388 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 19044 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15732 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 18860 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19320 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_3_
timestamp 1649977179
transform -1 0 18492 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_4_
timestamp 1649977179
transform -1 0 15916 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18860 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18492 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__282
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18952 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 19780 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19044 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20424 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 20792 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_4_
timestamp 1649977179
transform -1 0 19136 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_5_
timestamp 1649977179
transform -1 0 18860 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_6_
timestamp 1649977179
transform -1 0 19136 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_7__285
timestamp 1649977179
transform -1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_7_
timestamp 1649977179
transform 1 0 19780 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 20700 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 21344 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_2_
timestamp 1649977179
transform -1 0 20056 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_3_
timestamp 1649977179
transform 1 0 19688 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 20700 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 20056 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l5_in_0_
timestamp 1649977179
transform 1 0 20700 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17572 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 16744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 17388 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__286
timestamp 1649977179
transform -1 0 19136 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18584 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 18308 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 18952 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18492 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_2_
timestamp 1649977179
transform -1 0 18768 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_3__281
timestamp 1649977179
transform -1 0 19872 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18492 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_1_
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l4_in_0_
timestamp 1649977179
transform -1 0 20056 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20240 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 15272 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15824 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15180 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_2_
timestamp 1649977179
transform -1 0 16192 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l2_in_3__283
timestamp 1649977179
transform -1 0 16468 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 16008 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15180 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15364 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l4_in_0_
timestamp 1649977179
transform -1 0 15364 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20240 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16560 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17204 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15640 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_3_
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l1_in_3__284
timestamp 1649977179
transform -1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 16652 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16652 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16744 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5980 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7636 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_3_
timestamp 1649977179
transform 1 0 7176 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6900 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5980 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6900 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 7176 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 7728 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_3__287
timestamp 1649977179
transform -1 0 6900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7728 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 7268 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8280 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8004 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_3_
timestamp 1649977179
transform 1 0 7912 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_4_
timestamp 1649977179
transform 1 0 6900 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6900 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7452 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_3__289
timestamp 1649977179
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_3_
timestamp 1649977179
transform -1 0 6256 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6624 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5428 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 9200 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4232 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3680 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 3956 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2944 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_4_
timestamp 1649977179
transform 1 0 3956 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_5_
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_6_
timestamp 1649977179
transform 1 0 2760 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_7__292
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_7_
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3128 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_2_
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_3_
timestamp 1649977179
transform 1 0 2576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l4_in_1_
timestamp 1649977179
transform -1 0 2576 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l5_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4048 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5152 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9936 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_2_
timestamp 1649977179
transform -1 0 10028 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l2_in_3__293
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_3_
timestamp 1649977179
transform -1 0 10396 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_0_
timestamp 1649977179
transform -1 0 8832 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9384 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8280 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10580 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_2_
timestamp 1649977179
transform -1 0 11040 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_3__288
timestamp 1649977179
transform 1 0 11224 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10580 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10488 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11316 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12052 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13248 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12144 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 12328 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_1_
timestamp 1649977179
transform -1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_2_
timestamp 1649977179
transform -1 0 13156 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l2_in_3__290
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_3_
timestamp 1649977179
transform 1 0 13156 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l3_in_1_
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13524 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13800 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14628 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16284 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_32.mux_l1_in_3__291
timestamp 1649977179
transform 1 0 15824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l1_in_3_
timestamp 1649977179
transform -1 0 15364 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15824 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_32.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 16008 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform -1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform -1 0 2116 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform -1 0 2116 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform -1 0 2116 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform -1 0 2116 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform -1 0 2116 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform -1 0 2116 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output151
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output152
timestamp 1649977179
transform -1 0 19412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output153
timestamp 1649977179
transform -1 0 19136 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output154
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output155
timestamp 1649977179
transform 1 0 21252 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output156
timestamp 1649977179
transform 1 0 21252 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output157
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output158
timestamp 1649977179
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output159
timestamp 1649977179
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output160
timestamp 1649977179
transform 1 0 21252 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output161
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output162
timestamp 1649977179
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output163
timestamp 1649977179
transform -1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output164
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output165
timestamp 1649977179
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output166
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output167
timestamp 1649977179
transform 1 0 16928 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output168
timestamp 1649977179
transform 1 0 20148 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output169
timestamp 1649977179
transform 1 0 20056 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1649977179
transform 1 0 20424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1649977179
transform 1 0 20792 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1649977179
transform 1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1649977179
transform -1 0 13892 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1649977179
transform -1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1649977179
transform -1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1649977179
transform -1 0 17020 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1649977179
transform -1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1649977179
transform 1 0 10120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1649977179
transform 1 0 17020 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1649977179
transform 1 0 17756 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1649977179
transform -1 0 18492 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1649977179
transform 1 0 12052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1649977179
transform 1 0 11776 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1649977179
transform 1 0 12144 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1649977179
transform 1 0 12880 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1649977179
transform 1 0 13248 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1649977179
transform 1 0 13616 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1649977179
transform 1 0 20700 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1649977179
transform -1 0 2484 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1649977179
transform -1 0 16560 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1649977179
transform -1 0 2116 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1649977179
transform -1 0 15824 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1649977179
transform -1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1649977179
transform -1 0 19964 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1649977179
transform -1 0 2484 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output215
timestamp 1649977179
transform -1 0 16560 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output216
timestamp 1649977179
transform -1 0 21252 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output217
timestamp 1649977179
transform -1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output218
timestamp 1649977179
transform 1 0 9016 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1649977179
transform -1 0 20332 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1649977179
transform -1 0 15456 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1649977179
transform -1 0 2852 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_0_FTB00
timestamp 1649977179
transform 1 0 18952 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_E_FTB01
timestamp 1649977179
transform 1 0 19872 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_1_W_FTB01
timestamp 1649977179
transform 1 0 16100 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_E_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_N_FTB01
timestamp 1649977179
transform 1 0 20700 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_S_FTB01
timestamp 1649977179
transform 1 0 20700 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_2_W_FTB01
timestamp 1649977179
transform -1 0 19780 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_E_FTB01
timestamp 1649977179
transform -1 0 18308 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_N_FTB01
timestamp 1649977179
transform 1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_S_FTB01
timestamp 1649977179
transform 1 0 18860 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  prog_clk_3_W_FTB01
timestamp 1649977179
transform 1 0 18492 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater223
timestamp 1649977179
transform 1 0 4508 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater224
timestamp 1649977179
transform 1 0 5060 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater225
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater226
timestamp 1649977179
transform -1 0 9292 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater227
timestamp 1649977179
transform 1 0 20148 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater228
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater229
timestamp 1649977179
transform -1 0 17664 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater230
timestamp 1649977179
transform 1 0 17296 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater231
timestamp 1649977179
transform -1 0 3864 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater232
timestamp 1649977179
transform -1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater233
timestamp 1649977179
transform 1 0 4232 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater234
timestamp 1649977179
transform 1 0 6072 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater235
timestamp 1649977179
transform -1 0 11960 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater236
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater237
timestamp 1649977179
transform -1 0 14352 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater238
timestamp 1649977179
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater239
timestamp 1649977179
transform 1 0 2760 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater240
timestamp 1649977179
transform -1 0 4508 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater241
timestamp 1649977179
transform 1 0 3956 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater242
timestamp 1649977179
transform 1 0 7728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater243
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater244
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater245
timestamp 1649977179
transform 1 0 6716 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater246
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater247
timestamp 1649977179
transform -1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater248
timestamp 1649977179
transform 1 0 6716 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater249
timestamp 1649977179
transform 1 0 9200 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater250
timestamp 1649977179
transform 1 0 10304 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater251
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater252
timestamp 1649977179
transform -1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater253
timestamp 1649977179
transform 1 0 3680 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater254
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater255
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater256
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater257
timestamp 1649977179
transform 1 0 12604 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater258
timestamp 1649977179
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater259
timestamp 1649977179
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater260
timestamp 1649977179
transform 1 0 13248 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater261
timestamp 1649977179
transform 1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater262
timestamp 1649977179
transform 1 0 12420 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater263
timestamp 1649977179
transform 1 0 14720 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater264
timestamp 1649977179
transform 1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater265
timestamp 1649977179
transform 1 0 16652 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater266
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater267
timestamp 1649977179
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater268
timestamp 1649977179
transform -1 0 14812 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater269
timestamp 1649977179
transform 1 0 14260 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater270
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater271
timestamp 1649977179
transform -1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater272
timestamp 1649977179
transform -1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater273
timestamp 1649977179
transform -1 0 17848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater274
timestamp 1649977179
transform 1 0 19320 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater275
timestamp 1649977179
transform -1 0 17848 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  repeater276
timestamp 1649977179
transform 1 0 17296 0 1 15232
box -38 -48 314 592
<< labels >>
rlabel metal2 s 18602 22200 18658 23000 6 Test_en_N_out
port 0 nsew signal tristate
rlabel metal2 s 21086 0 21142 800 6 Test_en_S_in
port 1 nsew signal input
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 3 nsew power input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 4 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 5 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 6 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 bottom_left_grid_pin_45_
port 7 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 bottom_left_grid_pin_46_
port 8 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 bottom_left_grid_pin_47_
port 9 nsew signal input
rlabel metal2 s 2686 0 2742 800 6 bottom_left_grid_pin_48_
port 10 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 bottom_left_grid_pin_49_
port 11 nsew signal input
rlabel metal2 s 3514 0 3570 800 6 ccff_head
port 12 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 ccff_tail
port 13 nsew signal tristate
rlabel metal3 s 0 3544 800 3664 6 chanx_left_in[0]
port 14 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 chanx_left_in[10]
port 15 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 chanx_left_in[11]
port 16 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[12]
port 17 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[13]
port 18 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[14]
port 19 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 chanx_left_in[15]
port 20 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[16]
port 21 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 chanx_left_in[17]
port 22 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 chanx_left_in[18]
port 23 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 chanx_left_in[19]
port 24 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 chanx_left_in[1]
port 25 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[2]
port 26 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[3]
port 27 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[4]
port 28 nsew signal input
rlabel metal3 s 0 5584 800 5704 6 chanx_left_in[5]
port 29 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 chanx_left_in[6]
port 30 nsew signal input
rlabel metal3 s 0 6400 800 6520 6 chanx_left_in[7]
port 31 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 chanx_left_in[8]
port 32 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 chanx_left_in[9]
port 33 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 chanx_left_out[0]
port 34 nsew signal tristate
rlabel metal3 s 0 16192 800 16312 6 chanx_left_out[10]
port 35 nsew signal tristate
rlabel metal3 s 0 16736 800 16856 6 chanx_left_out[11]
port 36 nsew signal tristate
rlabel metal3 s 0 17144 800 17264 6 chanx_left_out[12]
port 37 nsew signal tristate
rlabel metal3 s 0 17552 800 17672 6 chanx_left_out[13]
port 38 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[14]
port 39 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[15]
port 40 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[16]
port 41 nsew signal tristate
rlabel metal3 s 0 19184 800 19304 6 chanx_left_out[17]
port 42 nsew signal tristate
rlabel metal3 s 0 19592 800 19712 6 chanx_left_out[18]
port 43 nsew signal tristate
rlabel metal3 s 0 20136 800 20256 6 chanx_left_out[19]
port 44 nsew signal tristate
rlabel metal3 s 0 12384 800 12504 6 chanx_left_out[1]
port 45 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 chanx_left_out[2]
port 46 nsew signal tristate
rlabel metal3 s 0 13336 800 13456 6 chanx_left_out[3]
port 47 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[4]
port 48 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[5]
port 49 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[6]
port 50 nsew signal tristate
rlabel metal3 s 0 14968 800 15088 6 chanx_left_out[7]
port 51 nsew signal tristate
rlabel metal3 s 0 15376 800 15496 6 chanx_left_out[8]
port 52 nsew signal tristate
rlabel metal3 s 0 15784 800 15904 6 chanx_left_out[9]
port 53 nsew signal tristate
rlabel metal3 s 22200 3544 23000 3664 6 chanx_right_in[0]
port 54 nsew signal input
rlabel metal3 s 22200 7760 23000 7880 6 chanx_right_in[10]
port 55 nsew signal input
rlabel metal3 s 22200 8168 23000 8288 6 chanx_right_in[11]
port 56 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[12]
port 57 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[13]
port 58 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[14]
port 59 nsew signal input
rlabel metal3 s 22200 9800 23000 9920 6 chanx_right_in[15]
port 60 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[16]
port 61 nsew signal input
rlabel metal3 s 22200 10752 23000 10872 6 chanx_right_in[17]
port 62 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[18]
port 63 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[19]
port 64 nsew signal input
rlabel metal3 s 22200 3952 23000 4072 6 chanx_right_in[1]
port 65 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[2]
port 66 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[3]
port 67 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[4]
port 68 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[5]
port 69 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[6]
port 70 nsew signal input
rlabel metal3 s 22200 6400 23000 6520 6 chanx_right_in[7]
port 71 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[8]
port 72 nsew signal input
rlabel metal3 s 22200 7352 23000 7472 6 chanx_right_in[9]
port 73 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_out[0]
port 74 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[10]
port 75 nsew signal tristate
rlabel metal3 s 22200 16736 23000 16856 6 chanx_right_out[11]
port 76 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[12]
port 77 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[13]
port 78 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[14]
port 79 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[15]
port 80 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[16]
port 81 nsew signal tristate
rlabel metal3 s 22200 19184 23000 19304 6 chanx_right_out[17]
port 82 nsew signal tristate
rlabel metal3 s 22200 19592 23000 19712 6 chanx_right_out[18]
port 83 nsew signal tristate
rlabel metal3 s 22200 20136 23000 20256 6 chanx_right_out[19]
port 84 nsew signal tristate
rlabel metal3 s 22200 12384 23000 12504 6 chanx_right_out[1]
port 85 nsew signal tristate
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_out[2]
port 86 nsew signal tristate
rlabel metal3 s 22200 13336 23000 13456 6 chanx_right_out[3]
port 87 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[4]
port 88 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[5]
port 89 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[6]
port 90 nsew signal tristate
rlabel metal3 s 22200 14968 23000 15088 6 chanx_right_out[7]
port 91 nsew signal tristate
rlabel metal3 s 22200 15376 23000 15496 6 chanx_right_out[8]
port 92 nsew signal tristate
rlabel metal3 s 22200 15784 23000 15904 6 chanx_right_out[9]
port 93 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_in[0]
port 94 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 chany_bottom_in[10]
port 95 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[11]
port 96 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[12]
port 97 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[13]
port 98 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[14]
port 99 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[15]
port 100 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[16]
port 101 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 102 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 103 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 chany_bottom_in[19]
port 104 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_in[1]
port 105 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_in[2]
port 106 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[3]
port 107 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[4]
port 108 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[5]
port 109 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_in[6]
port 110 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[7]
port 111 nsew signal input
rlabel metal2 s 7654 0 7710 800 6 chany_bottom_in[8]
port 112 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_in[9]
port 113 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[0]
port 114 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[10]
port 115 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[11]
port 116 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[12]
port 117 nsew signal tristate
rlabel metal2 s 18142 0 18198 800 6 chany_bottom_out[13]
port 118 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[14]
port 119 nsew signal tristate
rlabel metal2 s 18970 0 19026 800 6 chany_bottom_out[15]
port 120 nsew signal tristate
rlabel metal2 s 19430 0 19486 800 6 chany_bottom_out[16]
port 121 nsew signal tristate
rlabel metal2 s 19798 0 19854 800 6 chany_bottom_out[17]
port 122 nsew signal tristate
rlabel metal2 s 20258 0 20314 800 6 chany_bottom_out[18]
port 123 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 chany_bottom_out[19]
port 124 nsew signal tristate
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_out[1]
port 125 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_out[2]
port 126 nsew signal tristate
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_out[3]
port 127 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[4]
port 128 nsew signal tristate
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_out[5]
port 129 nsew signal tristate
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_out[6]
port 130 nsew signal tristate
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_out[7]
port 131 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[8]
port 132 nsew signal tristate
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_out[9]
port 133 nsew signal tristate
rlabel metal2 s 3238 22200 3294 23000 6 chany_top_in[0]
port 134 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[10]
port 135 nsew signal input
rlabel metal2 s 7470 22200 7526 23000 6 chany_top_in[11]
port 136 nsew signal input
rlabel metal2 s 7838 22200 7894 23000 6 chany_top_in[12]
port 137 nsew signal input
rlabel metal2 s 8206 22200 8262 23000 6 chany_top_in[13]
port 138 nsew signal input
rlabel metal2 s 8574 22200 8630 23000 6 chany_top_in[14]
port 139 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[15]
port 140 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[16]
port 141 nsew signal input
rlabel metal2 s 9770 22200 9826 23000 6 chany_top_in[17]
port 142 nsew signal input
rlabel metal2 s 10138 22200 10194 23000 6 chany_top_in[18]
port 143 nsew signal input
rlabel metal2 s 10506 22200 10562 23000 6 chany_top_in[19]
port 144 nsew signal input
rlabel metal2 s 3606 22200 3662 23000 6 chany_top_in[1]
port 145 nsew signal input
rlabel metal2 s 3974 22200 4030 23000 6 chany_top_in[2]
port 146 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[3]
port 147 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[4]
port 148 nsew signal input
rlabel metal2 s 5170 22200 5226 23000 6 chany_top_in[5]
port 149 nsew signal input
rlabel metal2 s 5538 22200 5594 23000 6 chany_top_in[6]
port 150 nsew signal input
rlabel metal2 s 5906 22200 5962 23000 6 chany_top_in[7]
port 151 nsew signal input
rlabel metal2 s 6274 22200 6330 23000 6 chany_top_in[8]
port 152 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[9]
port 153 nsew signal input
rlabel metal2 s 10874 22200 10930 23000 6 chany_top_out[0]
port 154 nsew signal tristate
rlabel metal2 s 14738 22200 14794 23000 6 chany_top_out[10]
port 155 nsew signal tristate
rlabel metal2 s 15106 22200 15162 23000 6 chany_top_out[11]
port 156 nsew signal tristate
rlabel metal2 s 15474 22200 15530 23000 6 chany_top_out[12]
port 157 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[13]
port 158 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[14]
port 159 nsew signal tristate
rlabel metal2 s 16670 22200 16726 23000 6 chany_top_out[15]
port 160 nsew signal tristate
rlabel metal2 s 17038 22200 17094 23000 6 chany_top_out[16]
port 161 nsew signal tristate
rlabel metal2 s 17406 22200 17462 23000 6 chany_top_out[17]
port 162 nsew signal tristate
rlabel metal2 s 17774 22200 17830 23000 6 chany_top_out[18]
port 163 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[19]
port 164 nsew signal tristate
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_out[1]
port 165 nsew signal tristate
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_out[2]
port 166 nsew signal tristate
rlabel metal2 s 12070 22200 12126 23000 6 chany_top_out[3]
port 167 nsew signal tristate
rlabel metal2 s 12438 22200 12494 23000 6 chany_top_out[4]
port 168 nsew signal tristate
rlabel metal2 s 12806 22200 12862 23000 6 chany_top_out[5]
port 169 nsew signal tristate
rlabel metal2 s 13174 22200 13230 23000 6 chany_top_out[6]
port 170 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[7]
port 171 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[8]
port 172 nsew signal tristate
rlabel metal2 s 14370 22200 14426 23000 6 chany_top_out[9]
port 173 nsew signal tristate
rlabel metal3 s 22200 20544 23000 20664 6 clk_1_E_out
port 174 nsew signal tristate
rlabel metal2 s 18970 22200 19026 23000 6 clk_1_N_in
port 175 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 clk_1_W_out
port 176 nsew signal tristate
rlabel metal3 s 22200 20952 23000 21072 6 clk_2_E_out
port 177 nsew signal tristate
rlabel metal2 s 19338 22200 19394 23000 6 clk_2_N_in
port 178 nsew signal input
rlabel metal2 s 21638 22200 21694 23000 6 clk_2_N_out
port 179 nsew signal tristate
rlabel metal2 s 21454 0 21510 800 6 clk_2_S_out
port 180 nsew signal tristate
rlabel metal3 s 0 20952 800 21072 6 clk_2_W_out
port 181 nsew signal tristate
rlabel metal3 s 22200 21360 23000 21480 6 clk_3_E_out
port 182 nsew signal tristate
rlabel metal2 s 19706 22200 19762 23000 6 clk_3_N_in
port 183 nsew signal input
rlabel metal2 s 22006 22200 22062 23000 6 clk_3_N_out
port 184 nsew signal tristate
rlabel metal2 s 21914 0 21970 800 6 clk_3_S_out
port 185 nsew signal tristate
rlabel metal3 s 0 21360 800 21480 6 clk_3_W_out
port 186 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 187 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 188 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 189 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 left_bottom_grid_pin_37_
port 190 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 left_bottom_grid_pin_38_
port 191 nsew signal input
rlabel metal3 s 0 2184 800 2304 6 left_bottom_grid_pin_39_
port 192 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 left_bottom_grid_pin_40_
port 193 nsew signal input
rlabel metal3 s 0 3000 800 3120 6 left_bottom_grid_pin_41_
port 194 nsew signal input
rlabel metal2 s 20074 22200 20130 23000 6 prog_clk_0_N_in
port 195 nsew signal input
rlabel metal3 s 22200 21768 23000 21888 6 prog_clk_1_E_out
port 196 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 prog_clk_1_N_in
port 197 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 prog_clk_1_W_out
port 198 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_2_E_out
port 199 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 prog_clk_2_N_in
port 200 nsew signal input
rlabel metal2 s 22374 22200 22430 23000 6 prog_clk_2_N_out
port 201 nsew signal tristate
rlabel metal2 s 22282 0 22338 800 6 prog_clk_2_S_out
port 202 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 prog_clk_2_W_out
port 203 nsew signal tristate
rlabel metal3 s 22200 22584 23000 22704 6 prog_clk_3_E_out
port 204 nsew signal tristate
rlabel metal2 s 21270 22200 21326 23000 6 prog_clk_3_N_in
port 205 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 prog_clk_3_N_out
port 206 nsew signal tristate
rlabel metal2 s 22742 0 22798 800 6 prog_clk_3_S_out
port 207 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 prog_clk_3_W_out
port 208 nsew signal tristate
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 209 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 210 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 211 nsew signal input
rlabel metal3 s 22200 1368 23000 1488 6 right_bottom_grid_pin_37_
port 212 nsew signal input
rlabel metal3 s 22200 1776 23000 1896 6 right_bottom_grid_pin_38_
port 213 nsew signal input
rlabel metal3 s 22200 2184 23000 2304 6 right_bottom_grid_pin_39_
port 214 nsew signal input
rlabel metal3 s 22200 2592 23000 2712 6 right_bottom_grid_pin_40_
port 215 nsew signal input
rlabel metal3 s 22200 3000 23000 3120 6 right_bottom_grid_pin_41_
port 216 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 217 nsew signal input
rlabel metal2 s 570 22200 626 23000 6 top_left_grid_pin_43_
port 218 nsew signal input
rlabel metal2 s 938 22200 994 23000 6 top_left_grid_pin_44_
port 219 nsew signal input
rlabel metal2 s 1306 22200 1362 23000 6 top_left_grid_pin_45_
port 220 nsew signal input
rlabel metal2 s 1674 22200 1730 23000 6 top_left_grid_pin_46_
port 221 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_47_
port 222 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_48_
port 223 nsew signal input
rlabel metal2 s 2870 22200 2926 23000 6 top_left_grid_pin_49_
port 224 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
