module sb_2__2_ (SC_IN_BOT,
    SC_OUT_BOT,
    VGND,
    VPWR,
    bottom_left_grid_pin_42_,
    bottom_left_grid_pin_43_,
    bottom_left_grid_pin_44_,
    bottom_left_grid_pin_45_,
    bottom_left_grid_pin_46_,
    bottom_left_grid_pin_47_,
    bottom_left_grid_pin_48_,
    bottom_left_grid_pin_49_,
    bottom_right_grid_pin_1_,
    ccff_head,
    ccff_tail,
    left_bottom_grid_pin_34_,
    left_bottom_grid_pin_35_,
    left_bottom_grid_pin_36_,
    left_bottom_grid_pin_37_,
    left_bottom_grid_pin_38_,
    left_bottom_grid_pin_39_,
    left_bottom_grid_pin_40_,
    left_bottom_grid_pin_41_,
    left_top_grid_pin_1_,
    prog_clk_0_S_in,
    chanx_left_in,
    chanx_left_out,
    chany_bottom_in,
    chany_bottom_out);
 inout SC_IN_BOT;
 output SC_OUT_BOT;
 inout VGND;
 inout VPWR;
 inout bottom_left_grid_pin_42_;
 inout bottom_left_grid_pin_43_;
 inout bottom_left_grid_pin_44_;
 inout bottom_left_grid_pin_45_;
 inout bottom_left_grid_pin_46_;
 inout bottom_left_grid_pin_47_;
 inout bottom_left_grid_pin_48_;
 inout bottom_left_grid_pin_49_;
 inout bottom_right_grid_pin_1_;
 inout ccff_head;
 output ccff_tail;
 inout left_bottom_grid_pin_34_;
 inout left_bottom_grid_pin_35_;
 inout left_bottom_grid_pin_36_;
 inout left_bottom_grid_pin_37_;
 inout left_bottom_grid_pin_38_;
 inout left_bottom_grid_pin_39_;
 inout left_bottom_grid_pin_40_;
 inout left_bottom_grid_pin_41_;
 inout left_top_grid_pin_1_;
 inout prog_clk_0_S_in;
 inout [19:0] chanx_left_in;
 output [19:0] chanx_left_out;
 inout [19:0] chany_bottom_in;
 output [19:0] chany_bottom_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire \clknet_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_1_0_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_1_1_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_0_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_1_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_2_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_2_3_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_0_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_1_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_2_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_3_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_4_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_5_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_6_0_mem_bottom_track_1.prog_clk ;
 wire \clknet_3_7_0_mem_bottom_track_1.prog_clk ;
 wire \mem_bottom_track_1.ccff_tail ;
 wire \mem_bottom_track_1.mem_out[0] ;
 wire \mem_bottom_track_1.mem_out[1] ;
 wire \mem_bottom_track_1.prog_clk ;
 wire \mem_bottom_track_11.ccff_head ;
 wire \mem_bottom_track_11.ccff_tail ;
 wire \mem_bottom_track_11.mem_out[0] ;
 wire \mem_bottom_track_13.ccff_tail ;
 wire \mem_bottom_track_13.mem_out[0] ;
 wire \mem_bottom_track_15.ccff_tail ;
 wire \mem_bottom_track_15.mem_out[0] ;
 wire \mem_bottom_track_17.ccff_tail ;
 wire \mem_bottom_track_17.mem_out[0] ;
 wire \mem_bottom_track_19.ccff_tail ;
 wire \mem_bottom_track_19.mem_out[0] ;
 wire \mem_bottom_track_21.ccff_tail ;
 wire \mem_bottom_track_21.mem_out[0] ;
 wire \mem_bottom_track_23.ccff_tail ;
 wire \mem_bottom_track_23.mem_out[0] ;
 wire \mem_bottom_track_25.ccff_tail ;
 wire \mem_bottom_track_25.mem_out[0] ;
 wire \mem_bottom_track_27.ccff_tail ;
 wire \mem_bottom_track_27.mem_out[0] ;
 wire \mem_bottom_track_29.ccff_tail ;
 wire \mem_bottom_track_29.mem_out[0] ;
 wire \mem_bottom_track_3.ccff_tail ;
 wire \mem_bottom_track_3.mem_out[0] ;
 wire \mem_bottom_track_3.mem_out[1] ;
 wire \mem_bottom_track_5.ccff_tail ;
 wire \mem_bottom_track_5.mem_out[0] ;
 wire \mem_bottom_track_5.mem_out[1] ;
 wire \mem_bottom_track_7.ccff_tail ;
 wire \mem_bottom_track_7.mem_out[0] ;
 wire \mem_bottom_track_7.mem_out[1] ;
 wire \mem_bottom_track_9.mem_out[0] ;
 wire \mem_left_track_1.ccff_tail ;
 wire \mem_left_track_1.mem_out[0] ;
 wire \mem_left_track_1.mem_out[1] ;
 wire \mem_left_track_11.ccff_head ;
 wire \mem_left_track_11.ccff_tail ;
 wire \mem_left_track_11.mem_out[0] ;
 wire \mem_left_track_13.ccff_tail ;
 wire \mem_left_track_13.mem_out[0] ;
 wire \mem_left_track_15.ccff_tail ;
 wire \mem_left_track_15.mem_out[0] ;
 wire \mem_left_track_17.ccff_tail ;
 wire \mem_left_track_17.mem_out[0] ;
 wire \mem_left_track_19.ccff_tail ;
 wire \mem_left_track_19.mem_out[0] ;
 wire \mem_left_track_21.ccff_tail ;
 wire \mem_left_track_21.mem_out[0] ;
 wire \mem_left_track_23.ccff_tail ;
 wire \mem_left_track_23.mem_out[0] ;
 wire \mem_left_track_25.ccff_tail ;
 wire \mem_left_track_25.mem_out[0] ;
 wire \mem_left_track_27.ccff_tail ;
 wire \mem_left_track_27.mem_out[0] ;
 wire \mem_left_track_29.ccff_tail ;
 wire \mem_left_track_29.mem_out[0] ;
 wire \mem_left_track_3.ccff_tail ;
 wire \mem_left_track_3.mem_out[0] ;
 wire \mem_left_track_3.mem_out[1] ;
 wire \mem_left_track_31.ccff_tail ;
 wire \mem_left_track_31.mem_out[0] ;
 wire \mem_left_track_33.ccff_tail ;
 wire \mem_left_track_33.mem_out[0] ;
 wire \mem_left_track_35.ccff_tail ;
 wire \mem_left_track_35.mem_out[0] ;
 wire \mem_left_track_37.ccff_tail ;
 wire \mem_left_track_37.mem_out[0] ;
 wire \mem_left_track_39.mem_out[0] ;
 wire \mem_left_track_5.ccff_tail ;
 wire \mem_left_track_5.mem_out[0] ;
 wire \mem_left_track_5.mem_out[1] ;
 wire \mem_left_track_7.ccff_tail ;
 wire \mem_left_track_7.mem_out[0] ;
 wire \mem_left_track_7.mem_out[1] ;
 wire \mem_left_track_9.mem_out[0] ;
 wire \mux_bottom_track_1.out ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_11.out ;
 wire \mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_13.out ;
 wire \mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_15.out ;
 wire \mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_17.out ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_19.out ;
 wire \mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_21.out ;
 wire \mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_23.out ;
 wire \mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_25.out ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_27.out ;
 wire \mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_29.out ;
 wire \mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_3.out ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_5.out ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_bottom_track_7.out ;
 wire \mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_bottom_track_9.out ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_1.out ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_11.out ;
 wire \mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_13.out ;
 wire \mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_15.out ;
 wire \mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_17.out ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_19.out ;
 wire \mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_21.out ;
 wire \mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_23.out ;
 wire \mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_25.out ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_27.out ;
 wire \mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_29.out ;
 wire \mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_3.out ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_31.out ;
 wire \mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_33.out ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_35.out ;
 wire \mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_37.out ;
 wire \mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_39.out ;
 wire \mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_5.out ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X ;
 wire \mux_left_track_7.out ;
 wire \mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X ;
 wire \mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X ;
 wire \mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X ;
 wire \mux_left_track_9.out ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X ;
 wire \mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 ANTENNA__106__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(bottom_right_grid_pin_1_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(ccff_head));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(chanx_left_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(chanx_left_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(chanx_left_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(chanx_left_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(chanx_left_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(chanx_left_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(chanx_left_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(chanx_left_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(SC_IN_BOT));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(chanx_left_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(chanx_left_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(chanx_left_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(chanx_left_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(chanx_left_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(chanx_left_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(chanx_left_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(chanx_left_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(chanx_left_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(chanx_left_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(bottom_left_grid_pin_42_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(chanx_left_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(chanx_left_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(chany_bottom_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(chany_bottom_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(chany_bottom_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(chany_bottom_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(chany_bottom_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(chany_bottom_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(chany_bottom_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(chany_bottom_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(bottom_left_grid_pin_43_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(chany_bottom_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(chany_bottom_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(chany_bottom_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(chany_bottom_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(chany_bottom_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(chany_bottom_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(chany_bottom_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(chany_bottom_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(chany_bottom_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(chany_bottom_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(bottom_left_grid_pin_44_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(chany_bottom_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(chany_bottom_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(left_bottom_grid_pin_34_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(left_bottom_grid_pin_35_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(left_bottom_grid_pin_36_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(left_bottom_grid_pin_37_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(left_bottom_grid_pin_38_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(left_bottom_grid_pin_39_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(left_bottom_grid_pin_40_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(left_bottom_grid_pin_41_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(bottom_left_grid_pin_45_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(left_top_grid_pin_1_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(bottom_left_grid_pin_46_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(bottom_left_grid_pin_47_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(bottom_left_grid_pin_48_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(bottom_left_grid_pin_49_));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1  (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0  (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_25.mux_l1_in_1__A1  (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_27.mux_l1_in_0__A1  (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1  (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1  (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_0__A0  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_1__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_1.mux_l1_in_2__A1  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_15.mux_l1_in_0__A0  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_17.mux_l1_in_0__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_19.mux_l1_in_0__A0  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_21.mux_l1_in_0__A0  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_23.mux_l1_in_0__A0  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_25.mux_l1_in_0__A0  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_1__A0  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l1_in_1__A1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_3.mux_l2_in_1__A1  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_31.mux_l1_in_0__A0  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_33.mux_l1_in_0__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_35.mux_l1_in_0__A0  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_37.mux_l1_in_0__A0  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_39.mux_l1_in_0__A0  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l1_in_0__A0  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l1_in_1__A0  (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_5.mux_l1_in_2__A1  (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_7.mux_l1_in_1__A0  (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_7.mux_l1_in_1__A1  (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_7.mux_l2_in_1__A1  (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 \ANTENNA_mux_left_track_9.mux_l1_in_0__A0  (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_prog_clk_0_FTB00_A (.DIODE(prog_clk_0_S_in));
 sky130_fd_sc_hd__fill_2 FILLER_0_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_177 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_189 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_162 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_174 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_198 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_133 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_131 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_189 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_193 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_10 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_107 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_120 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_132 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_18 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_199 ();
 sky130_fd_sc_hd__decap_12 FILLER_17_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_201 ();
 sky130_fd_sc_hd__decap_12 FILLER_18_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_6 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_10 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_139 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_163 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_19_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_31 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_5 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_150 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_98 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_20_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_108 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_163 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_18 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_21_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_90 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_112 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_20 ();
 sky130_fd_sc_hd__decap_12 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_163 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_18 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_110 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_9 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_120 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_18 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_25_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_137 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_16 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_126 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_170 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_19 ();
 sky130_fd_sc_hd__decap_12 FILLER_27_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_108 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_28_30 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_91 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_163 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_20 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_220 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_29_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_107 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_89 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_106 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_118 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_14 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_142 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_144 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_192 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_35 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_40 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_52 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_84 ();
 sky130_fd_sc_hd__decap_12 FILLER_30_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_106 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_115 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_127 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_14 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_163 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_19 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_196 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_24 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_53 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_9 ();
 sky130_fd_sc_hd__decap_12 FILLER_31_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_135 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_156 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_168 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_20 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_9 ();
 sky130_fd_sc_hd__decap_12 FILLER_32_99 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_112 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_117 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_141 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_170 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_175 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_199 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_56 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_33_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_12 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_143 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_148 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_172 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_190 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_184 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_188 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_84 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_19 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_199 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_160 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_199 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_5 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_115 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_174 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_186 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_198 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_5 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_87 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_99 ();
 sky130_fd_sc_hd__conb_1 _035_ (.HI(_034_));
 sky130_fd_sc_hd__conb_1 _036_ (.HI(_000_));
 sky130_fd_sc_hd__conb_1 _037_ (.HI(_001_));
 sky130_fd_sc_hd__conb_1 _038_ (.HI(_002_));
 sky130_fd_sc_hd__conb_1 _039_ (.HI(_003_));
 sky130_fd_sc_hd__conb_1 _040_ (.HI(_004_));
 sky130_fd_sc_hd__conb_1 _041_ (.HI(_005_));
 sky130_fd_sc_hd__conb_1 _042_ (.HI(_006_));
 sky130_fd_sc_hd__conb_1 _043_ (.HI(_007_));
 sky130_fd_sc_hd__conb_1 _044_ (.HI(_008_));
 sky130_fd_sc_hd__conb_1 _045_ (.HI(_009_));
 sky130_fd_sc_hd__conb_1 _046_ (.HI(_010_));
 sky130_fd_sc_hd__conb_1 _047_ (.HI(_011_));
 sky130_fd_sc_hd__conb_1 _048_ (.HI(_012_));
 sky130_fd_sc_hd__conb_1 _049_ (.HI(_013_));
 sky130_fd_sc_hd__conb_1 _050_ (.HI(_014_));
 sky130_fd_sc_hd__conb_1 _051_ (.HI(_015_));
 sky130_fd_sc_hd__conb_1 _052_ (.HI(_016_));
 sky130_fd_sc_hd__conb_1 _053_ (.HI(_017_));
 sky130_fd_sc_hd__conb_1 _054_ (.HI(_018_));
 sky130_fd_sc_hd__conb_1 _055_ (.HI(_019_));
 sky130_fd_sc_hd__conb_1 _056_ (.HI(_020_));
 sky130_fd_sc_hd__conb_1 _057_ (.HI(_021_));
 sky130_fd_sc_hd__conb_1 _058_ (.HI(_022_));
 sky130_fd_sc_hd__conb_1 _059_ (.HI(_023_));
 sky130_fd_sc_hd__conb_1 _060_ (.HI(_024_));
 sky130_fd_sc_hd__conb_1 _061_ (.HI(_025_));
 sky130_fd_sc_hd__conb_1 _062_ (.HI(_026_));
 sky130_fd_sc_hd__conb_1 _063_ (.HI(_027_));
 sky130_fd_sc_hd__conb_1 _064_ (.HI(_028_));
 sky130_fd_sc_hd__conb_1 _065_ (.HI(_029_));
 sky130_fd_sc_hd__conb_1 _066_ (.HI(_030_));
 sky130_fd_sc_hd__conb_1 _067_ (.HI(_031_));
 sky130_fd_sc_hd__conb_1 _068_ (.HI(_032_));
 sky130_fd_sc_hd__conb_1 _069_ (.HI(_033_));
 sky130_fd_sc_hd__clkbuf_1 _070_ (.A(net1),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _071_ (.A(\mux_left_track_1.out ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _072_ (.A(\mux_left_track_3.out ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_1 _073_ (.A(\mux_left_track_5.out ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _074_ (.A(\mux_left_track_7.out ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _075_ (.A(\mux_left_track_9.out ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _076_ (.A(\mux_left_track_11.out ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _077_ (.A(\mux_left_track_13.out ),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_1 _078_ (.A(\mux_left_track_15.out ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _079_ (.A(\mux_left_track_17.out ),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 _080_ (.A(\mux_left_track_19.out ),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 _081_ (.A(\mux_left_track_21.out ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _082_ (.A(\mux_left_track_23.out ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _083_ (.A(\mux_left_track_25.out ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _084_ (.A(\mux_left_track_27.out ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _085_ (.A(\mux_left_track_29.out ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _086_ (.A(\mux_left_track_31.out ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _087_ (.A(\mux_left_track_33.out ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _088_ (.A(\mux_left_track_35.out ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 _089_ (.A(\mux_left_track_37.out ),
    .X(net72));
 sky130_fd_sc_hd__buf_1 _090_ (.A(\mux_left_track_39.out ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_1 _091_ (.A(\mux_bottom_track_1.out ),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 _092_ (.A(\mux_bottom_track_3.out ),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_1 _093_ (.A(\mux_bottom_track_5.out ),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 _094_ (.A(\mux_bottom_track_7.out ),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 _095_ (.A(\mux_bottom_track_9.out ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_1 _096_ (.A(\mux_bottom_track_11.out ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_1 _097_ (.A(\mux_bottom_track_13.out ),
    .X(net99));
 sky130_fd_sc_hd__clkbuf_1 _098_ (.A(\mux_bottom_track_15.out ),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 _099_ (.A(\mux_bottom_track_17.out ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 _100_ (.A(\mux_bottom_track_19.out ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 _101_ (.A(\mux_bottom_track_21.out ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 _102_ (.A(\mux_bottom_track_23.out ),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 _103_ (.A(\mux_bottom_track_25.out ),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 _104_ (.A(\mux_bottom_track_27.out ),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_1 _105_ (.A(\mux_bottom_track_29.out ),
    .X(net88));
 sky130_fd_sc_hd__buf_1 _106_ (.A(net19),
    .X(net89));
 sky130_fd_sc_hd__buf_1 _107_ (.A(net20),
    .X(net90));
 sky130_fd_sc_hd__buf_1 _108_ (.A(net21),
    .X(net91));
 sky130_fd_sc_hd__buf_1 _109_ (.A(net22),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_1 _110_ (.A(net12),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_mem_bottom_track_1.prog_clk  (.A(\mem_bottom_track_1.prog_clk ),
    .X(\clknet_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_1_0_0_mem_bottom_track_1.prog_clk  (.A(\clknet_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_1_0_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_1_1_0_mem_bottom_track_1.prog_clk  (.A(\clknet_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_1_1_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_0_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_0_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_1_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_1_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_2_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_2_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_2_3_0_mem_bottom_track_1.prog_clk  (.A(\clknet_1_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_2_3_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_0_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_0_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_1_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_0_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_1_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_2_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_2_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_3_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_1_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_3_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_4_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_2_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_4_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_5_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_2_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_5_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_6_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_3_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_6_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 \clkbuf_3_7_0_mem_bottom_track_1.prog_clk  (.A(\clknet_2_3_0_mem_bottom_track_1.prog_clk ),
    .X(\clknet_3_7_0_mem_bottom_track_1.prog_clk ));
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(SC_IN_BOT),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(bottom_right_grid_pin_1_),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(ccff_head),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(chanx_left_in[0]),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(chanx_left_in[10]),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(chanx_left_in[11]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(chanx_left_in[12]),
    .X(net15));
 sky130_fd_sc_hd__buf_1 input16 (.A(chanx_left_in[13]),
    .X(net16));
 sky130_fd_sc_hd__buf_1 input17 (.A(chanx_left_in[14]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(chanx_left_in[15]),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(chanx_left_in[16]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(bottom_left_grid_pin_42_),
    .X(net2));
 sky130_fd_sc_hd__buf_1 input20 (.A(chanx_left_in[17]),
    .X(net20));
 sky130_fd_sc_hd__buf_1 input21 (.A(chanx_left_in[18]),
    .X(net21));
 sky130_fd_sc_hd__buf_1 input22 (.A(chanx_left_in[19]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(chanx_left_in[1]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(chanx_left_in[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(chanx_left_in[3]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(chanx_left_in[4]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(chanx_left_in[5]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(chanx_left_in[6]),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_1 input29 (.A(chanx_left_in[7]),
    .X(net29));
 sky130_fd_sc_hd__buf_1 input3 (.A(bottom_left_grid_pin_43_),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(chanx_left_in[8]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_1 input31 (.A(chanx_left_in[9]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(chany_bottom_in[0]),
    .X(net32));
 sky130_fd_sc_hd__buf_1 input33 (.A(chany_bottom_in[10]),
    .X(net33));
 sky130_fd_sc_hd__buf_1 input34 (.A(chany_bottom_in[11]),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 input35 (.A(chany_bottom_in[12]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(chany_bottom_in[13]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(chany_bottom_in[14]),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(chany_bottom_in[15]),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(chany_bottom_in[16]),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input4 (.A(bottom_left_grid_pin_44_),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input40 (.A(chany_bottom_in[17]),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(chany_bottom_in[18]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(chany_bottom_in[19]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(chany_bottom_in[1]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(chany_bottom_in[2]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(chany_bottom_in[3]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(chany_bottom_in[4]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(chany_bottom_in[5]),
    .X(net47));
 sky130_fd_sc_hd__buf_1 input48 (.A(chany_bottom_in[6]),
    .X(net48));
 sky130_fd_sc_hd__buf_1 input49 (.A(chany_bottom_in[7]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(bottom_left_grid_pin_45_),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input50 (.A(chany_bottom_in[8]),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(chany_bottom_in[9]),
    .X(net51));
 sky130_fd_sc_hd__buf_1 input52 (.A(left_bottom_grid_pin_34_),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 input53 (.A(left_bottom_grid_pin_35_),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_2 input54 (.A(left_bottom_grid_pin_36_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input55 (.A(left_bottom_grid_pin_37_),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_2 input56 (.A(left_bottom_grid_pin_38_),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_2 input57 (.A(left_bottom_grid_pin_39_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(left_bottom_grid_pin_40_),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_2 input59 (.A(left_bottom_grid_pin_41_),
    .X(net59));
 sky130_fd_sc_hd__buf_1 input6 (.A(bottom_left_grid_pin_46_),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(left_top_grid_pin_1_),
    .X(net60));
 sky130_fd_sc_hd__buf_1 input7 (.A(bottom_left_grid_pin_47_),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(bottom_left_grid_pin_48_),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(bottom_left_grid_pin_49_),
    .X(net9));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(net11),
    .Q(\mem_bottom_track_1.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.mem_out[0] ),
    .Q(\mem_bottom_track_1.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.mem_out[1] ),
    .Q(\mem_bottom_track_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_11.ccff_head ),
    .Q(\mem_bottom_track_11.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_11.mem_out[0] ),
    .Q(\mem_bottom_track_11.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_11.ccff_tail ),
    .Q(\mem_bottom_track_13.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_13.mem_out[0] ),
    .Q(\mem_bottom_track_13.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_13.ccff_tail ),
    .Q(\mem_bottom_track_15.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_15.mem_out[0] ),
    .Q(\mem_bottom_track_15.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_15.ccff_tail ),
    .Q(\mem_bottom_track_17.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.mem_out[0] ),
    .Q(\mem_bottom_track_17.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_17.ccff_tail ),
    .Q(\mem_bottom_track_19.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_19.mem_out[0] ),
    .Q(\mem_bottom_track_19.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_19.ccff_tail ),
    .Q(\mem_bottom_track_21.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_21.mem_out[0] ),
    .Q(\mem_bottom_track_21.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_21.ccff_tail ),
    .Q(\mem_bottom_track_23.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_23.mem_out[0] ),
    .Q(\mem_bottom_track_23.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_23.ccff_tail ),
    .Q(\mem_bottom_track_25.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_25.mem_out[0] ),
    .Q(\mem_bottom_track_25.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_25.ccff_tail ),
    .Q(\mem_bottom_track_27.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_27.mem_out[0] ),
    .Q(\mem_bottom_track_27.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_5_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_27.ccff_tail ),
    .Q(\mem_bottom_track_29.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_29.mem_out[0] ),
    .Q(\mem_bottom_track_29.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_1.ccff_tail ),
    .Q(\mem_bottom_track_3.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.mem_out[0] ),
    .Q(\mem_bottom_track_3.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.mem_out[1] ),
    .Q(\mem_bottom_track_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_3.ccff_tail ),
    .Q(\mem_bottom_track_5.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.mem_out[0] ),
    .Q(\mem_bottom_track_5.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.mem_out[1] ),
    .Q(\mem_bottom_track_5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_5.ccff_tail ),
    .Q(\mem_bottom_track_7.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_7.mem_out[0] ),
    .Q(\mem_bottom_track_7.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_7.mem_out[1] ),
    .Q(\mem_bottom_track_7.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_4_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_7.ccff_tail ),
    .Q(\mem_bottom_track_9.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_9.mem_out[0] ),
    .Q(\mem_bottom_track_11.ccff_head ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_bottom_track_29.ccff_tail ),
    .Q(\mem_left_track_1.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.mem_out[0] ),
    .Q(\mem_left_track_1.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.mem_out[1] ),
    .Q(\mem_left_track_1.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_11.ccff_head ),
    .Q(\mem_left_track_11.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_11.mem_out[0] ),
    .Q(\mem_left_track_11.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_11.ccff_tail ),
    .Q(\mem_left_track_13.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_13.mem_out[0] ),
    .Q(\mem_left_track_13.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_13.ccff_tail ),
    .Q(\mem_left_track_15.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_15.mem_out[0] ),
    .Q(\mem_left_track_15.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_15.ccff_tail ),
    .Q(\mem_left_track_17.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.mem_out[0] ),
    .Q(\mem_left_track_17.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_17.ccff_tail ),
    .Q(\mem_left_track_19.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_19.mem_out[0] ),
    .Q(\mem_left_track_19.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_19.ccff_tail ),
    .Q(\mem_left_track_21.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_21.mem_out[0] ),
    .Q(\mem_left_track_21.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_21.ccff_tail ),
    .Q(\mem_left_track_23.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_23.mem_out[0] ),
    .Q(\mem_left_track_23.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_23.ccff_tail ),
    .Q(\mem_left_track_25.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_25.mem_out[0] ),
    .Q(\mem_left_track_25.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_25.ccff_tail ),
    .Q(\mem_left_track_27.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_27.mem_out[0] ),
    .Q(\mem_left_track_27.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_27.ccff_tail ),
    .Q(\mem_left_track_29.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_29.mem_out[0] ),
    .Q(\mem_left_track_29.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_6_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_1.ccff_tail ),
    .Q(\mem_left_track_3.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.mem_out[0] ),
    .Q(\mem_left_track_3.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.mem_out[1] ),
    .Q(\mem_left_track_3.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_29.ccff_tail ),
    .Q(\mem_left_track_31.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_31.mem_out[0] ),
    .Q(\mem_left_track_31.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_31.ccff_tail ),
    .Q(\mem_left_track_33.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_33.mem_out[0] ),
    .Q(\mem_left_track_33.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_33.ccff_tail ),
    .Q(\mem_left_track_35.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_35.mem_out[0] ),
    .Q(\mem_left_track_35.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_35.ccff_tail ),
    .Q(\mem_left_track_37.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_37.mem_out[0] ),
    .Q(\mem_left_track_37.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_3_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_37.ccff_tail ),
    .Q(\mem_left_track_39.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_7_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_39.mem_out[0] ),
    .Q(net62));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_3.ccff_tail ),
    .Q(\mem_left_track_5.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.mem_out[0] ),
    .Q(\mem_left_track_5.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_0_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.mem_out[1] ),
    .Q(\mem_left_track_5.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_5.ccff_tail ),
    .Q(\mem_left_track_7.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_7.mem_out[0] ),
    .Q(\mem_left_track_7.mem_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_7.mem_out[1] ),
    .Q(\mem_left_track_7.ccff_tail ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_  (.CLK(\clknet_3_1_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_7.ccff_tail ),
    .Q(\mem_left_track_9.mem_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 \mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_  (.CLK(\clknet_3_2_0_mem_bottom_track_1.prog_clk ),
    .D(\mem_left_track_9.mem_out[0] ),
    .Q(\mem_left_track_11.ccff_head ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_0_  (.A0(net3),
    .A1(net10),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_1_  (.A0(net7),
    .A1(net5),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l1_in_2_  (.A0(net23),
    .A1(net9),
    .S(\mem_bottom_track_1.mem_out[0] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l2_in_0_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_1.mem_out[1] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l2_in_1_  (.A0(_022_),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_1.mem_out[1] ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_1.mux_l3_in_0_  (.A0(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_bottom_track_1.ccff_tail ),
    .X(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_1.sky130_fd_sc_hd__mux2_1_5_X ),
    .X(\mux_bottom_track_1.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_11.mux_l1_in_0_  (.A0(net28),
    .A1(net2),
    .S(\mem_bottom_track_11.mem_out[0] ),
    .X(\mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_11.mux_l2_in_0_  (.A0(_023_),
    .A1(\mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_11.ccff_tail ),
    .X(\mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_11.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_11.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_13.mux_l1_in_0_  (.A0(net29),
    .A1(net3),
    .S(\mem_bottom_track_13.mem_out[0] ),
    .X(\mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_13.mux_l2_in_0_  (.A0(_024_),
    .A1(\mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_13.ccff_tail ),
    .X(\mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_13.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_13.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_15.mux_l1_in_0_  (.A0(net30),
    .A1(net4),
    .S(\mem_bottom_track_15.mem_out[0] ),
    .X(\mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_15.mux_l2_in_0_  (.A0(_025_),
    .A1(\mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_15.ccff_tail ),
    .X(\mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_15.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_15.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l1_in_0_  (.A0(net31),
    .A1(net5),
    .S(\mem_bottom_track_17.mem_out[0] ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_17.mux_l2_in_0_  (.A0(_026_),
    .A1(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_17.ccff_tail ),
    .X(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_17.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_17.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_19.mux_l1_in_0_  (.A0(net13),
    .A1(net6),
    .S(\mem_bottom_track_19.mem_out[0] ),
    .X(\mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_19.mux_l2_in_0_  (.A0(_027_),
    .A1(\mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_19.ccff_tail ),
    .X(\mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_19.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_19.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_21.mux_l1_in_0_  (.A0(net14),
    .A1(net7),
    .S(\mem_bottom_track_21.mem_out[0] ),
    .X(\mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_21.mux_l2_in_0_  (.A0(_028_),
    .A1(\mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_21.ccff_tail ),
    .X(\mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_21.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_21.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_23.mux_l1_in_0_  (.A0(net15),
    .A1(net8),
    .S(\mem_bottom_track_23.mem_out[0] ),
    .X(\mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_23.mux_l2_in_0_  (.A0(_029_),
    .A1(\mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_23.ccff_tail ),
    .X(\mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_23.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_23.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l1_in_0_  (.A0(net9),
    .A1(net10),
    .S(\mem_bottom_track_25.mem_out[0] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l1_in_1_  (.A0(_030_),
    .A1(net16),
    .S(\mem_bottom_track_25.mem_out[0] ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_25.mux_l2_in_0_  (.A0(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_25.ccff_tail ),
    .X(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_25.sky130_fd_sc_hd__mux2_1_2_X ),
    .X(\mux_bottom_track_25.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_27.mux_l1_in_0_  (.A0(net17),
    .A1(net2),
    .S(\mem_bottom_track_27.mem_out[0] ),
    .X(\mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_27.mux_l2_in_0_  (.A0(_031_),
    .A1(\mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_27.ccff_tail ),
    .X(\mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_27.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_27.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_29.mux_l1_in_0_  (.A0(net18),
    .A1(net3),
    .S(\mem_bottom_track_29.mem_out[0] ),
    .X(\mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_29.mux_l2_in_0_  (.A0(_032_),
    .A1(\mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_29.ccff_tail ),
    .X(\mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_29.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_29.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_0_  (.A0(net4),
    .A1(net2),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l1_in_1_  (.A0(net8),
    .A1(net6),
    .S(\mem_bottom_track_3.mem_out[0] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l2_in_0_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_3.mem_out[1] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l2_in_1_  (.A0(_033_),
    .A1(net24),
    .S(\mem_bottom_track_3.mem_out[1] ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_3.mux_l3_in_0_  (.A0(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_3.ccff_tail ),
    .X(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_3.sky130_fd_sc_hd__mux2_1_4_X ),
    .X(\mux_bottom_track_3.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l1_in_0_  (.A0(net3),
    .A1(net10),
    .S(\mem_bottom_track_5.mem_out[0] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l1_in_1_  (.A0(net7),
    .A1(net5),
    .S(\mem_bottom_track_5.mem_out[0] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l1_in_2_  (.A0(net25),
    .A1(net9),
    .S(\mem_bottom_track_5.mem_out[0] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_0_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l2_in_1_  (.A0(_034_),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_5.mem_out[1] ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_5.mux_l3_in_0_  (.A0(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_bottom_track_5.ccff_tail ),
    .X(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_5.sky130_fd_sc_hd__mux2_1_5_X ),
    .X(\mux_bottom_track_5.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_7.mux_l1_in_0_  (.A0(net4),
    .A1(net2),
    .S(\mem_bottom_track_7.mem_out[0] ),
    .X(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_7.mux_l1_in_1_  (.A0(net8),
    .A1(net6),
    .S(\mem_bottom_track_7.mem_out[0] ),
    .X(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_7.mux_l2_in_0_  (.A0(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_7.mem_out[1] ),
    .X(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_7.mux_l2_in_1_  (.A0(_000_),
    .A1(net26),
    .S(\mem_bottom_track_7.mem_out[1] ),
    .X(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_7.mux_l3_in_0_  (.A0(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_bottom_track_7.ccff_tail ),
    .X(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_7.sky130_fd_sc_hd__mux2_1_4_X ),
    .X(\mux_bottom_track_7.out ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l1_in_0_  (.A0(net27),
    .A1(net10),
    .S(\mem_bottom_track_9.mem_out[0] ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_bottom_track_9.mux_l2_in_0_  (.A0(_001_),
    .A1(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_bottom_track_11.ccff_head ),
    .X(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_bottom_track_9.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_bottom_track_9.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_0_  (.A0(net60),
    .A1(net42),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_1_  (.A0(net55),
    .A1(net53),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l1_in_2_  (.A0(net59),
    .A1(net57),
    .S(\mem_left_track_1.mem_out[0] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l2_in_0_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_1.mem_out[1] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l2_in_1_  (.A0(_002_),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_1.mem_out[1] ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_1.mux_l3_in_0_  (.A0(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_left_track_1.ccff_tail ),
    .X(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_1.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_1.sky130_fd_sc_hd__mux2_1_5_X ),
    .X(\mux_left_track_1.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_11.mux_l1_in_0_  (.A0(net52),
    .A1(net46),
    .S(\mem_left_track_11.mem_out[0] ),
    .X(\mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_11.mux_l2_in_0_  (.A0(_003_),
    .A1(\mux_left_track_11.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_11.ccff_tail ),
    .X(\mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_11.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_11.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_11.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_13.mux_l1_in_0_  (.A0(net53),
    .A1(net47),
    .S(\mem_left_track_13.mem_out[0] ),
    .X(\mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_13.mux_l2_in_0_  (.A0(_004_),
    .A1(\mux_left_track_13.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_13.ccff_tail ),
    .X(\mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_13.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_13.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_13.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_15.mux_l1_in_0_  (.A0(net54),
    .A1(net48),
    .S(\mem_left_track_15.mem_out[0] ),
    .X(\mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_15.mux_l2_in_0_  (.A0(_005_),
    .A1(\mux_left_track_15.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_15.ccff_tail ),
    .X(\mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_15.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_15.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_15.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l1_in_0_  (.A0(net55),
    .A1(net49),
    .S(\mem_left_track_17.mem_out[0] ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_17.mux_l2_in_0_  (.A0(_006_),
    .A1(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_17.ccff_tail ),
    .X(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_17.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_17.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_17.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_19.mux_l1_in_0_  (.A0(net56),
    .A1(net50),
    .S(\mem_left_track_19.mem_out[0] ),
    .X(\mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_19.mux_l2_in_0_  (.A0(_007_),
    .A1(\mux_left_track_19.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_19.ccff_tail ),
    .X(\mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_19.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_19.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_19.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_21.mux_l1_in_0_  (.A0(net57),
    .A1(net51),
    .S(\mem_left_track_21.mem_out[0] ),
    .X(\mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_21.mux_l2_in_0_  (.A0(_008_),
    .A1(\mux_left_track_21.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_21.ccff_tail ),
    .X(\mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_21.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_21.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_21.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_23.mux_l1_in_0_  (.A0(net58),
    .A1(net33),
    .S(\mem_left_track_23.mem_out[0] ),
    .X(\mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_23.mux_l2_in_0_  (.A0(_009_),
    .A1(\mux_left_track_23.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_23.ccff_tail ),
    .X(\mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_23.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_23.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_23.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l1_in_0_  (.A0(net60),
    .A1(net34),
    .S(\mem_left_track_25.mem_out[0] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l1_in_1_  (.A0(_010_),
    .A1(net59),
    .S(\mem_left_track_25.mem_out[0] ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_25.mux_l2_in_0_  (.A0(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_25.ccff_tail ),
    .X(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_25.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_25.sky130_fd_sc_hd__mux2_1_2_X ),
    .X(\mux_left_track_25.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_27.mux_l1_in_0_  (.A0(net52),
    .A1(net35),
    .S(\mem_left_track_27.mem_out[0] ),
    .X(\mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_27.mux_l2_in_0_  (.A0(_011_),
    .A1(\mux_left_track_27.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_27.ccff_tail ),
    .X(\mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_27.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_27.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_27.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_29.mux_l1_in_0_  (.A0(net53),
    .A1(net36),
    .S(\mem_left_track_29.mem_out[0] ),
    .X(\mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_29.mux_l2_in_0_  (.A0(_012_),
    .A1(\mux_left_track_29.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_29.ccff_tail ),
    .X(\mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_29.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_29.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_29.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_0_  (.A0(net52),
    .A1(net32),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l1_in_1_  (.A0(net56),
    .A1(net54),
    .S(\mem_left_track_3.mem_out[0] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l2_in_0_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_3.mem_out[1] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l2_in_1_  (.A0(_013_),
    .A1(net58),
    .S(\mem_left_track_3.mem_out[1] ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_3.mux_l3_in_0_  (.A0(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_3.ccff_tail ),
    .X(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_3.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_3.sky130_fd_sc_hd__mux2_1_4_X ),
    .X(\mux_left_track_3.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_31.mux_l1_in_0_  (.A0(net54),
    .A1(net37),
    .S(\mem_left_track_31.mem_out[0] ),
    .X(\mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_31.mux_l2_in_0_  (.A0(_014_),
    .A1(\mux_left_track_31.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_31.ccff_tail ),
    .X(\mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_31.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_31.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_31.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l1_in_0_  (.A0(net55),
    .A1(net38),
    .S(\mem_left_track_33.mem_out[0] ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_33.mux_l2_in_0_  (.A0(_015_),
    .A1(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_33.ccff_tail ),
    .X(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_33.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_33.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_33.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_35.mux_l1_in_0_  (.A0(net56),
    .A1(net39),
    .S(\mem_left_track_35.mem_out[0] ),
    .X(\mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_35.mux_l2_in_0_  (.A0(_016_),
    .A1(\mux_left_track_35.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_35.ccff_tail ),
    .X(\mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_35.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_35.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_35.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_37.mux_l1_in_0_  (.A0(net57),
    .A1(net40),
    .S(\mem_left_track_37.mem_out[0] ),
    .X(\mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_37.mux_l2_in_0_  (.A0(_017_),
    .A1(\mux_left_track_37.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_37.ccff_tail ),
    .X(\mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_37.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_37.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_37.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_39.mux_l1_in_0_  (.A0(net58),
    .A1(net41),
    .S(\mem_left_track_39.mem_out[0] ),
    .X(\mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_39.mux_l2_in_0_  (.A0(_018_),
    .A1(\mux_left_track_39.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(net62),
    .X(\mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_39.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_39.sky130_fd_sc_hd__mux2_1_1_X ),
    .X(\mux_left_track_39.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l1_in_0_  (.A0(net60),
    .A1(net43),
    .S(\mem_left_track_5.mem_out[0] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l1_in_1_  (.A0(net55),
    .A1(net53),
    .S(\mem_left_track_5.mem_out[0] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l1_in_2_  (.A0(net59),
    .A1(net57),
    .S(\mem_left_track_5.mem_out[0] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_0_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l2_in_1_  (.A0(_019_),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_5.mem_out[1] ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_5.mux_l3_in_0_  (.A0(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_4_X ),
    .A1(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_3_X ),
    .S(\mem_left_track_5.ccff_tail ),
    .X(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_5.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_5.sky130_fd_sc_hd__mux2_1_5_X ),
    .X(\mux_left_track_5.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_7.mux_l1_in_0_  (.A0(net52),
    .A1(net44),
    .S(\mem_left_track_7.mem_out[0] ),
    .X(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_7.mux_l1_in_1_  (.A0(net56),
    .A1(net54),
    .S(\mem_left_track_7.mem_out[0] ),
    .X(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_7.mux_l2_in_0_  (.A0(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_7.mem_out[1] ),
    .X(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_7.mux_l2_in_1_  (.A0(_020_),
    .A1(net58),
    .S(\mem_left_track_7.mem_out[1] ),
    .X(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_7.mux_l3_in_0_  (.A0(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_3_X ),
    .A1(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_2_X ),
    .S(\mem_left_track_7.ccff_tail ),
    .X(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_7.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_7.sky130_fd_sc_hd__mux2_1_4_X ),
    .X(\mux_left_track_7.out ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l1_in_0_  (.A0(net60),
    .A1(net45),
    .S(\mem_left_track_9.mem_out[0] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l1_in_1_  (.A0(_021_),
    .A1(net59),
    .S(\mem_left_track_9.mem_out[0] ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X ));
 sky130_fd_sc_hd__mux2_1 \mux_left_track_9.mux_l2_in_0_  (.A0(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_1_X ),
    .A1(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_0_X ),
    .S(\mem_left_track_11.ccff_head ),
    .X(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X ));
 sky130_fd_sc_hd__clkbuf_1 \mux_left_track_9.sky130_fd_sc_hd__buf_4_0_  (.A(\mux_left_track_9.sky130_fd_sc_hd__mux2_1_2_X ),
    .X(\mux_left_track_9.out ));
 sky130_fd_sc_hd__clkbuf_2 output100 (.A(net100),
    .X(chany_bottom_out[7]));
 sky130_fd_sc_hd__clkbuf_2 output101 (.A(net101),
    .X(chany_bottom_out[8]));
 sky130_fd_sc_hd__clkbuf_2 output102 (.A(net102),
    .X(chany_bottom_out[9]));
 sky130_fd_sc_hd__clkbuf_2 output61 (.A(net61),
    .X(SC_OUT_BOT));
 sky130_fd_sc_hd__clkbuf_2 output62 (.A(net62),
    .X(ccff_tail));
 sky130_fd_sc_hd__clkbuf_2 output63 (.A(net63),
    .X(chanx_left_out[0]));
 sky130_fd_sc_hd__clkbuf_2 output64 (.A(net64),
    .X(chanx_left_out[10]));
 sky130_fd_sc_hd__clkbuf_2 output65 (.A(net65),
    .X(chanx_left_out[11]));
 sky130_fd_sc_hd__clkbuf_2 output66 (.A(net66),
    .X(chanx_left_out[12]));
 sky130_fd_sc_hd__clkbuf_2 output67 (.A(net67),
    .X(chanx_left_out[13]));
 sky130_fd_sc_hd__clkbuf_2 output68 (.A(net68),
    .X(chanx_left_out[14]));
 sky130_fd_sc_hd__clkbuf_2 output69 (.A(net69),
    .X(chanx_left_out[15]));
 sky130_fd_sc_hd__clkbuf_2 output70 (.A(net70),
    .X(chanx_left_out[16]));
 sky130_fd_sc_hd__clkbuf_2 output71 (.A(net71),
    .X(chanx_left_out[17]));
 sky130_fd_sc_hd__clkbuf_2 output72 (.A(net72),
    .X(chanx_left_out[18]));
 sky130_fd_sc_hd__clkbuf_2 output73 (.A(net73),
    .X(chanx_left_out[19]));
 sky130_fd_sc_hd__clkbuf_2 output74 (.A(net74),
    .X(chanx_left_out[1]));
 sky130_fd_sc_hd__clkbuf_2 output75 (.A(net75),
    .X(chanx_left_out[2]));
 sky130_fd_sc_hd__clkbuf_2 output76 (.A(net76),
    .X(chanx_left_out[3]));
 sky130_fd_sc_hd__clkbuf_2 output77 (.A(net77),
    .X(chanx_left_out[4]));
 sky130_fd_sc_hd__clkbuf_2 output78 (.A(net78),
    .X(chanx_left_out[5]));
 sky130_fd_sc_hd__clkbuf_2 output79 (.A(net79),
    .X(chanx_left_out[6]));
 sky130_fd_sc_hd__clkbuf_2 output80 (.A(net80),
    .X(chanx_left_out[7]));
 sky130_fd_sc_hd__clkbuf_2 output81 (.A(net81),
    .X(chanx_left_out[8]));
 sky130_fd_sc_hd__clkbuf_2 output82 (.A(net82),
    .X(chanx_left_out[9]));
 sky130_fd_sc_hd__clkbuf_2 output83 (.A(net83),
    .X(chany_bottom_out[0]));
 sky130_fd_sc_hd__clkbuf_2 output84 (.A(net84),
    .X(chany_bottom_out[10]));
 sky130_fd_sc_hd__clkbuf_2 output85 (.A(net85),
    .X(chany_bottom_out[11]));
 sky130_fd_sc_hd__clkbuf_2 output86 (.A(net86),
    .X(chany_bottom_out[12]));
 sky130_fd_sc_hd__clkbuf_2 output87 (.A(net87),
    .X(chany_bottom_out[13]));
 sky130_fd_sc_hd__clkbuf_2 output88 (.A(net88),
    .X(chany_bottom_out[14]));
 sky130_fd_sc_hd__clkbuf_2 output89 (.A(net89),
    .X(chany_bottom_out[15]));
 sky130_fd_sc_hd__clkbuf_2 output90 (.A(net90),
    .X(chany_bottom_out[16]));
 sky130_fd_sc_hd__clkbuf_2 output91 (.A(net91),
    .X(chany_bottom_out[17]));
 sky130_fd_sc_hd__clkbuf_2 output92 (.A(net92),
    .X(chany_bottom_out[18]));
 sky130_fd_sc_hd__clkbuf_2 output93 (.A(net93),
    .X(chany_bottom_out[19]));
 sky130_fd_sc_hd__clkbuf_2 output94 (.A(net94),
    .X(chany_bottom_out[1]));
 sky130_fd_sc_hd__clkbuf_2 output95 (.A(net95),
    .X(chany_bottom_out[2]));
 sky130_fd_sc_hd__clkbuf_2 output96 (.A(net96),
    .X(chany_bottom_out[3]));
 sky130_fd_sc_hd__clkbuf_2 output97 (.A(net97),
    .X(chany_bottom_out[4]));
 sky130_fd_sc_hd__clkbuf_2 output98 (.A(net98),
    .X(chany_bottom_out[5]));
 sky130_fd_sc_hd__clkbuf_2 output99 (.A(net99),
    .X(chany_bottom_out[6]));
 sky130_fd_sc_hd__buf_8 prog_clk_0_FTB00 (.A(prog_clk_0_S_in),
    .X(\mem_bottom_track_1.prog_clk ));
endmodule
