* NGSPICE file created from sb_2__2_.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

.subckt sb_2__2_ SC_IN_BOT SC_OUT_BOT VGND VPWR bottom_left_grid_pin_42_ bottom_left_grid_pin_43_
+ bottom_left_grid_pin_44_ bottom_left_grid_pin_45_ bottom_left_grid_pin_46_ bottom_left_grid_pin_47_
+ bottom_left_grid_pin_48_ bottom_left_grid_pin_49_ bottom_right_grid_pin_1_ ccff_head
+ ccff_tail chanx_left_in[0] chanx_left_in[10] chanx_left_in[11] chanx_left_in[12]
+ chanx_left_in[13] chanx_left_in[14] chanx_left_in[15] chanx_left_in[16] chanx_left_in[17]
+ chanx_left_in[18] chanx_left_in[19] chanx_left_in[1] chanx_left_in[2] chanx_left_in[3]
+ chanx_left_in[4] chanx_left_in[5] chanx_left_in[6] chanx_left_in[7] chanx_left_in[8]
+ chanx_left_in[9] chanx_left_out[0] chanx_left_out[10] chanx_left_out[11] chanx_left_out[12]
+ chanx_left_out[13] chanx_left_out[14] chanx_left_out[15] chanx_left_out[16] chanx_left_out[17]
+ chanx_left_out[18] chanx_left_out[19] chanx_left_out[1] chanx_left_out[2] chanx_left_out[3]
+ chanx_left_out[4] chanx_left_out[5] chanx_left_out[6] chanx_left_out[7] chanx_left_out[8]
+ chanx_left_out[9] chany_bottom_in[0] chany_bottom_in[10] chany_bottom_in[11] chany_bottom_in[12]
+ chany_bottom_in[13] chany_bottom_in[14] chany_bottom_in[15] chany_bottom_in[16]
+ chany_bottom_in[17] chany_bottom_in[18] chany_bottom_in[19] chany_bottom_in[1] chany_bottom_in[2]
+ chany_bottom_in[3] chany_bottom_in[4] chany_bottom_in[5] chany_bottom_in[6] chany_bottom_in[7]
+ chany_bottom_in[8] chany_bottom_in[9] chany_bottom_out[0] chany_bottom_out[10] chany_bottom_out[11]
+ chany_bottom_out[12] chany_bottom_out[13] chany_bottom_out[14] chany_bottom_out[15]
+ chany_bottom_out[16] chany_bottom_out[17] chany_bottom_out[18] chany_bottom_out[19]
+ chany_bottom_out[1] chany_bottom_out[2] chany_bottom_out[3] chany_bottom_out[4]
+ chany_bottom_out[5] chany_bottom_out[6] chany_bottom_out[7] chany_bottom_out[8]
+ chany_bottom_out[9] left_bottom_grid_pin_34_ left_bottom_grid_pin_35_ left_bottom_grid_pin_36_
+ left_bottom_grid_pin_37_ left_bottom_grid_pin_38_ left_bottom_grid_pin_39_ left_bottom_grid_pin_40_
+ left_bottom_grid_pin_41_ left_top_grid_pin_1_ prog_clk_0_S_in
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_1_ input8/X input6/X mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold46/X VGND VGND VPWR VPWR hold33/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_mux_left_track_35.mux_l1_in_0__A1 input39/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input55_A left_bottom_grid_pin_37_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_17.mux_l1_in_0_ input31/X input5/X hold13/A VGND VGND VPWR VPWR
+ mux_bottom_track_17.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_128 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_7.mux_l2_in_1__105 VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/A0
+ mux_bottom_track_7.mux_l2_in_1__105/LO sky130_fd_sc_hd__conb_1
XFILLER_20_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold41 hold41/A VGND VGND VPWR VPWR hold41/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold30 hold30/A VGND VGND VPWR VPWR hold30/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold52 hold52/A VGND VGND VPWR VPWR hold52/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_29.mux_l2_in_0_ mux_bottom_track_29.mux_l2_in_0_/A0 mux_bottom_track_29.mux_l1_in_0_/X
+ hold11/A VGND VGND VPWR VPWR mux_bottom_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input18_A chanx_left_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput75 _073_/X VGND VGND VPWR VPWR chanx_left_out[2] sky130_fd_sc_hd__buf_2
Xoutput64 _081_/X VGND VGND VPWR VPWR chanx_left_out[10] sky130_fd_sc_hd__buf_2
Xoutput97 _095_/X VGND VGND VPWR VPWR chany_bottom_out[4] sky130_fd_sc_hd__buf_2
Xoutput86 _103_/X VGND VGND VPWR VPWR chany_bottom_out[12] sky130_fd_sc_hd__buf_2
Xmux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_3.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _092_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_16_175 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l1_in_0_ input4/X input2/X mux_bottom_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input48_A chany_bottom_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.sky130_fd_sc_hd__buf_4_0_ mux_left_track_9.mux_l2_in_0_/X VGND VGND
+ VPWR VPWR _075_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR hold49/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_31.sky130_fd_sc_hd__buf_4_0_ mux_left_track_31.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _086_/A sky130_fd_sc_hd__clkbuf_1
Xhold20 hold20/A VGND VGND VPWR VPWR hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold42 hold42/A VGND VGND VPWR VPWR hold42/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold53 hold53/A VGND VGND VPWR VPWR hold53/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold31 hold31/A VGND VGND VPWR VPWR hold31/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold28/X VGND VGND VPWR VPWR hold4/A sky130_fd_sc_hd__dfxtp_1
XFILLER_15_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput87 _104_/X VGND VGND VPWR VPWR chany_bottom_out[13] sky130_fd_sc_hd__buf_2
Xoutput98 _096_/X VGND VGND VPWR VPWR chany_bottom_out[5] sky130_fd_sc_hd__buf_2
Xoutput76 _074_/X VGND VGND VPWR VPWR chanx_left_out[3] sky130_fd_sc_hd__buf_2
Xoutput65 _082_/X VGND VGND VPWR VPWR chanx_left_out[11] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A chanx_left_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_25.sky130_fd_sc_hd__buf_4_0_ mux_left_track_25.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _083_/A sky130_fd_sc_hd__clkbuf_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR hold32/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_29.mux_l1_in_0_ input18/X input3/X hold18/A VGND VGND VPWR VPWR
+ mux_bottom_track_29.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_26_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_19.sky130_fd_sc_hd__buf_4_0_ mux_left_track_19.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _080_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l3_in_0_ mux_left_track_7.mux_l2_in_1_/X mux_left_track_7.mux_l2_in_0_/X
+ hold38/A VGND VGND VPWR VPWR mux_left_track_7.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l2_in_1_ mux_left_track_7.mux_l2_in_1_/A0 input58/X mux_left_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input60_A left_top_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold41/X VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xhold32 hold32/A VGND VGND VPWR VPWR hold32/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold10 hold10/A VGND VGND VPWR VPWR hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold54 hold54/A VGND VGND VPWR VPWR hold54/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold43 hold43/A VGND VGND VPWR VPWR hold43/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold21 hold21/A VGND VGND VPWR VPWR hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold31/X VGND VGND VPWR VPWR hold28/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_17.mux_l2_in_0__131 VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/A0
+ mux_bottom_track_17.mux_l2_in_0__131/LO sky130_fd_sc_hd__conb_1
XFILLER_25_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput99 _097_/X VGND VGND VPWR VPWR chany_bottom_out[6] sky130_fd_sc_hd__buf_2
Xoutput88 _105_/X VGND VGND VPWR VPWR chany_bottom_out[14] sky130_fd_sc_hd__buf_2
Xoutput77 _075_/X VGND VGND VPWR VPWR chanx_left_out[4] sky130_fd_sc_hd__buf_2
Xoutput66 _083_/X VGND VGND VPWR VPWR chanx_left_out[12] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A chanx_left_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_15.mux_l2_in_0_ mux_left_track_15.mux_l2_in_0_/A0 mux_left_track_15.mux_l1_in_0_/X
+ hold46/A VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xprog_clk_0_FTB00 prog_clk_0_S_in VGND VGND VPWR VPWR prog_clk_0_FTB00/X sky130_fd_sc_hd__buf_8
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_7.mux_l2_in_0_ mux_left_track_7.mux_l1_in_1_/X mux_left_track_7.mux_l1_in_0_/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input53_A left_bottom_grid_pin_35_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_21.mux_l2_in_0__133 VGND VGND VPWR VPWR mux_bottom_track_21.mux_l2_in_0_/A0
+ mux_bottom_track_21.mux_l2_in_0__133/LO sky130_fd_sc_hd__conb_1
XFILLER_20_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold22 hold22/A VGND VGND VPWR VPWR hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold11 hold11/A VGND VGND VPWR VPWR hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold44 hold44/A VGND VGND VPWR VPWR hold44/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold33 hold33/A VGND VGND VPWR VPWR hold33/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold55 hold55/A VGND VGND VPWR VPWR hold55/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_131 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_7.mux_l1_in_1_ input56/X input54/X mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_134 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput89 _106_/X VGND VGND VPWR VPWR chany_bottom_out[15] sky130_fd_sc_hd__buf_2
Xoutput78 _076_/X VGND VGND VPWR VPWR chanx_left_out[5] sky130_fd_sc_hd__buf_2
Xoutput67 _084_/X VGND VGND VPWR VPWR chanx_left_out[13] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A chanx_left_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold9/X VGND VGND VPWR VPWR mux_bottom_track_3.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_input8_A bottom_left_grid_pin_48_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_1__A0 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold10/X VGND VGND VPWR VPWR hold16/A sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l1_in_0_ input54/X input48/X hold54/A VGND VGND VPWR VPWR mux_left_track_15.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
X_110_ _110_/A VGND VGND VPWR VPWR _110_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input46_A chany_bottom_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_27.mux_l2_in_0_ mux_left_track_27.mux_l2_in_0_/A0 mux_left_track_27.mux_l1_in_0_/X
+ hold3/A VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold12 hold12/A VGND VGND VPWR VPWR hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold34 hold34/A VGND VGND VPWR VPWR hold34/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A VGND VGND VPWR VPWR hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold45 hold45/A VGND VGND VPWR VPWR hold45/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold56 hold56/A VGND VGND VPWR VPWR hold56/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_143 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_11.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _096_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_7.mux_l1_in_0_ input52/X input44/X mux_left_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_146 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput79 _077_/X VGND VGND VPWR VPWR chanx_left_out[6] sky130_fd_sc_hd__buf_2
Xoutput68 _085_/X VGND VGND VPWR VPWR chanx_left_out[14] sky130_fd_sc_hd__buf_2
XFILLER_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_190 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_12_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold29/X VGND VGND VPWR VPWR hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold39/X VGND VGND VPWR VPWR hold36/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold20/X VGND VGND VPWR VPWR hold10/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_27.mux_l2_in_0__116 VGND VGND VPWR VPWR mux_left_track_27.mux_l2_in_0_/A0
+ mux_left_track_27.mux_l2_in_0__116/LO sky130_fd_sc_hd__conb_1
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input39_A chany_bottom_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold57 hold57/A VGND VGND VPWR VPWR hold57/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold13 hold13/A VGND VGND VPWR VPWR hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold24 hold24/A VGND VGND VPWR VPWR hold24/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold46 hold46/A VGND VGND VPWR VPWR hold46/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold35 hold35/A VGND VGND VPWR VPWR hold35/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_10_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_155 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_9.mux_l2_in_0__106 VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/A0
+ mux_bottom_track_9.mux_l2_in_0__106/LO sky130_fd_sc_hd__conb_1
XFILLER_15_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_27.mux_l1_in_0_ input52/X input35/X hold60/A VGND VGND VPWR VPWR mux_left_track_27.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput69 _086_/X VGND VGND VPWR VPWR chanx_left_out[15] sky130_fd_sc_hd__buf_2
XFILLER_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_39.mux_l2_in_0_ mux_left_track_39.mux_l2_in_0_/A0 mux_left_track_39.mux_l1_in_0_/X
+ output62/A VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_bottom_track_13.mux_l2_in_0_ mux_bottom_track_13.mux_l2_in_0_/A0 mux_bottom_track_13.mux_l1_in_0_/X
+ hold34/A VGND VGND VPWR VPWR mux_bottom_track_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input21_A chanx_left_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold16/X VGND VGND VPWR VPWR hold29/A sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold51/X VGND VGND VPWR VPWR hold39/A sky130_fd_sc_hd__dfxtp_1
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_27.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _104_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_23_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_0__A0 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold13/X VGND VGND VPWR VPWR hold27/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_099_ _099_/A VGND VGND VPWR VPWR _099_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold60/X VGND VGND VPWR VPWR hold3/A sky130_fd_sc_hd__dfxtp_1
Xhold25 hold25/A VGND VGND VPWR VPWR hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold14 hold14/A VGND VGND VPWR VPWR hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_5.mux_l2_in_1__104 VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/A0
+ mux_bottom_track_5.mux_l2_in_1__104/LO sky130_fd_sc_hd__conb_1
Xhold58 hold58/A VGND VGND VPWR VPWR hold58/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold47 hold47/A VGND VGND VPWR VPWR hold47/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold36 hold36/A VGND VGND VPWR VPWR hold36/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input51_A chany_bottom_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_mux_left_track_23.mux_l1_in_0__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input14_A chanx_left_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_184 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input6_A bottom_left_grid_pin_46_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_39.mux_l1_in_0_ input58/X input41/X hold35/A VGND VGND VPWR VPWR mux_left_track_39.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_31.mux_l2_in_0__119 VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/A0
+ mux_left_track_31.mux_l2_in_0__119/LO sky130_fd_sc_hd__conb_1
XFILLER_27_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_13.mux_l1_in_0_ input29/X input3/X hold19/A VGND VGND VPWR VPWR
+ mux_bottom_track_13.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l2_in_0_ mux_bottom_track_25.mux_l1_in_1_/X mux_bottom_track_25.mux_l1_in_0_/X
+ hold49/A VGND VGND VPWR VPWR mux_bottom_track_25.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_29_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold22/X VGND VGND VPWR VPWR hold13/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_098_ _098_/A VGND VGND VPWR VPWR _098_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold5/X VGND VGND VPWR VPWR hold60/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_25.mux_l1_in_1_ mux_bottom_track_25.mux_l1_in_1_/A0 input16/X mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xhold26 hold26/A VGND VGND VPWR VPWR hold26/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold15 hold15/A VGND VGND VPWR VPWR hold15/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold59 hold59/A VGND VGND VPWR VPWR hold59/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold37 hold37/A VGND VGND VPWR VPWR hold37/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold48 hold48/A VGND VGND VPWR VPWR hold48/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_9.mux_l2_in_0_ mux_bottom_track_9.mux_l2_in_0_/A0 mux_bottom_track_9.mux_l1_in_0_/X
+ hold16/A VGND VGND VPWR VPWR mux_bottom_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input44_A chany_bottom_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_38 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_3.mux_l2_in_1__A1 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_5.sky130_fd_sc_hd__buf_4_0_ mux_left_track_5.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _073_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold59/X VGND VGND VPWR VPWR hold15/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_39.mux_l2_in_0__123 VGND VGND VPWR VPWR mux_left_track_39.mux_l2_in_0_/A0
+ mux_left_track_39.mux_l2_in_0__123/LO sky130_fd_sc_hd__conb_1
XFILLER_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.sky130_fd_sc_hd__buf_4_0_ mux_left_track_21.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _081_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_097_ _097_/A VGND VGND VPWR VPWR _097_/X sky130_fd_sc_hd__clkbuf_1
Xhold16 hold16/A VGND VGND VPWR VPWR hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold27 hold27/A VGND VGND VPWR VPWR hold27/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold38 hold38/A VGND VGND VPWR VPWR hold38/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_25.mux_l1_in_0_ input9/X input10/X mux_bottom_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xhold49 hold49/A VGND VGND VPWR VPWR hold49/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_15.sky130_fd_sc_hd__buf_4_0_ mux_left_track_15.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _078_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input37_A chany_bottom_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_15.mux_l2_in_0__130 VGND VGND VPWR VPWR mux_bottom_track_15.mux_l2_in_0_/A0
+ mux_bottom_track_15.mux_l2_in_0__130/LO sky130_fd_sc_hd__conb_1
XFILLER_31_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_3.mux_l3_in_0_ mux_left_track_3.mux_l2_in_1_/X mux_left_track_3.mux_l2_in_0_/X
+ hold17/A VGND VGND VPWR VPWR mux_left_track_3.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_9.mux_l1_in_0_ input27/X input10/X hold10/A VGND VGND VPWR VPWR
+ mux_bottom_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_25.mux_l1_in_1__115 VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/A0
+ mux_left_track_25.mux_l1_in_1__115/LO sky130_fd_sc_hd__conb_1
XANTENNA_mux_left_track_7.mux_l1_in_1__A0 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_9.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _095_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_5_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR hold59/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_1_ mux_left_track_3.mux_l2_in_1_/A0 input58/X hold57/A
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_3.mux_l2_in_1__118 VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_1_/A0
+ mux_left_track_3.mux_l2_in_1__118/LO sky130_fd_sc_hd__conb_1
XFILLER_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_096_ _096_/A VGND VGND VPWR VPWR _096_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR hold38/A sky130_fd_sc_hd__dfxtp_1
Xhold17 hold17/A VGND VGND VPWR VPWR hold17/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold28 hold28/A VGND VGND VPWR VPWR hold28/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold39 hold39/A VGND VGND VPWR VPWR hold39/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_3_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_13.mux_l2_in_0__109 VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/A0
+ mux_left_track_13.mux_l2_in_0__109/LO sky130_fd_sc_hd__conb_1
XFILLER_19_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_079_ _079_/A VGND VGND VPWR VPWR _079_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_16_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_11.mux_l2_in_0_ mux_left_track_11.mux_l2_in_0_/A0 mux_left_track_11.mux_l1_in_0_/X
+ hold43/A VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_37.sky130_fd_sc_hd__buf_4_0_ mux_left_track_37.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _089_/A sky130_fd_sc_hd__clkbuf_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold2/X VGND VGND VPWR VPWR hold37/A sky130_fd_sc_hd__dfxtp_1
Xmem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold11/X VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_3.mux_l2_in_0_ mux_left_track_3.mux_l1_in_1_/X mux_left_track_3.mux_l1_in_0_/X
+ hold57/A VGND VGND VPWR VPWR mux_left_track_3.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input12_A chanx_left_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input4_A bottom_left_grid_pin_44_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_3.mux_l1_in_1_ input56/X input54/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_095_ _095_/A VGND VGND VPWR VPWR _095_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_7.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_27_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold29 hold29/A VGND VGND VPWR VPWR hold29/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold18 hold18/A VGND VGND VPWR VPWR hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_078_ _078_/A VGND VGND VPWR VPWR _078_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input42_A chany_bottom_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_8_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold43/X VGND VGND VPWR VPWR hold2/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_11.mux_l1_in_0_ input52/X input46/X hold53/A VGND VGND VPWR VPWR mux_left_track_11.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_23.mux_l2_in_0_ mux_left_track_23.mux_l2_in_0_/A0 mux_left_track_23.mux_l1_in_0_/X
+ hold55/A VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_27_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_3.mux_l1_in_0_ input52/X input32/X mux_left_track_3.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold47/X VGND VGND VPWR VPWR hold51/A sky130_fd_sc_hd__dfxtp_1
X_094_ _094_/A VGND VGND VPWR VPWR _094_/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold58/X VGND VGND VPWR VPWR mux_left_track_7.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xhold19 hold19/A VGND VGND VPWR VPWR hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_077_ _077_/A VGND VGND VPWR VPWR _077_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input35_A chany_bottom_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_204 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_23.mux_l1_in_0_ input58/X input33/X hold50/A VGND VGND VPWR VPWR mux_left_track_23.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold56/X VGND VGND VPWR VPWR hold47/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_093_ _093_/A VGND VGND VPWR VPWR _093_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.mux_l2_in_0_ mux_left_track_35.mux_l2_in_0_/A0 mux_left_track_35.mux_l1_in_0_/X
+ hold4/A VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold6/X VGND VGND VPWR VPWR hold30/A sky130_fd_sc_hd__dfxtp_1
Xinput1 SC_IN_BOT VGND VGND VPWR VPWR _070_/A sky130_fd_sc_hd__clkbuf_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_3.mux_l2_in_1__103 VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/A0
+ mux_bottom_track_3.mux_l2_in_1__103/LO sky130_fd_sc_hd__conb_1
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_23.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _102_/A sky130_fd_sc_hd__clkbuf_1
X_076_ _076_/A VGND VGND VPWR VPWR _076_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_32_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold42/X VGND VGND VPWR VPWR hold48/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_37.mux_l1_in_0__A0 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input28_A chanx_left_in[6] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_17.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _099_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_12_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_42 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_7_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l3_in_0_ mux_bottom_track_5.mux_l2_in_1_/X mux_bottom_track_5.mux_l2_in_0_/X
+ hold44/A VGND VGND VPWR VPWR mux_bottom_track_5.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_5.mux_l2_in_1_ mux_bottom_track_5.mux_l2_in_1_/A0 mux_bottom_track_5.mux_l1_in_2_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
XANTENNA_input10_A bottom_right_grid_pin_1_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input2_A bottom_left_grid_pin_42_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_092_ _092_/A VGND VGND VPWR VPWR _092_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input58_A left_bottom_grid_pin_40_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold12/X VGND VGND VPWR VPWR hold6/A sky130_fd_sc_hd__dfxtp_1
Xinput2 bottom_left_grid_pin_42_ VGND VGND VPWR VPWR input2/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.mux_l1_in_2_ input25/X input9/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_119 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_075_ _075_/A VGND VGND VPWR VPWR _075_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_25_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold45/X VGND VGND VPWR VPWR hold42/A sky130_fd_sc_hd__dfxtp_1
XFILLER_24_111 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_37.mux_l1_in_0__A1 input40/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_35.mux_l1_in_0_ input56/X input39/X hold28/A VGND VGND VPWR VPWR mux_left_track_35.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_19.mux_l2_in_0_ mux_bottom_track_19.mux_l2_in_0_/A0 mux_bottom_track_19.mux_l1_in_0_/X
+ hold12/A VGND VGND VPWR VPWR mux_bottom_track_19.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_21_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput60 left_top_grid_pin_1_ VGND VGND VPWR VPWR input60/X sky130_fd_sc_hd__clkbuf_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold23/X VGND VGND VPWR VPWR hold7/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_54 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input40_A chany_bottom_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_21.mux_l2_in_0_ mux_bottom_track_21.mux_l2_in_0_/A0 mux_bottom_track_21.mux_l1_in_0_/X
+ hold30/A VGND VGND VPWR VPWR mux_bottom_track_21.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold21/X VGND VGND VPWR VPWR hold40/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_37.mux_l2_in_0__122 VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/A0
+ mux_left_track_37.mux_l2_in_0__122/LO sky130_fd_sc_hd__conb_1
XFILLER_32_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_5.mux_l2_in_0_ mux_bottom_track_5.mux_l1_in_1_/X mux_bottom_track_5.mux_l1_in_0_/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR hold44/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.sky130_fd_sc_hd__buf_4_0_ mux_left_track_1.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _071_/A sky130_fd_sc_hd__clkbuf_1
X_091_ _091_/A VGND VGND VPWR VPWR _091_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 bottom_left_grid_pin_43_ VGND VGND VPWR VPWR input3/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_1_ input7/X input5/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_074_ _074_/A VGND VGND VPWR VPWR _074_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_123 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput50 chany_bottom_in[8] VGND VGND VPWR VPWR input50/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_prog_clk_0_FTB00_A prog_clk_0_S_in VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_mux_left_track_1.mux_l1_in_0__A0 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold49/X VGND VGND VPWR VPWR hold23/A sky130_fd_sc_hd__dfxtp_1
XFILLER_32_66 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_input33_A chany_bottom_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ _109_/A VGND VGND VPWR VPWR _109_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_11.sky130_fd_sc_hd__buf_4_0_ mux_left_track_11.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _076_/A sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold4/X VGND VGND VPWR VPWR hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_27_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_19.mux_l1_in_0_ input13/X input6/X hold26/A VGND VGND VPWR VPWR
+ mux_bottom_track_19.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_bottom_track_21.mux_l1_in_0_ input14/X input7/X hold6/A VGND VGND VPWR VPWR mux_bottom_track_21.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_29.mux_l2_in_0__137 VGND VGND VPWR VPWR mux_bottom_track_29.mux_l2_in_0_/A0
+ mux_bottom_track_29.mux_l2_in_0__137/LO sky130_fd_sc_hd__conb_1
XFILLER_24_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_090_ _090_/A VGND VGND VPWR VPWR _090_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_5.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _093_/A sky130_fd_sc_hd__clkbuf_1
Xinput4 bottom_left_grid_pin_44_ VGND VGND VPWR VPWR input4/X sky130_fd_sc_hd__clkbuf_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_bottom_track_5.mux_l1_in_0_ input3/X input10/X mux_bottom_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_11.mux_l2_in_0__108 VGND VGND VPWR VPWR mux_left_track_11.mux_l2_in_0_/A0
+ mux_left_track_11.mux_l2_in_0__108/LO sky130_fd_sc_hd__conb_1
XFILLER_27_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_073_ _073_/A VGND VGND VPWR VPWR _073_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_105 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput51 chany_bottom_in[9] VGND VGND VPWR VPWR input51/X sky130_fd_sc_hd__clkbuf_1
Xinput40 chany_bottom_in[17] VGND VGND VPWR VPWR input40/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input26_A chanx_left_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_108_ _108_/A VGND VGND VPWR VPWR _108_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_1__107 VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/A0
+ mux_left_track_1.mux_l2_in_1__107/LO sky130_fd_sc_hd__conb_1
XFILLER_1_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_33.sky130_fd_sc_hd__buf_4_0_ mux_left_track_33.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _087_/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold32/X VGND VGND VPWR VPWR mux_bottom_track_5.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_24_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput5 bottom_left_grid_pin_45_ VGND VGND VPWR VPWR input5/X sky130_fd_sc_hd__clkbuf_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_27.sky130_fd_sc_hd__buf_4_0_ mux_left_track_27.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _084_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_19.mux_l2_in_0__112 VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/A0
+ mux_left_track_19.mux_l2_in_0__112/LO sky130_fd_sc_hd__conb_1
XFILLER_2_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_072_ _072_/A VGND VGND VPWR VPWR _072_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input56_A left_bottom_grid_pin_38_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_18_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_117 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput41 chany_bottom_in[18] VGND VGND VPWR VPWR input41/X sky130_fd_sc_hd__clkbuf_1
Xinput52 left_bottom_grid_pin_34_ VGND VGND VPWR VPWR input52/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput30 chanx_left_in[8] VGND VGND VPWR VPWR input30/X sky130_fd_sc_hd__clkbuf_1
XFILLER_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input19_A chanx_left_in[16] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_107_ _107_/A VGND VGND VPWR VPWR _107_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_23.mux_l2_in_0__114 VGND VGND VPWR VPWR mux_left_track_23.mux_l2_in_0_/A0
+ mux_left_track_23.mux_l2_in_0__114/LO sky130_fd_sc_hd__conb_1
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold19/X VGND VGND VPWR VPWR hold34/A sky130_fd_sc_hd__dfxtp_1
XFILLER_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput6 bottom_left_grid_pin_46_ VGND VGND VPWR VPWR input6/X sky130_fd_sc_hd__clkbuf_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_3.mux_l1_in_1__A0 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold50/X VGND VGND VPWR VPWR hold55/A sky130_fd_sc_hd__dfxtp_1
X_071_ _071_/A VGND VGND VPWR VPWR _071_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input49_A chany_bottom_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l2_in_0_ mux_left_track_17.mux_l2_in_0_/A0 mux_left_track_17.mux_l1_in_0_/X
+ hold56/A VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput31 chanx_left_in[9] VGND VGND VPWR VPWR input31/X sky130_fd_sc_hd__clkbuf_1
Xinput20 chanx_left_in[17] VGND VGND VPWR VPWR _107_/A sky130_fd_sc_hd__clkbuf_1
Xinput53 left_bottom_grid_pin_35_ VGND VGND VPWR VPWR input53/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 chany_bottom_in[19] VGND VGND VPWR VPWR input42/X sky130_fd_sc_hd__clkbuf_1
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_106_ _106_/A VGND VGND VPWR VPWR _106_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_9.mux_l2_in_0_ mux_left_track_9.mux_l1_in_1_/X mux_left_track_9.mux_l1_in_0_/X
+ hold1/A VGND VGND VPWR VPWR mux_left_track_9.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input31_A chanx_left_in[9] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_1_ mux_left_track_9.mux_l1_in_1_/A0 input59/X mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold8/X VGND VGND VPWR VPWR hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput7 bottom_left_grid_pin_47_ VGND VGND VPWR VPWR input7/X sky130_fd_sc_hd__clkbuf_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold36/X VGND VGND VPWR VPWR hold50/A sky130_fd_sc_hd__dfxtp_1
X_070_ _070_/A VGND VGND VPWR VPWR _070_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold26/X VGND VGND VPWR VPWR hold12/A sky130_fd_sc_hd__dfxtp_1
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput32 chany_bottom_in[0] VGND VGND VPWR VPWR input32/X sky130_fd_sc_hd__clkbuf_1
Xinput54 left_bottom_grid_pin_36_ VGND VGND VPWR VPWR input54/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput10 bottom_right_grid_pin_1_ VGND VGND VPWR VPWR input10/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput43 chany_bottom_in[1] VGND VGND VPWR VPWR input43/X sky130_fd_sc_hd__clkbuf_1
Xinput21 chanx_left_in[18] VGND VGND VPWR VPWR _108_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_105_ _105_/A VGND VGND VPWR VPWR _105_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold24/X VGND VGND VPWR VPWR hold45/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.mux_l1_in_0_ input55/X input49/X hold33/A VGND VGND VPWR VPWR mux_left_track_17.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_29.mux_l2_in_0_ mux_left_track_29.mux_l2_in_0_/A0 mux_left_track_29.mux_l1_in_0_/X
+ hold45/A VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_input24_A chanx_left_in[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_200 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_17_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_31.mux_l2_in_0_ mux_left_track_31.mux_l2_in_0_/A0 mux_left_track_31.mux_l1_in_0_/X
+ hold48/A VGND VGND VPWR VPWR mux_left_track_31.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_9.mux_l1_in_0_ input60/X input45/X mux_left_track_9.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_13.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _097_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_24_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_14_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 bottom_left_grid_pin_48_ VGND VGND VPWR VPWR input8/X sky130_fd_sc_hd__clkbuf_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_25_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l3_in_0_ mux_bottom_track_1.mux_l2_in_1_/X mux_bottom_track_1.mux_l2_in_0_/X
+ hold9/A VGND VGND VPWR VPWR mux_bottom_track_1.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_17.mux_l1_in_0__A0 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input54_A left_bottom_grid_pin_36_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold27/X VGND VGND VPWR VPWR hold26/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput33 chany_bottom_in[10] VGND VGND VPWR VPWR input33/X sky130_fd_sc_hd__clkbuf_1
Xinput55 left_bottom_grid_pin_37_ VGND VGND VPWR VPWR input55/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput44 chany_bottom_in[2] VGND VGND VPWR VPWR input44/X sky130_fd_sc_hd__clkbuf_1
Xinput11 ccff_head VGND VGND VPWR VPWR input11/X sky130_fd_sc_hd__clkbuf_1
Xinput22 chanx_left_in[19] VGND VGND VPWR VPWR _109_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold3/X VGND VGND VPWR VPWR hold24/A sky130_fd_sc_hd__dfxtp_1
XFILLER_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_1.mux_l2_in_1_ mux_bottom_track_1.mux_l2_in_1_/A0 mux_bottom_track_1.mux_l1_in_2_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
X_104_ _104_/A VGND VGND VPWR VPWR _104_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_35.mux_l2_in_0__121 VGND VGND VPWR VPWR mux_left_track_35.mux_l2_in_0_/A0
+ mux_left_track_35.mux_l2_in_0__121/LO sky130_fd_sc_hd__conb_1
XFILLER_4_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input17_A chanx_left_in[14] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_1.mux_l1_in_2_ input23/X input9/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input9_A bottom_left_grid_pin_49_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_29.mux_l1_in_0_ input53/X input36/X hold24/A VGND VGND VPWR VPWR mux_left_track_29.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_31.mux_l1_in_0_ input54/X input37/X hold42/A VGND VGND VPWR VPWR mux_left_track_31.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput9 bottom_left_grid_pin_49_ VGND VGND VPWR VPWR input9/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold57/X VGND VGND VPWR VPWR hold17/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_25.mux_l1_in_0__A0 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_15.mux_l2_in_0_ mux_bottom_track_15.mux_l2_in_0_/A0 mux_bottom_track_15.mux_l1_in_0_/X
+ hold22/A VGND VGND VPWR VPWR mux_bottom_track_15.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input47_A chany_bottom_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput56 left_bottom_grid_pin_38_ VGND VGND VPWR VPWR input56/X sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 chany_bottom_in[11] VGND VGND VPWR VPWR input34/X sky130_fd_sc_hd__clkbuf_1
Xinput45 chany_bottom_in[3] VGND VGND VPWR VPWR input45/X sky130_fd_sc_hd__clkbuf_1
Xinput12 chanx_left_in[0] VGND VGND VPWR VPWR _110_/A sky130_fd_sc_hd__clkbuf_1
Xinput23 chanx_left_in[1] VGND VGND VPWR VPWR input23/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_29.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_29.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _105_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_20_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_103_ _103_/A VGND VGND VPWR VPWR _103_/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_1.mux_l2_in_0_ mux_bottom_track_1.mux_l1_in_1_/X mux_bottom_track_1.mux_l1_in_0_/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_22_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xhold1 hold1/A VGND VGND VPWR VPWR hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_mux_left_track_5.mux_l1_in_2__A1 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_1__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xmux_bottom_track_1.mux_l1_in_1_ input7/X input5/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_33.mux_l1_in_0__A0 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_27.mux_l2_in_0__136 VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/A0
+ mux_bottom_track_27.mux_l2_in_0__136/LO sky130_fd_sc_hd__conb_1
XFILLER_30_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_3.mux_l1_in_1_/S VGND VGND VPWR VPWR hold57/A sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_1.mux_l2_in_1__127 VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/A0
+ mux_bottom_track_1.mux_l2_in_1__127/LO sky130_fd_sc_hd__conb_1
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput100 _098_/X VGND VGND VPWR VPWR chany_bottom_out[7] sky130_fd_sc_hd__buf_2
XFILLER_11_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput13 chanx_left_in[10] VGND VGND VPWR VPWR input13/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_15.mux_l1_in_0_ input30/X input4/X hold14/A VGND VGND VPWR VPWR
+ mux_bottom_track_15.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xinput24 chanx_left_in[2] VGND VGND VPWR VPWR input24/X sky130_fd_sc_hd__clkbuf_1
Xinput57 left_bottom_grid_pin_39_ VGND VGND VPWR VPWR input57/X sky130_fd_sc_hd__clkbuf_2
Xinput46 chany_bottom_in[4] VGND VGND VPWR VPWR input46/X sky130_fd_sc_hd__clkbuf_1
Xinput35 chany_bottom_in[12] VGND VGND VPWR VPWR input35/X sky130_fd_sc_hd__clkbuf_1
Xmux_bottom_track_27.mux_l2_in_0_ mux_bottom_track_27.mux_l2_in_0_/A0 mux_bottom_track_27.mux_l1_in_0_/X
+ hold7/A VGND VGND VPWR VPWR mux_bottom_track_27.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_122 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_20_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_1.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _091_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_11_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_102_ _102_/A VGND VGND VPWR VPWR _102_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold2 hold2/A VGND VGND VPWR VPWR hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_1.mux_l1_in_0_ input3/X input10/X mux_bottom_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input22_A chanx_left_in[19] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold54/X VGND VGND VPWR VPWR hold46/A sky130_fd_sc_hd__dfxtp_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold15/X VGND VGND VPWR VPWR mux_left_track_3.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_7.sky130_fd_sc_hd__buf_4_0_ mux_left_track_7.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _074_/A sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_17.mux_l2_in_0__111 VGND VGND VPWR VPWR mux_left_track_17.mux_l2_in_0_/A0
+ mux_left_track_17.mux_l2_in_0__111/LO sky130_fd_sc_hd__conb_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput101 _099_/X VGND VGND VPWR VPWR chany_bottom_out[8] sky130_fd_sc_hd__buf_2
Xclkbuf_0_mem_bottom_track_1.prog_clk prog_clk_0_FTB00/X VGND VGND VPWR VPWR clkbuf_0_mem_bottom_track_1.prog_clk/X
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput36 chany_bottom_in[13] VGND VGND VPWR VPWR input36/X sky130_fd_sc_hd__clkbuf_1
Xinput25 chanx_left_in[3] VGND VGND VPWR VPWR input25/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput14 chanx_left_in[11] VGND VGND VPWR VPWR input14/X sky130_fd_sc_hd__clkbuf_1
Xinput47 chany_bottom_in[5] VGND VGND VPWR VPWR input47/X sky130_fd_sc_hd__clkbuf_1
Xinput58 left_bottom_grid_pin_40_ VGND VGND VPWR VPWR input58/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_9.mux_l1_in_1_/S VGND VGND VPWR VPWR hold1/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_101_ _101_/A VGND VGND VPWR VPWR _101_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_2__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_input52_A left_bottom_grid_pin_34_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_23.sky130_fd_sc_hd__buf_4_0_ mux_left_track_23.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _082_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_27.mux_l1_in_0_ input17/X input2/X hold23/A VGND VGND VPWR VPWR
+ mux_bottom_track_27.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold3 hold3/A VGND VGND VPWR VPWR hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_13_207 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_17.sky130_fd_sc_hd__buf_4_0_ mux_left_track_17.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _079_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input15_A chanx_left_in[12] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.mux_l2_in_0__113 VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/A0
+ mux_left_track_21.mux_l2_in_0__113/LO sky130_fd_sc_hd__conb_1
XFILLER_8_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_left_track_5.mux_l3_in_0_ mux_left_track_5.mux_l2_in_1_/X mux_left_track_5.mux_l2_in_0_/X
+ hold58/A VGND VGND VPWR VPWR mux_left_track_5.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input7_A bottom_left_grid_pin_47_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold37/X VGND VGND VPWR VPWR hold54/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_29_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_27_129 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_121 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_1_ mux_left_track_5.mux_l2_in_1_/A0 mux_left_track_5.mux_l1_in_2_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput102 _100_/X VGND VGND VPWR VPWR chany_bottom_out[9] sky130_fd_sc_hd__buf_2
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 chanx_left_in[4] VGND VGND VPWR VPWR input26/X sky130_fd_sc_hd__clkbuf_1
Xinput59 left_bottom_grid_pin_41_ VGND VGND VPWR VPWR input59/X sky130_fd_sc_hd__clkbuf_2
Xinput37 chany_bottom_in[14] VGND VGND VPWR VPWR input37/X sky130_fd_sc_hd__clkbuf_1
Xinput48 chany_bottom_in[6] VGND VGND VPWR VPWR input48/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput15 chanx_left_in[12] VGND VGND VPWR VPWR input15/X sky130_fd_sc_hd__clkbuf_1
Xmem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold38/X VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_100_ _100_/A VGND VGND VPWR VPWR _100_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input45_A chany_bottom_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_2_ input59/X input57/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_41 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_33_85 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold4 hold4/A VGND VGND VPWR VPWR hold4/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_13_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_13.mux_l2_in_0_ mux_left_track_13.mux_l2_in_0_/A0 mux_left_track_13.mux_l1_in_0_/X
+ hold37/A VGND VGND VPWR VPWR mux_left_track_13.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_64 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_39.sky130_fd_sc_hd__buf_4_0_ mux_left_track_39.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _090_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_29_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_32_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_5.mux_l2_in_0_ mux_left_track_5.mux_l1_in_1_/X mux_left_track_5.mux_l1_in_0_/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_11_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xinput38 chany_bottom_in[15] VGND VGND VPWR VPWR input38/X sky130_fd_sc_hd__clkbuf_1
Xinput27 chanx_left_in[5] VGND VGND VPWR VPWR input27/X sky130_fd_sc_hd__clkbuf_1
Xinput16 chanx_left_in[13] VGND VGND VPWR VPWR input16/X sky130_fd_sc_hd__clkbuf_1
Xinput49 chany_bottom_in[7] VGND VGND VPWR VPWR input49/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input38_A chany_bottom_in[15] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_5.mux_l1_in_1_ input55/X input53/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold25/X VGND VGND VPWR VPWR hold41/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_25.mux_l1_in_1__135 VGND VGND VPWR VPWR mux_bottom_track_25.mux_l1_in_1_/A0
+ mux_bottom_track_25.mux_l1_in_1__135/LO sky130_fd_sc_hd__conb_1
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold52/X VGND VGND VPWR VPWR hold31/A sky130_fd_sc_hd__dfxtp_1
XFILLER_33_97 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold5 hold5/A VGND VGND VPWR VPWR hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_22_209 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l2_in_1_/S VGND VGND VPWR VPWR hold9/A sky130_fd_sc_hd__dfxtp_1
XFILLER_14_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_input20_A chanx_left_in[17] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_13.mux_l2_in_0__129 VGND VGND VPWR VPWR mux_bottom_track_13.mux_l2_in_0_/A0
+ mux_bottom_track_13.mux_l2_in_0__129/LO sky130_fd_sc_hd__conb_1
Xmux_left_track_13.mux_l1_in_0_ input53/X input47/X hold2/A VGND VGND VPWR VPWR mux_left_track_13.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_142 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmux_left_track_25.mux_l2_in_0_ mux_left_track_25.mux_l1_in_1_/X mux_left_track_25.mux_l1_in_0_/X
+ hold5/A VGND VGND VPWR VPWR mux_left_track_25.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput39 chany_bottom_in[16] VGND VGND VPWR VPWR input39/X sky130_fd_sc_hd__clkbuf_1
Xinput28 chanx_left_in[6] VGND VGND VPWR VPWR input28/X sky130_fd_sc_hd__clkbuf_1
Xinput17 chanx_left_in[14] VGND VGND VPWR VPWR input17/X sky130_fd_sc_hd__clkbuf_1
XFILLER_9_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold30/X VGND VGND VPWR VPWR hold25/A sky130_fd_sc_hd__dfxtp_1
Xmux_left_track_5.mux_l1_in_0_ input60/X input43/X mux_left_track_5.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_1_ mux_left_track_25.mux_l1_in_1_/A0 input59/X mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
X_089_ _089_/A VGND VGND VPWR VPWR _089_/X sky130_fd_sc_hd__clkbuf_1
Xmux_left_track_33.mux_l2_in_0__120 VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/A0
+ mux_left_track_33.mux_l2_in_0__120/LO sky130_fd_sc_hd__conb_1
XFILLER_17_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold48/X VGND VGND VPWR VPWR hold52/A sky130_fd_sc_hd__dfxtp_1
XFILLER_3_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input50_A chany_bottom_in[8] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold6 hold6/A VGND VGND VPWR VPWR hold6/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_30_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_1.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_bottom_track_1.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
Xmem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X
+ hold18/X VGND VGND VPWR VPWR hold11/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_39.mux_l1_in_0__A0 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_4__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_input13_A chanx_left_in[10] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_140 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold35/X VGND VGND VPWR VPWR output62/A sky130_fd_sc_hd__dfxtp_1
XANTENNA_input5_A bottom_left_grid_pin_45_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_154 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR hold20/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_113 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 chanx_left_in[15] VGND VGND VPWR VPWR input18/X sky130_fd_sc_hd__clkbuf_1
XFILLER_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput29 chanx_left_in[7] VGND VGND VPWR VPWR input29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_25.mux_l1_in_0_ input60/X input34/X mux_left_track_25.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
X_088_ _088_/A VGND VGND VPWR VPWR _088_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_6_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_left_track_37.mux_l2_in_0_ mux_left_track_37.mux_l2_in_0_/A0 mux_left_track_37.mux_l1_in_0_/X
+ hold40/A VGND VGND VPWR VPWR mux_left_track_37.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
Xmux_left_track_7.mux_l2_in_1__125 VGND VGND VPWR VPWR mux_left_track_7.mux_l2_in_1_/A0
+ mux_left_track_7.mux_l2_in_1__125/LO sky130_fd_sc_hd__conb_1
XFILLER_3_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input43_A chany_bottom_in[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold7 hold7/A VGND VGND VPWR VPWR hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xmux_bottom_track_11.mux_l2_in_0_ mux_bottom_track_11.mux_l2_in_0_/A0 mux_bottom_track_11.mux_l1_in_0_/X
+ hold8/A VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ input11/X VGND VGND VPWR VPWR mux_bottom_track_1.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
Xmux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_25.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _103_/A sky130_fd_sc_hd__clkbuf_1
Xmem_bottom_track_29.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X
+ hold7/X VGND VGND VPWR VPWR hold18/A sky130_fd_sc_hd__dfxtp_1
XFILLER_5_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_152 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ hold40/X VGND VGND VPWR VPWR hold35/A sky130_fd_sc_hd__dfxtp_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_7.mux_l3_in_0_ mux_bottom_track_7.mux_l2_in_1_/X mux_bottom_track_7.mux_l2_in_0_/X
+ hold20/A VGND VGND VPWR VPWR mux_bottom_track_7.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_177 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_19.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _100_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_1_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ mux_bottom_track_7.mux_l1_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_23_125 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput19 chanx_left_in[16] VGND VGND VPWR VPWR _106_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_1_ mux_bottom_track_7.mux_l2_in_1_/A0 input26/X mux_bottom_track_7.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_22_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_087_ _087_/A VGND VGND VPWR VPWR _087_/X sky130_fd_sc_hd__clkbuf_1
Xhold8 hold8/A VGND VGND VPWR VPWR hold8/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xclkbuf_3_5__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_5__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XANTENNA_input36_A chany_bottom_in[13] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_37.mux_l1_in_0_ input57/X input40/X hold21/A VGND VGND VPWR VPWR mux_left_track_37.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_14_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmux_bottom_track_11.mux_l1_in_0_ input28/X input2/X hold29/A VGND VGND VPWR VPWR
+ mux_bottom_track_11.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_6_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_15.mux_l2_in_0__110 VGND VGND VPWR VPWR mux_left_track_15.mux_l2_in_0_/A0
+ mux_left_track_15.mux_l2_in_0__110/LO sky130_fd_sc_hd__conb_1
XFILLER_6_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_23.mux_l2_in_0_ mux_bottom_track_23.mux_l2_in_0_/A0 mux_bottom_track_23.mux_l1_in_0_/X
+ hold41/A VGND VGND VPWR VPWR mux_bottom_track_23.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ hold44/X VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
XFILLER_23_137 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.mux_l2_in_0_ mux_bottom_track_7.mux_l1_in_1_/X mux_bottom_track_7.mux_l1_in_0_/X
+ mux_bottom_track_7.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_7.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_8_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_086_ _086_/A VGND VGND VPWR VPWR _086_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_3.sky130_fd_sc_hd__buf_4_0_ mux_left_track_3.mux_l3_in_0_/X VGND VGND
+ VPWR VPWR _072_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_21.mux_l1_in_0__A0 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_57 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold9 hold9/A VGND VGND VPWR VPWR hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input29_A chanx_left_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_7.mux_l1_in_1_ input8/X input6/X mux_bottom_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input11_A ccff_head VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput90 _107_/X VGND VGND VPWR VPWR chany_bottom_out[16] sky130_fd_sc_hd__buf_2
XFILLER_23_149 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mux_left_track_1.mux_l1_in_2__A1 input57/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input3_A bottom_left_grid_pin_43_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_13.sky130_fd_sc_hd__buf_4_0_ mux_left_track_13.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _077_/A sky130_fd_sc_hd__clkbuf_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input59_A left_bottom_grid_pin_41_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_23.mux_l1_in_0_ input15/X input8/X hold25/A VGND VGND VPWR VPWR
+ mux_bottom_track_23.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold14/X VGND VGND VPWR VPWR hold22/A sky130_fd_sc_hd__dfxtp_1
XFILLER_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_171 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_9.mux_l1_in_1__126 VGND VGND VPWR VPWR mux_left_track_9.mux_l1_in_1_/A0
+ mux_left_track_9.mux_l1_in_1__126/LO sky130_fd_sc_hd__conb_1
XFILLER_9_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_6__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_3__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_25.mux_l1_in_1_/S VGND VGND VPWR VPWR hold5/A sky130_fd_sc_hd__dfxtp_1
X_085_ _085_/A VGND VGND VPWR VPWR _085_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_26_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_21.mux_l1_in_0__A1 input51/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_69 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.mux_l3_in_0_ mux_left_track_1.mux_l2_in_1_/X mux_left_track_1.mux_l2_in_0_/X
+ hold15/A VGND VGND VPWR VPWR mux_left_track_1.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_33_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_bottom_track_7.mux_l1_in_0_ input4/X input2/X mux_bottom_track_7.mux_l1_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_7.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_7.mux_l3_in_0_/X VGND
+ VGND VPWR VPWR _094_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_input41_A chany_bottom_in[18] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_1.mux_l2_in_1_ mux_left_track_1.mux_l2_in_1_/A0 mux_left_track_1.mux_l1_in_2_/X
+ hold59/A VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_1.mux_l1_in_2_ input59/X input57/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_2_/X sky130_fd_sc_hd__mux2_1
Xoutput91 _108_/X VGND VGND VPWR VPWR chany_bottom_out[17] sky130_fd_sc_hd__buf_2
Xoutput80 _078_/X VGND VGND VPWR VPWR chanx_left_out[7] sky130_fd_sc_hd__buf_2
XFILLER_31_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_6__f_mem_bottom_track_1.prog_clk/X
+ hold34/X VGND VGND VPWR VPWR hold14/A sky130_fd_sc_hd__dfxtp_1
XFILLER_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_183 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmux_left_track_35.sky130_fd_sc_hd__buf_4_0_ mux_left_track_35.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _088_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold55/X VGND VGND VPWR VPWR mux_left_track_25.mux_l1_in_1_/S sky130_fd_sc_hd__dfxtp_1
X_084_ _084_/A VGND VGND VPWR VPWR _084_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_5.mux_l1_in_1__A0 input55/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_29.sky130_fd_sc_hd__buf_4_0_ mux_left_track_29.mux_l2_in_0_/X VGND
+ VGND VPWR VPWR _085_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_28_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_input34_A chany_bottom_in[11] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l2_in_0_ mux_left_track_1.mux_l1_in_1_/X mux_left_track_1.mux_l1_in_0_/X
+ hold59/A VGND VGND VPWR VPWR mux_left_track_1.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_4_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_7__f_mem_bottom_track_1.prog_clk clkbuf_0_mem_bottom_track_1.prog_clk/X
+ VGND VGND VPWR VPWR clkbuf_3_7__f_mem_bottom_track_1.prog_clk/X sky130_fd_sc_hd__clkbuf_16
Xmux_bottom_track_11.mux_l2_in_0__128 VGND VGND VPWR VPWR mux_bottom_track_11.mux_l2_in_0_/A0
+ mux_bottom_track_11.mux_l2_in_0__128/LO sky130_fd_sc_hd__conb_1
XFILLER_17_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_1.mux_l1_in_1_ input55/X input53/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_1_/X sky130_fd_sc_hd__mux2_1
XFILLER_25_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_81 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput70 _087_/X VGND VGND VPWR VPWR chanx_left_out[16] sky130_fd_sc_hd__buf_2
Xoutput92 _109_/X VGND VGND VPWR VPWR chany_bottom_out[18] sky130_fd_sc_hd__buf_2
Xoutput81 _079_/X VGND VGND VPWR VPWR chanx_left_out[8] sky130_fd_sc_hd__buf_2
XFILLER_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_195 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_083_ _083_/A VGND VGND VPWR VPWR _083_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_15_202 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_23_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_205 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_19.mux_l2_in_0_ mux_left_track_19.mux_l2_in_0_/A0 mux_left_track_19.mux_l1_in_0_/X
+ hold51/A VGND VGND VPWR VPWR mux_left_track_19.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_input27_A chanx_left_in[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_21.mux_l2_in_0_ mux_left_track_21.mux_l2_in_0_/A0 mux_left_track_21.mux_l1_in_0_/X
+ hold36/A VGND VGND VPWR VPWR mux_left_track_21.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmux_bottom_track_19.mux_l2_in_0__132 VGND VGND VPWR VPWR mux_bottom_track_19.mux_l2_in_0_/A0
+ mux_bottom_track_19.mux_l2_in_0__132/LO sky130_fd_sc_hd__conb_1
XFILLER_17_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_left_track_1.mux_l1_in_0_ input60/X input42/X mux_left_track_1.mux_l1_in_2_/S
+ VGND VGND VPWR VPWR mux_left_track_1.mux_l1_in_0_/X sky130_fd_sc_hd__mux2_1
Xoutput93 _110_/X VGND VGND VPWR VPWR chany_bottom_out[19] sky130_fd_sc_hd__buf_2
Xoutput82 _080_/X VGND VGND VPWR VPWR chanx_left_out[9] sky130_fd_sc_hd__buf_2
Xoutput71 _088_/X VGND VGND VPWR VPWR chanx_left_out[17] sky130_fd_sc_hd__buf_2
XFILLER_31_93 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_141 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input1_A SC_IN_BOT VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l2_in_1_/S VGND VGND VPWR VPWR hold58/A sky130_fd_sc_hd__dfxtp_1
XFILLER_10_199 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
X_082_ _082_/A VGND VGND VPWR VPWR _082_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_input57_A left_bottom_grid_pin_39_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_5.mux_l2_in_1__124 VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/A0
+ mux_left_track_5.mux_l2_in_1__124/LO sky130_fd_sc_hd__conb_1
XFILLER_15_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_23.mux_l2_in_0__134 VGND VGND VPWR VPWR mux_bottom_track_23.mux_l2_in_0_/A0
+ mux_bottom_track_23.mux_l2_in_0__134/LO sky130_fd_sc_hd__conb_1
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_mux_left_track_19.mux_l1_in_0__A0 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_169 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_1__f_mem_bottom_track_1.prog_clk/X
+ hold53/X VGND VGND VPWR VPWR hold43/A sky130_fd_sc_hd__dfxtp_1
Xhold60 hold60/A VGND VGND VPWR VPWR hold60/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmux_left_track_19.mux_l1_in_0_ input56/X input50/X hold47/A VGND VGND VPWR VPWR mux_left_track_19.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_17_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_109 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_mux_left_track_9.mux_l1_in_0__A0 input60/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput61 _070_/X VGND VGND VPWR VPWR SC_OUT_BOT sky130_fd_sc_hd__buf_2
Xoutput83 _091_/X VGND VGND VPWR VPWR chany_bottom_out[0] sky130_fd_sc_hd__buf_2
Xoutput94 _092_/X VGND VGND VPWR VPWR chany_bottom_out[1] sky130_fd_sc_hd__buf_2
Xmux_left_track_21.mux_l1_in_0_ input57/X input51/X hold39/A VGND VGND VPWR VPWR mux_left_track_21.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
Xoutput72 _089_/X VGND VGND VPWR VPWR chanx_left_out[18] sky130_fd_sc_hd__buf_2
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmux_left_track_33.mux_l2_in_0_ mux_left_track_33.mux_l2_in_0_/A0 mux_left_track_33.mux_l1_in_0_/X
+ hold31/A VGND VGND VPWR VPWR mux_left_track_33.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_153 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_22_197 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
Xmux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_21.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _101_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_13_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_0__f_mem_bottom_track_1.prog_clk/X
+ mux_left_track_5.mux_l1_in_2_/S VGND VGND VPWR VPWR mux_left_track_5.mux_l2_in_1_/S
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_10_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_081_ _081_/A VGND VGND VPWR VPWR _081_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_18_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_ mux_bottom_track_15.mux_l2_in_0_/X
+ VGND VGND VPWR VPWR _098_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_17_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l3_in_0_ mux_bottom_track_3.mux_l2_in_1_/X mux_bottom_track_3.mux_l2_in_0_/X
+ hold32/A VGND VGND VPWR VPWR mux_bottom_track_3.mux_l3_in_0_/X sky130_fd_sc_hd__mux2_1
XANTENNA_mux_left_track_19.mux_l1_in_0__A1 input50/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold1/X VGND VGND VPWR VPWR hold53/A sky130_fd_sc_hd__dfxtp_1
XFILLER_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_input32_A chany_bottom_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold50 hold50/A VGND VGND VPWR VPWR hold50/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l2_in_1_ mux_bottom_track_3.mux_l2_in_1_/A0 input24/X mux_bottom_track_3.mux_l2_in_1_/S
+ VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_1_/X sky130_fd_sc_hd__mux2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_181 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_1_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput73 _090_/X VGND VGND VPWR VPWR chanx_left_out[19] sky130_fd_sc_hd__buf_2
Xoutput95 _093_/X VGND VGND VPWR VPWR chany_bottom_out[2] sky130_fd_sc_hd__buf_2
Xoutput84 _101_/X VGND VGND VPWR VPWR chany_bottom_out[10] sky130_fd_sc_hd__buf_2
Xoutput62 output62/A VGND VGND VPWR VPWR ccff_tail sky130_fd_sc_hd__buf_2
XFILLER_16_151 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_165 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_ clkbuf_3_2__f_mem_bottom_track_1.prog_clk/X
+ hold33/X VGND VGND VPWR VPWR hold56/A sky130_fd_sc_hd__dfxtp_1
XFILLER_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_ clkbuf_3_4__f_mem_bottom_track_1.prog_clk/X
+ hold17/X VGND VGND VPWR VPWR mux_left_track_5.mux_l1_in_2_/S sky130_fd_sc_hd__dfxtp_1
XANTENNA_mux_left_track_35.mux_l1_in_0__A0 input56/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_080_ _080_/A VGND VGND VPWR VPWR _080_/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__108__A _108_/A VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_left_track_33.mux_l1_in_0_ input55/X input38/X hold52/A VGND VGND VPWR VPWR mux_left_track_33.mux_l1_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_5_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_mux_left_track_7.mux_l2_in_1__A1 input58/X VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmux_bottom_track_17.mux_l2_in_0_ mux_bottom_track_17.mux_l2_in_0_/A0 mux_bottom_track_17.mux_l1_in_0_/X
+ hold27/A VGND VGND VPWR VPWR mux_bottom_track_17.mux_l2_in_0_/X sky130_fd_sc_hd__mux2_1
XFILLER_2_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_left_track_29.mux_l2_in_0__117 VGND VGND VPWR VPWR mux_left_track_29.mux_l2_in_0_/A0
+ mux_left_track_29.mux_l2_in_0__117/LO sky130_fd_sc_hd__conb_1
XFILLER_7_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_116 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_4_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold40 hold40/A VGND VGND VPWR VPWR hold40/X sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA_input25_A chanx_left_in[3] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold51 hold51/A VGND VGND VPWR VPWR hold51/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xmux_bottom_track_3.mux_l2_in_0_ mux_bottom_track_3.mux_l1_in_1_/X mux_bottom_track_3.mux_l1_in_0_/X
+ mux_bottom_track_3.mux_l2_in_1_/S VGND VGND VPWR VPWR mux_bottom_track_3.mux_l2_in_0_/X
+ sky130_fd_sc_hd__mux2_1
XFILLER_19_193 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_15_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput96 _094_/X VGND VGND VPWR VPWR chany_bottom_out[3] sky130_fd_sc_hd__buf_2
Xoutput85 _102_/X VGND VGND VPWR VPWR chany_bottom_out[11] sky130_fd_sc_hd__buf_2
Xoutput63 _071_/X VGND VGND VPWR VPWR chanx_left_out[0] sky130_fd_sc_hd__buf_2
Xoutput74 _072_/X VGND VGND VPWR VPWR chanx_left_out[1] sky130_fd_sc_hd__buf_2
XFILLER_16_163 VGND VPWR VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_31_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

