magic
tech sky130A
magscale 1 2
timestamp 1650891882
<< viali >>
rect 1593 17289 1627 17323
rect 1961 17289 1995 17323
rect 2329 17289 2363 17323
rect 2697 17289 2731 17323
rect 3157 17289 3191 17323
rect 4169 17289 4203 17323
rect 4997 17289 5031 17323
rect 6101 17289 6135 17323
rect 7481 17289 7515 17323
rect 7849 17289 7883 17323
rect 9965 17221 9999 17255
rect 11713 17221 11747 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 2973 17153 3007 17187
rect 3617 17153 3651 17187
rect 3793 17153 3827 17187
rect 4353 17153 4387 17187
rect 4445 17153 4479 17187
rect 4813 17153 4847 17187
rect 5181 17153 5215 17187
rect 5549 17153 5583 17187
rect 5917 17153 5951 17187
rect 6401 17153 6435 17187
rect 6929 17153 6963 17187
rect 7389 17153 7423 17187
rect 8217 17153 8251 17187
rect 9597 17153 9631 17187
rect 10057 17153 10091 17187
rect 11897 17153 11931 17187
rect 13093 17153 13127 17187
rect 14372 17153 14406 17187
rect 7573 17085 7607 17119
rect 8309 17085 8343 17119
rect 8401 17085 8435 17119
rect 9781 17085 9815 17119
rect 11069 17085 11103 17119
rect 11345 17085 11379 17119
rect 11529 17085 11563 17119
rect 12173 17085 12207 17119
rect 12449 17085 12483 17119
rect 13369 17085 13403 17119
rect 14105 17085 14139 17119
rect 3433 17017 3467 17051
rect 4629 17017 4663 17051
rect 6561 17017 6595 17051
rect 8769 17017 8803 17051
rect 15485 17017 15519 17051
rect 3985 16949 4019 16983
rect 5365 16949 5399 16983
rect 5733 16949 5767 16983
rect 6745 16949 6779 16983
rect 7021 16949 7055 16983
rect 8953 16949 8987 16983
rect 10425 16949 10459 16983
rect 12081 16949 12115 16983
rect 15577 16949 15611 16983
rect 1869 16745 1903 16779
rect 2237 16745 2271 16779
rect 4169 16745 4203 16779
rect 4445 16745 4479 16779
rect 4905 16745 4939 16779
rect 8309 16745 8343 16779
rect 10701 16745 10735 16779
rect 15577 16745 15611 16779
rect 1501 16677 1535 16711
rect 2881 16677 2915 16711
rect 3617 16677 3651 16711
rect 3893 16677 3927 16711
rect 6561 16609 6595 16643
rect 6653 16609 6687 16643
rect 8953 16609 8987 16643
rect 11437 16609 11471 16643
rect 11621 16609 11655 16643
rect 13461 16609 13495 16643
rect 14105 16609 14139 16643
rect 1685 16541 1719 16575
rect 2053 16541 2087 16575
rect 2421 16541 2455 16575
rect 2513 16541 2547 16575
rect 3065 16541 3099 16575
rect 3157 16541 3191 16575
rect 3433 16541 3467 16575
rect 3985 16541 4019 16575
rect 4629 16541 4663 16575
rect 4721 16541 4755 16575
rect 4997 16541 5031 16575
rect 5365 16541 5399 16575
rect 6929 16541 6963 16575
rect 9321 16541 9355 16575
rect 11161 16541 11195 16575
rect 13645 16541 13679 16575
rect 6009 16473 6043 16507
rect 7174 16473 7208 16507
rect 8677 16473 8711 16507
rect 9137 16473 9171 16507
rect 9588 16473 9622 16507
rect 11805 16473 11839 16507
rect 13194 16473 13228 16507
rect 14372 16473 14406 16507
rect 2697 16405 2731 16439
rect 3341 16405 3375 16439
rect 5181 16405 5215 16439
rect 6101 16405 6135 16439
rect 6469 16405 6503 16439
rect 8585 16405 8619 16439
rect 10793 16405 10827 16439
rect 11253 16405 11287 16439
rect 12081 16405 12115 16439
rect 13737 16405 13771 16439
rect 15485 16405 15519 16439
rect 1961 16201 1995 16235
rect 2513 16201 2547 16235
rect 2881 16201 2915 16235
rect 4077 16201 4111 16235
rect 4353 16201 4387 16235
rect 4905 16201 4939 16235
rect 5641 16201 5675 16235
rect 6377 16201 6411 16235
rect 7849 16201 7883 16235
rect 8217 16201 8251 16235
rect 9873 16201 9907 16235
rect 10425 16201 10459 16235
rect 11529 16201 11563 16235
rect 12817 16201 12851 16235
rect 8668 16133 8702 16167
rect 11253 16133 11287 16167
rect 15669 16133 15703 16167
rect 1685 16065 1719 16099
rect 1777 16065 1811 16099
rect 2421 16065 2455 16099
rect 2697 16065 2731 16099
rect 3065 16065 3099 16099
rect 3341 16065 3375 16099
rect 3433 16065 3467 16099
rect 3893 16065 3927 16099
rect 4261 16065 4295 16099
rect 4537 16065 4571 16099
rect 4629 16065 4663 16099
rect 5089 16065 5123 16099
rect 5181 16065 5215 16099
rect 5465 16065 5499 16099
rect 5733 16065 5767 16099
rect 7490 16065 7524 16099
rect 7757 16065 7791 16099
rect 8033 16065 8067 16099
rect 8401 16065 8435 16099
rect 11897 16065 11931 16099
rect 12541 16065 12575 16099
rect 13737 16065 13771 16099
rect 10241 15997 10275 16031
rect 10333 15997 10367 16031
rect 10977 15997 11011 16031
rect 11989 15997 12023 16031
rect 12081 15997 12115 16031
rect 13461 15997 13495 16031
rect 13829 15997 13863 16031
rect 14013 15997 14047 16031
rect 2237 15929 2271 15963
rect 3157 15929 3191 15963
rect 3709 15929 3743 15963
rect 4813 15929 4847 15963
rect 5917 15929 5951 15963
rect 11069 15929 11103 15963
rect 12357 15929 12391 15963
rect 1501 15861 1535 15895
rect 3617 15861 3651 15895
rect 5365 15861 5399 15895
rect 6101 15861 6135 15895
rect 9781 15861 9815 15895
rect 10793 15861 10827 15895
rect 1501 15657 1535 15691
rect 1777 15657 1811 15691
rect 2145 15657 2179 15691
rect 2421 15657 2455 15691
rect 2697 15657 2731 15691
rect 2973 15657 3007 15691
rect 3617 15657 3651 15691
rect 3893 15657 3927 15691
rect 6285 15657 6319 15691
rect 7205 15657 7239 15691
rect 9965 15657 9999 15691
rect 10977 15657 11011 15691
rect 3249 15589 3283 15623
rect 4077 15589 4111 15623
rect 12725 15589 12759 15623
rect 6653 15521 6687 15555
rect 8585 15521 8619 15555
rect 9413 15521 9447 15555
rect 10517 15521 10551 15555
rect 10701 15521 10735 15555
rect 11529 15521 11563 15555
rect 12541 15521 12575 15555
rect 13369 15521 13403 15555
rect 14105 15521 14139 15555
rect 1685 15453 1719 15487
rect 1961 15453 1995 15487
rect 2329 15453 2363 15487
rect 2605 15453 2639 15487
rect 2881 15453 2915 15487
rect 3157 15453 3191 15487
rect 3433 15453 3467 15487
rect 4169 15453 4203 15487
rect 4905 15453 4939 15487
rect 6837 15453 6871 15487
rect 7297 15453 7331 15487
rect 7573 15453 7607 15487
rect 9137 15453 9171 15487
rect 12265 15453 12299 15487
rect 14381 15453 14415 15487
rect 15025 15453 15059 15487
rect 5172 15385 5206 15419
rect 8217 15385 8251 15419
rect 8401 15385 8435 15419
rect 9597 15385 9631 15419
rect 13737 15385 13771 15419
rect 15669 15385 15703 15419
rect 4813 15317 4847 15351
rect 6745 15317 6779 15351
rect 8953 15317 8987 15351
rect 9505 15317 9539 15351
rect 10057 15317 10091 15351
rect 10425 15317 10459 15351
rect 11345 15317 11379 15351
rect 11437 15317 11471 15351
rect 11897 15317 11931 15351
rect 12357 15317 12391 15351
rect 13093 15317 13127 15351
rect 13185 15317 13219 15351
rect 13645 15317 13679 15351
rect 5457 15113 5491 15147
rect 5825 15113 5859 15147
rect 5917 15113 5951 15147
rect 6377 15113 6411 15147
rect 7205 15113 7239 15147
rect 8493 15113 8527 15147
rect 9505 15113 9539 15147
rect 11345 15113 11379 15147
rect 12265 15113 12299 15147
rect 12357 15113 12391 15147
rect 13001 15113 13035 15147
rect 15577 15113 15611 15147
rect 7573 15045 7607 15079
rect 8309 15045 8343 15079
rect 10232 15045 10266 15079
rect 14013 15045 14047 15079
rect 2706 14977 2740 15011
rect 2973 14977 3007 15011
rect 3065 14977 3099 15011
rect 3332 14977 3366 15011
rect 4905 14977 4939 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 8677 14977 8711 15011
rect 9137 14977 9171 15011
rect 9597 14977 9631 15011
rect 11713 14977 11747 15011
rect 12909 14977 12943 15011
rect 13369 14977 13403 15011
rect 14197 14977 14231 15011
rect 15117 14977 15151 15011
rect 4997 14909 5031 14943
rect 5089 14909 5123 14943
rect 6101 14909 6135 14943
rect 7021 14909 7055 14943
rect 7665 14909 7699 14943
rect 7849 14909 7883 14943
rect 8861 14909 8895 14943
rect 9045 14909 9079 14943
rect 9965 14909 9999 14943
rect 12449 14909 12483 14943
rect 13461 14909 13495 14943
rect 13645 14909 13679 14943
rect 14473 14909 14507 14943
rect 1501 14841 1535 14875
rect 11529 14841 11563 14875
rect 1593 14773 1627 14807
rect 4445 14773 4479 14807
rect 4537 14773 4571 14807
rect 8217 14773 8251 14807
rect 9781 14773 9815 14807
rect 11897 14773 11931 14807
rect 12725 14773 12759 14807
rect 13921 14773 13955 14807
rect 15393 14773 15427 14807
rect 1501 14569 1535 14603
rect 7757 14569 7791 14603
rect 9229 14569 9263 14603
rect 12633 14569 12667 14603
rect 2881 14501 2915 14535
rect 12357 14501 12391 14535
rect 15577 14501 15611 14535
rect 2145 14433 2179 14467
rect 3433 14433 3467 14467
rect 3985 14433 4019 14467
rect 5917 14433 5951 14467
rect 8401 14433 8435 14467
rect 9781 14433 9815 14467
rect 10333 14433 10367 14467
rect 13093 14433 13127 14467
rect 1685 14365 1719 14399
rect 1961 14365 1995 14399
rect 4445 14365 4479 14399
rect 6193 14365 6227 14399
rect 8125 14365 8159 14399
rect 9689 14365 9723 14399
rect 10517 14365 10551 14399
rect 10977 14365 11011 14399
rect 11244 14365 11278 14399
rect 12449 14365 12483 14399
rect 13369 14365 13403 14399
rect 14105 14365 14139 14399
rect 2421 14297 2455 14331
rect 3341 14297 3375 14331
rect 4712 14297 4746 14331
rect 6460 14297 6494 14331
rect 8217 14297 8251 14331
rect 8953 14297 8987 14331
rect 9597 14297 9631 14331
rect 12725 14297 12759 14331
rect 12909 14297 12943 14331
rect 14350 14297 14384 14331
rect 1777 14229 1811 14263
rect 2329 14229 2363 14263
rect 2789 14229 2823 14263
rect 3249 14229 3283 14263
rect 3893 14229 3927 14263
rect 4169 14229 4203 14263
rect 5825 14229 5859 14263
rect 7573 14229 7607 14263
rect 8677 14229 8711 14263
rect 10425 14229 10459 14263
rect 10885 14229 10919 14263
rect 15485 14229 15519 14263
rect 1777 14025 1811 14059
rect 2513 14025 2547 14059
rect 2973 14025 3007 14059
rect 3801 14025 3835 14059
rect 4169 14025 4203 14059
rect 4997 14025 5031 14059
rect 5365 14025 5399 14059
rect 5733 14025 5767 14059
rect 6193 14025 6227 14059
rect 6745 14025 6779 14059
rect 7389 14025 7423 14059
rect 11345 14025 11379 14059
rect 11989 14025 12023 14059
rect 12357 14025 12391 14059
rect 12817 14025 12851 14059
rect 2421 13957 2455 13991
rect 3341 13957 3375 13991
rect 4905 13957 4939 13991
rect 6837 13957 6871 13991
rect 7297 13957 7331 13991
rect 11529 13957 11563 13991
rect 1685 13889 1719 13923
rect 1961 13889 1995 13923
rect 3433 13889 3467 13923
rect 5825 13889 5859 13923
rect 7757 13889 7791 13923
rect 8024 13889 8058 13923
rect 9229 13889 9263 13923
rect 9485 13889 9519 13923
rect 10701 13889 10735 13923
rect 12449 13889 12483 13923
rect 13185 13889 13219 13923
rect 13277 13889 13311 13923
rect 13645 13889 13679 13923
rect 2329 13821 2363 13855
rect 3525 13821 3559 13855
rect 4261 13821 4295 13855
rect 4445 13821 4479 13855
rect 4813 13821 4847 13855
rect 5549 13821 5583 13855
rect 7021 13821 7055 13855
rect 11897 13821 11931 13855
rect 12541 13821 12575 13855
rect 13369 13821 13403 13855
rect 13921 13821 13955 13855
rect 15485 13821 15519 13855
rect 15669 13821 15703 13855
rect 1501 13753 1535 13787
rect 2881 13753 2915 13787
rect 7573 13753 7607 13787
rect 9137 13753 9171 13787
rect 10609 13753 10643 13787
rect 6377 13685 6411 13719
rect 2697 13481 2731 13515
rect 5181 13481 5215 13515
rect 5733 13481 5767 13515
rect 7389 13481 7423 13515
rect 8953 13481 8987 13515
rect 9597 13481 9631 13515
rect 11897 13481 11931 13515
rect 14105 13481 14139 13515
rect 3801 13413 3835 13447
rect 4261 13413 4295 13447
rect 9505 13413 9539 13447
rect 12265 13413 12299 13447
rect 3341 13345 3375 13379
rect 4629 13345 4663 13379
rect 4721 13345 4755 13379
rect 8769 13345 8803 13379
rect 10149 13345 10183 13379
rect 14657 13345 14691 13379
rect 15577 13345 15611 13379
rect 1685 13277 1719 13311
rect 2605 13277 2639 13311
rect 3065 13277 3099 13311
rect 3525 13277 3559 13311
rect 3985 13277 4019 13311
rect 8513 13277 8547 13311
rect 9321 13277 9355 13311
rect 13645 13277 13679 13311
rect 15393 13277 15427 13311
rect 1777 13209 1811 13243
rect 4813 13209 4847 13243
rect 7021 13209 7055 13243
rect 10057 13209 10091 13243
rect 10425 13209 10459 13243
rect 13378 13209 13412 13243
rect 15301 13209 15335 13243
rect 1501 13141 1535 13175
rect 1961 13141 1995 13175
rect 3157 13141 3191 13175
rect 4169 13141 4203 13175
rect 7205 13141 7239 13175
rect 9965 13141 9999 13175
rect 13737 13141 13771 13175
rect 14473 13141 14507 13175
rect 14565 13141 14599 13175
rect 14933 13141 14967 13175
rect 3249 12937 3283 12971
rect 4721 12937 4755 12971
rect 4997 12937 5031 12971
rect 5365 12937 5399 12971
rect 5825 12937 5859 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 7665 12937 7699 12971
rect 9781 12937 9815 12971
rect 10333 12937 10367 12971
rect 10977 12937 11011 12971
rect 11161 12937 11195 12971
rect 11529 12937 11563 12971
rect 14473 12937 14507 12971
rect 15025 12937 15059 12971
rect 3586 12869 3620 12903
rect 5273 12869 5307 12903
rect 5733 12869 5767 12903
rect 7757 12869 7791 12903
rect 8861 12869 8895 12903
rect 13001 12869 13035 12903
rect 1869 12801 1903 12835
rect 2136 12801 2170 12835
rect 3341 12801 3375 12835
rect 8125 12801 8159 12835
rect 9137 12801 9171 12835
rect 10425 12801 10459 12835
rect 11897 12801 11931 12835
rect 12357 12801 12391 12835
rect 13921 12801 13955 12835
rect 14565 12801 14599 12835
rect 15669 12801 15703 12835
rect 6009 12733 6043 12767
rect 6837 12733 6871 12767
rect 6929 12733 6963 12767
rect 7849 12733 7883 12767
rect 10609 12733 10643 12767
rect 11345 12733 11379 12767
rect 11989 12733 12023 12767
rect 12173 12733 12207 12767
rect 12817 12733 12851 12767
rect 13277 12733 13311 12767
rect 14289 12733 14323 12767
rect 8769 12665 8803 12699
rect 14933 12665 14967 12699
rect 1593 12597 1627 12631
rect 1777 12597 1811 12631
rect 7297 12597 7331 12631
rect 9965 12597 9999 12631
rect 2145 12393 2179 12427
rect 3157 12393 3191 12427
rect 3801 12393 3835 12427
rect 8677 12393 8711 12427
rect 10701 12393 10735 12427
rect 10977 12393 11011 12427
rect 12633 12393 12667 12427
rect 15669 12393 15703 12427
rect 2973 12325 3007 12359
rect 4813 12325 4847 12359
rect 10333 12325 10367 12359
rect 10885 12325 10919 12359
rect 4353 12257 4387 12291
rect 5273 12257 5307 12291
rect 5457 12257 5491 12291
rect 13185 12257 13219 12291
rect 14197 12257 14231 12291
rect 15117 12257 15151 12291
rect 1501 12189 1535 12223
rect 2513 12189 2547 12223
rect 2789 12189 2823 12223
rect 5641 12189 5675 12223
rect 5825 12189 5859 12223
rect 7297 12189 7331 12223
rect 8953 12189 8987 12223
rect 11161 12189 11195 12223
rect 13001 12189 13035 12223
rect 14473 12189 14507 12223
rect 15301 12189 15335 12223
rect 3341 12121 3375 12155
rect 3617 12121 3651 12155
rect 4169 12121 4203 12155
rect 6092 12121 6126 12155
rect 7542 12121 7576 12155
rect 9220 12121 9254 12155
rect 11428 12121 11462 12155
rect 13737 12121 13771 12155
rect 2329 12053 2363 12087
rect 2605 12053 2639 12087
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 5181 12053 5215 12087
rect 7205 12053 7239 12087
rect 12541 12053 12575 12087
rect 13093 12053 13127 12087
rect 13645 12053 13679 12087
rect 14381 12053 14415 12087
rect 14841 12053 14875 12087
rect 15209 12053 15243 12087
rect 3801 11849 3835 11883
rect 4353 11849 4387 11883
rect 4721 11849 4755 11883
rect 5181 11849 5215 11883
rect 6009 11849 6043 11883
rect 6929 11849 6963 11883
rect 7297 11849 7331 11883
rect 7757 11849 7791 11883
rect 9321 11849 9355 11883
rect 9873 11849 9907 11883
rect 10333 11849 10367 11883
rect 11529 11849 11563 11883
rect 12909 11849 12943 11883
rect 13553 11849 13587 11883
rect 14013 11849 14047 11883
rect 14197 11849 14231 11883
rect 14749 11849 14783 11883
rect 15025 11849 15059 11883
rect 6837 11781 6871 11815
rect 13461 11781 13495 11815
rect 14381 11781 14415 11815
rect 15393 11781 15427 11815
rect 2533 11713 2567 11747
rect 2789 11713 2823 11747
rect 3249 11713 3283 11747
rect 4261 11713 4295 11747
rect 5089 11713 5123 11747
rect 5825 11713 5859 11747
rect 7665 11713 7699 11747
rect 8125 11713 8159 11747
rect 8677 11713 8711 11747
rect 10241 11713 10275 11747
rect 11897 11713 11931 11747
rect 11989 11713 12023 11747
rect 13829 11713 13863 11747
rect 14841 11713 14875 11747
rect 15117 11713 15151 11747
rect 3341 11645 3375 11679
rect 3433 11645 3467 11679
rect 4445 11645 4479 11679
rect 5273 11645 5307 11679
rect 7021 11645 7055 11679
rect 7849 11645 7883 11679
rect 10517 11645 10551 11679
rect 12081 11645 12115 11679
rect 14473 11645 14507 11679
rect 6469 11577 6503 11611
rect 13001 11577 13035 11611
rect 1409 11509 1443 11543
rect 2881 11509 2915 11543
rect 3893 11509 3927 11543
rect 5549 11509 5583 11543
rect 9505 11509 9539 11543
rect 12449 11509 12483 11543
rect 12725 11509 12759 11543
rect 13277 11509 13311 11543
rect 2697 11305 2731 11339
rect 3617 11305 3651 11339
rect 3801 11305 3835 11339
rect 5273 11305 5307 11339
rect 6469 11305 6503 11339
rect 10149 11305 10183 11339
rect 13645 11305 13679 11339
rect 15209 11305 15243 11339
rect 15531 11305 15565 11339
rect 8953 11237 8987 11271
rect 13921 11237 13955 11271
rect 2053 11169 2087 11203
rect 2237 11169 2271 11203
rect 2973 11169 3007 11203
rect 3157 11169 3191 11203
rect 5825 11169 5859 11203
rect 7205 11169 7239 11203
rect 7389 11169 7423 11203
rect 8401 11169 8435 11203
rect 8585 11169 8619 11203
rect 9505 11169 9539 11203
rect 10793 11169 10827 11203
rect 13461 11169 13495 11203
rect 14197 11169 14231 11203
rect 15301 11169 15335 11203
rect 1685 11101 1719 11135
rect 2329 11101 2363 11135
rect 5181 11101 5215 11135
rect 9321 11101 9355 11135
rect 10517 11101 10551 11135
rect 10609 11101 10643 11135
rect 11621 11101 11655 11135
rect 11713 11101 11747 11135
rect 14381 11101 14415 11135
rect 15602 11101 15636 11135
rect 4914 11033 4948 11067
rect 5641 11033 5675 11067
rect 6101 11033 6135 11067
rect 7113 11033 7147 11067
rect 8309 11033 8343 11067
rect 9781 11033 9815 11067
rect 10977 11033 11011 11067
rect 11958 11033 11992 11067
rect 14473 11033 14507 11067
rect 15025 11033 15059 11067
rect 1501 10965 1535 10999
rect 3249 10965 3283 10999
rect 5733 10965 5767 10999
rect 6745 10965 6779 10999
rect 7941 10965 7975 10999
rect 9413 10965 9447 10999
rect 13093 10965 13127 10999
rect 13185 10965 13219 10999
rect 14841 10965 14875 10999
rect 1501 10761 1535 10795
rect 3065 10761 3099 10795
rect 7757 10761 7791 10795
rect 11713 10761 11747 10795
rect 4353 10693 4387 10727
rect 9689 10693 9723 10727
rect 1685 10625 1719 10659
rect 5558 10625 5592 10659
rect 5825 10625 5859 10659
rect 6377 10625 6411 10659
rect 6644 10625 6678 10659
rect 11078 10625 11112 10659
rect 11345 10625 11379 10659
rect 12837 10625 12871 10659
rect 13093 10625 13127 10659
rect 13185 10625 13219 10659
rect 13452 10625 13486 10659
rect 15025 10625 15059 10659
rect 6101 10557 6135 10591
rect 15117 10557 15151 10591
rect 15209 10557 15243 10591
rect 4445 10489 4479 10523
rect 8401 10489 8435 10523
rect 14657 10489 14691 10523
rect 15485 10489 15519 10523
rect 5917 10421 5951 10455
rect 9965 10421 9999 10455
rect 14565 10421 14599 10455
rect 3249 10217 3283 10251
rect 3617 10217 3651 10251
rect 5641 10217 5675 10251
rect 7297 10217 7331 10251
rect 9505 10217 9539 10251
rect 11713 10217 11747 10251
rect 7389 10149 7423 10183
rect 2697 10081 2731 10115
rect 4445 10081 4479 10115
rect 8769 10081 8803 10115
rect 10149 10081 10183 10115
rect 12817 10081 12851 10115
rect 13645 10081 13679 10115
rect 14565 10081 14599 10115
rect 14657 10081 14691 10115
rect 15117 10081 15151 10115
rect 1685 10013 1719 10047
rect 1961 10013 1995 10047
rect 2421 10013 2455 10047
rect 2881 10013 2915 10047
rect 4169 10013 4203 10047
rect 4997 10013 5031 10047
rect 7113 10013 7147 10047
rect 8513 10013 8547 10047
rect 9873 10013 9907 10047
rect 12633 10013 12667 10047
rect 14473 10013 14507 10047
rect 15393 10013 15427 10047
rect 2789 9945 2823 9979
rect 4261 9945 4295 9979
rect 6868 9945 6902 9979
rect 10425 9945 10459 9979
rect 12725 9945 12759 9979
rect 1501 9877 1535 9911
rect 1777 9877 1811 9911
rect 2053 9877 2087 9911
rect 3341 9877 3375 9911
rect 3801 9877 3835 9911
rect 4629 9877 4663 9911
rect 4905 9877 4939 9911
rect 5733 9877 5767 9911
rect 9965 9877 9999 9911
rect 12265 9877 12299 9911
rect 13093 9877 13127 9911
rect 13461 9877 13495 9911
rect 13553 9877 13587 9911
rect 14105 9877 14139 9911
rect 15577 9877 15611 9911
rect 4353 9673 4387 9707
rect 9873 9673 9907 9707
rect 10241 9673 10275 9707
rect 10333 9673 10367 9707
rect 11529 9673 11563 9707
rect 12817 9673 12851 9707
rect 13185 9673 13219 9707
rect 2789 9605 2823 9639
rect 5917 9605 5951 9639
rect 6745 9605 6779 9639
rect 8401 9605 8435 9639
rect 8953 9605 8987 9639
rect 9781 9605 9815 9639
rect 10793 9605 10827 9639
rect 11989 9605 12023 9639
rect 12725 9605 12759 9639
rect 1685 9537 1719 9571
rect 1961 9537 1995 9571
rect 2237 9537 2271 9571
rect 3157 9537 3191 9571
rect 4261 9537 4295 9571
rect 5181 9537 5215 9571
rect 5273 9537 5307 9571
rect 6101 9537 6135 9571
rect 7573 9537 7607 9571
rect 8493 9537 8527 9571
rect 10701 9537 10735 9571
rect 11897 9537 11931 9571
rect 13553 9537 13587 9571
rect 14381 9537 14415 9571
rect 3065 9469 3099 9503
rect 4445 9469 4479 9503
rect 5365 9469 5399 9503
rect 5641 9469 5675 9503
rect 6561 9469 6595 9503
rect 6653 9469 6687 9503
rect 7665 9469 7699 9503
rect 7849 9469 7883 9503
rect 8677 9469 8711 9503
rect 9597 9469 9631 9503
rect 10885 9469 10919 9503
rect 12081 9469 12115 9503
rect 12909 9469 12943 9503
rect 13645 9469 13679 9503
rect 13829 9469 13863 9503
rect 14473 9469 14507 9503
rect 14565 9469 14599 9503
rect 3893 9401 3927 9435
rect 7113 9401 7147 9435
rect 8033 9401 8067 9435
rect 9229 9401 9263 9435
rect 12357 9401 12391 9435
rect 15025 9401 15059 9435
rect 1501 9333 1535 9367
rect 1777 9333 1811 9367
rect 2053 9333 2087 9367
rect 2421 9333 2455 9367
rect 2605 9333 2639 9367
rect 3801 9333 3835 9367
rect 4813 9333 4847 9367
rect 7205 9333 7239 9367
rect 9045 9333 9079 9367
rect 11253 9333 11287 9367
rect 14013 9333 14047 9367
rect 14933 9333 14967 9367
rect 15301 9333 15335 9367
rect 3801 9129 3835 9163
rect 3985 9129 4019 9163
rect 4169 9129 4203 9163
rect 8953 9129 8987 9163
rect 3617 9061 3651 9095
rect 4629 8993 4663 9027
rect 4721 8993 4755 9027
rect 6469 8993 6503 9027
rect 8217 8993 8251 9027
rect 9505 8993 9539 9027
rect 12357 8993 12391 9027
rect 14565 8993 14599 9027
rect 1685 8925 1719 8959
rect 1777 8925 1811 8959
rect 2237 8925 2271 8959
rect 4997 8925 5031 8959
rect 7941 8925 7975 8959
rect 10149 8925 10183 8959
rect 10885 8925 10919 8959
rect 12541 8925 12575 8959
rect 14105 8925 14139 8959
rect 14841 8925 14875 8959
rect 15485 8925 15519 8959
rect 2504 8857 2538 8891
rect 5242 8857 5276 8891
rect 6714 8857 6748 8891
rect 10793 8857 10827 8891
rect 11130 8857 11164 8891
rect 12808 8857 12842 8891
rect 15301 8857 15335 8891
rect 1501 8789 1535 8823
rect 1961 8789 1995 8823
rect 2145 8789 2179 8823
rect 4537 8789 4571 8823
rect 6377 8789 6411 8823
rect 7849 8789 7883 8823
rect 9321 8789 9355 8823
rect 9413 8789 9447 8823
rect 9781 8789 9815 8823
rect 12265 8789 12299 8823
rect 13921 8789 13955 8823
rect 14381 8789 14415 8823
rect 14657 8789 14691 8823
rect 15025 8789 15059 8823
rect 15669 8789 15703 8823
rect 1777 8585 1811 8619
rect 3249 8585 3283 8619
rect 4721 8585 4755 8619
rect 5733 8585 5767 8619
rect 5825 8585 5859 8619
rect 8125 8585 8159 8619
rect 8953 8585 8987 8619
rect 9321 8585 9355 8619
rect 9873 8585 9907 8619
rect 9965 8585 9999 8619
rect 12173 8585 12207 8619
rect 12541 8585 12575 8619
rect 12909 8585 12943 8619
rect 13369 8585 13403 8619
rect 7113 8517 7147 8551
rect 1685 8449 1719 8483
rect 1961 8449 1995 8483
rect 2237 8449 2271 8483
rect 2513 8449 2547 8483
rect 2789 8449 2823 8483
rect 3065 8449 3099 8483
rect 4362 8449 4396 8483
rect 4629 8449 4663 8483
rect 5365 8449 5399 8483
rect 6377 8449 6411 8483
rect 8493 8449 8527 8483
rect 11089 8449 11123 8483
rect 11345 8449 11379 8483
rect 12081 8449 12115 8483
rect 13001 8449 13035 8483
rect 13461 8449 13495 8483
rect 13921 8449 13955 8483
rect 5641 8381 5675 8415
rect 7205 8381 7239 8415
rect 7297 8381 7331 8415
rect 7573 8381 7607 8415
rect 8585 8381 8619 8415
rect 8677 8381 8711 8415
rect 9413 8381 9447 8415
rect 9505 8381 9539 8415
rect 11713 8381 11747 8415
rect 11989 8381 12023 8415
rect 12817 8381 12851 8415
rect 1501 8313 1535 8347
rect 2053 8313 2087 8347
rect 2605 8313 2639 8347
rect 2881 8313 2915 8347
rect 6193 8313 6227 8347
rect 6745 8313 6779 8347
rect 7757 8313 7791 8347
rect 13829 8313 13863 8347
rect 2329 8245 2363 8279
rect 6561 8245 6595 8279
rect 7941 8245 7975 8279
rect 15393 8245 15427 8279
rect 2513 8041 2547 8075
rect 5273 8041 5307 8075
rect 6101 8041 6135 8075
rect 8309 8041 8343 8075
rect 8953 8041 8987 8075
rect 9781 8041 9815 8075
rect 11253 8041 11287 8075
rect 14105 8041 14139 8075
rect 15117 8041 15151 8075
rect 1501 7973 1535 8007
rect 3801 7973 3835 8007
rect 9965 7973 9999 8007
rect 13829 7973 13863 8007
rect 5181 7905 5215 7939
rect 5825 7905 5859 7939
rect 6561 7905 6595 7939
rect 6745 7905 6779 7939
rect 6929 7905 6963 7939
rect 8493 7905 8527 7939
rect 9413 7905 9447 7939
rect 9505 7905 9539 7939
rect 10885 7905 10919 7939
rect 11989 7905 12023 7939
rect 14657 7905 14691 7939
rect 1685 7837 1719 7871
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 2329 7837 2363 7871
rect 3433 7837 3467 7871
rect 5641 7837 5675 7871
rect 5733 7837 5767 7871
rect 7185 7837 7219 7871
rect 10241 7837 10275 7871
rect 12265 7837 12299 7871
rect 13001 7837 13035 7871
rect 14473 7837 14507 7871
rect 2697 7769 2731 7803
rect 4936 7769 4970 7803
rect 6469 7769 6503 7803
rect 9321 7769 9355 7803
rect 10701 7769 10735 7803
rect 11805 7769 11839 7803
rect 13553 7769 13587 7803
rect 14565 7769 14599 7803
rect 15393 7769 15427 7803
rect 1777 7701 1811 7735
rect 2053 7701 2087 7735
rect 2789 7701 2823 7735
rect 3525 7701 3559 7735
rect 8769 7701 8803 7735
rect 10333 7701 10367 7735
rect 10793 7701 10827 7735
rect 11437 7701 11471 7735
rect 11897 7701 11931 7735
rect 12909 7701 12943 7735
rect 13369 7701 13403 7735
rect 13645 7701 13679 7735
rect 14933 7701 14967 7735
rect 15577 7701 15611 7735
rect 3065 7497 3099 7531
rect 4997 7497 5031 7531
rect 6377 7497 6411 7531
rect 7665 7497 7699 7531
rect 7849 7497 7883 7531
rect 10425 7497 10459 7531
rect 13461 7497 13495 7531
rect 15025 7497 15059 7531
rect 15669 7497 15703 7531
rect 4353 7429 4387 7463
rect 4537 7429 4571 7463
rect 6837 7429 6871 7463
rect 8962 7429 8996 7463
rect 12642 7429 12676 7463
rect 14841 7429 14875 7463
rect 1685 7361 1719 7395
rect 2053 7361 2087 7395
rect 2513 7361 2547 7395
rect 5825 7361 5859 7395
rect 5917 7361 5951 7395
rect 6745 7361 6779 7395
rect 7389 7361 7423 7395
rect 7573 7361 7607 7395
rect 9229 7361 9263 7395
rect 10057 7361 10091 7395
rect 12909 7361 12943 7395
rect 14749 7361 14783 7395
rect 5089 7293 5123 7327
rect 5273 7293 5307 7327
rect 6101 7293 6135 7327
rect 6929 7293 6963 7327
rect 9781 7293 9815 7327
rect 9965 7293 9999 7327
rect 10517 7293 10551 7327
rect 15393 7293 15427 7327
rect 9505 7225 9539 7259
rect 11529 7225 11563 7259
rect 1501 7157 1535 7191
rect 1869 7157 1903 7191
rect 2329 7157 2363 7191
rect 4629 7157 4663 7191
rect 5457 7157 5491 7191
rect 7205 7157 7239 7191
rect 9413 7157 9447 7191
rect 10747 7157 10781 7191
rect 15301 7157 15335 7191
rect 3617 6953 3651 6987
rect 6009 6953 6043 6987
rect 11253 6953 11287 6987
rect 12909 6953 12943 6987
rect 14933 6953 14967 6987
rect 4077 6885 4111 6919
rect 11161 6885 11195 6919
rect 14565 6885 14599 6919
rect 15393 6885 15427 6919
rect 1593 6817 1627 6851
rect 4537 6817 4571 6851
rect 4721 6817 4755 6851
rect 5365 6817 5399 6851
rect 5549 6817 5583 6851
rect 6653 6817 6687 6851
rect 7481 6817 7515 6851
rect 7665 6817 7699 6851
rect 9045 6817 9079 6851
rect 11805 6817 11839 6851
rect 12541 6817 12575 6851
rect 12633 6817 12667 6851
rect 13461 6817 13495 6851
rect 2237 6749 2271 6783
rect 3893 6749 3927 6783
rect 4353 6749 4387 6783
rect 6469 6749 6503 6783
rect 6561 6749 6595 6783
rect 8125 6749 8159 6783
rect 9321 6749 9355 6783
rect 9781 6749 9815 6783
rect 13277 6749 13311 6783
rect 14197 6749 14231 6783
rect 14749 6749 14783 6783
rect 1685 6681 1719 6715
rect 2504 6681 2538 6715
rect 4813 6681 4847 6715
rect 7389 6681 7423 6715
rect 8769 6681 8803 6715
rect 10026 6681 10060 6715
rect 15025 6681 15059 6715
rect 15209 6681 15243 6715
rect 15577 6681 15611 6715
rect 1777 6613 1811 6647
rect 2145 6613 2179 6647
rect 4169 6613 4203 6647
rect 5181 6613 5215 6647
rect 5641 6613 5675 6647
rect 6101 6613 6135 6647
rect 7021 6613 7055 6647
rect 7941 6613 7975 6647
rect 9229 6613 9263 6647
rect 9689 6613 9723 6647
rect 11621 6613 11655 6647
rect 11713 6613 11747 6647
rect 12081 6613 12115 6647
rect 12449 6613 12483 6647
rect 13369 6613 13403 6647
rect 13737 6613 13771 6647
rect 14381 6613 14415 6647
rect 2053 6409 2087 6443
rect 4261 6409 4295 6443
rect 4629 6409 4663 6443
rect 4997 6409 5031 6443
rect 8585 6409 8619 6443
rect 11161 6409 11195 6443
rect 11713 6409 11747 6443
rect 11897 6409 11931 6443
rect 12265 6409 12299 6443
rect 14289 6409 14323 6443
rect 14473 6409 14507 6443
rect 8156 6341 8190 6375
rect 9720 6341 9754 6375
rect 13093 6341 13127 6375
rect 13921 6341 13955 6375
rect 1685 6273 1719 6307
rect 1777 6273 1811 6307
rect 3166 6273 3200 6307
rect 3709 6273 3743 6307
rect 4169 6273 4203 6307
rect 5825 6273 5859 6307
rect 6377 6273 6411 6307
rect 9965 6273 9999 6307
rect 11529 6273 11563 6307
rect 12357 6273 12391 6307
rect 14841 6273 14875 6307
rect 15393 6273 15427 6307
rect 3433 6205 3467 6239
rect 4353 6205 4387 6239
rect 5089 6205 5123 6239
rect 5181 6205 5215 6239
rect 5917 6205 5951 6239
rect 6101 6205 6135 6239
rect 6929 6205 6963 6239
rect 8401 6205 8435 6239
rect 10241 6205 10275 6239
rect 10517 6205 10551 6239
rect 12541 6205 12575 6239
rect 12909 6205 12943 6239
rect 13001 6205 13035 6239
rect 13737 6205 13771 6239
rect 13829 6205 13863 6239
rect 14933 6205 14967 6239
rect 15025 6205 15059 6239
rect 1501 6137 1535 6171
rect 5457 6137 5491 6171
rect 13461 6137 13495 6171
rect 1961 6069 1995 6103
rect 3525 6069 3559 6103
rect 3801 6069 3835 6103
rect 7021 6069 7055 6103
rect 10057 6069 10091 6103
rect 15577 6069 15611 6103
rect 3893 5865 3927 5899
rect 8953 5865 8987 5899
rect 9229 5865 9263 5899
rect 11713 5865 11747 5899
rect 14841 5865 14875 5899
rect 2789 5797 2823 5831
rect 2881 5797 2915 5831
rect 6929 5797 6963 5831
rect 13829 5797 13863 5831
rect 3525 5729 3559 5763
rect 6285 5729 6319 5763
rect 7665 5729 7699 5763
rect 8401 5729 8435 5763
rect 8677 5729 8711 5763
rect 10149 5729 10183 5763
rect 12817 5729 12851 5763
rect 13277 5729 13311 5763
rect 14289 5729 14323 5763
rect 15485 5729 15519 5763
rect 1409 5661 1443 5695
rect 3249 5661 3283 5695
rect 5365 5661 5399 5695
rect 6101 5661 6135 5695
rect 6469 5661 6503 5695
rect 7389 5661 7423 5695
rect 7481 5661 7515 5695
rect 9137 5637 9171 5671
rect 9413 5661 9447 5695
rect 12633 5661 12667 5695
rect 14473 5661 14507 5695
rect 15393 5661 15427 5695
rect 1676 5593 1710 5627
rect 3341 5593 3375 5627
rect 5098 5593 5132 5627
rect 6561 5593 6595 5627
rect 8309 5593 8343 5627
rect 10425 5593 10459 5627
rect 13461 5593 13495 5627
rect 3985 5525 4019 5559
rect 5457 5525 5491 5559
rect 7021 5525 7055 5559
rect 7849 5525 7883 5559
rect 8217 5525 8251 5559
rect 9597 5525 9631 5559
rect 9965 5525 9999 5559
rect 10057 5525 10091 5559
rect 12265 5525 12299 5559
rect 12725 5525 12759 5559
rect 13369 5525 13403 5559
rect 14381 5525 14415 5559
rect 14933 5525 14967 5559
rect 15301 5525 15335 5559
rect 1501 5321 1535 5355
rect 1777 5321 1811 5355
rect 3065 5321 3099 5355
rect 6469 5321 6503 5355
rect 7113 5321 7147 5355
rect 7941 5321 7975 5355
rect 8401 5321 8435 5355
rect 9965 5321 9999 5355
rect 11529 5321 11563 5355
rect 13001 5321 13035 5355
rect 13461 5321 13495 5355
rect 14381 5321 14415 5355
rect 11100 5253 11134 5287
rect 15669 5253 15703 5287
rect 1685 5185 1719 5219
rect 2145 5185 2179 5219
rect 4353 5185 4387 5219
rect 4445 5185 4479 5219
rect 4813 5185 4847 5219
rect 5080 5185 5114 5219
rect 6653 5185 6687 5219
rect 9514 5185 9548 5219
rect 9781 5185 9815 5219
rect 11345 5185 11379 5219
rect 12653 5185 12687 5219
rect 13369 5185 13403 5219
rect 2237 5117 2271 5151
rect 2421 5117 2455 5151
rect 7205 5117 7239 5151
rect 7297 5117 7331 5151
rect 7665 5117 7699 5151
rect 7849 5117 7883 5151
rect 12909 5117 12943 5151
rect 13553 5117 13587 5151
rect 6745 5049 6779 5083
rect 4629 4981 4663 5015
rect 6193 4981 6227 5015
rect 8309 4981 8343 5015
rect 2881 4777 2915 4811
rect 7941 4777 7975 4811
rect 12449 4777 12483 4811
rect 13921 4777 13955 4811
rect 14749 4777 14783 4811
rect 5181 4709 5215 4743
rect 7757 4709 7791 4743
rect 11345 4709 11379 4743
rect 2513 4641 2547 4675
rect 2697 4641 2731 4675
rect 3525 4641 3559 4675
rect 3801 4641 3835 4675
rect 5917 4641 5951 4675
rect 8401 4641 8435 4675
rect 8493 4641 8527 4675
rect 9137 4641 9171 4675
rect 9781 4641 9815 4675
rect 10701 4641 10735 4675
rect 11897 4641 11931 4675
rect 11989 4641 12023 4675
rect 15669 4641 15703 4675
rect 1685 4573 1719 4607
rect 2421 4573 2455 4607
rect 3341 4573 3375 4607
rect 5273 4573 5307 4607
rect 5825 4573 5859 4607
rect 6173 4573 6207 4607
rect 7665 4573 7699 4607
rect 9413 4573 9447 4607
rect 9873 4573 9907 4607
rect 10425 4573 10459 4607
rect 11529 4573 11563 4607
rect 12541 4573 12575 4607
rect 14105 4573 14139 4607
rect 15393 4573 15427 4607
rect 1961 4505 1995 4539
rect 4068 4505 4102 4539
rect 12081 4505 12115 4539
rect 12808 4505 12842 4539
rect 1501 4437 1535 4471
rect 2053 4437 2087 4471
rect 3249 4437 3283 4471
rect 5457 4437 5491 4471
rect 5641 4437 5675 4471
rect 7297 4437 7331 4471
rect 7481 4437 7515 4471
rect 8309 4437 8343 4471
rect 9229 4437 9263 4471
rect 9965 4437 9999 4471
rect 10333 4437 10367 4471
rect 1777 4233 1811 4267
rect 4445 4233 4479 4267
rect 6837 4233 6871 4267
rect 10057 4233 10091 4267
rect 12081 4233 12115 4267
rect 12449 4233 12483 4267
rect 14933 4233 14967 4267
rect 15301 4233 15335 4267
rect 6745 4165 6779 4199
rect 2504 4097 2538 4131
rect 3709 4097 3743 4131
rect 4353 4097 4387 4131
rect 5558 4097 5592 4131
rect 5825 4097 5859 4131
rect 6193 4097 6227 4131
rect 7297 4097 7331 4131
rect 8217 4097 8251 4131
rect 8953 4097 8987 4131
rect 9413 4097 9447 4131
rect 9873 4097 9907 4131
rect 10517 4097 10551 4131
rect 10609 4097 10643 4131
rect 11069 4097 11103 4131
rect 11989 4097 12023 4131
rect 12808 4097 12842 4131
rect 14841 4097 14875 4131
rect 15393 4097 15427 4131
rect 1593 4029 1627 4063
rect 1685 4029 1719 4063
rect 2237 4029 2271 4063
rect 6929 4029 6963 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 10701 4029 10735 4063
rect 11253 4029 11287 4063
rect 11897 4029 11931 4063
rect 12541 4029 12575 4063
rect 14565 4029 14599 4063
rect 15577 4029 15611 4063
rect 8033 3961 8067 3995
rect 10149 3961 10183 3995
rect 11529 3961 11563 3995
rect 13921 3961 13955 3995
rect 2145 3893 2179 3927
rect 3617 3893 3651 3927
rect 6009 3893 6043 3927
rect 6377 3893 6411 3927
rect 7941 3893 7975 3927
rect 8309 3893 8343 3927
rect 9781 3893 9815 3927
rect 1961 3689 1995 3723
rect 7389 3689 7423 3723
rect 9137 3689 9171 3723
rect 9597 3689 9631 3723
rect 1685 3621 1719 3655
rect 2881 3621 2915 3655
rect 2421 3553 2455 3587
rect 2513 3553 2547 3587
rect 3525 3553 3559 3587
rect 4537 3553 4571 3587
rect 5089 3553 5123 3587
rect 6377 3553 6411 3587
rect 7021 3553 7055 3587
rect 7205 3553 7239 3587
rect 8769 3553 8803 3587
rect 10149 3553 10183 3587
rect 12817 3553 12851 3587
rect 13921 3553 13955 3587
rect 14565 3553 14599 3587
rect 14841 3553 14875 3587
rect 15485 3553 15519 3587
rect 1869 3485 1903 3519
rect 2329 3485 2363 3519
rect 3341 3485 3375 3519
rect 5181 3485 5215 3519
rect 6101 3485 6135 3519
rect 8502 3485 8536 3519
rect 8953 3485 8987 3519
rect 9505 3485 9539 3519
rect 10057 3485 10091 3519
rect 10425 3485 10459 3519
rect 12725 3485 12759 3519
rect 13645 3485 13679 3519
rect 14105 3485 14139 3519
rect 14289 3485 14323 3519
rect 3249 3417 3283 3451
rect 1501 3349 1535 3383
rect 3893 3349 3927 3383
rect 3985 3349 4019 3383
rect 4353 3349 4387 3383
rect 4445 3349 4479 3383
rect 5273 3349 5307 3383
rect 5641 3349 5675 3383
rect 5733 3349 5767 3383
rect 6193 3349 6227 3383
rect 6561 3349 6595 3383
rect 6929 3349 6963 3383
rect 9321 3349 9355 3383
rect 9965 3349 9999 3383
rect 11713 3349 11747 3383
rect 12265 3349 12299 3383
rect 12633 3349 12667 3383
rect 3893 3145 3927 3179
rect 4353 3145 4387 3179
rect 4721 3145 4755 3179
rect 5181 3145 5215 3179
rect 5549 3145 5583 3179
rect 5641 3145 5675 3179
rect 11897 3145 11931 3179
rect 11989 3145 12023 3179
rect 14473 3145 14507 3179
rect 2320 3077 2354 3111
rect 6377 3077 6411 3111
rect 7674 3077 7708 3111
rect 12725 3077 12759 3111
rect 13338 3077 13372 3111
rect 1409 3009 1443 3043
rect 1961 3009 1995 3043
rect 2053 3009 2087 3043
rect 3709 3009 3743 3043
rect 4261 3009 4295 3043
rect 6193 3009 6227 3043
rect 7941 3009 7975 3043
rect 8033 3009 8067 3043
rect 8217 3009 8251 3043
rect 9525 3009 9559 3043
rect 9781 3009 9815 3043
rect 10986 3009 11020 3043
rect 11253 3009 11287 3043
rect 12541 3009 12575 3043
rect 12909 3009 12943 3043
rect 13093 3009 13127 3043
rect 14841 3009 14875 3043
rect 15485 3009 15519 3043
rect 4813 2941 4847 2975
rect 4905 2941 4939 2975
rect 5733 2941 5767 2975
rect 12081 2941 12115 2975
rect 12357 2941 12391 2975
rect 14565 2941 14599 2975
rect 1593 2873 1627 2907
rect 3525 2873 3559 2907
rect 4077 2873 4111 2907
rect 6561 2873 6595 2907
rect 9873 2873 9907 2907
rect 1777 2805 1811 2839
rect 3433 2805 3467 2839
rect 6009 2805 6043 2839
rect 8401 2805 8435 2839
rect 11529 2805 11563 2839
rect 15669 2805 15703 2839
rect 1593 2601 1627 2635
rect 4537 2601 4571 2635
rect 5641 2601 5675 2635
rect 8125 2601 8159 2635
rect 9045 2601 9079 2635
rect 10425 2601 10459 2635
rect 15485 2601 15519 2635
rect 2053 2533 2087 2567
rect 2697 2533 2731 2567
rect 4261 2533 4295 2567
rect 8217 2533 8251 2567
rect 8493 2533 8527 2567
rect 10517 2533 10551 2567
rect 5181 2465 5215 2499
rect 9597 2465 9631 2499
rect 11069 2465 11103 2499
rect 11529 2465 11563 2499
rect 11805 2465 11839 2499
rect 13277 2465 13311 2499
rect 13737 2465 13771 2499
rect 1777 2397 1811 2431
rect 1869 2397 1903 2431
rect 2513 2397 2547 2431
rect 2881 2397 2915 2431
rect 3249 2397 3283 2431
rect 3617 2397 3651 2431
rect 4077 2397 4111 2431
rect 4445 2397 4479 2431
rect 5825 2397 5859 2431
rect 6193 2397 6227 2431
rect 6965 2397 6999 2431
rect 7492 2397 7526 2431
rect 8401 2397 8435 2431
rect 9413 2397 9447 2431
rect 9505 2397 9539 2431
rect 10057 2397 10091 2431
rect 10241 2397 10275 2431
rect 10885 2397 10919 2431
rect 13001 2397 13035 2431
rect 13921 2397 13955 2431
rect 14565 2397 14599 2431
rect 14841 2397 14875 2431
rect 4997 2329 5031 2363
rect 6561 2329 6595 2363
rect 7205 2329 7239 2363
rect 8677 2329 8711 2363
rect 10977 2329 11011 2363
rect 14289 2329 14323 2363
rect 2329 2261 2363 2295
rect 3065 2261 3099 2295
rect 3433 2261 3467 2295
rect 3893 2261 3927 2295
rect 4905 2261 4939 2295
rect 5457 2261 5491 2295
rect 6009 2261 6043 2295
rect 6469 2261 6503 2295
rect 6837 2261 6871 2295
rect 7297 2261 7331 2295
rect 9965 2261 9999 2295
rect 14197 2261 14231 2295
<< metal1 >>
rect 6454 17620 6460 17672
rect 6512 17660 6518 17672
rect 8386 17660 8392 17672
rect 6512 17632 8392 17660
rect 6512 17620 6518 17632
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 5534 17552 5540 17604
rect 5592 17592 5598 17604
rect 6730 17592 6736 17604
rect 5592 17564 6736 17592
rect 5592 17552 5598 17564
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 7282 17552 7288 17604
rect 7340 17592 7346 17604
rect 12526 17592 12532 17604
rect 7340 17564 12532 17592
rect 7340 17552 7346 17564
rect 12526 17552 12532 17564
rect 12584 17552 12590 17604
rect 198 17484 204 17536
rect 256 17524 262 17536
rect 3786 17524 3792 17536
rect 256 17496 3792 17524
rect 256 17484 262 17496
rect 3786 17484 3792 17496
rect 3844 17484 3850 17536
rect 9030 17484 9036 17536
rect 9088 17524 9094 17536
rect 11422 17524 11428 17536
rect 9088 17496 11428 17524
rect 9088 17484 9094 17496
rect 11422 17484 11428 17496
rect 11480 17484 11486 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 1581 17323 1639 17329
rect 1581 17289 1593 17323
rect 1627 17320 1639 17323
rect 1762 17320 1768 17332
rect 1627 17292 1768 17320
rect 1627 17289 1639 17292
rect 1581 17283 1639 17289
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 1949 17323 2007 17329
rect 1949 17289 1961 17323
rect 1995 17320 2007 17323
rect 2222 17320 2228 17332
rect 1995 17292 2228 17320
rect 1995 17289 2007 17292
rect 1949 17283 2007 17289
rect 2222 17280 2228 17292
rect 2280 17280 2286 17332
rect 2317 17323 2375 17329
rect 2317 17289 2329 17323
rect 2363 17320 2375 17323
rect 2590 17320 2596 17332
rect 2363 17292 2596 17320
rect 2363 17289 2375 17292
rect 2317 17283 2375 17289
rect 2590 17280 2596 17292
rect 2648 17280 2654 17332
rect 2685 17323 2743 17329
rect 2685 17289 2697 17323
rect 2731 17320 2743 17323
rect 3050 17320 3056 17332
rect 2731 17292 3056 17320
rect 2731 17289 2743 17292
rect 2685 17283 2743 17289
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3145 17323 3203 17329
rect 3145 17289 3157 17323
rect 3191 17320 3203 17323
rect 3418 17320 3424 17332
rect 3191 17292 3424 17320
rect 3191 17289 3203 17292
rect 3145 17283 3203 17289
rect 3418 17280 3424 17292
rect 3476 17280 3482 17332
rect 4157 17323 4215 17329
rect 4157 17289 4169 17323
rect 4203 17320 4215 17323
rect 4614 17320 4620 17332
rect 4203 17292 4620 17320
rect 4203 17289 4215 17292
rect 4157 17283 4215 17289
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 4985 17323 5043 17329
rect 4985 17289 4997 17323
rect 5031 17320 5043 17323
rect 5902 17320 5908 17332
rect 5031 17292 5908 17320
rect 5031 17289 5043 17292
rect 4985 17283 5043 17289
rect 5902 17280 5908 17292
rect 5960 17280 5966 17332
rect 6089 17323 6147 17329
rect 6089 17289 6101 17323
rect 6135 17320 6147 17323
rect 7469 17323 7527 17329
rect 6135 17292 7236 17320
rect 6135 17289 6147 17292
rect 6089 17283 6147 17289
rect 3694 17252 3700 17264
rect 2884 17224 3700 17252
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 1765 17147 1823 17153
rect 1780 17048 1808 17147
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2884 17193 2912 17224
rect 3694 17212 3700 17224
rect 3752 17212 3758 17264
rect 5626 17212 5632 17264
rect 5684 17212 5690 17264
rect 7098 17252 7104 17264
rect 5736 17224 7104 17252
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2869 17187 2927 17193
rect 2869 17153 2881 17187
rect 2915 17153 2927 17187
rect 2869 17147 2927 17153
rect 2961 17187 3019 17193
rect 2961 17153 2973 17187
rect 3007 17184 3019 17187
rect 3142 17184 3148 17196
rect 3007 17156 3148 17184
rect 3007 17153 3019 17156
rect 2961 17147 3019 17153
rect 2516 17116 2544 17147
rect 3142 17144 3148 17156
rect 3200 17144 3206 17196
rect 3602 17184 3608 17196
rect 3563 17156 3608 17184
rect 3602 17144 3608 17156
rect 3660 17144 3666 17196
rect 3786 17193 3792 17196
rect 3781 17184 3792 17193
rect 3747 17156 3792 17184
rect 3781 17147 3792 17156
rect 3844 17184 3850 17196
rect 4338 17184 4344 17196
rect 3844 17156 4200 17184
rect 4299 17156 4344 17184
rect 3786 17144 3792 17147
rect 3844 17144 3850 17156
rect 3234 17116 3240 17128
rect 2516 17088 3240 17116
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 4172 17116 4200 17156
rect 4338 17144 4344 17156
rect 4396 17144 4402 17196
rect 4430 17144 4436 17196
rect 4488 17184 4494 17196
rect 4488 17156 4533 17184
rect 4488 17144 4494 17156
rect 4614 17144 4620 17196
rect 4672 17184 4678 17196
rect 4801 17187 4859 17193
rect 4801 17184 4813 17187
rect 4672 17156 4813 17184
rect 4672 17144 4678 17156
rect 4801 17153 4813 17156
rect 4847 17153 4859 17187
rect 5166 17184 5172 17196
rect 5127 17156 5172 17184
rect 4801 17147 4859 17153
rect 5166 17144 5172 17156
rect 5224 17144 5230 17196
rect 5537 17187 5595 17193
rect 5537 17153 5549 17187
rect 5583 17184 5595 17187
rect 5644 17184 5672 17212
rect 5583 17156 5672 17184
rect 5583 17153 5595 17156
rect 5537 17147 5595 17153
rect 5626 17116 5632 17128
rect 4172 17088 5632 17116
rect 5626 17076 5632 17088
rect 5684 17076 5690 17128
rect 3326 17048 3332 17060
rect 1780 17020 3332 17048
rect 3326 17008 3332 17020
rect 3384 17008 3390 17060
rect 3421 17051 3479 17057
rect 3421 17017 3433 17051
rect 3467 17048 3479 17051
rect 4246 17048 4252 17060
rect 3467 17020 4252 17048
rect 3467 17017 3479 17020
rect 3421 17011 3479 17017
rect 4246 17008 4252 17020
rect 4304 17008 4310 17060
rect 4617 17051 4675 17057
rect 4617 17017 4629 17051
rect 4663 17048 4675 17051
rect 5442 17048 5448 17060
rect 4663 17020 5448 17048
rect 4663 17017 4675 17020
rect 4617 17011 4675 17017
rect 5442 17008 5448 17020
rect 5500 17008 5506 17060
rect 3970 16980 3976 16992
rect 3931 16952 3976 16980
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 5353 16983 5411 16989
rect 5353 16949 5365 16983
rect 5399 16980 5411 16983
rect 5534 16980 5540 16992
rect 5399 16952 5540 16980
rect 5399 16949 5411 16952
rect 5353 16943 5411 16949
rect 5534 16940 5540 16952
rect 5592 16940 5598 16992
rect 5736 16989 5764 17224
rect 7098 17212 7104 17224
rect 7156 17212 7162 17264
rect 7208 17252 7236 17292
rect 7469 17289 7481 17323
rect 7515 17320 7527 17323
rect 7837 17323 7895 17329
rect 7837 17320 7849 17323
rect 7515 17292 7849 17320
rect 7515 17289 7527 17292
rect 7469 17283 7527 17289
rect 7837 17289 7849 17292
rect 7883 17289 7895 17323
rect 7837 17283 7895 17289
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 8904 17292 11744 17320
rect 8904 17280 8910 17292
rect 11716 17264 11744 17292
rect 7558 17252 7564 17264
rect 7208 17224 7564 17252
rect 7558 17212 7564 17224
rect 7616 17212 7622 17264
rect 9953 17255 10011 17261
rect 9953 17221 9965 17255
rect 9999 17252 10011 17255
rect 11514 17252 11520 17264
rect 9999 17224 11520 17252
rect 9999 17221 10011 17224
rect 9953 17215 10011 17221
rect 11514 17212 11520 17224
rect 11572 17212 11578 17264
rect 11698 17252 11704 17264
rect 11659 17224 11704 17252
rect 11698 17212 11704 17224
rect 11756 17212 11762 17264
rect 15746 17252 15752 17264
rect 13188 17224 15752 17252
rect 5902 17184 5908 17196
rect 5863 17156 5908 17184
rect 5902 17144 5908 17156
rect 5960 17144 5966 17196
rect 5994 17144 6000 17196
rect 6052 17184 6058 17196
rect 6389 17187 6447 17193
rect 6389 17184 6401 17187
rect 6052 17156 6401 17184
rect 6052 17144 6058 17156
rect 6389 17153 6401 17156
rect 6435 17184 6447 17187
rect 6917 17187 6975 17193
rect 6435 17156 6868 17184
rect 6435 17153 6447 17156
rect 6389 17147 6447 17153
rect 6840 17116 6868 17156
rect 6917 17153 6929 17187
rect 6963 17184 6975 17187
rect 7190 17184 7196 17196
rect 6963 17156 7196 17184
rect 6963 17153 6975 17156
rect 6917 17147 6975 17153
rect 7190 17144 7196 17156
rect 7248 17144 7254 17196
rect 7374 17184 7380 17196
rect 7335 17156 7380 17184
rect 7374 17144 7380 17156
rect 7432 17144 7438 17196
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 7668 17156 8217 17184
rect 6840 17088 6960 17116
rect 6549 17051 6607 17057
rect 6549 17017 6561 17051
rect 6595 17048 6607 17051
rect 6822 17048 6828 17060
rect 6595 17020 6828 17048
rect 6595 17017 6607 17020
rect 6549 17011 6607 17017
rect 6822 17008 6828 17020
rect 6880 17008 6886 17060
rect 6932 17048 6960 17088
rect 7466 17076 7472 17128
rect 7524 17116 7530 17128
rect 7561 17119 7619 17125
rect 7561 17116 7573 17119
rect 7524 17088 7573 17116
rect 7524 17076 7530 17088
rect 7561 17085 7573 17088
rect 7607 17085 7619 17119
rect 7561 17079 7619 17085
rect 7668 17048 7696 17156
rect 8205 17153 8217 17156
rect 8251 17184 8263 17187
rect 9306 17184 9312 17196
rect 8251 17156 9312 17184
rect 8251 17153 8263 17156
rect 8205 17147 8263 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 9582 17184 9588 17196
rect 9543 17156 9588 17184
rect 9582 17144 9588 17156
rect 9640 17144 9646 17196
rect 10042 17184 10048 17196
rect 10003 17156 10048 17184
rect 10042 17144 10048 17156
rect 10100 17144 10106 17196
rect 11882 17184 11888 17196
rect 11843 17156 11888 17184
rect 11882 17144 11888 17156
rect 11940 17144 11946 17196
rect 12618 17144 12624 17196
rect 12676 17184 12682 17196
rect 13081 17187 13139 17193
rect 13081 17184 13093 17187
rect 12676 17156 13093 17184
rect 12676 17144 12682 17156
rect 13081 17153 13093 17156
rect 13127 17153 13139 17187
rect 13081 17147 13139 17153
rect 8110 17076 8116 17128
rect 8168 17116 8174 17128
rect 8297 17119 8355 17125
rect 8297 17116 8309 17119
rect 8168 17088 8309 17116
rect 8168 17076 8174 17088
rect 8297 17085 8309 17088
rect 8343 17085 8355 17119
rect 8297 17079 8355 17085
rect 8389 17119 8447 17125
rect 8389 17085 8401 17119
rect 8435 17085 8447 17119
rect 9769 17119 9827 17125
rect 8389 17079 8447 17085
rect 8496 17088 9674 17116
rect 6932 17020 7696 17048
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 8404 17048 8432 17079
rect 8260 17020 8432 17048
rect 8260 17008 8266 17020
rect 5721 16983 5779 16989
rect 5721 16949 5733 16983
rect 5767 16949 5779 16983
rect 5721 16943 5779 16949
rect 6454 16940 6460 16992
rect 6512 16980 6518 16992
rect 6733 16983 6791 16989
rect 6733 16980 6745 16983
rect 6512 16952 6745 16980
rect 6512 16940 6518 16952
rect 6733 16949 6745 16952
rect 6779 16949 6791 16983
rect 6733 16943 6791 16949
rect 7009 16983 7067 16989
rect 7009 16949 7021 16983
rect 7055 16980 7067 16983
rect 7098 16980 7104 16992
rect 7055 16952 7104 16980
rect 7055 16949 7067 16952
rect 7009 16943 7067 16949
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 8018 16940 8024 16992
rect 8076 16980 8082 16992
rect 8496 16980 8524 17088
rect 8757 17051 8815 17057
rect 8757 17017 8769 17051
rect 8803 17048 8815 17051
rect 9214 17048 9220 17060
rect 8803 17020 9220 17048
rect 8803 17017 8815 17020
rect 8757 17011 8815 17017
rect 9214 17008 9220 17020
rect 9272 17008 9278 17060
rect 8938 16980 8944 16992
rect 8076 16952 8524 16980
rect 8899 16952 8944 16980
rect 8076 16940 8082 16952
rect 8938 16940 8944 16952
rect 8996 16940 9002 16992
rect 9646 16980 9674 17088
rect 9769 17085 9781 17119
rect 9815 17085 9827 17119
rect 11054 17116 11060 17128
rect 11015 17088 11060 17116
rect 9769 17079 9827 17085
rect 9784 17048 9812 17079
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17085 11391 17119
rect 11333 17079 11391 17085
rect 10686 17048 10692 17060
rect 9784 17020 10692 17048
rect 10686 17008 10692 17020
rect 10744 17008 10750 17060
rect 11146 17008 11152 17060
rect 11204 17048 11210 17060
rect 11348 17048 11376 17079
rect 11422 17076 11428 17128
rect 11480 17116 11486 17128
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 11480 17088 11529 17116
rect 11480 17076 11486 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 11698 17076 11704 17128
rect 11756 17116 11762 17128
rect 12066 17116 12072 17128
rect 11756 17088 12072 17116
rect 11756 17076 11762 17088
rect 12066 17076 12072 17088
rect 12124 17116 12130 17128
rect 12161 17119 12219 17125
rect 12161 17116 12173 17119
rect 12124 17088 12173 17116
rect 12124 17076 12130 17088
rect 12161 17085 12173 17088
rect 12207 17085 12219 17119
rect 12161 17079 12219 17085
rect 12434 17076 12440 17128
rect 12492 17116 12498 17128
rect 12492 17088 12537 17116
rect 12492 17076 12498 17088
rect 13188 17048 13216 17224
rect 15746 17212 15752 17224
rect 15804 17212 15810 17264
rect 14360 17187 14418 17193
rect 14360 17153 14372 17187
rect 14406 17184 14418 17187
rect 14826 17184 14832 17196
rect 14406 17156 14832 17184
rect 14406 17153 14418 17156
rect 14360 17147 14418 17153
rect 14826 17144 14832 17156
rect 14884 17144 14890 17196
rect 13357 17119 13415 17125
rect 13357 17085 13369 17119
rect 13403 17116 13415 17119
rect 13446 17116 13452 17128
rect 13403 17088 13452 17116
rect 13403 17085 13415 17088
rect 13357 17079 13415 17085
rect 13446 17076 13452 17088
rect 13504 17076 13510 17128
rect 13814 17076 13820 17128
rect 13872 17116 13878 17128
rect 14093 17119 14151 17125
rect 14093 17116 14105 17119
rect 13872 17088 14105 17116
rect 13872 17076 13878 17088
rect 14093 17085 14105 17088
rect 14139 17085 14151 17119
rect 14093 17079 14151 17085
rect 11204 17020 13216 17048
rect 15473 17051 15531 17057
rect 11204 17008 11210 17020
rect 15473 17017 15485 17051
rect 15519 17048 15531 17051
rect 15838 17048 15844 17060
rect 15519 17020 15844 17048
rect 15519 17017 15531 17020
rect 15473 17011 15531 17017
rect 15838 17008 15844 17020
rect 15896 17008 15902 17060
rect 10134 16980 10140 16992
rect 9646 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10413 16983 10471 16989
rect 10413 16980 10425 16983
rect 10284 16952 10425 16980
rect 10284 16940 10290 16952
rect 10413 16949 10425 16952
rect 10459 16949 10471 16983
rect 10413 16943 10471 16949
rect 10778 16940 10784 16992
rect 10836 16980 10842 16992
rect 11882 16980 11888 16992
rect 10836 16952 11888 16980
rect 10836 16940 10842 16952
rect 11882 16940 11888 16952
rect 11940 16940 11946 16992
rect 12069 16983 12127 16989
rect 12069 16949 12081 16983
rect 12115 16980 12127 16983
rect 12526 16980 12532 16992
rect 12115 16952 12532 16980
rect 12115 16949 12127 16952
rect 12069 16943 12127 16949
rect 12526 16940 12532 16952
rect 12584 16980 12590 16992
rect 13078 16980 13084 16992
rect 12584 16952 13084 16980
rect 12584 16940 12590 16952
rect 13078 16940 13084 16952
rect 13136 16940 13142 16992
rect 15378 16940 15384 16992
rect 15436 16980 15442 16992
rect 15565 16983 15623 16989
rect 15565 16980 15577 16983
rect 15436 16952 15577 16980
rect 15436 16940 15442 16952
rect 15565 16949 15577 16952
rect 15611 16949 15623 16983
rect 15565 16943 15623 16949
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 1854 16776 1860 16788
rect 1815 16748 1860 16776
rect 1854 16736 1860 16748
rect 1912 16736 1918 16788
rect 2225 16779 2283 16785
rect 2225 16745 2237 16779
rect 2271 16776 2283 16779
rect 2682 16776 2688 16788
rect 2271 16748 2688 16776
rect 2271 16745 2283 16748
rect 2225 16739 2283 16745
rect 2682 16736 2688 16748
rect 2740 16736 2746 16788
rect 3786 16736 3792 16788
rect 3844 16776 3850 16788
rect 4157 16779 4215 16785
rect 4157 16776 4169 16779
rect 3844 16748 4169 16776
rect 3844 16736 3850 16748
rect 4157 16745 4169 16748
rect 4203 16745 4215 16779
rect 4430 16776 4436 16788
rect 4391 16748 4436 16776
rect 4157 16739 4215 16745
rect 4430 16736 4436 16748
rect 4488 16736 4494 16788
rect 4893 16779 4951 16785
rect 4893 16745 4905 16779
rect 4939 16776 4951 16779
rect 5166 16776 5172 16788
rect 4939 16748 5172 16776
rect 4939 16745 4951 16748
rect 4893 16739 4951 16745
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 5810 16736 5816 16788
rect 5868 16776 5874 16788
rect 7098 16776 7104 16788
rect 5868 16748 7104 16776
rect 5868 16736 5874 16748
rect 7098 16736 7104 16748
rect 7156 16736 7162 16788
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 8846 16776 8852 16788
rect 8343 16748 8852 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 8846 16736 8852 16748
rect 8904 16776 8910 16788
rect 9582 16776 9588 16788
rect 8904 16748 9588 16776
rect 8904 16736 8910 16748
rect 9582 16736 9588 16748
rect 9640 16736 9646 16788
rect 10686 16776 10692 16788
rect 10647 16748 10692 16776
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11054 16736 11060 16788
rect 11112 16776 11118 16788
rect 15565 16779 15623 16785
rect 15565 16776 15577 16779
rect 11112 16748 15577 16776
rect 11112 16736 11118 16748
rect 1486 16708 1492 16720
rect 1447 16680 1492 16708
rect 1486 16668 1492 16680
rect 1544 16668 1550 16720
rect 2869 16711 2927 16717
rect 2869 16677 2881 16711
rect 2915 16708 2927 16711
rect 3142 16708 3148 16720
rect 2915 16680 3148 16708
rect 2915 16677 2927 16680
rect 2869 16671 2927 16677
rect 3142 16668 3148 16680
rect 3200 16668 3206 16720
rect 3605 16711 3663 16717
rect 3605 16677 3617 16711
rect 3651 16677 3663 16711
rect 3605 16671 3663 16677
rect 3881 16711 3939 16717
rect 3881 16677 3893 16711
rect 3927 16708 3939 16711
rect 5994 16708 6000 16720
rect 3927 16680 6000 16708
rect 3927 16677 3939 16680
rect 3881 16671 3939 16677
rect 3620 16640 3648 16671
rect 5994 16668 6000 16680
rect 6052 16668 6058 16720
rect 6914 16708 6920 16720
rect 6564 16680 6920 16708
rect 3252 16612 3556 16640
rect 3620 16612 4108 16640
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 1946 16572 1952 16584
rect 1719 16544 1952 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2041 16575 2099 16581
rect 2041 16541 2053 16575
rect 2087 16541 2099 16575
rect 2406 16572 2412 16584
rect 2367 16544 2412 16572
rect 2041 16535 2099 16541
rect 2056 16504 2084 16535
rect 2406 16532 2412 16544
rect 2464 16532 2470 16584
rect 2498 16532 2504 16584
rect 2556 16572 2562 16584
rect 2556 16544 2601 16572
rect 2556 16532 2562 16544
rect 2958 16532 2964 16584
rect 3016 16572 3022 16584
rect 3053 16575 3111 16581
rect 3053 16572 3065 16575
rect 3016 16544 3065 16572
rect 3016 16532 3022 16544
rect 3053 16541 3065 16544
rect 3099 16541 3111 16575
rect 3053 16535 3111 16541
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3252 16572 3280 16612
rect 3528 16584 3556 16612
rect 3191 16544 3280 16572
rect 3421 16575 3479 16581
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 3421 16541 3433 16575
rect 3467 16541 3479 16575
rect 3421 16535 3479 16541
rect 2590 16504 2596 16516
rect 2056 16476 2596 16504
rect 2590 16464 2596 16476
rect 2648 16464 2654 16516
rect 3436 16504 3464 16535
rect 3510 16532 3516 16584
rect 3568 16532 3574 16584
rect 3973 16575 4031 16581
rect 3973 16572 3985 16575
rect 3896 16544 3985 16572
rect 3786 16504 3792 16516
rect 3436 16476 3792 16504
rect 3786 16464 3792 16476
rect 3844 16464 3850 16516
rect 934 16396 940 16448
rect 992 16436 998 16448
rect 2685 16439 2743 16445
rect 2685 16436 2697 16439
rect 992 16408 2697 16436
rect 992 16396 998 16408
rect 2685 16405 2697 16408
rect 2731 16405 2743 16439
rect 2685 16399 2743 16405
rect 3329 16439 3387 16445
rect 3329 16405 3341 16439
rect 3375 16436 3387 16439
rect 3896 16436 3924 16544
rect 3973 16541 3985 16544
rect 4019 16541 4031 16575
rect 3973 16535 4031 16541
rect 4080 16504 4108 16612
rect 4908 16612 5120 16640
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 4617 16575 4675 16581
rect 4617 16572 4629 16575
rect 4580 16544 4629 16572
rect 4580 16532 4586 16544
rect 4617 16541 4629 16544
rect 4663 16541 4675 16575
rect 4617 16535 4675 16541
rect 4709 16575 4767 16581
rect 4709 16541 4721 16575
rect 4755 16572 4767 16575
rect 4908 16572 4936 16612
rect 4755 16544 4936 16572
rect 4985 16575 5043 16581
rect 4755 16541 4767 16544
rect 4709 16535 4767 16541
rect 4985 16541 4997 16575
rect 5031 16541 5043 16575
rect 5092 16572 5120 16612
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 6564 16649 6592 16680
rect 6914 16668 6920 16680
rect 6972 16668 6978 16720
rect 11330 16668 11336 16720
rect 11388 16668 11394 16720
rect 6549 16643 6607 16649
rect 6236 16612 6500 16640
rect 6236 16600 6242 16612
rect 5166 16572 5172 16584
rect 5092 16544 5172 16572
rect 4985 16535 5043 16541
rect 5000 16504 5028 16535
rect 5166 16532 5172 16544
rect 5224 16532 5230 16584
rect 5353 16575 5411 16581
rect 5353 16541 5365 16575
rect 5399 16572 5411 16575
rect 6362 16572 6368 16584
rect 5399 16544 6368 16572
rect 5399 16541 5411 16544
rect 5353 16535 5411 16541
rect 6362 16532 6368 16544
rect 6420 16532 6426 16584
rect 6472 16572 6500 16612
rect 6549 16609 6561 16643
rect 6595 16609 6607 16643
rect 6549 16603 6607 16609
rect 6641 16643 6699 16649
rect 6641 16609 6653 16643
rect 6687 16609 6699 16643
rect 6641 16603 6699 16609
rect 6656 16572 6684 16603
rect 8110 16600 8116 16652
rect 8168 16640 8174 16652
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8168 16612 8953 16640
rect 8168 16600 8174 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 11348 16640 11376 16668
rect 11425 16643 11483 16649
rect 11425 16640 11437 16643
rect 8941 16603 8999 16609
rect 10888 16612 11437 16640
rect 6472 16544 6684 16572
rect 6917 16575 6975 16581
rect 6917 16541 6929 16575
rect 6963 16572 6975 16575
rect 7742 16572 7748 16584
rect 6963 16544 7748 16572
rect 6963 16541 6975 16544
rect 6917 16535 6975 16541
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8294 16532 8300 16584
rect 8352 16572 8358 16584
rect 9309 16575 9367 16581
rect 9309 16572 9321 16575
rect 8352 16544 9321 16572
rect 8352 16532 8358 16544
rect 9309 16541 9321 16544
rect 9355 16541 9367 16575
rect 10888 16572 10916 16612
rect 11425 16609 11437 16612
rect 11471 16609 11483 16643
rect 11425 16603 11483 16609
rect 11609 16643 11667 16649
rect 11609 16609 11621 16643
rect 11655 16640 11667 16643
rect 11790 16640 11796 16652
rect 11655 16612 11796 16640
rect 11655 16609 11667 16612
rect 11609 16603 11667 16609
rect 11790 16600 11796 16612
rect 11848 16600 11854 16652
rect 9309 16535 9367 16541
rect 9600 16544 10916 16572
rect 9600 16516 9628 16544
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 11149 16575 11207 16581
rect 11149 16572 11161 16575
rect 11112 16544 11161 16572
rect 11112 16532 11118 16544
rect 11149 16541 11161 16544
rect 11195 16541 11207 16575
rect 12084 16572 12112 16748
rect 15565 16745 15577 16748
rect 15611 16745 15623 16779
rect 15565 16739 15623 16745
rect 13449 16643 13507 16649
rect 13449 16609 13461 16643
rect 13495 16640 13507 16643
rect 13814 16640 13820 16652
rect 13495 16612 13820 16640
rect 13495 16609 13507 16612
rect 13449 16603 13507 16609
rect 13814 16600 13820 16612
rect 13872 16640 13878 16652
rect 14093 16643 14151 16649
rect 14093 16640 14105 16643
rect 13872 16612 14105 16640
rect 13872 16600 13878 16612
rect 14093 16609 14105 16612
rect 14139 16609 14151 16643
rect 14093 16603 14151 16609
rect 13633 16575 13691 16581
rect 13633 16572 13645 16575
rect 11149 16535 11207 16541
rect 11808 16544 12112 16572
rect 12820 16544 13645 16572
rect 4080 16476 5028 16504
rect 5997 16507 6055 16513
rect 5997 16473 6009 16507
rect 6043 16504 6055 16507
rect 7162 16507 7220 16513
rect 7162 16504 7174 16507
rect 6043 16476 7174 16504
rect 6043 16473 6055 16476
rect 5997 16467 6055 16473
rect 7162 16473 7174 16476
rect 7208 16473 7220 16507
rect 7162 16467 7220 16473
rect 7834 16464 7840 16516
rect 7892 16504 7898 16516
rect 8665 16507 8723 16513
rect 8665 16504 8677 16507
rect 7892 16476 8677 16504
rect 7892 16464 7898 16476
rect 8665 16473 8677 16476
rect 8711 16473 8723 16507
rect 8665 16467 8723 16473
rect 9125 16507 9183 16513
rect 9125 16473 9137 16507
rect 9171 16504 9183 16507
rect 9214 16504 9220 16516
rect 9171 16476 9220 16504
rect 9171 16473 9183 16476
rect 9125 16467 9183 16473
rect 3375 16408 3924 16436
rect 3375 16405 3387 16408
rect 3329 16399 3387 16405
rect 5074 16396 5080 16448
rect 5132 16436 5138 16448
rect 5169 16439 5227 16445
rect 5169 16436 5181 16439
rect 5132 16408 5181 16436
rect 5132 16396 5138 16408
rect 5169 16405 5181 16408
rect 5215 16405 5227 16439
rect 6086 16436 6092 16448
rect 6047 16408 6092 16436
rect 5169 16399 5227 16405
rect 6086 16396 6092 16408
rect 6144 16396 6150 16448
rect 6454 16436 6460 16448
rect 6415 16408 6460 16436
rect 6454 16396 6460 16408
rect 6512 16396 6518 16448
rect 8018 16396 8024 16448
rect 8076 16436 8082 16448
rect 8573 16439 8631 16445
rect 8573 16436 8585 16439
rect 8076 16408 8585 16436
rect 8076 16396 8082 16408
rect 8573 16405 8585 16408
rect 8619 16405 8631 16439
rect 8680 16436 8708 16467
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 9582 16513 9588 16516
rect 9576 16504 9588 16513
rect 9543 16476 9588 16504
rect 9576 16467 9588 16476
rect 9582 16464 9588 16467
rect 9640 16464 9646 16516
rect 10134 16464 10140 16516
rect 10192 16504 10198 16516
rect 11808 16513 11836 16544
rect 11793 16507 11851 16513
rect 10192 16476 11100 16504
rect 10192 16464 10198 16476
rect 11072 16448 11100 16476
rect 11793 16473 11805 16507
rect 11839 16473 11851 16507
rect 11793 16467 11851 16473
rect 11882 16464 11888 16516
rect 11940 16504 11946 16516
rect 12820 16504 12848 16544
rect 13633 16541 13645 16544
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 11940 16476 12848 16504
rect 11940 16464 11946 16476
rect 13170 16464 13176 16516
rect 13228 16513 13234 16516
rect 13228 16504 13240 16513
rect 13228 16476 13273 16504
rect 13228 16467 13240 16476
rect 13228 16464 13234 16467
rect 13538 16464 13544 16516
rect 13596 16504 13602 16516
rect 14360 16507 14418 16513
rect 14360 16504 14372 16507
rect 13596 16476 14372 16504
rect 13596 16464 13602 16476
rect 14360 16473 14372 16476
rect 14406 16504 14418 16507
rect 16022 16504 16028 16516
rect 14406 16476 16028 16504
rect 14406 16473 14418 16476
rect 14360 16467 14418 16473
rect 16022 16464 16028 16476
rect 16080 16464 16086 16516
rect 9950 16436 9956 16448
rect 8680 16408 9956 16436
rect 8573 16399 8631 16405
rect 9950 16396 9956 16408
rect 10008 16396 10014 16448
rect 10778 16396 10784 16448
rect 10836 16436 10842 16448
rect 10836 16408 10881 16436
rect 10836 16396 10842 16408
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11241 16439 11299 16445
rect 11241 16436 11253 16439
rect 11112 16408 11253 16436
rect 11112 16396 11118 16408
rect 11241 16405 11253 16408
rect 11287 16405 11299 16439
rect 11241 16399 11299 16405
rect 11422 16396 11428 16448
rect 11480 16436 11486 16448
rect 12069 16439 12127 16445
rect 12069 16436 12081 16439
rect 11480 16408 12081 16436
rect 11480 16396 11486 16408
rect 12069 16405 12081 16408
rect 12115 16436 12127 16439
rect 12526 16436 12532 16448
rect 12115 16408 12532 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 12526 16396 12532 16408
rect 12584 16396 12590 16448
rect 13354 16396 13360 16448
rect 13412 16436 13418 16448
rect 13725 16439 13783 16445
rect 13725 16436 13737 16439
rect 13412 16408 13737 16436
rect 13412 16396 13418 16408
rect 13725 16405 13737 16408
rect 13771 16405 13783 16439
rect 15470 16436 15476 16448
rect 15431 16408 15476 16436
rect 13725 16399 13783 16405
rect 15470 16396 15476 16408
rect 15528 16396 15534 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 566 16192 572 16244
rect 624 16232 630 16244
rect 1949 16235 2007 16241
rect 1949 16232 1961 16235
rect 624 16204 1961 16232
rect 624 16192 630 16204
rect 1949 16201 1961 16204
rect 1995 16201 2007 16235
rect 1949 16195 2007 16201
rect 2130 16192 2136 16244
rect 2188 16232 2194 16244
rect 2501 16235 2559 16241
rect 2501 16232 2513 16235
rect 2188 16204 2513 16232
rect 2188 16192 2194 16204
rect 2501 16201 2513 16204
rect 2547 16201 2559 16235
rect 2501 16195 2559 16201
rect 2869 16235 2927 16241
rect 2869 16201 2881 16235
rect 2915 16232 2927 16235
rect 3234 16232 3240 16244
rect 2915 16204 3240 16232
rect 2915 16201 2927 16204
rect 2869 16195 2927 16201
rect 3234 16192 3240 16204
rect 3292 16192 3298 16244
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 4065 16235 4123 16241
rect 4065 16232 4077 16235
rect 3660 16204 4077 16232
rect 3660 16192 3666 16204
rect 4065 16201 4077 16204
rect 4111 16201 4123 16235
rect 4338 16232 4344 16244
rect 4299 16204 4344 16232
rect 4065 16195 4123 16201
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 4614 16192 4620 16244
rect 4672 16232 4678 16244
rect 4893 16235 4951 16241
rect 4893 16232 4905 16235
rect 4672 16204 4905 16232
rect 4672 16192 4678 16204
rect 4893 16201 4905 16204
rect 4939 16201 4951 16235
rect 4893 16195 4951 16201
rect 5534 16192 5540 16244
rect 5592 16192 5598 16244
rect 5629 16235 5687 16241
rect 5629 16201 5641 16235
rect 5675 16232 5687 16235
rect 5902 16232 5908 16244
rect 5675 16204 5908 16232
rect 5675 16201 5687 16204
rect 5629 16195 5687 16201
rect 5902 16192 5908 16204
rect 5960 16192 5966 16244
rect 6362 16232 6368 16244
rect 6323 16204 6368 16232
rect 6362 16192 6368 16204
rect 6420 16192 6426 16244
rect 7006 16192 7012 16244
rect 7064 16232 7070 16244
rect 7834 16232 7840 16244
rect 7064 16204 7696 16232
rect 7795 16204 7840 16232
rect 7064 16192 7070 16204
rect 2222 16124 2228 16176
rect 2280 16164 2286 16176
rect 2280 16136 3372 16164
rect 2280 16124 2286 16136
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1636 16068 1685 16096
rect 1636 16056 1642 16068
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 2409 16099 2467 16105
rect 1820 16068 1865 16096
rect 1820 16056 1826 16068
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 2590 16096 2596 16108
rect 2455 16068 2596 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2590 16056 2596 16068
rect 2648 16056 2654 16108
rect 2685 16099 2743 16105
rect 2685 16065 2697 16099
rect 2731 16065 2743 16099
rect 2685 16059 2743 16065
rect 3053 16099 3111 16105
rect 3053 16065 3065 16099
rect 3099 16096 3111 16099
rect 3234 16096 3240 16108
rect 3099 16068 3240 16096
rect 3099 16065 3111 16068
rect 3053 16059 3111 16065
rect 2314 15988 2320 16040
rect 2372 16028 2378 16040
rect 2700 16028 2728 16059
rect 3234 16056 3240 16068
rect 3292 16056 3298 16108
rect 3344 16105 3372 16136
rect 4430 16124 4436 16176
rect 4488 16164 4494 16176
rect 4488 16136 5203 16164
rect 4488 16124 4494 16136
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16065 3387 16099
rect 3329 16059 3387 16065
rect 3418 16056 3424 16108
rect 3476 16096 3482 16108
rect 3786 16096 3792 16108
rect 3476 16068 3792 16096
rect 3476 16056 3482 16068
rect 3786 16056 3792 16068
rect 3844 16056 3850 16108
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16096 3939 16099
rect 3970 16096 3976 16108
rect 3927 16068 3976 16096
rect 3927 16065 3939 16068
rect 3881 16059 3939 16065
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4246 16096 4252 16108
rect 4207 16068 4252 16096
rect 4246 16056 4252 16068
rect 4304 16056 4310 16108
rect 4525 16099 4583 16105
rect 4525 16065 4537 16099
rect 4571 16065 4583 16099
rect 4525 16059 4583 16065
rect 4617 16099 4675 16105
rect 4617 16065 4629 16099
rect 4663 16096 4675 16099
rect 4982 16096 4988 16108
rect 4663 16068 4988 16096
rect 4663 16065 4675 16068
rect 4617 16059 4675 16065
rect 2372 16000 2728 16028
rect 2372 15988 2378 16000
rect 2958 15988 2964 16040
rect 3016 16028 3022 16040
rect 4540 16028 4568 16059
rect 4982 16056 4988 16068
rect 5040 16056 5046 16108
rect 5175 16105 5203 16136
rect 5077 16099 5135 16105
rect 5077 16065 5089 16099
rect 5123 16065 5135 16099
rect 5077 16059 5135 16065
rect 5169 16099 5227 16105
rect 5169 16065 5181 16099
rect 5215 16096 5227 16099
rect 5350 16096 5356 16108
rect 5215 16068 5356 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 4706 16028 4712 16040
rect 3016 16000 3924 16028
rect 4540 16000 4712 16028
rect 3016 15988 3022 16000
rect 3896 15972 3924 16000
rect 4706 15988 4712 16000
rect 4764 15988 4770 16040
rect 5092 16028 5120 16059
rect 5350 16056 5356 16068
rect 5408 16056 5414 16108
rect 5453 16099 5511 16105
rect 5453 16065 5465 16099
rect 5499 16096 5511 16099
rect 5552 16096 5580 16192
rect 7668 16164 7696 16204
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 7926 16192 7932 16244
rect 7984 16232 7990 16244
rect 8205 16235 8263 16241
rect 8205 16232 8217 16235
rect 7984 16204 8217 16232
rect 7984 16192 7990 16204
rect 8205 16201 8217 16204
rect 8251 16201 8263 16235
rect 8205 16195 8263 16201
rect 9122 16192 9128 16244
rect 9180 16232 9186 16244
rect 9861 16235 9919 16241
rect 9861 16232 9873 16235
rect 9180 16204 9873 16232
rect 9180 16192 9186 16204
rect 9861 16201 9873 16204
rect 9907 16201 9919 16235
rect 9861 16195 9919 16201
rect 10413 16235 10471 16241
rect 10413 16201 10425 16235
rect 10459 16232 10471 16235
rect 10778 16232 10784 16244
rect 10459 16204 10784 16232
rect 10459 16201 10471 16204
rect 10413 16195 10471 16201
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11514 16232 11520 16244
rect 11475 16204 11520 16232
rect 11514 16192 11520 16204
rect 11572 16192 11578 16244
rect 12526 16192 12532 16244
rect 12584 16232 12590 16244
rect 12805 16235 12863 16241
rect 12805 16232 12817 16235
rect 12584 16204 12817 16232
rect 12584 16192 12590 16204
rect 12805 16201 12817 16204
rect 12851 16232 12863 16235
rect 14550 16232 14556 16244
rect 12851 16204 14556 16232
rect 12851 16201 12863 16204
rect 12805 16195 12863 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 16574 16232 16580 16244
rect 14660 16204 16580 16232
rect 8656 16167 8714 16173
rect 7668 16136 8064 16164
rect 5499 16068 5580 16096
rect 5721 16100 5779 16105
rect 5721 16099 5856 16100
rect 5499 16065 5511 16068
rect 5453 16059 5511 16065
rect 5721 16065 5733 16099
rect 5767 16072 5856 16099
rect 5767 16065 5779 16072
rect 5721 16059 5779 16065
rect 5534 16028 5540 16040
rect 5092 16000 5540 16028
rect 5534 15988 5540 16000
rect 5592 15988 5598 16040
rect 1394 15920 1400 15972
rect 1452 15960 1458 15972
rect 2225 15963 2283 15969
rect 2225 15960 2237 15963
rect 1452 15932 2237 15960
rect 1452 15920 1458 15932
rect 2225 15929 2237 15932
rect 2271 15929 2283 15963
rect 2225 15923 2283 15929
rect 2406 15920 2412 15972
rect 2464 15960 2470 15972
rect 3145 15963 3203 15969
rect 3145 15960 3157 15963
rect 2464 15932 3157 15960
rect 2464 15920 2470 15932
rect 3145 15929 3157 15932
rect 3191 15929 3203 15963
rect 3694 15960 3700 15972
rect 3655 15932 3700 15960
rect 3145 15923 3203 15929
rect 3694 15920 3700 15932
rect 3752 15920 3758 15972
rect 3878 15920 3884 15972
rect 3936 15920 3942 15972
rect 4801 15963 4859 15969
rect 4801 15929 4813 15963
rect 4847 15960 4859 15963
rect 5828 15960 5856 16072
rect 6178 16056 6184 16108
rect 6236 16096 6242 16108
rect 7466 16096 7472 16108
rect 7524 16105 7530 16108
rect 6236 16068 7472 16096
rect 6236 16056 6242 16068
rect 7466 16056 7472 16068
rect 7524 16059 7536 16105
rect 7742 16096 7748 16108
rect 7703 16068 7748 16096
rect 7524 16056 7530 16059
rect 7742 16056 7748 16068
rect 7800 16056 7806 16108
rect 8036 16105 8064 16136
rect 8656 16133 8668 16167
rect 8702 16164 8714 16167
rect 8938 16164 8944 16176
rect 8702 16136 8944 16164
rect 8702 16133 8714 16136
rect 8656 16127 8714 16133
rect 8938 16124 8944 16136
rect 8996 16124 9002 16176
rect 9214 16124 9220 16176
rect 9272 16164 9278 16176
rect 11238 16164 11244 16176
rect 9272 16136 10824 16164
rect 11199 16136 11244 16164
rect 9272 16124 9278 16136
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16065 8079 16099
rect 8021 16059 8079 16065
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 8352 16068 8401 16096
rect 8352 16056 8358 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 10686 16096 10692 16108
rect 8389 16059 8447 16065
rect 10244 16068 10692 16096
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10244 16037 10272 16068
rect 10686 16056 10692 16068
rect 10744 16056 10750 16108
rect 10796 16096 10824 16136
rect 11238 16124 11244 16136
rect 11296 16124 11302 16176
rect 12894 16164 12900 16176
rect 11348 16136 12900 16164
rect 11348 16096 11376 16136
rect 12894 16124 12900 16136
rect 12952 16124 12958 16176
rect 14660 16164 14688 16204
rect 16574 16192 16580 16204
rect 16632 16192 16638 16244
rect 15654 16164 15660 16176
rect 13188 16136 14688 16164
rect 15615 16136 15660 16164
rect 13188 16108 13216 16136
rect 15654 16124 15660 16136
rect 15712 16124 15718 16176
rect 11882 16096 11888 16108
rect 10796 16068 11376 16096
rect 11843 16068 11888 16096
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 12529 16099 12587 16105
rect 11992 16068 12434 16096
rect 11992 16040 12020 16068
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 10192 16000 10241 16028
rect 10192 15988 10198 16000
rect 10229 15997 10241 16000
rect 10275 15997 10287 16031
rect 10229 15991 10287 15997
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 15997 10379 16031
rect 10321 15991 10379 15997
rect 10965 16031 11023 16037
rect 10965 15997 10977 16031
rect 11011 16028 11023 16031
rect 11514 16028 11520 16040
rect 11011 16000 11520 16028
rect 11011 15997 11023 16000
rect 10965 15991 11023 15997
rect 4847 15932 5856 15960
rect 5905 15963 5963 15969
rect 4847 15929 4859 15932
rect 4801 15923 4859 15929
rect 5905 15929 5917 15963
rect 5951 15960 5963 15963
rect 6270 15960 6276 15972
rect 5951 15932 6276 15960
rect 5951 15929 5963 15932
rect 5905 15923 5963 15929
rect 6270 15920 6276 15932
rect 6328 15920 6334 15972
rect 9950 15920 9956 15972
rect 10008 15960 10014 15972
rect 10336 15960 10364 15991
rect 11514 15988 11520 16000
rect 11572 15988 11578 16040
rect 11974 16028 11980 16040
rect 11935 16000 11980 16028
rect 11974 15988 11980 16000
rect 12032 15988 12038 16040
rect 12069 16031 12127 16037
rect 12069 15997 12081 16031
rect 12115 15997 12127 16031
rect 12406 16028 12434 16068
rect 12529 16065 12541 16099
rect 12575 16096 12587 16099
rect 13170 16096 13176 16108
rect 12575 16068 13176 16096
rect 12575 16065 12587 16068
rect 12529 16059 12587 16065
rect 13170 16056 13176 16068
rect 13228 16056 13234 16108
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13538 16096 13544 16108
rect 13320 16068 13544 16096
rect 13320 16056 13326 16068
rect 13538 16056 13544 16068
rect 13596 16096 13602 16108
rect 13725 16099 13783 16105
rect 13725 16096 13737 16099
rect 13596 16068 13737 16096
rect 13596 16056 13602 16068
rect 13725 16065 13737 16068
rect 13771 16065 13783 16099
rect 13725 16059 13783 16065
rect 13449 16031 13507 16037
rect 13449 16028 13461 16031
rect 12406 16000 13461 16028
rect 12069 15991 12127 15997
rect 13449 15997 13461 16000
rect 13495 15997 13507 16031
rect 13449 15991 13507 15997
rect 13817 16031 13875 16037
rect 13817 15997 13829 16031
rect 13863 15997 13875 16031
rect 13817 15991 13875 15997
rect 14001 16031 14059 16037
rect 14001 15997 14013 16031
rect 14047 16028 14059 16031
rect 15562 16028 15568 16040
rect 14047 16000 15568 16028
rect 14047 15997 14059 16000
rect 14001 15991 14059 15997
rect 11054 15960 11060 15972
rect 10008 15932 10364 15960
rect 11015 15932 11060 15960
rect 10008 15920 10014 15932
rect 11054 15920 11060 15932
rect 11112 15920 11118 15972
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 12084 15960 12112 15991
rect 11388 15932 12112 15960
rect 12345 15963 12403 15969
rect 11388 15920 11394 15932
rect 12345 15929 12357 15963
rect 12391 15929 12403 15963
rect 13832 15960 13860 15991
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 13906 15960 13912 15972
rect 13832 15932 13912 15960
rect 12345 15923 12403 15929
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 3602 15892 3608 15904
rect 3563 15864 3608 15892
rect 3602 15852 3608 15864
rect 3660 15852 3666 15904
rect 5353 15895 5411 15901
rect 5353 15861 5365 15895
rect 5399 15892 5411 15895
rect 5718 15892 5724 15904
rect 5399 15864 5724 15892
rect 5399 15861 5411 15864
rect 5353 15855 5411 15861
rect 5718 15852 5724 15864
rect 5776 15852 5782 15904
rect 5994 15852 6000 15904
rect 6052 15892 6058 15904
rect 6089 15895 6147 15901
rect 6089 15892 6101 15895
rect 6052 15864 6101 15892
rect 6052 15852 6058 15864
rect 6089 15861 6101 15864
rect 6135 15892 6147 15895
rect 8110 15892 8116 15904
rect 6135 15864 8116 15892
rect 6135 15861 6147 15864
rect 6089 15855 6147 15861
rect 8110 15852 8116 15864
rect 8168 15852 8174 15904
rect 9582 15852 9588 15904
rect 9640 15892 9646 15904
rect 9766 15892 9772 15904
rect 9640 15864 9772 15892
rect 9640 15852 9646 15864
rect 9766 15852 9772 15864
rect 9824 15852 9830 15904
rect 10778 15892 10784 15904
rect 10739 15864 10784 15892
rect 10778 15852 10784 15864
rect 10836 15852 10842 15904
rect 11514 15852 11520 15904
rect 11572 15892 11578 15904
rect 12360 15892 12388 15923
rect 13906 15920 13912 15932
rect 13964 15920 13970 15972
rect 11572 15864 12388 15892
rect 11572 15852 11578 15864
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 1489 15691 1547 15697
rect 1489 15657 1501 15691
rect 1535 15688 1547 15691
rect 1578 15688 1584 15700
rect 1535 15660 1584 15688
rect 1535 15657 1547 15660
rect 1489 15651 1547 15657
rect 1578 15648 1584 15660
rect 1636 15648 1642 15700
rect 1762 15688 1768 15700
rect 1723 15660 1768 15688
rect 1762 15648 1768 15660
rect 1820 15648 1826 15700
rect 1946 15648 1952 15700
rect 2004 15688 2010 15700
rect 2133 15691 2191 15697
rect 2133 15688 2145 15691
rect 2004 15660 2145 15688
rect 2004 15648 2010 15660
rect 2133 15657 2145 15660
rect 2179 15657 2191 15691
rect 2133 15651 2191 15657
rect 2409 15691 2467 15697
rect 2409 15657 2421 15691
rect 2455 15688 2467 15691
rect 2498 15688 2504 15700
rect 2455 15660 2504 15688
rect 2455 15657 2467 15660
rect 2409 15651 2467 15657
rect 2498 15648 2504 15660
rect 2556 15648 2562 15700
rect 2682 15688 2688 15700
rect 2643 15660 2688 15688
rect 2682 15648 2688 15660
rect 2740 15648 2746 15700
rect 2961 15691 3019 15697
rect 2961 15657 2973 15691
rect 3007 15688 3019 15691
rect 3326 15688 3332 15700
rect 3007 15660 3332 15688
rect 3007 15657 3019 15660
rect 2961 15651 3019 15657
rect 3326 15648 3332 15660
rect 3384 15648 3390 15700
rect 3602 15688 3608 15700
rect 3563 15660 3608 15688
rect 3602 15648 3608 15660
rect 3660 15648 3666 15700
rect 3881 15691 3939 15697
rect 3881 15657 3893 15691
rect 3927 15688 3939 15691
rect 4430 15688 4436 15700
rect 3927 15660 4436 15688
rect 3927 15657 3939 15660
rect 3881 15651 3939 15657
rect 4430 15648 4436 15660
rect 4488 15648 4494 15700
rect 4522 15648 4528 15700
rect 4580 15688 4586 15700
rect 5258 15688 5264 15700
rect 4580 15660 5264 15688
rect 4580 15648 4586 15660
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 6178 15648 6184 15700
rect 6236 15688 6242 15700
rect 6273 15691 6331 15697
rect 6273 15688 6285 15691
rect 6236 15660 6285 15688
rect 6236 15648 6242 15660
rect 6273 15657 6285 15660
rect 6319 15657 6331 15691
rect 6273 15651 6331 15657
rect 7193 15691 7251 15697
rect 7193 15657 7205 15691
rect 7239 15688 7251 15691
rect 7374 15688 7380 15700
rect 7239 15660 7380 15688
rect 7239 15657 7251 15660
rect 7193 15651 7251 15657
rect 7374 15648 7380 15660
rect 7432 15648 7438 15700
rect 9950 15688 9956 15700
rect 9911 15660 9956 15688
rect 9950 15648 9956 15660
rect 10008 15648 10014 15700
rect 10042 15648 10048 15700
rect 10100 15688 10106 15700
rect 10965 15691 11023 15697
rect 10965 15688 10977 15691
rect 10100 15660 10977 15688
rect 10100 15648 10106 15660
rect 10965 15657 10977 15660
rect 11011 15657 11023 15691
rect 10965 15651 11023 15657
rect 13262 15648 13268 15700
rect 13320 15688 13326 15700
rect 15378 15688 15384 15700
rect 13320 15660 15384 15688
rect 13320 15648 13326 15660
rect 15378 15648 15384 15660
rect 15436 15648 15442 15700
rect 2590 15580 2596 15632
rect 2648 15620 2654 15632
rect 3237 15623 3295 15629
rect 3237 15620 3249 15623
rect 2648 15592 3249 15620
rect 2648 15580 2654 15592
rect 3237 15589 3249 15592
rect 3283 15589 3295 15623
rect 4062 15620 4068 15632
rect 4023 15592 4068 15620
rect 3237 15583 3295 15589
rect 4062 15580 4068 15592
rect 4120 15580 4126 15632
rect 7006 15620 7012 15632
rect 6656 15592 7012 15620
rect 4522 15552 4528 15564
rect 1688 15524 4528 15552
rect 1688 15493 1716 15524
rect 4522 15512 4528 15524
rect 4580 15512 4586 15564
rect 6656 15561 6684 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 10778 15620 10784 15632
rect 10520 15592 10784 15620
rect 6641 15555 6699 15561
rect 6641 15521 6653 15555
rect 6687 15521 6699 15555
rect 8573 15555 8631 15561
rect 8573 15552 8585 15555
rect 6641 15515 6699 15521
rect 6840 15524 8585 15552
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1946 15484 1952 15496
rect 1907 15456 1952 15484
rect 1673 15447 1731 15453
rect 1946 15444 1952 15456
rect 2004 15444 2010 15496
rect 2314 15484 2320 15496
rect 2275 15456 2320 15484
rect 2314 15444 2320 15456
rect 2372 15444 2378 15496
rect 2498 15444 2504 15496
rect 2556 15484 2562 15496
rect 2593 15487 2651 15493
rect 2593 15484 2605 15487
rect 2556 15456 2605 15484
rect 2556 15444 2562 15456
rect 2593 15453 2605 15456
rect 2639 15453 2651 15487
rect 2593 15447 2651 15453
rect 2869 15487 2927 15493
rect 2869 15453 2881 15487
rect 2915 15453 2927 15487
rect 3142 15484 3148 15496
rect 3103 15456 3148 15484
rect 2869 15447 2927 15453
rect 2884 15348 2912 15447
rect 3142 15444 3148 15456
rect 3200 15444 3206 15496
rect 3421 15487 3479 15493
rect 3421 15453 3433 15487
rect 3467 15453 3479 15487
rect 3421 15447 3479 15453
rect 4157 15487 4215 15493
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4430 15484 4436 15496
rect 4203 15456 4436 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 3436 15416 3464 15447
rect 4430 15444 4436 15456
rect 4488 15444 4494 15496
rect 4893 15487 4951 15493
rect 4893 15453 4905 15487
rect 4939 15484 4951 15487
rect 5718 15484 5724 15496
rect 4939 15456 5724 15484
rect 4939 15453 4951 15456
rect 4893 15447 4951 15453
rect 5718 15444 5724 15456
rect 5776 15444 5782 15496
rect 5160 15419 5218 15425
rect 3436 15388 5120 15416
rect 3418 15348 3424 15360
rect 2884 15320 3424 15348
rect 3418 15308 3424 15320
rect 3476 15308 3482 15360
rect 4338 15308 4344 15360
rect 4396 15348 4402 15360
rect 4801 15351 4859 15357
rect 4801 15348 4813 15351
rect 4396 15320 4813 15348
rect 4396 15308 4402 15320
rect 4801 15317 4813 15320
rect 4847 15317 4859 15351
rect 5092 15348 5120 15388
rect 5160 15385 5172 15419
rect 5206 15416 5218 15419
rect 6656 15416 6684 15515
rect 6840 15493 6868 15524
rect 8573 15521 8585 15524
rect 8619 15521 8631 15555
rect 8573 15515 8631 15521
rect 9401 15555 9459 15561
rect 9401 15521 9413 15555
rect 9447 15552 9459 15555
rect 9766 15552 9772 15564
rect 9447 15524 9772 15552
rect 9447 15521 9459 15524
rect 9401 15515 9459 15521
rect 9766 15512 9772 15524
rect 9824 15512 9830 15564
rect 9950 15512 9956 15564
rect 10008 15552 10014 15564
rect 10520 15561 10548 15592
rect 10778 15580 10784 15592
rect 10836 15580 10842 15632
rect 12713 15623 12771 15629
rect 12713 15620 12725 15623
rect 12268 15592 12725 15620
rect 10505 15555 10563 15561
rect 10008 15524 10456 15552
rect 10008 15512 10014 15524
rect 6825 15487 6883 15493
rect 6825 15453 6837 15487
rect 6871 15453 6883 15487
rect 6825 15447 6883 15453
rect 7098 15444 7104 15496
rect 7156 15484 7162 15496
rect 7282 15484 7288 15496
rect 7156 15456 7288 15484
rect 7156 15444 7162 15456
rect 7282 15444 7288 15456
rect 7340 15444 7346 15496
rect 7558 15484 7564 15496
rect 7519 15456 7564 15484
rect 7558 15444 7564 15456
rect 7616 15444 7622 15496
rect 9122 15484 9128 15496
rect 9083 15456 9128 15484
rect 9122 15444 9128 15456
rect 9180 15444 9186 15496
rect 10428 15484 10456 15524
rect 10505 15521 10517 15555
rect 10551 15521 10563 15555
rect 10505 15515 10563 15521
rect 10689 15555 10747 15561
rect 10689 15521 10701 15555
rect 10735 15552 10747 15555
rect 10962 15552 10968 15564
rect 10735 15524 10968 15552
rect 10735 15521 10747 15524
rect 10689 15515 10747 15521
rect 10962 15512 10968 15524
rect 11020 15512 11026 15564
rect 11330 15512 11336 15564
rect 11388 15552 11394 15564
rect 11517 15555 11575 15561
rect 11517 15552 11529 15555
rect 11388 15524 11529 15552
rect 11388 15512 11394 15524
rect 11517 15521 11529 15524
rect 11563 15521 11575 15555
rect 11517 15515 11575 15521
rect 11698 15512 11704 15564
rect 11756 15512 11762 15564
rect 11716 15484 11744 15512
rect 12268 15493 12296 15592
rect 12713 15589 12725 15592
rect 12759 15589 12771 15623
rect 13722 15620 13728 15632
rect 12713 15583 12771 15589
rect 13372 15592 13728 15620
rect 13372 15561 13400 15592
rect 13722 15580 13728 15592
rect 13780 15580 13786 15632
rect 12529 15555 12587 15561
rect 12529 15521 12541 15555
rect 12575 15521 12587 15555
rect 12529 15515 12587 15521
rect 13357 15555 13415 15561
rect 13357 15521 13369 15555
rect 13403 15521 13415 15555
rect 13357 15515 13415 15521
rect 10428 15456 11744 15484
rect 12253 15487 12311 15493
rect 12253 15453 12265 15487
rect 12299 15453 12311 15487
rect 12544 15484 12572 15515
rect 13630 15512 13636 15564
rect 13688 15552 13694 15564
rect 14093 15555 14151 15561
rect 14093 15552 14105 15555
rect 13688 15524 14105 15552
rect 13688 15512 13694 15524
rect 14093 15521 14105 15524
rect 14139 15552 14151 15555
rect 14918 15552 14924 15564
rect 14139 15524 14924 15552
rect 14139 15521 14151 15524
rect 14093 15515 14151 15521
rect 14918 15512 14924 15524
rect 14976 15512 14982 15564
rect 12986 15484 12992 15496
rect 12544 15456 12992 15484
rect 12253 15447 12311 15453
rect 12986 15444 12992 15456
rect 13044 15484 13050 15496
rect 14182 15484 14188 15496
rect 13044 15456 14188 15484
rect 13044 15444 13050 15456
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 14369 15487 14427 15493
rect 14369 15453 14381 15487
rect 14415 15484 14427 15487
rect 14458 15484 14464 15496
rect 14415 15456 14464 15484
rect 14415 15453 14427 15456
rect 14369 15447 14427 15453
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15010 15484 15016 15496
rect 14971 15456 15016 15484
rect 15010 15444 15016 15456
rect 15068 15444 15074 15496
rect 15930 15484 15936 15496
rect 15304 15456 15936 15484
rect 5206 15388 6684 15416
rect 5206 15385 5218 15388
rect 5160 15379 5218 15385
rect 8110 15376 8116 15428
rect 8168 15416 8174 15428
rect 8205 15419 8263 15425
rect 8205 15416 8217 15419
rect 8168 15388 8217 15416
rect 8168 15376 8174 15388
rect 8205 15385 8217 15388
rect 8251 15385 8263 15419
rect 8205 15379 8263 15385
rect 8389 15419 8447 15425
rect 8389 15385 8401 15419
rect 8435 15416 8447 15419
rect 9030 15416 9036 15428
rect 8435 15388 9036 15416
rect 8435 15385 8447 15388
rect 8389 15379 8447 15385
rect 9030 15376 9036 15388
rect 9088 15376 9094 15428
rect 9585 15419 9643 15425
rect 9585 15385 9597 15419
rect 9631 15416 9643 15419
rect 9631 15388 10640 15416
rect 9631 15385 9643 15388
rect 9585 15379 9643 15385
rect 5442 15348 5448 15360
rect 5092 15320 5448 15348
rect 4801 15311 4859 15317
rect 5442 15308 5448 15320
rect 5500 15308 5506 15360
rect 6733 15351 6791 15357
rect 6733 15317 6745 15351
rect 6779 15348 6791 15351
rect 7374 15348 7380 15360
rect 6779 15320 7380 15348
rect 6779 15317 6791 15320
rect 6733 15311 6791 15317
rect 7374 15308 7380 15320
rect 7432 15308 7438 15360
rect 8938 15348 8944 15360
rect 8899 15320 8944 15348
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 9490 15348 9496 15360
rect 9451 15320 9496 15348
rect 9490 15308 9496 15320
rect 9548 15308 9554 15360
rect 10042 15348 10048 15360
rect 10003 15320 10048 15348
rect 10042 15308 10048 15320
rect 10100 15308 10106 15360
rect 10226 15308 10232 15360
rect 10284 15348 10290 15360
rect 10413 15351 10471 15357
rect 10413 15348 10425 15351
rect 10284 15320 10425 15348
rect 10284 15308 10290 15320
rect 10413 15317 10425 15320
rect 10459 15317 10471 15351
rect 10612 15348 10640 15388
rect 10686 15376 10692 15428
rect 10744 15416 10750 15428
rect 13725 15419 13783 15425
rect 10744 15388 11928 15416
rect 10744 15376 10750 15388
rect 10778 15348 10784 15360
rect 10612 15320 10784 15348
rect 10413 15311 10471 15317
rect 10778 15308 10784 15320
rect 10836 15308 10842 15360
rect 11330 15348 11336 15360
rect 11291 15320 11336 15348
rect 11330 15308 11336 15320
rect 11388 15308 11394 15360
rect 11425 15351 11483 15357
rect 11425 15317 11437 15351
rect 11471 15348 11483 15351
rect 11514 15348 11520 15360
rect 11471 15320 11520 15348
rect 11471 15317 11483 15320
rect 11425 15311 11483 15317
rect 11514 15308 11520 15320
rect 11572 15308 11578 15360
rect 11900 15357 11928 15388
rect 13725 15385 13737 15419
rect 13771 15416 13783 15419
rect 15304 15416 15332 15456
rect 15930 15444 15936 15456
rect 15988 15484 15994 15496
rect 16114 15484 16120 15496
rect 15988 15456 16120 15484
rect 15988 15444 15994 15456
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 15654 15416 15660 15428
rect 13771 15388 15332 15416
rect 15615 15388 15660 15416
rect 13771 15385 13783 15388
rect 13725 15379 13783 15385
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 11885 15351 11943 15357
rect 11885 15317 11897 15351
rect 11931 15317 11943 15351
rect 11885 15311 11943 15317
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15348 12403 15351
rect 12894 15348 12900 15360
rect 12391 15320 12900 15348
rect 12391 15317 12403 15320
rect 12345 15311 12403 15317
rect 12894 15308 12900 15320
rect 12952 15308 12958 15360
rect 13078 15348 13084 15360
rect 13039 15320 13084 15348
rect 13078 15308 13084 15320
rect 13136 15308 13142 15360
rect 13173 15351 13231 15357
rect 13173 15317 13185 15351
rect 13219 15348 13231 15351
rect 13262 15348 13268 15360
rect 13219 15320 13268 15348
rect 13219 15317 13231 15320
rect 13173 15311 13231 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 13630 15348 13636 15360
rect 13591 15320 13636 15348
rect 13630 15308 13636 15320
rect 13688 15308 13694 15360
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 4522 15104 4528 15156
rect 4580 15144 4586 15156
rect 5445 15147 5503 15153
rect 5445 15144 5457 15147
rect 4580 15116 5457 15144
rect 4580 15104 4586 15116
rect 5445 15113 5457 15116
rect 5491 15113 5503 15147
rect 5810 15144 5816 15156
rect 5771 15116 5816 15144
rect 5445 15107 5503 15113
rect 5810 15104 5816 15116
rect 5868 15104 5874 15156
rect 5905 15147 5963 15153
rect 5905 15113 5917 15147
rect 5951 15144 5963 15147
rect 6086 15144 6092 15156
rect 5951 15116 6092 15144
rect 5951 15113 5963 15116
rect 5905 15107 5963 15113
rect 6086 15104 6092 15116
rect 6144 15104 6150 15156
rect 6365 15147 6423 15153
rect 6365 15113 6377 15147
rect 6411 15144 6423 15147
rect 6454 15144 6460 15156
rect 6411 15116 6460 15144
rect 6411 15113 6423 15116
rect 6365 15107 6423 15113
rect 6454 15104 6460 15116
rect 6512 15104 6518 15156
rect 6914 15104 6920 15156
rect 6972 15144 6978 15156
rect 7193 15147 7251 15153
rect 7193 15144 7205 15147
rect 6972 15116 7205 15144
rect 6972 15104 6978 15116
rect 7193 15113 7205 15116
rect 7239 15113 7251 15147
rect 7193 15107 7251 15113
rect 7282 15104 7288 15156
rect 7340 15144 7346 15156
rect 8481 15147 8539 15153
rect 8481 15144 8493 15147
rect 7340 15116 8493 15144
rect 7340 15104 7346 15116
rect 8481 15113 8493 15116
rect 8527 15113 8539 15147
rect 9490 15144 9496 15156
rect 9451 15116 9496 15144
rect 8481 15107 8539 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 10042 15104 10048 15156
rect 10100 15144 10106 15156
rect 10870 15144 10876 15156
rect 10100 15116 10876 15144
rect 10100 15104 10106 15116
rect 10870 15104 10876 15116
rect 10928 15104 10934 15156
rect 10962 15104 10968 15156
rect 11020 15144 11026 15156
rect 11333 15147 11391 15153
rect 11333 15144 11345 15147
rect 11020 15116 11345 15144
rect 11020 15104 11026 15116
rect 11333 15113 11345 15116
rect 11379 15144 11391 15147
rect 11974 15144 11980 15156
rect 11379 15116 11980 15144
rect 11379 15113 11391 15116
rect 11333 15107 11391 15113
rect 11974 15104 11980 15116
rect 12032 15104 12038 15156
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15113 12311 15147
rect 12253 15107 12311 15113
rect 12345 15147 12403 15153
rect 12345 15113 12357 15147
rect 12391 15144 12403 15147
rect 12802 15144 12808 15156
rect 12391 15116 12808 15144
rect 12391 15113 12403 15116
rect 12345 15107 12403 15113
rect 5718 15076 5724 15088
rect 3068 15048 5724 15076
rect 2682 15008 2688 15020
rect 2740 15017 2746 15020
rect 3068 15017 3096 15048
rect 5718 15036 5724 15048
rect 5776 15036 5782 15088
rect 7561 15079 7619 15085
rect 7561 15076 7573 15079
rect 6012 15048 7573 15076
rect 3326 15017 3332 15020
rect 2652 14980 2688 15008
rect 2682 14968 2688 14980
rect 2740 14971 2752 15017
rect 2961 15011 3019 15017
rect 2961 14977 2973 15011
rect 3007 15008 3019 15011
rect 3053 15011 3111 15017
rect 3053 15008 3065 15011
rect 3007 14980 3065 15008
rect 3007 14977 3019 14980
rect 2961 14971 3019 14977
rect 3053 14977 3065 14980
rect 3099 14977 3111 15011
rect 3320 15008 3332 15017
rect 3287 14980 3332 15008
rect 3053 14971 3111 14977
rect 3320 14971 3332 14980
rect 2740 14968 2746 14971
rect 3326 14968 3332 14971
rect 3384 14968 3390 15020
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 4893 15011 4951 15017
rect 4893 15008 4905 15011
rect 4304 14980 4905 15008
rect 4304 14968 4310 14980
rect 4893 14977 4905 14980
rect 4939 15008 4951 15011
rect 5166 15008 5172 15020
rect 4939 14980 5172 15008
rect 4939 14977 4951 14980
rect 4893 14971 4951 14977
rect 5166 14968 5172 14980
rect 5224 15008 5230 15020
rect 5350 15008 5356 15020
rect 5224 14980 5356 15008
rect 5224 14968 5230 14980
rect 5350 14968 5356 14980
rect 5408 14968 5414 15020
rect 5442 14968 5448 15020
rect 5500 15008 5506 15020
rect 6012 15008 6040 15048
rect 7208 15020 7236 15048
rect 7561 15045 7573 15048
rect 7607 15045 7619 15079
rect 7561 15039 7619 15045
rect 8297 15079 8355 15085
rect 8297 15045 8309 15079
rect 8343 15076 8355 15079
rect 9030 15076 9036 15088
rect 8343 15048 9036 15076
rect 8343 15045 8355 15048
rect 8297 15039 8355 15045
rect 9030 15036 9036 15048
rect 9088 15036 9094 15088
rect 10226 15085 10232 15088
rect 10220 15076 10232 15085
rect 10187 15048 10232 15076
rect 10220 15039 10232 15048
rect 10226 15036 10232 15039
rect 10284 15036 10290 15088
rect 12158 15036 12164 15088
rect 12216 15076 12222 15088
rect 12268 15076 12296 15107
rect 12802 15104 12808 15116
rect 12860 15104 12866 15156
rect 12894 15104 12900 15156
rect 12952 15144 12958 15156
rect 12989 15147 13047 15153
rect 12989 15144 13001 15147
rect 12952 15116 13001 15144
rect 12952 15104 12958 15116
rect 12989 15113 13001 15116
rect 13035 15113 13047 15147
rect 12989 15107 13047 15113
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 15562 15144 15568 15156
rect 15252 15116 15568 15144
rect 15252 15104 15258 15116
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 12216 15048 12296 15076
rect 14001 15079 14059 15085
rect 12216 15036 12222 15048
rect 14001 15045 14013 15079
rect 14047 15076 14059 15079
rect 15010 15076 15016 15088
rect 14047 15048 15016 15076
rect 14047 15045 14059 15048
rect 14001 15039 14059 15045
rect 15010 15036 15016 15048
rect 15068 15076 15074 15088
rect 15286 15076 15292 15088
rect 15068 15048 15292 15076
rect 15068 15036 15074 15048
rect 15286 15036 15292 15048
rect 15344 15036 15350 15088
rect 6730 15008 6736 15020
rect 5500 14980 6040 15008
rect 6643 14980 6736 15008
rect 5500 14968 5506 14980
rect 6730 14968 6736 14980
rect 6788 14968 6794 15020
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 7098 15008 7104 15020
rect 6871 14980 7104 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 7190 14968 7196 15020
rect 7248 14968 7254 15020
rect 8665 15011 8723 15017
rect 8665 14977 8677 15011
rect 8711 15008 8723 15011
rect 8754 15008 8760 15020
rect 8711 14980 8760 15008
rect 8711 14977 8723 14980
rect 8665 14971 8723 14977
rect 8754 14968 8760 14980
rect 8812 14968 8818 15020
rect 8938 14968 8944 15020
rect 8996 15008 9002 15020
rect 9125 15011 9183 15017
rect 9125 15008 9137 15011
rect 8996 14980 9137 15008
rect 8996 14968 9002 14980
rect 9125 14977 9137 14980
rect 9171 15008 9183 15011
rect 9585 15011 9643 15017
rect 9585 15008 9597 15011
rect 9171 14980 9597 15008
rect 9171 14977 9183 14980
rect 9125 14971 9183 14977
rect 9585 14977 9597 14980
rect 9631 14977 9643 15011
rect 9585 14971 9643 14977
rect 11701 15011 11759 15017
rect 11701 14977 11713 15011
rect 11747 15008 11759 15011
rect 11747 15006 12204 15008
rect 12250 15006 12256 15020
rect 11747 14980 12256 15006
rect 11747 14977 11759 14980
rect 12176 14978 12256 14980
rect 11701 14971 11759 14977
rect 12250 14968 12256 14978
rect 12308 14968 12314 15020
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 12897 15011 12955 15017
rect 12897 15008 12909 15011
rect 12676 14980 12909 15008
rect 12676 14968 12682 14980
rect 12897 14977 12909 14980
rect 12943 14977 12955 15011
rect 12897 14971 12955 14977
rect 13357 15011 13415 15017
rect 13357 14977 13369 15011
rect 13403 15008 13415 15011
rect 13906 15008 13912 15020
rect 13403 14980 13912 15008
rect 13403 14977 13415 14980
rect 13357 14971 13415 14977
rect 13906 14968 13912 14980
rect 13964 14968 13970 15020
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 15008 14243 15011
rect 14366 15008 14372 15020
rect 14231 14980 14372 15008
rect 14231 14977 14243 14980
rect 14185 14971 14243 14977
rect 14366 14968 14372 14980
rect 14424 15008 14430 15020
rect 14642 15008 14648 15020
rect 14424 14980 14648 15008
rect 14424 14968 14430 14980
rect 14642 14968 14648 14980
rect 14700 14968 14706 15020
rect 15102 15008 15108 15020
rect 15063 14980 15108 15008
rect 15102 14968 15108 14980
rect 15160 14968 15166 15020
rect 4062 14900 4068 14952
rect 4120 14940 4126 14952
rect 4985 14943 5043 14949
rect 4985 14940 4997 14943
rect 4120 14912 4997 14940
rect 4120 14900 4126 14912
rect 4985 14909 4997 14912
rect 5031 14909 5043 14943
rect 4985 14903 5043 14909
rect 5077 14943 5135 14949
rect 5077 14909 5089 14943
rect 5123 14909 5135 14943
rect 5077 14903 5135 14909
rect 6089 14943 6147 14949
rect 6089 14909 6101 14943
rect 6135 14940 6147 14943
rect 6362 14940 6368 14952
rect 6135 14912 6368 14940
rect 6135 14909 6147 14912
rect 6089 14903 6147 14909
rect 1489 14875 1547 14881
rect 1489 14841 1501 14875
rect 1535 14872 1547 14875
rect 1535 14844 2084 14872
rect 1535 14841 1547 14844
rect 1489 14835 1547 14841
rect 1578 14804 1584 14816
rect 1539 14776 1584 14804
rect 1578 14764 1584 14776
rect 1636 14764 1642 14816
rect 2056 14804 2084 14844
rect 4614 14832 4620 14884
rect 4672 14872 4678 14884
rect 5092 14872 5120 14903
rect 6362 14900 6368 14912
rect 6420 14900 6426 14952
rect 6748 14940 6776 14968
rect 6914 14940 6920 14952
rect 6748 14912 6920 14940
rect 6914 14900 6920 14912
rect 6972 14900 6978 14952
rect 7006 14900 7012 14952
rect 7064 14940 7070 14952
rect 7650 14940 7656 14952
rect 7064 14912 7157 14940
rect 7611 14912 7656 14940
rect 7064 14900 7070 14912
rect 7650 14900 7656 14912
rect 7708 14900 7714 14952
rect 7837 14943 7895 14949
rect 7837 14909 7849 14943
rect 7883 14940 7895 14943
rect 8202 14940 8208 14952
rect 7883 14912 8208 14940
rect 7883 14909 7895 14912
rect 7837 14903 7895 14909
rect 4672 14844 5120 14872
rect 7024 14872 7052 14900
rect 7282 14872 7288 14884
rect 7024 14844 7288 14872
rect 4672 14832 4678 14844
rect 7282 14832 7288 14844
rect 7340 14872 7346 14884
rect 7852 14872 7880 14903
rect 8202 14900 8208 14912
rect 8260 14900 8266 14952
rect 8846 14940 8852 14952
rect 8807 14912 8852 14940
rect 8846 14900 8852 14912
rect 8904 14900 8910 14952
rect 9033 14943 9091 14949
rect 9033 14909 9045 14943
rect 9079 14940 9091 14943
rect 9766 14940 9772 14952
rect 9079 14912 9772 14940
rect 9079 14909 9091 14912
rect 9033 14903 9091 14909
rect 9766 14900 9772 14912
rect 9824 14900 9830 14952
rect 9953 14943 10011 14949
rect 9953 14909 9965 14943
rect 9999 14909 10011 14943
rect 9953 14903 10011 14909
rect 7340 14844 7880 14872
rect 7340 14832 7346 14844
rect 4246 14804 4252 14816
rect 2056 14776 4252 14804
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4430 14804 4436 14816
rect 4391 14776 4436 14804
rect 4430 14764 4436 14776
rect 4488 14764 4494 14816
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4580 14776 4625 14804
rect 4580 14764 4586 14776
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 8205 14807 8263 14813
rect 8205 14804 8217 14807
rect 5224 14776 8217 14804
rect 5224 14764 5230 14776
rect 8205 14773 8217 14776
rect 8251 14773 8263 14807
rect 8205 14767 8263 14773
rect 8846 14764 8852 14816
rect 8904 14804 8910 14816
rect 9306 14804 9312 14816
rect 8904 14776 9312 14804
rect 8904 14764 8910 14776
rect 9306 14764 9312 14776
rect 9364 14764 9370 14816
rect 9769 14807 9827 14813
rect 9769 14773 9781 14807
rect 9815 14804 9827 14807
rect 9858 14804 9864 14816
rect 9815 14776 9864 14804
rect 9815 14773 9827 14776
rect 9769 14767 9827 14773
rect 9858 14764 9864 14776
rect 9916 14764 9922 14816
rect 9968 14804 9996 14903
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 12434 14940 12440 14952
rect 11020 14912 11652 14940
rect 12395 14912 12440 14940
rect 11020 14900 11026 14912
rect 11514 14872 11520 14884
rect 11475 14844 11520 14872
rect 11514 14832 11520 14844
rect 11572 14832 11578 14884
rect 11624 14872 11652 14912
rect 12434 14900 12440 14912
rect 12492 14900 12498 14952
rect 13078 14900 13084 14952
rect 13136 14940 13142 14952
rect 13449 14943 13507 14949
rect 13449 14940 13461 14943
rect 13136 14912 13461 14940
rect 13136 14900 13142 14912
rect 13449 14909 13461 14912
rect 13495 14909 13507 14943
rect 13449 14903 13507 14909
rect 13633 14943 13691 14949
rect 13633 14909 13645 14943
rect 13679 14940 13691 14943
rect 13722 14940 13728 14952
rect 13679 14912 13728 14940
rect 13679 14909 13691 14912
rect 13633 14903 13691 14909
rect 13722 14900 13728 14912
rect 13780 14900 13786 14952
rect 14461 14943 14519 14949
rect 14461 14909 14473 14943
rect 14507 14940 14519 14943
rect 14550 14940 14556 14952
rect 14507 14912 14556 14940
rect 14507 14909 14519 14912
rect 14461 14903 14519 14909
rect 14550 14900 14556 14912
rect 14608 14900 14614 14952
rect 14734 14900 14740 14952
rect 14792 14900 14798 14952
rect 11624 14844 12434 14872
rect 10962 14804 10968 14816
rect 9968 14776 10968 14804
rect 10962 14764 10968 14776
rect 11020 14764 11026 14816
rect 11882 14804 11888 14816
rect 11843 14776 11888 14804
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 12406 14804 12434 14844
rect 12894 14832 12900 14884
rect 12952 14872 12958 14884
rect 14752 14872 14780 14900
rect 15102 14872 15108 14884
rect 12952 14844 15108 14872
rect 12952 14832 12958 14844
rect 15102 14832 15108 14844
rect 15160 14832 15166 14884
rect 15838 14872 15844 14884
rect 15396 14844 15844 14872
rect 12713 14807 12771 14813
rect 12713 14804 12725 14807
rect 12406 14776 12725 14804
rect 12713 14773 12725 14776
rect 12759 14773 12771 14807
rect 12713 14767 12771 14773
rect 13909 14807 13967 14813
rect 13909 14773 13921 14807
rect 13955 14804 13967 14807
rect 14734 14804 14740 14816
rect 13955 14776 14740 14804
rect 13955 14773 13967 14776
rect 13909 14767 13967 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 15396 14813 15424 14844
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 15381 14807 15439 14813
rect 15381 14773 15393 14807
rect 15427 14773 15439 14807
rect 15381 14767 15439 14773
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1486 14600 1492 14612
rect 1447 14572 1492 14600
rect 1486 14560 1492 14572
rect 1544 14560 1550 14612
rect 4356 14572 7144 14600
rect 2866 14532 2872 14544
rect 2827 14504 2872 14532
rect 2866 14492 2872 14504
rect 2924 14492 2930 14544
rect 1578 14424 1584 14476
rect 1636 14464 1642 14476
rect 2133 14467 2191 14473
rect 2133 14464 2145 14467
rect 1636 14436 2145 14464
rect 1636 14424 1642 14436
rect 2133 14433 2145 14436
rect 2179 14464 2191 14467
rect 3326 14464 3332 14476
rect 2179 14436 3332 14464
rect 2179 14433 2191 14436
rect 2133 14427 2191 14433
rect 3326 14424 3332 14436
rect 3384 14464 3390 14476
rect 3421 14467 3479 14473
rect 3421 14464 3433 14467
rect 3384 14436 3433 14464
rect 3384 14424 3390 14436
rect 3421 14433 3433 14436
rect 3467 14433 3479 14467
rect 3421 14427 3479 14433
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 3973 14467 4031 14473
rect 3973 14464 3985 14467
rect 3752 14436 3985 14464
rect 3752 14424 3758 14436
rect 3973 14433 3985 14436
rect 4019 14464 4031 14467
rect 4062 14464 4068 14476
rect 4019 14436 4068 14464
rect 4019 14433 4031 14436
rect 3973 14427 4031 14433
rect 4062 14424 4068 14436
rect 4120 14424 4126 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1949 14399 2007 14405
rect 1719 14368 1808 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 1780 14269 1808 14368
rect 1949 14365 1961 14399
rect 1995 14396 2007 14399
rect 4356 14396 4384 14572
rect 5626 14492 5632 14544
rect 5684 14532 5690 14544
rect 6086 14532 6092 14544
rect 5684 14504 6092 14532
rect 5684 14492 5690 14504
rect 6086 14492 6092 14504
rect 6144 14492 6150 14544
rect 7116 14532 7144 14572
rect 7650 14560 7656 14612
rect 7708 14600 7714 14612
rect 7745 14603 7803 14609
rect 7745 14600 7757 14603
rect 7708 14572 7757 14600
rect 7708 14560 7714 14572
rect 7745 14569 7757 14572
rect 7791 14569 7803 14603
rect 9217 14603 9275 14609
rect 9217 14600 9229 14603
rect 7745 14563 7803 14569
rect 7852 14572 9229 14600
rect 7852 14532 7880 14572
rect 9217 14569 9229 14572
rect 9263 14569 9275 14603
rect 11882 14600 11888 14612
rect 9217 14563 9275 14569
rect 10704 14572 11888 14600
rect 10502 14532 10508 14544
rect 7116 14504 7880 14532
rect 8404 14504 10508 14532
rect 8404 14473 8432 14504
rect 10502 14492 10508 14504
rect 10560 14492 10566 14544
rect 5905 14467 5963 14473
rect 5905 14464 5917 14467
rect 5460 14436 5917 14464
rect 1995 14368 4384 14396
rect 4433 14399 4491 14405
rect 1995 14365 2007 14368
rect 1949 14359 2007 14365
rect 4433 14365 4445 14399
rect 4479 14396 4491 14399
rect 4479 14368 4660 14396
rect 4479 14365 4491 14368
rect 4433 14359 4491 14365
rect 2409 14331 2467 14337
rect 2409 14297 2421 14331
rect 2455 14328 2467 14331
rect 2958 14328 2964 14340
rect 2455 14300 2964 14328
rect 2455 14297 2467 14300
rect 2409 14291 2467 14297
rect 2958 14288 2964 14300
rect 3016 14288 3022 14340
rect 3329 14331 3387 14337
rect 3329 14297 3341 14331
rect 3375 14328 3387 14331
rect 4522 14328 4528 14340
rect 3375 14300 4528 14328
rect 3375 14297 3387 14300
rect 3329 14291 3387 14297
rect 4522 14288 4528 14300
rect 4580 14288 4586 14340
rect 1765 14263 1823 14269
rect 1765 14229 1777 14263
rect 1811 14229 1823 14263
rect 2314 14260 2320 14272
rect 2275 14232 2320 14260
rect 1765 14223 1823 14229
rect 2314 14220 2320 14232
rect 2372 14220 2378 14272
rect 2774 14220 2780 14272
rect 2832 14260 2838 14272
rect 3237 14263 3295 14269
rect 2832 14232 2877 14260
rect 2832 14220 2838 14232
rect 3237 14229 3249 14263
rect 3283 14260 3295 14263
rect 3602 14260 3608 14272
rect 3283 14232 3608 14260
rect 3283 14229 3295 14232
rect 3237 14223 3295 14229
rect 3602 14220 3608 14232
rect 3660 14220 3666 14272
rect 3878 14260 3884 14272
rect 3839 14232 3884 14260
rect 3878 14220 3884 14232
rect 3936 14220 3942 14272
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4632 14260 4660 14368
rect 4706 14337 4712 14340
rect 4700 14291 4712 14337
rect 4764 14328 4770 14340
rect 4764 14300 4800 14328
rect 4706 14288 4712 14291
rect 4764 14288 4770 14300
rect 5350 14288 5356 14340
rect 5408 14328 5414 14340
rect 5460 14328 5488 14436
rect 5905 14433 5917 14436
rect 5951 14433 5963 14467
rect 5905 14427 5963 14433
rect 8389 14467 8447 14473
rect 8389 14433 8401 14467
rect 8435 14433 8447 14467
rect 8389 14427 8447 14433
rect 9214 14424 9220 14476
rect 9272 14464 9278 14476
rect 9769 14467 9827 14473
rect 9769 14464 9781 14467
rect 9272 14436 9781 14464
rect 9272 14424 9278 14436
rect 9769 14433 9781 14436
rect 9815 14433 9827 14467
rect 10318 14464 10324 14476
rect 10279 14436 10324 14464
rect 9769 14427 9827 14433
rect 10318 14424 10324 14436
rect 10376 14424 10382 14476
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 6181 14399 6239 14405
rect 6181 14396 6193 14399
rect 5776 14368 6193 14396
rect 5776 14356 5782 14368
rect 6181 14365 6193 14368
rect 6227 14396 6239 14399
rect 7742 14396 7748 14408
rect 6227 14368 7748 14396
rect 6227 14365 6239 14368
rect 6181 14359 6239 14365
rect 7742 14356 7748 14368
rect 7800 14356 7806 14408
rect 8110 14396 8116 14408
rect 8023 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14396 8174 14408
rect 9677 14399 9735 14405
rect 9677 14396 9689 14399
rect 8168 14368 9076 14396
rect 8168 14356 8174 14368
rect 5736 14328 5764 14356
rect 6454 14337 6460 14340
rect 6448 14328 6460 14337
rect 5408 14300 5488 14328
rect 5552 14300 5764 14328
rect 5828 14300 6460 14328
rect 5408 14288 5414 14300
rect 5552 14260 5580 14300
rect 4632 14232 5580 14260
rect 5626 14220 5632 14272
rect 5684 14260 5690 14272
rect 5828 14269 5856 14300
rect 6448 14291 6460 14300
rect 6454 14288 6460 14291
rect 6512 14288 6518 14340
rect 6822 14288 6828 14340
rect 6880 14328 6886 14340
rect 8205 14331 8263 14337
rect 8205 14328 8217 14331
rect 6880 14300 8217 14328
rect 6880 14288 6886 14300
rect 8205 14297 8217 14300
rect 8251 14297 8263 14331
rect 8754 14328 8760 14340
rect 8205 14291 8263 14297
rect 8588 14300 8760 14328
rect 5813 14263 5871 14269
rect 5813 14260 5825 14263
rect 5684 14232 5825 14260
rect 5684 14220 5690 14232
rect 5813 14229 5825 14232
rect 5859 14229 5871 14263
rect 5813 14223 5871 14229
rect 7006 14220 7012 14272
rect 7064 14260 7070 14272
rect 7561 14263 7619 14269
rect 7561 14260 7573 14263
rect 7064 14232 7573 14260
rect 7064 14220 7070 14232
rect 7561 14229 7573 14232
rect 7607 14229 7619 14263
rect 7561 14223 7619 14229
rect 8110 14220 8116 14272
rect 8168 14260 8174 14272
rect 8588 14260 8616 14300
rect 8754 14288 8760 14300
rect 8812 14328 8818 14340
rect 8941 14331 8999 14337
rect 8941 14328 8953 14331
rect 8812 14300 8953 14328
rect 8812 14288 8818 14300
rect 8941 14297 8953 14300
rect 8987 14297 8999 14331
rect 8941 14291 8999 14297
rect 8168 14232 8616 14260
rect 8665 14263 8723 14269
rect 8168 14220 8174 14232
rect 8665 14229 8677 14263
rect 8711 14260 8723 14263
rect 8846 14260 8852 14272
rect 8711 14232 8852 14260
rect 8711 14229 8723 14232
rect 8665 14223 8723 14229
rect 8846 14220 8852 14232
rect 8904 14220 8910 14272
rect 9048 14260 9076 14368
rect 9508 14368 9689 14396
rect 9122 14288 9128 14340
rect 9180 14328 9186 14340
rect 9508 14328 9536 14368
rect 9677 14365 9689 14368
rect 9723 14365 9735 14399
rect 9677 14359 9735 14365
rect 10505 14399 10563 14405
rect 10505 14365 10517 14399
rect 10551 14396 10563 14399
rect 10704 14396 10732 14572
rect 11882 14560 11888 14572
rect 11940 14560 11946 14612
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 16942 14600 16948 14612
rect 12667 14572 16948 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 16942 14560 16948 14572
rect 17000 14560 17006 14612
rect 12345 14535 12403 14541
rect 12345 14501 12357 14535
rect 12391 14532 12403 14535
rect 13722 14532 13728 14544
rect 12391 14504 13728 14532
rect 12391 14501 12403 14504
rect 12345 14495 12403 14501
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 15102 14492 15108 14544
rect 15160 14532 15166 14544
rect 15565 14535 15623 14541
rect 15565 14532 15577 14535
rect 15160 14504 15577 14532
rect 15160 14492 15166 14504
rect 15565 14501 15577 14504
rect 15611 14501 15623 14535
rect 15565 14495 15623 14501
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 12710 14464 12716 14476
rect 12584 14436 12716 14464
rect 12584 14424 12590 14436
rect 12710 14424 12716 14436
rect 12768 14424 12774 14476
rect 12986 14424 12992 14476
rect 13044 14464 13050 14476
rect 13081 14467 13139 14473
rect 13081 14464 13093 14467
rect 13044 14436 13093 14464
rect 13044 14424 13050 14436
rect 13081 14433 13093 14436
rect 13127 14433 13139 14467
rect 13081 14427 13139 14433
rect 10962 14396 10968 14408
rect 10551 14368 10732 14396
rect 10923 14368 10968 14396
rect 10551 14365 10563 14368
rect 10505 14359 10563 14365
rect 10962 14356 10968 14368
rect 11020 14356 11026 14408
rect 11232 14399 11290 14405
rect 11232 14365 11244 14399
rect 11278 14396 11290 14399
rect 11698 14396 11704 14408
rect 11278 14368 11704 14396
rect 11278 14365 11290 14368
rect 11232 14359 11290 14365
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 12437 14399 12495 14405
rect 12437 14365 12449 14399
rect 12483 14396 12495 14399
rect 12483 14368 13032 14396
rect 12483 14365 12495 14368
rect 12437 14359 12495 14365
rect 9180 14300 9536 14328
rect 9585 14331 9643 14337
rect 9180 14288 9186 14300
rect 9585 14297 9597 14331
rect 9631 14328 9643 14331
rect 12710 14328 12716 14340
rect 9631 14300 11100 14328
rect 12671 14300 12716 14328
rect 9631 14297 9643 14300
rect 9585 14291 9643 14297
rect 9490 14260 9496 14272
rect 9048 14232 9496 14260
rect 9490 14220 9496 14232
rect 9548 14220 9554 14272
rect 9674 14220 9680 14272
rect 9732 14260 9738 14272
rect 10318 14260 10324 14272
rect 9732 14232 10324 14260
rect 9732 14220 9738 14232
rect 10318 14220 10324 14232
rect 10376 14220 10382 14272
rect 10413 14263 10471 14269
rect 10413 14229 10425 14263
rect 10459 14260 10471 14263
rect 10686 14260 10692 14272
rect 10459 14232 10692 14260
rect 10459 14229 10471 14232
rect 10413 14223 10471 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 10870 14260 10876 14272
rect 10831 14232 10876 14260
rect 10870 14220 10876 14232
rect 10928 14220 10934 14272
rect 11072 14260 11100 14300
rect 12710 14288 12716 14300
rect 12768 14288 12774 14340
rect 12894 14328 12900 14340
rect 12855 14300 12900 14328
rect 12894 14288 12900 14300
rect 12952 14288 12958 14340
rect 11974 14260 11980 14272
rect 11072 14232 11980 14260
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 13004 14260 13032 14368
rect 13170 14356 13176 14408
rect 13228 14396 13234 14408
rect 13357 14399 13415 14405
rect 13357 14396 13369 14399
rect 13228 14368 13369 14396
rect 13228 14356 13234 14368
rect 13357 14365 13369 14368
rect 13403 14365 13415 14399
rect 13357 14359 13415 14365
rect 13814 14356 13820 14408
rect 13872 14396 13878 14408
rect 14093 14399 14151 14405
rect 14093 14396 14105 14399
rect 13872 14368 14105 14396
rect 13872 14356 13878 14368
rect 14093 14365 14105 14368
rect 14139 14365 14151 14399
rect 14093 14359 14151 14365
rect 13722 14288 13728 14340
rect 13780 14328 13786 14340
rect 14338 14331 14396 14337
rect 14338 14328 14350 14331
rect 13780 14300 14350 14328
rect 13780 14288 13786 14300
rect 14338 14297 14350 14300
rect 14384 14297 14396 14331
rect 14338 14291 14396 14297
rect 15286 14288 15292 14340
rect 15344 14328 15350 14340
rect 15344 14300 15516 14328
rect 15344 14288 15350 14300
rect 15378 14260 15384 14272
rect 13004 14232 15384 14260
rect 15378 14220 15384 14232
rect 15436 14220 15442 14272
rect 15488 14269 15516 14300
rect 15473 14263 15531 14269
rect 15473 14229 15485 14263
rect 15519 14229 15531 14263
rect 15473 14223 15531 14229
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 1765 14059 1823 14065
rect 1765 14025 1777 14059
rect 1811 14025 1823 14059
rect 1765 14019 1823 14025
rect 2501 14059 2559 14065
rect 2501 14025 2513 14059
rect 2547 14056 2559 14059
rect 2866 14056 2872 14068
rect 2547 14028 2872 14056
rect 2547 14025 2559 14028
rect 2501 14019 2559 14025
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13920 1731 13923
rect 1780 13920 1808 14019
rect 2866 14016 2872 14028
rect 2924 14016 2930 14068
rect 2958 14016 2964 14068
rect 3016 14056 3022 14068
rect 3016 14028 3061 14056
rect 3016 14016 3022 14028
rect 3602 14016 3608 14068
rect 3660 14056 3666 14068
rect 3789 14059 3847 14065
rect 3789 14056 3801 14059
rect 3660 14028 3801 14056
rect 3660 14016 3666 14028
rect 3789 14025 3801 14028
rect 3835 14025 3847 14059
rect 4154 14056 4160 14068
rect 4115 14028 4160 14056
rect 3789 14019 3847 14025
rect 4154 14016 4160 14028
rect 4212 14016 4218 14068
rect 4246 14016 4252 14068
rect 4304 14056 4310 14068
rect 4985 14059 5043 14065
rect 4985 14056 4997 14059
rect 4304 14028 4997 14056
rect 4304 14016 4310 14028
rect 4985 14025 4997 14028
rect 5031 14056 5043 14059
rect 5166 14056 5172 14068
rect 5031 14028 5172 14056
rect 5031 14025 5043 14028
rect 4985 14019 5043 14025
rect 5166 14016 5172 14028
rect 5224 14016 5230 14068
rect 5353 14059 5411 14065
rect 5353 14025 5365 14059
rect 5399 14025 5411 14059
rect 5353 14019 5411 14025
rect 2409 13991 2467 13997
rect 2409 13957 2421 13991
rect 2455 13988 2467 13991
rect 2774 13988 2780 14000
rect 2455 13960 2780 13988
rect 2455 13957 2467 13960
rect 2409 13951 2467 13957
rect 2774 13948 2780 13960
rect 2832 13948 2838 14000
rect 3234 13948 3240 14000
rect 3292 13988 3298 14000
rect 3329 13991 3387 13997
rect 3329 13988 3341 13991
rect 3292 13960 3341 13988
rect 3292 13948 3298 13960
rect 3329 13957 3341 13960
rect 3375 13957 3387 13991
rect 3329 13951 3387 13957
rect 4522 13948 4528 14000
rect 4580 13988 4586 14000
rect 4893 13991 4951 13997
rect 4893 13988 4905 13991
rect 4580 13960 4905 13988
rect 4580 13948 4586 13960
rect 4893 13957 4905 13960
rect 4939 13957 4951 13991
rect 5368 13988 5396 14019
rect 5442 14016 5448 14068
rect 5500 14056 5506 14068
rect 5721 14059 5779 14065
rect 5721 14056 5733 14059
rect 5500 14028 5733 14056
rect 5500 14016 5506 14028
rect 5721 14025 5733 14028
rect 5767 14025 5779 14059
rect 5721 14019 5779 14025
rect 6181 14059 6239 14065
rect 6181 14025 6193 14059
rect 6227 14056 6239 14059
rect 6733 14059 6791 14065
rect 6733 14056 6745 14059
rect 6227 14028 6745 14056
rect 6227 14025 6239 14028
rect 6181 14019 6239 14025
rect 6733 14025 6745 14028
rect 6779 14025 6791 14059
rect 7374 14056 7380 14068
rect 7335 14028 7380 14056
rect 6733 14019 6791 14025
rect 7374 14016 7380 14028
rect 7432 14056 7438 14068
rect 7650 14056 7656 14068
rect 7432 14028 7656 14056
rect 7432 14016 7438 14028
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 10134 14056 10140 14068
rect 7760 14028 10140 14056
rect 6825 13991 6883 13997
rect 6825 13988 6837 13991
rect 5368 13960 6837 13988
rect 4893 13951 4951 13957
rect 6825 13957 6837 13960
rect 6871 13957 6883 13991
rect 6825 13951 6883 13957
rect 1719 13892 1808 13920
rect 1949 13923 2007 13929
rect 1719 13889 1731 13892
rect 1673 13883 1731 13889
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 2590 13920 2596 13932
rect 1995 13892 2596 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2590 13880 2596 13892
rect 2648 13880 2654 13932
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13920 3479 13923
rect 4338 13920 4344 13932
rect 3467 13892 4344 13920
rect 3467 13889 3479 13892
rect 3421 13883 3479 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 4908 13920 4936 13951
rect 6914 13948 6920 14000
rect 6972 13988 6978 14000
rect 7285 13991 7343 13997
rect 7285 13988 7297 13991
rect 6972 13960 7297 13988
rect 6972 13948 6978 13960
rect 7285 13957 7297 13960
rect 7331 13988 7343 13991
rect 7760 13988 7788 14028
rect 10134 14016 10140 14028
rect 10192 14016 10198 14068
rect 10318 14016 10324 14068
rect 10376 14056 10382 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 10376 14028 11345 14056
rect 10376 14016 10382 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11974 14056 11980 14068
rect 11935 14028 11980 14056
rect 11333 14019 11391 14025
rect 11974 14016 11980 14028
rect 12032 14016 12038 14068
rect 12345 14059 12403 14065
rect 12345 14025 12357 14059
rect 12391 14056 12403 14059
rect 12802 14056 12808 14068
rect 12391 14028 12572 14056
rect 12763 14028 12808 14056
rect 12391 14025 12403 14028
rect 12345 14019 12403 14025
rect 7331 13960 7788 13988
rect 7331 13957 7343 13960
rect 7285 13951 7343 13957
rect 9573 13948 9579 14000
rect 9631 13988 9637 14000
rect 10962 13988 10968 14000
rect 9631 13960 10968 13988
rect 9631 13948 9637 13960
rect 10962 13948 10968 13960
rect 11020 13948 11026 14000
rect 11238 13948 11244 14000
rect 11296 13988 11302 14000
rect 11517 13991 11575 13997
rect 11517 13988 11529 13991
rect 11296 13960 11529 13988
rect 11296 13948 11302 13960
rect 11517 13957 11529 13960
rect 11563 13957 11575 13991
rect 12544 13988 12572 14028
rect 12802 14016 12808 14028
rect 12860 14016 12866 14068
rect 12894 14016 12900 14068
rect 12952 14056 12958 14068
rect 13262 14056 13268 14068
rect 12952 14028 13268 14056
rect 12952 14016 12958 14028
rect 13262 14016 13268 14028
rect 13320 14016 13326 14068
rect 13354 14016 13360 14068
rect 13412 14056 13418 14068
rect 13722 14056 13728 14068
rect 13412 14028 13728 14056
rect 13412 14016 13418 14028
rect 13722 14016 13728 14028
rect 13780 14016 13786 14068
rect 12618 13988 12624 14000
rect 12544 13960 12624 13988
rect 11517 13951 11575 13957
rect 12618 13948 12624 13960
rect 12676 13948 12682 14000
rect 13998 13988 14004 14000
rect 13096 13960 14004 13988
rect 5813 13923 5871 13929
rect 4908 13892 5764 13920
rect 2317 13855 2375 13861
rect 2317 13821 2329 13855
rect 2363 13821 2375 13855
rect 2317 13815 2375 13821
rect 1486 13784 1492 13796
rect 1447 13756 1492 13784
rect 1486 13744 1492 13756
rect 1544 13744 1550 13796
rect 2332 13716 2360 13815
rect 2682 13812 2688 13864
rect 2740 13852 2746 13864
rect 3513 13855 3571 13861
rect 3513 13852 3525 13855
rect 2740 13824 3525 13852
rect 2740 13812 2746 13824
rect 3513 13821 3525 13824
rect 3559 13852 3571 13855
rect 3878 13852 3884 13864
rect 3559 13824 3884 13852
rect 3559 13821 3571 13824
rect 3513 13815 3571 13821
rect 3878 13812 3884 13824
rect 3936 13852 3942 13864
rect 3936 13824 4108 13852
rect 3936 13812 3942 13824
rect 2869 13787 2927 13793
rect 2869 13753 2881 13787
rect 2915 13784 2927 13787
rect 3970 13784 3976 13796
rect 2915 13756 3976 13784
rect 2915 13753 2927 13756
rect 2869 13747 2927 13753
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 4080 13784 4108 13824
rect 4154 13812 4160 13864
rect 4212 13852 4218 13864
rect 4249 13855 4307 13861
rect 4249 13852 4261 13855
rect 4212 13824 4261 13852
rect 4212 13812 4218 13824
rect 4249 13821 4261 13824
rect 4295 13821 4307 13855
rect 4249 13815 4307 13821
rect 4433 13855 4491 13861
rect 4433 13821 4445 13855
rect 4479 13852 4491 13855
rect 4614 13852 4620 13864
rect 4479 13824 4620 13852
rect 4479 13821 4491 13824
rect 4433 13815 4491 13821
rect 4448 13784 4476 13815
rect 4614 13812 4620 13824
rect 4672 13812 4678 13864
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 5537 13855 5595 13861
rect 5537 13821 5549 13855
rect 5583 13821 5595 13855
rect 5736 13852 5764 13892
rect 5813 13889 5825 13923
rect 5859 13920 5871 13923
rect 5902 13920 5908 13932
rect 5859 13892 5908 13920
rect 5859 13889 5871 13892
rect 5813 13883 5871 13889
rect 5902 13880 5908 13892
rect 5960 13920 5966 13932
rect 7558 13920 7564 13932
rect 5960 13892 7564 13920
rect 5960 13880 5966 13892
rect 7558 13880 7564 13892
rect 7616 13880 7622 13932
rect 7742 13920 7748 13932
rect 7703 13892 7748 13920
rect 7742 13880 7748 13892
rect 7800 13880 7806 13932
rect 8018 13929 8024 13932
rect 8012 13883 8024 13929
rect 8076 13920 8082 13932
rect 8076 13892 8112 13920
rect 8018 13880 8024 13883
rect 8076 13880 8082 13892
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 8754 13920 8760 13932
rect 8352 13892 8760 13920
rect 8352 13880 8358 13892
rect 8754 13880 8760 13892
rect 8812 13920 8818 13932
rect 9217 13923 9275 13929
rect 9217 13920 9229 13923
rect 8812 13892 9229 13920
rect 8812 13880 8818 13892
rect 9217 13889 9229 13892
rect 9263 13889 9275 13923
rect 9217 13883 9275 13889
rect 9306 13880 9312 13932
rect 9364 13920 9370 13932
rect 9473 13923 9531 13929
rect 9473 13920 9485 13923
rect 9364 13892 9485 13920
rect 9364 13880 9370 13892
rect 9473 13889 9485 13892
rect 9519 13889 9531 13923
rect 9473 13883 9531 13889
rect 10502 13880 10508 13932
rect 10560 13920 10566 13932
rect 10689 13923 10747 13929
rect 10689 13920 10701 13923
rect 10560 13892 10701 13920
rect 10560 13880 10566 13892
rect 10689 13889 10701 13892
rect 10735 13889 10747 13923
rect 10689 13883 10747 13889
rect 12437 13923 12495 13929
rect 12437 13889 12449 13923
rect 12483 13920 12495 13923
rect 13096 13920 13124 13960
rect 13998 13948 14004 13960
rect 14056 13948 14062 14000
rect 12483 13892 13124 13920
rect 13173 13923 13231 13929
rect 12483 13889 12495 13892
rect 12437 13883 12495 13889
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 6822 13852 6828 13864
rect 5736 13824 6828 13852
rect 5537 13815 5595 13821
rect 4080 13756 4476 13784
rect 4816 13784 4844 13815
rect 5552 13784 5580 13815
rect 6822 13812 6828 13824
rect 6880 13812 6886 13864
rect 7006 13852 7012 13864
rect 6967 13824 7012 13852
rect 7006 13812 7012 13824
rect 7064 13812 7070 13864
rect 11885 13855 11943 13861
rect 11885 13821 11897 13855
rect 11931 13852 11943 13855
rect 11931 13824 12388 13852
rect 11931 13821 11943 13824
rect 11885 13815 11943 13821
rect 5626 13784 5632 13796
rect 4816 13756 5632 13784
rect 5626 13744 5632 13756
rect 5684 13744 5690 13796
rect 6178 13744 6184 13796
rect 6236 13784 6242 13796
rect 7561 13787 7619 13793
rect 7561 13784 7573 13787
rect 6236 13756 7573 13784
rect 6236 13744 6242 13756
rect 7561 13753 7573 13756
rect 7607 13753 7619 13787
rect 7561 13747 7619 13753
rect 9125 13787 9183 13793
rect 9125 13753 9137 13787
rect 9171 13784 9183 13787
rect 9214 13784 9220 13796
rect 9171 13756 9220 13784
rect 9171 13753 9183 13756
rect 9125 13747 9183 13753
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 10502 13744 10508 13796
rect 10560 13784 10566 13796
rect 10597 13787 10655 13793
rect 10597 13784 10609 13787
rect 10560 13756 10609 13784
rect 10560 13744 10566 13756
rect 10597 13753 10609 13756
rect 10643 13753 10655 13787
rect 10597 13747 10655 13753
rect 11698 13744 11704 13796
rect 11756 13784 11762 13796
rect 12158 13784 12164 13796
rect 11756 13756 12164 13784
rect 11756 13744 11762 13756
rect 12158 13744 12164 13756
rect 12216 13744 12222 13796
rect 4430 13716 4436 13728
rect 2332 13688 4436 13716
rect 4430 13676 4436 13688
rect 4488 13676 4494 13728
rect 6362 13676 6368 13728
rect 6420 13716 6426 13728
rect 6420 13688 6465 13716
rect 6420 13676 6426 13688
rect 8018 13676 8024 13728
rect 8076 13716 8082 13728
rect 10134 13716 10140 13728
rect 8076 13688 10140 13716
rect 8076 13676 8082 13688
rect 10134 13676 10140 13688
rect 10192 13676 10198 13728
rect 11238 13676 11244 13728
rect 11296 13716 11302 13728
rect 11882 13716 11888 13728
rect 11296 13688 11888 13716
rect 11296 13676 11302 13688
rect 11882 13676 11888 13688
rect 11940 13676 11946 13728
rect 12360 13716 12388 13824
rect 12526 13812 12532 13864
rect 12584 13852 12590 13864
rect 12584 13824 12629 13852
rect 12584 13812 12590 13824
rect 12986 13812 12992 13864
rect 13044 13852 13050 13864
rect 13188 13852 13216 13883
rect 13262 13880 13268 13932
rect 13320 13920 13326 13932
rect 13633 13923 13691 13929
rect 13633 13920 13645 13923
rect 13320 13892 13645 13920
rect 13320 13880 13326 13892
rect 13633 13889 13645 13892
rect 13679 13889 13691 13923
rect 13633 13883 13691 13889
rect 13354 13852 13360 13864
rect 13044 13824 13216 13852
rect 13315 13824 13360 13852
rect 13044 13812 13050 13824
rect 13354 13812 13360 13824
rect 13412 13812 13418 13864
rect 13906 13852 13912 13864
rect 13867 13824 13912 13852
rect 13906 13812 13912 13824
rect 13964 13812 13970 13864
rect 15470 13852 15476 13864
rect 15431 13824 15476 13852
rect 15470 13812 15476 13824
rect 15528 13812 15534 13864
rect 15657 13855 15715 13861
rect 15657 13821 15669 13855
rect 15703 13852 15715 13855
rect 15746 13852 15752 13864
rect 15703 13824 15752 13852
rect 15703 13821 15715 13824
rect 15657 13815 15715 13821
rect 15746 13812 15752 13824
rect 15804 13812 15810 13864
rect 15010 13716 15016 13728
rect 12360 13688 15016 13716
rect 15010 13676 15016 13688
rect 15068 13676 15074 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 2314 13472 2320 13524
rect 2372 13512 2378 13524
rect 2685 13515 2743 13521
rect 2685 13512 2697 13515
rect 2372 13484 2697 13512
rect 2372 13472 2378 13484
rect 2685 13481 2697 13484
rect 2731 13481 2743 13515
rect 5166 13512 5172 13524
rect 5127 13484 5172 13512
rect 2685 13475 2743 13481
rect 5166 13472 5172 13484
rect 5224 13472 5230 13524
rect 5718 13512 5724 13524
rect 5679 13484 5724 13512
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 7282 13472 7288 13524
rect 7340 13512 7346 13524
rect 7377 13515 7435 13521
rect 7377 13512 7389 13515
rect 7340 13484 7389 13512
rect 7340 13472 7346 13484
rect 7377 13481 7389 13484
rect 7423 13481 7435 13515
rect 7377 13475 7435 13481
rect 7466 13472 7472 13524
rect 7524 13512 7530 13524
rect 8846 13512 8852 13524
rect 7524 13484 8852 13512
rect 7524 13472 7530 13484
rect 8846 13472 8852 13484
rect 8904 13512 8910 13524
rect 8941 13515 8999 13521
rect 8941 13512 8953 13515
rect 8904 13484 8953 13512
rect 8904 13472 8910 13484
rect 8941 13481 8953 13484
rect 8987 13481 8999 13515
rect 9582 13512 9588 13524
rect 9543 13484 9588 13512
rect 8941 13475 8999 13481
rect 9582 13472 9588 13484
rect 9640 13472 9646 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11885 13515 11943 13521
rect 11885 13512 11897 13515
rect 11020 13484 11897 13512
rect 11020 13472 11026 13484
rect 11885 13481 11897 13484
rect 11931 13512 11943 13515
rect 13814 13512 13820 13524
rect 11931 13484 13820 13512
rect 11931 13481 11943 13484
rect 11885 13475 11943 13481
rect 13814 13472 13820 13484
rect 13872 13472 13878 13524
rect 13906 13472 13912 13524
rect 13964 13512 13970 13524
rect 14093 13515 14151 13521
rect 14093 13512 14105 13515
rect 13964 13484 14105 13512
rect 13964 13472 13970 13484
rect 14093 13481 14105 13484
rect 14139 13481 14151 13515
rect 14093 13475 14151 13481
rect 3789 13447 3847 13453
rect 3789 13444 3801 13447
rect 1688 13416 3801 13444
rect 1688 13317 1716 13416
rect 3789 13413 3801 13416
rect 3835 13413 3847 13447
rect 3789 13407 3847 13413
rect 4154 13404 4160 13456
rect 4212 13444 4218 13456
rect 4249 13447 4307 13453
rect 4249 13444 4261 13447
rect 4212 13416 4261 13444
rect 4212 13404 4218 13416
rect 4249 13413 4261 13416
rect 4295 13444 4307 13447
rect 5810 13444 5816 13456
rect 4295 13416 5816 13444
rect 4295 13413 4307 13416
rect 4249 13407 4307 13413
rect 5810 13404 5816 13416
rect 5868 13404 5874 13456
rect 9493 13447 9551 13453
rect 9493 13413 9505 13447
rect 9539 13444 9551 13447
rect 9950 13444 9956 13456
rect 9539 13416 9956 13444
rect 9539 13413 9551 13416
rect 9493 13407 9551 13413
rect 9950 13404 9956 13416
rect 10008 13404 10014 13456
rect 10870 13404 10876 13456
rect 10928 13444 10934 13456
rect 12066 13444 12072 13456
rect 10928 13416 12072 13444
rect 10928 13404 10934 13416
rect 12066 13404 12072 13416
rect 12124 13404 12130 13456
rect 12250 13444 12256 13456
rect 12163 13416 12256 13444
rect 12250 13404 12256 13416
rect 12308 13404 12314 13456
rect 14274 13404 14280 13456
rect 14332 13444 14338 13456
rect 15286 13444 15292 13456
rect 14332 13416 15292 13444
rect 14332 13404 14338 13416
rect 15286 13404 15292 13416
rect 15344 13404 15350 13456
rect 2866 13336 2872 13388
rect 2924 13376 2930 13388
rect 3234 13376 3240 13388
rect 2924 13348 3240 13376
rect 2924 13336 2930 13348
rect 3234 13336 3240 13348
rect 3292 13336 3298 13388
rect 3329 13379 3387 13385
rect 3329 13345 3341 13379
rect 3375 13376 3387 13379
rect 3878 13376 3884 13388
rect 3375 13348 3884 13376
rect 3375 13345 3387 13348
rect 3329 13339 3387 13345
rect 3878 13336 3884 13348
rect 3936 13336 3942 13388
rect 4617 13379 4675 13385
rect 4617 13345 4629 13379
rect 4663 13345 4675 13379
rect 4617 13339 4675 13345
rect 4709 13379 4767 13385
rect 4709 13345 4721 13379
rect 4755 13376 4767 13379
rect 6362 13376 6368 13388
rect 4755 13348 6368 13376
rect 4755 13345 4767 13348
rect 4709 13339 4767 13345
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 2593 13311 2651 13317
rect 2593 13277 2605 13311
rect 2639 13308 2651 13311
rect 3053 13311 3111 13317
rect 2639 13280 2774 13308
rect 2639 13277 2651 13280
rect 2593 13271 2651 13277
rect 1302 13200 1308 13252
rect 1360 13240 1366 13252
rect 1765 13243 1823 13249
rect 1765 13240 1777 13243
rect 1360 13212 1777 13240
rect 1360 13200 1366 13212
rect 1765 13209 1777 13212
rect 1811 13240 1823 13243
rect 2222 13240 2228 13252
rect 1811 13212 2228 13240
rect 1811 13209 1823 13212
rect 1765 13203 1823 13209
rect 2222 13200 2228 13212
rect 2280 13200 2286 13252
rect 2746 13240 2774 13280
rect 3053 13277 3065 13311
rect 3099 13308 3111 13311
rect 3142 13308 3148 13320
rect 3099 13280 3148 13308
rect 3099 13277 3111 13280
rect 3053 13271 3111 13277
rect 3142 13268 3148 13280
rect 3200 13308 3206 13320
rect 3510 13308 3516 13320
rect 3200 13280 3516 13308
rect 3200 13268 3206 13280
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 3970 13308 3976 13320
rect 3931 13280 3976 13308
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 4632 13308 4660 13339
rect 6362 13336 6368 13348
rect 6420 13336 6426 13388
rect 8754 13376 8760 13388
rect 8715 13348 8760 13376
rect 8754 13336 8760 13348
rect 8812 13336 8818 13388
rect 10134 13376 10140 13388
rect 10095 13348 10140 13376
rect 10134 13336 10140 13348
rect 10192 13376 10198 13388
rect 12268 13376 12296 13404
rect 10192 13348 12296 13376
rect 10192 13336 10198 13348
rect 14366 13336 14372 13388
rect 14424 13376 14430 13388
rect 14645 13379 14703 13385
rect 14645 13376 14657 13379
rect 14424 13348 14657 13376
rect 14424 13336 14430 13348
rect 14645 13345 14657 13348
rect 14691 13345 14703 13379
rect 15562 13376 15568 13388
rect 15523 13348 15568 13376
rect 14645 13339 14703 13345
rect 15562 13336 15568 13348
rect 15620 13336 15626 13388
rect 6270 13308 6276 13320
rect 4632 13280 6276 13308
rect 6270 13268 6276 13280
rect 6328 13268 6334 13320
rect 8501 13311 8559 13317
rect 8501 13277 8513 13311
rect 8547 13308 8559 13311
rect 9122 13308 9128 13320
rect 8547 13280 9128 13308
rect 8547 13277 8559 13280
rect 8501 13271 8559 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9309 13311 9367 13317
rect 9309 13277 9321 13311
rect 9355 13308 9367 13311
rect 9355 13280 12112 13308
rect 9355 13277 9367 13280
rect 9309 13271 9367 13277
rect 3234 13240 3240 13252
rect 2746 13212 3240 13240
rect 3234 13200 3240 13212
rect 3292 13200 3298 13252
rect 4801 13243 4859 13249
rect 4801 13209 4813 13243
rect 4847 13240 4859 13243
rect 5350 13240 5356 13252
rect 4847 13212 5356 13240
rect 4847 13209 4859 13212
rect 4801 13203 4859 13209
rect 5350 13200 5356 13212
rect 5408 13200 5414 13252
rect 7006 13240 7012 13252
rect 6967 13212 7012 13240
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 8662 13200 8668 13252
rect 8720 13240 8726 13252
rect 9582 13240 9588 13252
rect 8720 13212 9588 13240
rect 8720 13200 8726 13212
rect 9582 13200 9588 13212
rect 9640 13200 9646 13252
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 10045 13243 10103 13249
rect 10045 13240 10057 13243
rect 9732 13212 10057 13240
rect 9732 13200 9738 13212
rect 10045 13209 10057 13212
rect 10091 13209 10103 13243
rect 10045 13203 10103 13209
rect 10226 13200 10232 13252
rect 10284 13240 10290 13252
rect 10413 13243 10471 13249
rect 10413 13240 10425 13243
rect 10284 13212 10425 13240
rect 10284 13200 10290 13212
rect 10413 13209 10425 13212
rect 10459 13209 10471 13243
rect 10413 13203 10471 13209
rect 11330 13200 11336 13252
rect 11388 13240 11394 13252
rect 12084 13240 12112 13280
rect 12802 13268 12808 13320
rect 12860 13308 12866 13320
rect 13633 13311 13691 13317
rect 12860 13280 13483 13308
rect 12860 13268 12866 13280
rect 12434 13240 12440 13252
rect 11388 13212 12020 13240
rect 12084 13212 12440 13240
rect 11388 13200 11394 13212
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1946 13172 1952 13184
rect 1907 13144 1952 13172
rect 1946 13132 1952 13144
rect 2004 13132 2010 13184
rect 3145 13175 3203 13181
rect 3145 13141 3157 13175
rect 3191 13172 3203 13175
rect 3418 13172 3424 13184
rect 3191 13144 3424 13172
rect 3191 13141 3203 13144
rect 3145 13135 3203 13141
rect 3418 13132 3424 13144
rect 3476 13132 3482 13184
rect 4157 13175 4215 13181
rect 4157 13141 4169 13175
rect 4203 13172 4215 13175
rect 6822 13172 6828 13184
rect 4203 13144 6828 13172
rect 4203 13141 4215 13144
rect 4157 13135 4215 13141
rect 6822 13132 6828 13144
rect 6880 13132 6886 13184
rect 6914 13132 6920 13184
rect 6972 13172 6978 13184
rect 7193 13175 7251 13181
rect 7193 13172 7205 13175
rect 6972 13144 7205 13172
rect 6972 13132 6978 13144
rect 7193 13141 7205 13144
rect 7239 13172 7251 13175
rect 8018 13172 8024 13184
rect 7239 13144 8024 13172
rect 7239 13141 7251 13144
rect 7193 13135 7251 13141
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 9953 13175 10011 13181
rect 9953 13141 9965 13175
rect 9999 13172 10011 13175
rect 11514 13172 11520 13184
rect 9999 13144 11520 13172
rect 9999 13141 10011 13144
rect 9953 13135 10011 13141
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 11992 13172 12020 13212
rect 12434 13200 12440 13212
rect 12492 13200 12498 13252
rect 12618 13200 12624 13252
rect 12676 13240 12682 13252
rect 13262 13240 13268 13252
rect 12676 13212 13268 13240
rect 12676 13200 12682 13212
rect 13262 13200 13268 13212
rect 13320 13240 13326 13252
rect 13366 13243 13424 13249
rect 13366 13240 13378 13243
rect 13320 13212 13378 13240
rect 13320 13200 13326 13212
rect 13366 13209 13378 13212
rect 13412 13209 13424 13243
rect 13455 13240 13483 13280
rect 13633 13277 13645 13311
rect 13679 13277 13691 13311
rect 13633 13271 13691 13277
rect 13648 13240 13676 13271
rect 14090 13268 14096 13320
rect 14148 13308 14154 13320
rect 15381 13311 15439 13317
rect 15381 13308 15393 13311
rect 14148 13280 15393 13308
rect 14148 13268 14154 13280
rect 15381 13277 15393 13280
rect 15427 13277 15439 13311
rect 15381 13271 15439 13277
rect 13455 13212 13676 13240
rect 13366 13203 13424 13209
rect 13906 13200 13912 13252
rect 13964 13240 13970 13252
rect 15289 13243 15347 13249
rect 13964 13212 14964 13240
rect 13964 13200 13970 13212
rect 13725 13175 13783 13181
rect 13725 13172 13737 13175
rect 11992 13144 13737 13172
rect 13725 13141 13737 13144
rect 13771 13141 13783 13175
rect 13725 13135 13783 13141
rect 14182 13132 14188 13184
rect 14240 13172 14246 13184
rect 14461 13175 14519 13181
rect 14461 13172 14473 13175
rect 14240 13144 14473 13172
rect 14240 13132 14246 13144
rect 14461 13141 14473 13144
rect 14507 13141 14519 13175
rect 14461 13135 14519 13141
rect 14550 13132 14556 13184
rect 14608 13172 14614 13184
rect 14936 13181 14964 13212
rect 15289 13209 15301 13243
rect 15335 13240 15347 13243
rect 15654 13240 15660 13252
rect 15335 13212 15660 13240
rect 15335 13209 15347 13212
rect 15289 13203 15347 13209
rect 15654 13200 15660 13212
rect 15712 13200 15718 13252
rect 14921 13175 14979 13181
rect 14608 13144 14653 13172
rect 14608 13132 14614 13144
rect 14921 13141 14933 13175
rect 14967 13141 14979 13175
rect 14921 13135 14979 13141
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 1946 12928 1952 12980
rect 2004 12968 2010 12980
rect 2004 12940 3188 12968
rect 2004 12928 2010 12940
rect 3160 12900 3188 12940
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 3292 12940 3337 12968
rect 3292 12928 3298 12940
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 4709 12971 4767 12977
rect 4709 12968 4721 12971
rect 4672 12940 4721 12968
rect 4672 12928 4678 12940
rect 4709 12937 4721 12940
rect 4755 12937 4767 12971
rect 4709 12931 4767 12937
rect 4985 12971 5043 12977
rect 4985 12937 4997 12971
rect 5031 12968 5043 12971
rect 5074 12968 5080 12980
rect 5031 12940 5080 12968
rect 5031 12937 5043 12940
rect 4985 12931 5043 12937
rect 5074 12928 5080 12940
rect 5132 12928 5138 12980
rect 5350 12968 5356 12980
rect 5311 12940 5356 12968
rect 5350 12928 5356 12940
rect 5408 12928 5414 12980
rect 5813 12971 5871 12977
rect 5813 12937 5825 12971
rect 5859 12968 5871 12971
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 5859 12940 6377 12968
rect 5859 12937 5871 12940
rect 5813 12931 5871 12937
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6730 12968 6736 12980
rect 6691 12940 6736 12968
rect 6365 12931 6423 12937
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7466 12928 7472 12980
rect 7524 12968 7530 12980
rect 7653 12971 7711 12977
rect 7653 12968 7665 12971
rect 7524 12940 7665 12968
rect 7524 12928 7530 12940
rect 7653 12937 7665 12940
rect 7699 12937 7711 12971
rect 7653 12931 7711 12937
rect 8110 12928 8116 12980
rect 8168 12968 8174 12980
rect 8168 12940 8984 12968
rect 8168 12928 8174 12940
rect 3574 12903 3632 12909
rect 3574 12900 3586 12903
rect 1872 12872 3096 12900
rect 3160 12872 3586 12900
rect 1872 12841 1900 12872
rect 2130 12841 2136 12844
rect 1857 12835 1915 12841
rect 1857 12801 1869 12835
rect 1903 12801 1915 12835
rect 1857 12795 1915 12801
rect 2124 12795 2136 12841
rect 2188 12832 2194 12844
rect 3068 12832 3096 12872
rect 3574 12869 3586 12872
rect 3620 12869 3632 12903
rect 5258 12900 5264 12912
rect 5219 12872 5264 12900
rect 3574 12863 3632 12869
rect 5258 12860 5264 12872
rect 5316 12900 5322 12912
rect 5721 12903 5779 12909
rect 5721 12900 5733 12903
rect 5316 12872 5733 12900
rect 5316 12860 5322 12872
rect 5721 12869 5733 12872
rect 5767 12900 5779 12903
rect 6178 12900 6184 12912
rect 5767 12872 6184 12900
rect 5767 12869 5779 12872
rect 5721 12863 5779 12869
rect 6178 12860 6184 12872
rect 6236 12860 6242 12912
rect 7745 12903 7803 12909
rect 7745 12869 7757 12903
rect 7791 12900 7803 12903
rect 8849 12903 8907 12909
rect 8849 12900 8861 12903
rect 7791 12872 8861 12900
rect 7791 12869 7803 12872
rect 7745 12863 7803 12869
rect 8849 12869 8861 12872
rect 8895 12869 8907 12903
rect 8956 12900 8984 12940
rect 9306 12928 9312 12980
rect 9364 12968 9370 12980
rect 9769 12971 9827 12977
rect 9769 12968 9781 12971
rect 9364 12940 9781 12968
rect 9364 12928 9370 12940
rect 9769 12937 9781 12940
rect 9815 12937 9827 12971
rect 9769 12931 9827 12937
rect 9858 12928 9864 12980
rect 9916 12968 9922 12980
rect 10321 12971 10379 12977
rect 10321 12968 10333 12971
rect 9916 12940 10333 12968
rect 9916 12928 9922 12940
rect 10321 12937 10333 12940
rect 10367 12937 10379 12971
rect 10962 12968 10968 12980
rect 10923 12940 10968 12968
rect 10321 12931 10379 12937
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 11149 12971 11207 12977
rect 11149 12937 11161 12971
rect 11195 12968 11207 12971
rect 11238 12968 11244 12980
rect 11195 12940 11244 12968
rect 11195 12937 11207 12940
rect 11149 12931 11207 12937
rect 11164 12900 11192 12931
rect 11238 12928 11244 12940
rect 11296 12928 11302 12980
rect 11514 12968 11520 12980
rect 11475 12940 11520 12968
rect 11514 12928 11520 12940
rect 11572 12928 11578 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 14090 12968 14096 12980
rect 12124 12940 14096 12968
rect 12124 12928 12130 12940
rect 14090 12928 14096 12940
rect 14148 12928 14154 12980
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 14734 12968 14740 12980
rect 14507 12940 14740 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 14826 12928 14832 12980
rect 14884 12968 14890 12980
rect 15013 12971 15071 12977
rect 15013 12968 15025 12971
rect 14884 12940 15025 12968
rect 14884 12928 14890 12940
rect 15013 12937 15025 12940
rect 15059 12937 15071 12971
rect 15013 12931 15071 12937
rect 12986 12900 12992 12912
rect 8956 12872 11192 12900
rect 12899 12872 12992 12900
rect 8849 12863 8907 12869
rect 3142 12832 3148 12844
rect 2188 12804 2224 12832
rect 3055 12804 3148 12832
rect 2130 12792 2136 12795
rect 2188 12792 2194 12804
rect 3142 12792 3148 12804
rect 3200 12832 3206 12844
rect 3329 12835 3387 12841
rect 3329 12832 3341 12835
rect 3200 12804 3341 12832
rect 3200 12792 3206 12804
rect 3329 12801 3341 12804
rect 3375 12801 3387 12835
rect 3329 12795 3387 12801
rect 4062 12792 4068 12844
rect 4120 12832 4126 12844
rect 4120 12804 6123 12832
rect 4120 12792 4126 12804
rect 5997 12767 6055 12773
rect 5997 12733 6009 12767
rect 6043 12733 6055 12767
rect 6095 12764 6123 12804
rect 6454 12792 6460 12844
rect 6512 12832 6518 12844
rect 8110 12832 8116 12844
rect 6512 12804 6960 12832
rect 8071 12804 8116 12832
rect 6512 12792 6518 12804
rect 6822 12764 6828 12776
rect 6095 12736 6828 12764
rect 5997 12727 6055 12733
rect 2866 12656 2872 12708
rect 2924 12656 2930 12708
rect 6012 12696 6040 12727
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6932 12773 6960 12804
rect 8110 12792 8116 12804
rect 8168 12792 8174 12844
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 7834 12764 7840 12776
rect 7156 12736 7840 12764
rect 7156 12724 7162 12736
rect 7834 12724 7840 12736
rect 7892 12724 7898 12776
rect 8864 12764 8892 12863
rect 12986 12860 12992 12872
rect 13044 12900 13050 12912
rect 14752 12900 14780 12928
rect 13044 12872 14412 12900
rect 14752 12872 15148 12900
rect 13044 12860 13050 12872
rect 9125 12835 9183 12841
rect 9125 12801 9137 12835
rect 9171 12832 9183 12835
rect 9214 12832 9220 12844
rect 9171 12804 9220 12832
rect 9171 12801 9183 12804
rect 9125 12795 9183 12801
rect 9214 12792 9220 12804
rect 9272 12792 9278 12844
rect 9766 12792 9772 12844
rect 9824 12832 9830 12844
rect 9950 12832 9956 12844
rect 9824 12804 9956 12832
rect 9824 12792 9830 12804
rect 9950 12792 9956 12804
rect 10008 12832 10014 12844
rect 10413 12835 10471 12841
rect 10413 12832 10425 12835
rect 10008 12804 10425 12832
rect 10008 12792 10014 12804
rect 10413 12801 10425 12804
rect 10459 12801 10471 12835
rect 10413 12795 10471 12801
rect 10502 12792 10508 12844
rect 10560 12832 10566 12844
rect 11514 12832 11520 12844
rect 10560 12804 11520 12832
rect 10560 12792 10566 12804
rect 11514 12792 11520 12804
rect 11572 12832 11578 12844
rect 11885 12835 11943 12841
rect 11885 12832 11897 12835
rect 11572 12804 11897 12832
rect 11572 12792 11578 12804
rect 11885 12801 11897 12804
rect 11931 12832 11943 12835
rect 12345 12835 12403 12841
rect 12345 12832 12357 12835
rect 11931 12804 12357 12832
rect 11931 12801 11943 12804
rect 11885 12795 11943 12801
rect 12345 12801 12357 12804
rect 12391 12801 12403 12835
rect 13906 12832 13912 12844
rect 13867 12804 13912 12832
rect 12345 12795 12403 12801
rect 13906 12792 13912 12804
rect 13964 12792 13970 12844
rect 10597 12767 10655 12773
rect 8864 12736 9168 12764
rect 7116 12696 7144 12724
rect 6012 12668 7144 12696
rect 8757 12699 8815 12705
rect 1578 12628 1584 12640
rect 1539 12600 1584 12628
rect 1578 12588 1584 12600
rect 1636 12588 1642 12640
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 2222 12628 2228 12640
rect 1811 12600 2228 12628
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 2222 12588 2228 12600
rect 2280 12628 2286 12640
rect 2884 12628 2912 12656
rect 6104 12640 6132 12668
rect 8757 12665 8769 12699
rect 8803 12696 8815 12699
rect 9030 12696 9036 12708
rect 8803 12668 9036 12696
rect 8803 12665 8815 12668
rect 8757 12659 8815 12665
rect 9030 12656 9036 12668
rect 9088 12656 9094 12708
rect 9140 12640 9168 12736
rect 10597 12733 10609 12767
rect 10643 12764 10655 12767
rect 10778 12764 10784 12776
rect 10643 12736 10784 12764
rect 10643 12733 10655 12736
rect 10597 12727 10655 12733
rect 10778 12724 10784 12736
rect 10836 12724 10842 12776
rect 11333 12767 11391 12773
rect 11333 12733 11345 12767
rect 11379 12764 11391 12767
rect 11698 12764 11704 12776
rect 11379 12736 11704 12764
rect 11379 12733 11391 12736
rect 11333 12727 11391 12733
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 11974 12764 11980 12776
rect 11935 12736 11980 12764
rect 11974 12724 11980 12736
rect 12032 12724 12038 12776
rect 12161 12767 12219 12773
rect 12161 12733 12173 12767
rect 12207 12733 12219 12767
rect 12802 12764 12808 12776
rect 12763 12736 12808 12764
rect 12161 12727 12219 12733
rect 9766 12656 9772 12708
rect 9824 12696 9830 12708
rect 10042 12696 10048 12708
rect 9824 12668 10048 12696
rect 9824 12656 9830 12668
rect 10042 12656 10048 12668
rect 10100 12656 10106 12708
rect 12176 12696 12204 12727
rect 12802 12724 12808 12736
rect 12860 12724 12866 12776
rect 13262 12764 13268 12776
rect 13223 12736 13268 12764
rect 13262 12724 13268 12736
rect 13320 12724 13326 12776
rect 13814 12724 13820 12776
rect 13872 12764 13878 12776
rect 14274 12764 14280 12776
rect 13872 12736 14280 12764
rect 13872 12724 13878 12736
rect 14274 12724 14280 12736
rect 14332 12724 14338 12776
rect 14384 12764 14412 12872
rect 15120 12844 15148 12872
rect 14553 12835 14611 12841
rect 14553 12801 14565 12835
rect 14599 12832 14611 12835
rect 15010 12832 15016 12844
rect 14599 12804 15016 12832
rect 14599 12801 14611 12804
rect 14553 12795 14611 12801
rect 15010 12792 15016 12804
rect 15068 12792 15074 12844
rect 15102 12792 15108 12844
rect 15160 12792 15166 12844
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15620 12804 15669 12832
rect 15620 12792 15626 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 16298 12764 16304 12776
rect 14384 12736 16304 12764
rect 16298 12724 16304 12736
rect 16356 12724 16362 12776
rect 12526 12696 12532 12708
rect 12176 12668 12532 12696
rect 12526 12656 12532 12668
rect 12584 12656 12590 12708
rect 14921 12699 14979 12705
rect 14921 12665 14933 12699
rect 14967 12696 14979 12699
rect 15286 12696 15292 12708
rect 14967 12668 15292 12696
rect 14967 12665 14979 12668
rect 14921 12659 14979 12665
rect 15286 12656 15292 12668
rect 15344 12656 15350 12708
rect 2280 12600 2912 12628
rect 2280 12588 2286 12600
rect 6086 12588 6092 12640
rect 6144 12588 6150 12640
rect 6454 12588 6460 12640
rect 6512 12628 6518 12640
rect 7285 12631 7343 12637
rect 7285 12628 7297 12631
rect 6512 12600 7297 12628
rect 6512 12588 6518 12600
rect 7285 12597 7297 12600
rect 7331 12597 7343 12631
rect 7285 12591 7343 12597
rect 9122 12588 9128 12640
rect 9180 12588 9186 12640
rect 9953 12631 10011 12637
rect 9953 12597 9965 12631
rect 9999 12628 10011 12631
rect 10134 12628 10140 12640
rect 9999 12600 10140 12628
rect 9999 12597 10011 12600
rect 9953 12591 10011 12597
rect 10134 12588 10140 12600
rect 10192 12588 10198 12640
rect 10962 12588 10968 12640
rect 11020 12628 11026 12640
rect 11146 12628 11152 12640
rect 11020 12600 11152 12628
rect 11020 12588 11026 12600
rect 11146 12588 11152 12600
rect 11204 12588 11210 12640
rect 13630 12588 13636 12640
rect 13688 12628 13694 12640
rect 15010 12628 15016 12640
rect 13688 12600 15016 12628
rect 13688 12588 13694 12600
rect 15010 12588 15016 12600
rect 15068 12588 15074 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 2130 12424 2136 12436
rect 2091 12396 2136 12424
rect 2130 12384 2136 12396
rect 2188 12384 2194 12436
rect 3145 12427 3203 12433
rect 3145 12393 3157 12427
rect 3191 12424 3203 12427
rect 3326 12424 3332 12436
rect 3191 12396 3332 12424
rect 3191 12393 3203 12396
rect 3145 12387 3203 12393
rect 3326 12384 3332 12396
rect 3384 12384 3390 12436
rect 3418 12384 3424 12436
rect 3476 12424 3482 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3476 12396 3801 12424
rect 3476 12384 3482 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 5074 12384 5080 12436
rect 5132 12424 5138 12436
rect 5258 12424 5264 12436
rect 5132 12396 5264 12424
rect 5132 12384 5138 12396
rect 5258 12384 5264 12396
rect 5316 12384 5322 12436
rect 8294 12424 8300 12436
rect 5460 12396 8300 12424
rect 2498 12316 2504 12368
rect 2556 12316 2562 12368
rect 2590 12316 2596 12368
rect 2648 12356 2654 12368
rect 2961 12359 3019 12365
rect 2648 12328 2912 12356
rect 2648 12316 2654 12328
rect 2516 12288 2544 12316
rect 2516 12260 2728 12288
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 1489 12223 1547 12229
rect 1489 12220 1501 12223
rect 1452 12192 1501 12220
rect 1452 12180 1458 12192
rect 1489 12189 1501 12192
rect 1535 12189 1547 12223
rect 1489 12183 1547 12189
rect 2501 12223 2559 12229
rect 2501 12189 2513 12223
rect 2547 12220 2559 12223
rect 2547 12192 2636 12220
rect 2547 12189 2559 12192
rect 2501 12183 2559 12189
rect 2314 12084 2320 12096
rect 2275 12056 2320 12084
rect 2314 12044 2320 12056
rect 2372 12044 2378 12096
rect 2608 12093 2636 12192
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12053 2651 12087
rect 2700 12084 2728 12260
rect 2777 12223 2835 12229
rect 2777 12189 2789 12223
rect 2823 12189 2835 12223
rect 2884 12220 2912 12328
rect 2961 12325 2973 12359
rect 3007 12356 3019 12359
rect 3602 12356 3608 12368
rect 3007 12328 3608 12356
rect 3007 12325 3019 12328
rect 2961 12319 3019 12325
rect 3602 12316 3608 12328
rect 3660 12316 3666 12368
rect 4801 12359 4859 12365
rect 4801 12325 4813 12359
rect 4847 12325 4859 12359
rect 4801 12319 4859 12325
rect 3234 12248 3240 12300
rect 3292 12288 3298 12300
rect 4341 12291 4399 12297
rect 4341 12288 4353 12291
rect 3292 12260 4353 12288
rect 3292 12248 3298 12260
rect 4341 12257 4353 12260
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 4816 12220 4844 12319
rect 5166 12248 5172 12300
rect 5224 12288 5230 12300
rect 5460 12297 5488 12396
rect 8294 12384 8300 12396
rect 8352 12424 8358 12436
rect 8665 12427 8723 12433
rect 8665 12424 8677 12427
rect 8352 12396 8677 12424
rect 8352 12384 8358 12396
rect 8665 12393 8677 12396
rect 8711 12393 8723 12427
rect 10686 12424 10692 12436
rect 10647 12396 10692 12424
rect 8665 12387 8723 12393
rect 10686 12384 10692 12396
rect 10744 12384 10750 12436
rect 10962 12424 10968 12436
rect 10923 12396 10968 12424
rect 10962 12384 10968 12396
rect 11020 12384 11026 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 12492 12396 12633 12424
rect 12492 12384 12498 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 15654 12424 15660 12436
rect 15615 12396 15660 12424
rect 12621 12387 12679 12393
rect 15654 12384 15660 12396
rect 15712 12384 15718 12436
rect 10321 12359 10379 12365
rect 10321 12325 10333 12359
rect 10367 12356 10379 12359
rect 10778 12356 10784 12368
rect 10367 12328 10784 12356
rect 10367 12325 10379 12328
rect 10321 12319 10379 12325
rect 10778 12316 10784 12328
rect 10836 12316 10842 12368
rect 10873 12359 10931 12365
rect 10873 12325 10885 12359
rect 10919 12356 10931 12359
rect 11054 12356 11060 12368
rect 10919 12328 11060 12356
rect 10919 12325 10931 12328
rect 10873 12319 10931 12325
rect 11054 12316 11060 12328
rect 11112 12316 11118 12368
rect 5261 12291 5319 12297
rect 5261 12288 5273 12291
rect 5224 12260 5273 12288
rect 5224 12248 5230 12260
rect 5261 12257 5273 12260
rect 5307 12257 5319 12291
rect 5261 12251 5319 12257
rect 5445 12291 5503 12297
rect 5445 12257 5457 12291
rect 5491 12257 5503 12291
rect 5445 12251 5503 12257
rect 12526 12248 12532 12300
rect 12584 12288 12590 12300
rect 13173 12291 13231 12297
rect 13173 12288 13185 12291
rect 12584 12260 13185 12288
rect 12584 12248 12590 12260
rect 13173 12257 13185 12260
rect 13219 12257 13231 12291
rect 13173 12251 13231 12257
rect 13446 12248 13452 12300
rect 13504 12288 13510 12300
rect 13630 12288 13636 12300
rect 13504 12260 13636 12288
rect 13504 12248 13510 12260
rect 13630 12248 13636 12260
rect 13688 12248 13694 12300
rect 14090 12248 14096 12300
rect 14148 12288 14154 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 14148 12260 14197 12288
rect 14148 12248 14154 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 15105 12291 15163 12297
rect 15105 12257 15117 12291
rect 15151 12288 15163 12291
rect 16022 12288 16028 12300
rect 15151 12260 16028 12288
rect 15151 12257 15163 12260
rect 15105 12251 15163 12257
rect 16022 12248 16028 12260
rect 16080 12248 16086 12300
rect 2884 12192 4844 12220
rect 2777 12183 2835 12189
rect 2792 12152 2820 12183
rect 5534 12180 5540 12232
rect 5592 12220 5598 12232
rect 5629 12223 5687 12229
rect 5629 12220 5641 12223
rect 5592 12192 5641 12220
rect 5592 12180 5598 12192
rect 5629 12189 5641 12192
rect 5675 12189 5687 12223
rect 5810 12220 5816 12232
rect 5771 12192 5816 12220
rect 5629 12183 5687 12189
rect 5810 12180 5816 12192
rect 5868 12220 5874 12232
rect 7285 12223 7343 12229
rect 7285 12220 7297 12223
rect 5868 12192 6745 12220
rect 5868 12180 5874 12192
rect 2866 12152 2872 12164
rect 2792 12124 2872 12152
rect 2866 12112 2872 12124
rect 2924 12112 2930 12164
rect 3329 12155 3387 12161
rect 3329 12121 3341 12155
rect 3375 12152 3387 12155
rect 3510 12152 3516 12164
rect 3375 12124 3516 12152
rect 3375 12121 3387 12124
rect 3329 12115 3387 12121
rect 3510 12112 3516 12124
rect 3568 12112 3574 12164
rect 3605 12155 3663 12161
rect 3605 12121 3617 12155
rect 3651 12152 3663 12155
rect 4062 12152 4068 12164
rect 3651 12124 4068 12152
rect 3651 12121 3663 12124
rect 3605 12115 3663 12121
rect 4062 12112 4068 12124
rect 4120 12112 4126 12164
rect 4157 12155 4215 12161
rect 4157 12121 4169 12155
rect 4203 12152 4215 12155
rect 4982 12152 4988 12164
rect 4203 12124 4988 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 4982 12112 4988 12124
rect 5040 12112 5046 12164
rect 6086 12161 6092 12164
rect 6080 12115 6092 12161
rect 6144 12152 6150 12164
rect 6717 12152 6745 12192
rect 6932 12192 7297 12220
rect 6932 12152 6960 12192
rect 7285 12189 7297 12192
rect 7331 12189 7343 12223
rect 8938 12220 8944 12232
rect 8899 12192 8944 12220
rect 7285 12183 7343 12189
rect 8938 12180 8944 12192
rect 8996 12220 9002 12232
rect 11149 12223 11207 12229
rect 11149 12220 11161 12223
rect 8996 12192 11161 12220
rect 8996 12180 9002 12192
rect 11149 12189 11161 12192
rect 11195 12220 11207 12223
rect 11238 12220 11244 12232
rect 11195 12192 11244 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 12989 12223 13047 12229
rect 12989 12220 13001 12223
rect 12860 12192 13001 12220
rect 12860 12180 12866 12192
rect 12989 12189 13001 12192
rect 13035 12189 13047 12223
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 12989 12183 13047 12189
rect 13372 12192 14473 12220
rect 7530 12155 7588 12161
rect 7530 12152 7542 12155
rect 6144 12124 6180 12152
rect 6717 12124 6960 12152
rect 7208 12124 7542 12152
rect 6086 12112 6092 12115
rect 6144 12112 6150 12124
rect 4249 12087 4307 12093
rect 4249 12084 4261 12087
rect 2700 12056 4261 12084
rect 2593 12047 2651 12053
rect 4249 12053 4261 12056
rect 4295 12084 4307 12087
rect 4614 12084 4620 12096
rect 4295 12056 4620 12084
rect 4295 12053 4307 12056
rect 4249 12047 4307 12053
rect 4614 12044 4620 12056
rect 4672 12044 4678 12096
rect 4709 12087 4767 12093
rect 4709 12053 4721 12087
rect 4755 12084 4767 12087
rect 5074 12084 5080 12096
rect 4755 12056 5080 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 5074 12044 5080 12056
rect 5132 12044 5138 12096
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5442 12084 5448 12096
rect 5215 12056 5448 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5442 12044 5448 12056
rect 5500 12044 5506 12096
rect 6362 12044 6368 12096
rect 6420 12084 6426 12096
rect 6822 12084 6828 12096
rect 6420 12056 6828 12084
rect 6420 12044 6426 12056
rect 6822 12044 6828 12056
rect 6880 12084 6886 12096
rect 7208 12093 7236 12124
rect 7530 12121 7542 12124
rect 7576 12121 7588 12155
rect 7530 12115 7588 12121
rect 9208 12155 9266 12161
rect 9208 12121 9220 12155
rect 9254 12152 9266 12155
rect 9306 12152 9312 12164
rect 9254 12124 9312 12152
rect 9254 12121 9266 12124
rect 9208 12115 9266 12121
rect 9306 12112 9312 12124
rect 9364 12112 9370 12164
rect 10778 12112 10784 12164
rect 10836 12152 10842 12164
rect 11422 12161 11428 12164
rect 11416 12152 11428 12161
rect 10836 12124 11428 12152
rect 10836 12112 10842 12124
rect 11416 12115 11428 12124
rect 11422 12112 11428 12115
rect 11480 12112 11486 12164
rect 13372 12152 13400 12192
rect 14461 12189 14473 12192
rect 14507 12220 14519 12223
rect 14734 12220 14740 12232
rect 14507 12192 14740 12220
rect 14507 12189 14519 12192
rect 14461 12183 14519 12189
rect 14734 12180 14740 12192
rect 14792 12180 14798 12232
rect 15286 12220 15292 12232
rect 15247 12192 15292 12220
rect 15286 12180 15292 12192
rect 15344 12180 15350 12232
rect 12406 12124 13400 12152
rect 7193 12087 7251 12093
rect 7193 12084 7205 12087
rect 6880 12056 7205 12084
rect 6880 12044 6886 12056
rect 7193 12053 7205 12056
rect 7239 12053 7251 12087
rect 7193 12047 7251 12053
rect 8846 12044 8852 12096
rect 8904 12084 8910 12096
rect 12406 12084 12434 12124
rect 13446 12112 13452 12164
rect 13504 12152 13510 12164
rect 13725 12155 13783 12161
rect 13725 12152 13737 12155
rect 13504 12124 13737 12152
rect 13504 12112 13510 12124
rect 13725 12121 13737 12124
rect 13771 12121 13783 12155
rect 13725 12115 13783 12121
rect 15102 12112 15108 12164
rect 15160 12152 15166 12164
rect 15160 12124 15332 12152
rect 15160 12112 15166 12124
rect 15304 12096 15332 12124
rect 12526 12084 12532 12096
rect 8904 12056 12434 12084
rect 12487 12056 12532 12084
rect 8904 12044 8910 12056
rect 12526 12044 12532 12056
rect 12584 12044 12590 12096
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 13081 12087 13139 12093
rect 13081 12084 13093 12087
rect 12676 12056 13093 12084
rect 12676 12044 12682 12056
rect 13081 12053 13093 12056
rect 13127 12053 13139 12087
rect 13081 12047 13139 12053
rect 13170 12044 13176 12096
rect 13228 12084 13234 12096
rect 13633 12087 13691 12093
rect 13633 12084 13645 12087
rect 13228 12056 13645 12084
rect 13228 12044 13234 12056
rect 13633 12053 13645 12056
rect 13679 12053 13691 12087
rect 13633 12047 13691 12053
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 14369 12087 14427 12093
rect 14369 12084 14381 12087
rect 14148 12056 14381 12084
rect 14148 12044 14154 12056
rect 14369 12053 14381 12056
rect 14415 12053 14427 12087
rect 14369 12047 14427 12053
rect 14829 12087 14887 12093
rect 14829 12053 14841 12087
rect 14875 12084 14887 12087
rect 15197 12087 15255 12093
rect 15197 12084 15209 12087
rect 14875 12056 15209 12084
rect 14875 12053 14887 12056
rect 14829 12047 14887 12053
rect 15197 12053 15209 12056
rect 15243 12053 15255 12087
rect 15197 12047 15255 12053
rect 15286 12044 15292 12096
rect 15344 12044 15350 12096
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 3234 11840 3240 11892
rect 3292 11880 3298 11892
rect 3789 11883 3847 11889
rect 3789 11880 3801 11883
rect 3292 11852 3801 11880
rect 3292 11840 3298 11852
rect 3789 11849 3801 11852
rect 3835 11880 3847 11883
rect 4062 11880 4068 11892
rect 3835 11852 4068 11880
rect 3835 11849 3847 11852
rect 3789 11843 3847 11849
rect 4062 11840 4068 11852
rect 4120 11840 4126 11892
rect 4341 11883 4399 11889
rect 4341 11849 4353 11883
rect 4387 11880 4399 11883
rect 4709 11883 4767 11889
rect 4709 11880 4721 11883
rect 4387 11852 4721 11880
rect 4387 11849 4399 11852
rect 4341 11843 4399 11849
rect 4709 11849 4721 11852
rect 4755 11849 4767 11883
rect 5166 11880 5172 11892
rect 5127 11852 5172 11880
rect 4709 11843 4767 11849
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 5994 11880 6000 11892
rect 5955 11852 6000 11880
rect 5994 11840 6000 11852
rect 6052 11840 6058 11892
rect 6454 11840 6460 11892
rect 6512 11880 6518 11892
rect 6917 11883 6975 11889
rect 6917 11880 6929 11883
rect 6512 11852 6929 11880
rect 6512 11840 6518 11852
rect 6917 11849 6929 11852
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 7285 11883 7343 11889
rect 7285 11849 7297 11883
rect 7331 11849 7343 11883
rect 7742 11880 7748 11892
rect 7703 11852 7748 11880
rect 7285 11843 7343 11849
rect 3418 11772 3424 11824
rect 3476 11812 3482 11824
rect 5902 11812 5908 11824
rect 3476 11784 5908 11812
rect 3476 11772 3482 11784
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 6825 11815 6883 11821
rect 6825 11781 6837 11815
rect 6871 11812 6883 11815
rect 7300 11812 7328 11843
rect 7742 11840 7748 11852
rect 7800 11840 7806 11892
rect 9306 11880 9312 11892
rect 9267 11852 9312 11880
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 9674 11840 9680 11892
rect 9732 11880 9738 11892
rect 9861 11883 9919 11889
rect 9861 11880 9873 11883
rect 9732 11852 9873 11880
rect 9732 11840 9738 11852
rect 9861 11849 9873 11852
rect 9907 11849 9919 11883
rect 9861 11843 9919 11849
rect 10134 11840 10140 11892
rect 10192 11880 10198 11892
rect 10321 11883 10379 11889
rect 10321 11880 10333 11883
rect 10192 11852 10333 11880
rect 10192 11840 10198 11852
rect 10321 11849 10333 11852
rect 10367 11849 10379 11883
rect 10321 11843 10379 11849
rect 11517 11883 11575 11889
rect 11517 11849 11529 11883
rect 11563 11880 11575 11883
rect 11882 11880 11888 11892
rect 11563 11852 11888 11880
rect 11563 11849 11575 11852
rect 11517 11843 11575 11849
rect 11882 11840 11888 11852
rect 11940 11840 11946 11892
rect 12897 11883 12955 11889
rect 12897 11880 12909 11883
rect 11992 11852 12909 11880
rect 11330 11812 11336 11824
rect 6871 11784 7328 11812
rect 7392 11784 11336 11812
rect 6871 11781 6883 11784
rect 6825 11775 6883 11781
rect 2521 11747 2579 11753
rect 2521 11713 2533 11747
rect 2567 11744 2579 11747
rect 2777 11747 2835 11753
rect 2567 11716 2728 11744
rect 2567 11713 2579 11716
rect 2521 11707 2579 11713
rect 2700 11676 2728 11716
rect 2777 11713 2789 11747
rect 2823 11744 2835 11747
rect 3142 11744 3148 11756
rect 2823 11716 3148 11744
rect 2823 11713 2835 11716
rect 2777 11707 2835 11713
rect 3142 11704 3148 11716
rect 3200 11704 3206 11756
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3602 11744 3608 11756
rect 3283 11716 3608 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3602 11704 3608 11716
rect 3660 11704 3666 11756
rect 4246 11744 4252 11756
rect 4207 11716 4252 11744
rect 4246 11704 4252 11716
rect 4304 11704 4310 11756
rect 4982 11704 4988 11756
rect 5040 11744 5046 11756
rect 5077 11747 5135 11753
rect 5077 11744 5089 11747
rect 5040 11716 5089 11744
rect 5040 11704 5046 11716
rect 5077 11713 5089 11716
rect 5123 11713 5135 11747
rect 5077 11707 5135 11713
rect 5626 11704 5632 11756
rect 5684 11744 5690 11756
rect 5813 11747 5871 11753
rect 5813 11744 5825 11747
rect 5684 11716 5825 11744
rect 5684 11704 5690 11716
rect 5813 11713 5825 11716
rect 5859 11744 5871 11747
rect 5994 11744 6000 11756
rect 5859 11716 6000 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 6454 11704 6460 11756
rect 6512 11744 6518 11756
rect 7392 11744 7420 11784
rect 6512 11716 7420 11744
rect 7653 11747 7711 11753
rect 6512 11704 6518 11716
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 8113 11747 8171 11753
rect 8113 11744 8125 11747
rect 7699 11716 8125 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 8113 11713 8125 11716
rect 8159 11713 8171 11747
rect 8113 11707 8171 11713
rect 3326 11676 3332 11688
rect 2700 11648 3188 11676
rect 3287 11648 3332 11676
rect 3160 11608 3188 11648
rect 3326 11636 3332 11648
rect 3384 11636 3390 11688
rect 3421 11679 3479 11685
rect 3421 11645 3433 11679
rect 3467 11676 3479 11679
rect 3786 11676 3792 11688
rect 3467 11648 3792 11676
rect 3467 11645 3479 11648
rect 3421 11639 3479 11645
rect 3436 11608 3464 11639
rect 3786 11636 3792 11648
rect 3844 11676 3850 11688
rect 4433 11679 4491 11685
rect 4433 11676 4445 11679
rect 3844 11648 4445 11676
rect 3844 11636 3850 11648
rect 4433 11645 4445 11648
rect 4479 11645 4491 11679
rect 4433 11639 4491 11645
rect 4890 11636 4896 11688
rect 4948 11676 4954 11688
rect 5261 11679 5319 11685
rect 5261 11676 5273 11679
rect 4948 11648 5273 11676
rect 4948 11636 4954 11648
rect 5261 11645 5273 11648
rect 5307 11645 5319 11679
rect 5261 11639 5319 11645
rect 5368 11648 6776 11676
rect 3160 11580 3464 11608
rect 3510 11568 3516 11620
rect 3568 11608 3574 11620
rect 5368 11608 5396 11648
rect 3568 11580 5396 11608
rect 3568 11568 3574 11580
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 6457 11611 6515 11617
rect 6457 11608 6469 11611
rect 5500 11580 6469 11608
rect 5500 11568 5506 11580
rect 6457 11577 6469 11580
rect 6503 11577 6515 11611
rect 6748 11608 6776 11648
rect 6822 11636 6828 11688
rect 6880 11676 6886 11688
rect 7009 11679 7067 11685
rect 7009 11676 7021 11679
rect 6880 11648 7021 11676
rect 6880 11636 6886 11648
rect 7009 11645 7021 11648
rect 7055 11645 7067 11679
rect 7834 11676 7840 11688
rect 7795 11648 7840 11676
rect 7009 11639 7067 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 7374 11608 7380 11620
rect 6748 11580 7380 11608
rect 6457 11571 6515 11577
rect 7374 11568 7380 11580
rect 7432 11568 7438 11620
rect 8220 11608 8248 11784
rect 11330 11772 11336 11784
rect 11388 11772 11394 11824
rect 11992 11812 12020 11852
rect 12897 11849 12909 11852
rect 12943 11880 12955 11883
rect 13170 11880 13176 11892
rect 12943 11852 13176 11880
rect 12943 11849 12955 11852
rect 12897 11843 12955 11849
rect 13170 11840 13176 11852
rect 13228 11840 13234 11892
rect 13354 11840 13360 11892
rect 13412 11880 13418 11892
rect 13541 11883 13599 11889
rect 13541 11880 13553 11883
rect 13412 11852 13553 11880
rect 13412 11840 13418 11852
rect 13541 11849 13553 11852
rect 13587 11849 13599 11883
rect 13541 11843 13599 11849
rect 14001 11883 14059 11889
rect 14001 11849 14013 11883
rect 14047 11880 14059 11883
rect 14090 11880 14096 11892
rect 14047 11852 14096 11880
rect 14047 11849 14059 11852
rect 14001 11843 14059 11849
rect 14090 11840 14096 11852
rect 14148 11840 14154 11892
rect 14185 11883 14243 11889
rect 14185 11849 14197 11883
rect 14231 11880 14243 11883
rect 14458 11880 14464 11892
rect 14231 11852 14464 11880
rect 14231 11849 14243 11852
rect 14185 11843 14243 11849
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 14734 11880 14740 11892
rect 14695 11852 14740 11880
rect 14734 11840 14740 11852
rect 14792 11840 14798 11892
rect 14826 11840 14832 11892
rect 14884 11840 14890 11892
rect 15013 11883 15071 11889
rect 15013 11849 15025 11883
rect 15059 11880 15071 11883
rect 15746 11880 15752 11892
rect 15059 11852 15752 11880
rect 15059 11849 15071 11852
rect 15013 11843 15071 11849
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 12802 11812 12808 11824
rect 11900 11784 12020 11812
rect 12406 11784 12808 11812
rect 11900 11756 11928 11784
rect 8294 11704 8300 11756
rect 8352 11744 8358 11756
rect 8665 11747 8723 11753
rect 8665 11744 8677 11747
rect 8352 11716 8677 11744
rect 8352 11704 8358 11716
rect 8665 11713 8677 11716
rect 8711 11713 8723 11747
rect 8665 11707 8723 11713
rect 10134 11704 10140 11756
rect 10192 11744 10198 11756
rect 10229 11747 10287 11753
rect 10229 11744 10241 11747
rect 10192 11716 10241 11744
rect 10192 11704 10198 11716
rect 10229 11713 10241 11716
rect 10275 11713 10287 11747
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 10229 11707 10287 11713
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 11974 11704 11980 11756
rect 12032 11744 12038 11756
rect 12406 11744 12434 11784
rect 12802 11772 12808 11784
rect 12860 11772 12866 11824
rect 13446 11812 13452 11824
rect 12912 11784 13452 11812
rect 12032 11716 12434 11744
rect 12032 11704 12038 11716
rect 10505 11679 10563 11685
rect 10505 11645 10517 11679
rect 10551 11645 10563 11679
rect 10505 11639 10563 11645
rect 8294 11608 8300 11620
rect 8220 11580 8300 11608
rect 8294 11568 8300 11580
rect 8352 11568 8358 11620
rect 10520 11608 10548 11639
rect 11422 11636 11428 11688
rect 11480 11676 11486 11688
rect 12069 11679 12127 11685
rect 12069 11676 12081 11679
rect 11480 11648 12081 11676
rect 11480 11636 11486 11648
rect 12069 11645 12081 11648
rect 12115 11645 12127 11679
rect 12069 11639 12127 11645
rect 12342 11636 12348 11688
rect 12400 11676 12406 11688
rect 12912 11676 12940 11784
rect 13446 11772 13452 11784
rect 13504 11772 13510 11824
rect 14369 11815 14427 11821
rect 14369 11781 14381 11815
rect 14415 11812 14427 11815
rect 14844 11812 14872 11840
rect 15378 11812 15384 11824
rect 14415 11784 14872 11812
rect 15339 11784 15384 11812
rect 14415 11781 14427 11784
rect 14369 11775 14427 11781
rect 15378 11772 15384 11784
rect 15436 11772 15442 11824
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11744 13875 11747
rect 14642 11744 14648 11756
rect 13863 11716 14648 11744
rect 13863 11713 13875 11716
rect 13817 11707 13875 11713
rect 14642 11704 14648 11716
rect 14700 11704 14706 11756
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11713 14887 11747
rect 15102 11744 15108 11756
rect 15063 11716 15108 11744
rect 14829 11707 14887 11713
rect 12400 11648 12940 11676
rect 12400 11636 12406 11648
rect 13722 11636 13728 11688
rect 13780 11676 13786 11688
rect 14458 11676 14464 11688
rect 13780 11648 14464 11676
rect 13780 11636 13786 11648
rect 14458 11636 14464 11648
rect 14516 11636 14522 11688
rect 14844 11676 14872 11707
rect 15102 11704 15108 11716
rect 15160 11704 15166 11756
rect 15378 11676 15384 11688
rect 14844 11648 15384 11676
rect 15378 11636 15384 11648
rect 15436 11676 15442 11688
rect 16114 11676 16120 11688
rect 15436 11648 16120 11676
rect 15436 11636 15442 11648
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 12526 11608 12532 11620
rect 10520 11580 12532 11608
rect 12526 11568 12532 11580
rect 12584 11568 12590 11620
rect 12986 11608 12992 11620
rect 12899 11580 12992 11608
rect 12986 11568 12992 11580
rect 13044 11608 13050 11620
rect 13044 11580 16160 11608
rect 13044 11568 13050 11580
rect 16132 11552 16160 11580
rect 1394 11540 1400 11552
rect 1355 11512 1400 11540
rect 1394 11500 1400 11512
rect 1452 11500 1458 11552
rect 2406 11500 2412 11552
rect 2464 11540 2470 11552
rect 2869 11543 2927 11549
rect 2869 11540 2881 11543
rect 2464 11512 2881 11540
rect 2464 11500 2470 11512
rect 2869 11509 2881 11512
rect 2915 11509 2927 11543
rect 3878 11540 3884 11552
rect 3839 11512 3884 11540
rect 2869 11503 2927 11509
rect 3878 11500 3884 11512
rect 3936 11500 3942 11552
rect 4338 11500 4344 11552
rect 4396 11540 4402 11552
rect 4982 11540 4988 11552
rect 4396 11512 4988 11540
rect 4396 11500 4402 11512
rect 4982 11500 4988 11512
rect 5040 11540 5046 11552
rect 5258 11540 5264 11552
rect 5040 11512 5264 11540
rect 5040 11500 5046 11512
rect 5258 11500 5264 11512
rect 5316 11540 5322 11552
rect 5537 11543 5595 11549
rect 5537 11540 5549 11543
rect 5316 11512 5549 11540
rect 5316 11500 5322 11512
rect 5537 11509 5549 11512
rect 5583 11509 5595 11543
rect 5537 11503 5595 11509
rect 8386 11500 8392 11552
rect 8444 11540 8450 11552
rect 9493 11543 9551 11549
rect 9493 11540 9505 11543
rect 8444 11512 9505 11540
rect 8444 11500 8450 11512
rect 9493 11509 9505 11512
rect 9539 11540 9551 11543
rect 10962 11540 10968 11552
rect 9539 11512 10968 11540
rect 9539 11509 9551 11512
rect 9493 11503 9551 11509
rect 10962 11500 10968 11512
rect 11020 11500 11026 11552
rect 11606 11500 11612 11552
rect 11664 11540 11670 11552
rect 12342 11540 12348 11552
rect 11664 11512 12348 11540
rect 11664 11500 11670 11512
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 12434 11500 12440 11552
rect 12492 11540 12498 11552
rect 12713 11543 12771 11549
rect 12492 11512 12537 11540
rect 12492 11500 12498 11512
rect 12713 11509 12725 11543
rect 12759 11540 12771 11543
rect 12802 11540 12808 11552
rect 12759 11512 12808 11540
rect 12759 11509 12771 11512
rect 12713 11503 12771 11509
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13078 11500 13084 11552
rect 13136 11540 13142 11552
rect 13265 11543 13323 11549
rect 13265 11540 13277 11543
rect 13136 11512 13277 11540
rect 13136 11500 13142 11512
rect 13265 11509 13277 11512
rect 13311 11540 13323 11543
rect 13354 11540 13360 11552
rect 13311 11512 13360 11540
rect 13311 11509 13323 11512
rect 13265 11503 13323 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 16114 11500 16120 11552
rect 16172 11500 16178 11552
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 2682 11336 2688 11348
rect 2643 11308 2688 11336
rect 2682 11296 2688 11308
rect 2740 11296 2746 11348
rect 3602 11336 3608 11348
rect 3563 11308 3608 11336
rect 3602 11296 3608 11308
rect 3660 11296 3666 11348
rect 3786 11336 3792 11348
rect 3747 11308 3792 11336
rect 3786 11296 3792 11308
rect 3844 11296 3850 11348
rect 4246 11296 4252 11348
rect 4304 11336 4310 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4304 11308 5273 11336
rect 4304 11296 4310 11308
rect 5261 11305 5273 11308
rect 5307 11305 5319 11339
rect 6454 11336 6460 11348
rect 6415 11308 6460 11336
rect 5261 11299 5319 11305
rect 6454 11296 6460 11308
rect 6512 11296 6518 11348
rect 8846 11296 8852 11348
rect 8904 11336 8910 11348
rect 10134 11336 10140 11348
rect 8904 11308 9674 11336
rect 10095 11308 10140 11336
rect 8904 11296 8910 11308
rect 2866 11228 2872 11280
rect 2924 11268 2930 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 2924 11240 3188 11268
rect 2924 11228 2930 11240
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 2041 11203 2099 11209
rect 2041 11200 2053 11203
rect 1452 11172 2053 11200
rect 1452 11160 1458 11172
rect 2041 11169 2053 11172
rect 2087 11169 2099 11203
rect 2041 11163 2099 11169
rect 2225 11203 2283 11209
rect 2225 11169 2237 11203
rect 2271 11200 2283 11203
rect 2406 11200 2412 11212
rect 2271 11172 2412 11200
rect 2271 11169 2283 11172
rect 2225 11163 2283 11169
rect 2406 11160 2412 11172
rect 2464 11160 2470 11212
rect 2774 11160 2780 11212
rect 2832 11200 2838 11212
rect 3160 11209 3188 11240
rect 7208 11240 8953 11268
rect 2961 11203 3019 11209
rect 2961 11200 2973 11203
rect 2832 11172 2973 11200
rect 2832 11160 2838 11172
rect 2961 11169 2973 11172
rect 3007 11169 3019 11203
rect 2961 11163 3019 11169
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 3418 11200 3424 11212
rect 3191 11172 3424 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 5718 11200 5724 11212
rect 5184 11172 5724 11200
rect 1670 11132 1676 11144
rect 1631 11104 1676 11132
rect 1670 11092 1676 11104
rect 1728 11092 1734 11144
rect 2317 11135 2375 11141
rect 2317 11101 2329 11135
rect 2363 11132 2375 11135
rect 2363 11104 3004 11132
rect 2363 11101 2375 11104
rect 2317 11095 2375 11101
rect 2038 11024 2044 11076
rect 2096 11064 2102 11076
rect 2866 11064 2872 11076
rect 2096 11036 2872 11064
rect 2096 11024 2102 11036
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 2976 11064 3004 11104
rect 3050 11092 3056 11144
rect 3108 11132 3114 11144
rect 5184 11141 5212 11172
rect 5718 11160 5724 11172
rect 5776 11160 5782 11212
rect 7208 11209 7236 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 9646 11268 9674 11308
rect 10134 11296 10140 11308
rect 10192 11296 10198 11348
rect 10428 11308 13308 11336
rect 10428 11268 10456 11308
rect 11146 11268 11152 11280
rect 9646 11240 10456 11268
rect 10520 11240 11152 11268
rect 8941 11231 8999 11237
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 7377 11203 7435 11209
rect 7377 11169 7389 11203
rect 7423 11200 7435 11203
rect 7742 11200 7748 11212
rect 7423 11172 7748 11200
rect 7423 11169 7435 11172
rect 7377 11163 7435 11169
rect 5169 11135 5227 11141
rect 5169 11132 5181 11135
rect 3108 11104 5181 11132
rect 3108 11092 3114 11104
rect 5169 11101 5181 11104
rect 5215 11101 5227 11135
rect 5828 11132 5856 11163
rect 7742 11160 7748 11172
rect 7800 11200 7806 11212
rect 8110 11200 8116 11212
rect 7800 11172 8116 11200
rect 7800 11160 7806 11172
rect 8110 11160 8116 11172
rect 8168 11160 8174 11212
rect 8386 11200 8392 11212
rect 8347 11172 8392 11200
rect 8386 11160 8392 11172
rect 8444 11160 8450 11212
rect 8573 11203 8631 11209
rect 8573 11169 8585 11203
rect 8619 11200 8631 11203
rect 9030 11200 9036 11212
rect 8619 11172 9036 11200
rect 8619 11169 8631 11172
rect 8573 11163 8631 11169
rect 9030 11160 9036 11172
rect 9088 11160 9094 11212
rect 9493 11203 9551 11209
rect 9493 11200 9505 11203
rect 9140 11172 9505 11200
rect 5169 11095 5227 11101
rect 5552 11104 5856 11132
rect 3878 11064 3884 11076
rect 2976 11036 3884 11064
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4430 11024 4436 11076
rect 4488 11064 4494 11076
rect 4890 11064 4896 11076
rect 4948 11073 4954 11076
rect 4488 11036 4896 11064
rect 4488 11024 4494 11036
rect 4890 11024 4896 11036
rect 4948 11064 4960 11073
rect 5552 11064 5580 11104
rect 6914 11092 6920 11144
rect 6972 11132 6978 11144
rect 7466 11132 7472 11144
rect 6972 11104 7472 11132
rect 6972 11092 6978 11104
rect 7466 11092 7472 11104
rect 7524 11132 7530 11144
rect 9140 11132 9168 11172
rect 9493 11169 9505 11172
rect 9539 11169 9551 11203
rect 9493 11163 9551 11169
rect 9766 11160 9772 11212
rect 9824 11200 9830 11212
rect 10520 11200 10548 11240
rect 11146 11228 11152 11240
rect 11204 11228 11210 11280
rect 10778 11200 10784 11212
rect 9824 11172 10548 11200
rect 10739 11172 10784 11200
rect 9824 11160 9830 11172
rect 7524 11104 9168 11132
rect 9309 11135 9367 11141
rect 7524 11092 7530 11104
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 10134 11132 10140 11144
rect 9355 11104 10140 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 10134 11092 10140 11104
rect 10192 11092 10198 11144
rect 10520 11141 10548 11172
rect 10778 11160 10784 11172
rect 10836 11160 10842 11212
rect 11238 11160 11244 11212
rect 11296 11200 11302 11212
rect 11296 11172 11744 11200
rect 11296 11160 11302 11172
rect 10505 11135 10563 11141
rect 10505 11101 10517 11135
rect 10551 11101 10563 11135
rect 10505 11095 10563 11101
rect 10597 11135 10655 11141
rect 10597 11101 10609 11135
rect 10643 11132 10655 11135
rect 10870 11132 10876 11144
rect 10643 11104 10876 11132
rect 10643 11101 10655 11104
rect 10597 11095 10655 11101
rect 10870 11092 10876 11104
rect 10928 11132 10934 11144
rect 11422 11132 11428 11144
rect 10928 11104 11428 11132
rect 10928 11092 10934 11104
rect 11422 11092 11428 11104
rect 11480 11092 11486 11144
rect 11606 11132 11612 11144
rect 11567 11104 11612 11132
rect 11606 11092 11612 11104
rect 11664 11092 11670 11144
rect 11716 11141 11744 11172
rect 11701 11135 11759 11141
rect 11701 11101 11713 11135
rect 11747 11132 11759 11135
rect 12894 11132 12900 11144
rect 11747 11104 12900 11132
rect 11747 11101 11759 11104
rect 11701 11095 11759 11101
rect 12894 11092 12900 11104
rect 12952 11092 12958 11144
rect 13280 11132 13308 11308
rect 13538 11296 13544 11348
rect 13596 11336 13602 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 13596 11308 13645 11336
rect 13596 11296 13602 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 15197 11339 15255 11345
rect 15197 11305 15209 11339
rect 15243 11336 15255 11339
rect 15378 11336 15384 11348
rect 15243 11308 15384 11336
rect 15243 11305 15255 11308
rect 15197 11299 15255 11305
rect 15378 11296 15384 11308
rect 15436 11296 15442 11348
rect 15470 11296 15476 11348
rect 15528 11345 15534 11348
rect 15528 11339 15577 11345
rect 15528 11305 15531 11339
rect 15565 11305 15577 11339
rect 15528 11299 15577 11305
rect 15528 11296 15534 11299
rect 13909 11271 13967 11277
rect 13909 11237 13921 11271
rect 13955 11268 13967 11271
rect 15930 11268 15936 11280
rect 13955 11240 15936 11268
rect 13955 11237 13967 11240
rect 13909 11231 13967 11237
rect 15930 11228 15936 11240
rect 15988 11228 15994 11280
rect 13446 11200 13452 11212
rect 13359 11172 13452 11200
rect 13446 11160 13452 11172
rect 13504 11200 13510 11212
rect 13630 11200 13636 11212
rect 13504 11172 13636 11200
rect 13504 11160 13510 11172
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13814 11160 13820 11212
rect 13872 11200 13878 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 13872 11172 14197 11200
rect 13872 11160 13878 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14550 11200 14556 11212
rect 14185 11163 14243 11169
rect 14384 11172 14556 11200
rect 14384 11141 14412 11172
rect 14550 11160 14556 11172
rect 14608 11200 14614 11212
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 14608 11172 15301 11200
rect 14608 11160 14614 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 14369 11135 14427 11141
rect 14369 11132 14381 11135
rect 13280 11104 14381 11132
rect 14369 11101 14381 11104
rect 14415 11101 14427 11135
rect 14369 11095 14427 11101
rect 15194 11092 15200 11144
rect 15252 11132 15258 11144
rect 15590 11135 15648 11141
rect 15590 11132 15602 11135
rect 15252 11104 15602 11132
rect 15252 11092 15258 11104
rect 15590 11101 15602 11104
rect 15636 11101 15648 11135
rect 15590 11095 15648 11101
rect 4948 11036 5580 11064
rect 5629 11067 5687 11073
rect 4948 11027 4960 11036
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 6089 11067 6147 11073
rect 6089 11064 6101 11067
rect 5675 11036 6101 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 6089 11033 6101 11036
rect 6135 11033 6147 11067
rect 6454 11064 6460 11076
rect 6089 11027 6147 11033
rect 6196 11036 6460 11064
rect 4948 11024 4954 11027
rect 1486 10996 1492 11008
rect 1447 10968 1492 10996
rect 1486 10956 1492 10968
rect 1544 10956 1550 11008
rect 3234 10956 3240 11008
rect 3292 10996 3298 11008
rect 5718 10996 5724 11008
rect 3292 10968 3337 10996
rect 5631 10968 5724 10996
rect 3292 10956 3298 10968
rect 5718 10956 5724 10968
rect 5776 10996 5782 11008
rect 6196 10996 6224 11036
rect 6454 11024 6460 11036
rect 6512 11024 6518 11076
rect 7098 11064 7104 11076
rect 7059 11036 7104 11064
rect 7098 11024 7104 11036
rect 7156 11024 7162 11076
rect 8297 11067 8355 11073
rect 8297 11033 8309 11067
rect 8343 11064 8355 11067
rect 9769 11067 9827 11073
rect 9769 11064 9781 11067
rect 8343 11036 9781 11064
rect 8343 11033 8355 11036
rect 8297 11027 8355 11033
rect 9769 11033 9781 11036
rect 9815 11033 9827 11067
rect 9769 11027 9827 11033
rect 10965 11067 11023 11073
rect 10965 11033 10977 11067
rect 11011 11064 11023 11067
rect 11946 11067 12004 11073
rect 11946 11064 11958 11067
rect 11011 11036 11958 11064
rect 11011 11033 11023 11036
rect 10965 11027 11023 11033
rect 11946 11033 11958 11036
rect 11992 11033 12004 11067
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 11946 11027 12004 11033
rect 12406 11036 14473 11064
rect 6730 10996 6736 11008
rect 5776 10968 6224 10996
rect 6691 10968 6736 10996
rect 5776 10956 5782 10968
rect 6730 10956 6736 10968
rect 6788 10956 6794 11008
rect 7926 10996 7932 11008
rect 7887 10968 7932 10996
rect 7926 10956 7932 10968
rect 7984 10956 7990 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 9456 10968 9501 10996
rect 9456 10956 9462 10968
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 12406 10996 12434 11036
rect 14461 11033 14473 11036
rect 14507 11064 14519 11067
rect 15013 11067 15071 11073
rect 15013 11064 15025 11067
rect 14507 11036 15025 11064
rect 14507 11033 14519 11036
rect 14461 11027 14519 11033
rect 15013 11033 15025 11036
rect 15059 11064 15071 11067
rect 15378 11064 15384 11076
rect 15059 11036 15384 11064
rect 15059 11033 15071 11036
rect 15013 11027 15071 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 9640 10968 12434 10996
rect 9640 10956 9646 10968
rect 12894 10956 12900 11008
rect 12952 10996 12958 11008
rect 13081 10999 13139 11005
rect 13081 10996 13093 10999
rect 12952 10968 13093 10996
rect 12952 10956 12958 10968
rect 13081 10965 13093 10968
rect 13127 10965 13139 10999
rect 13081 10959 13139 10965
rect 13170 10956 13176 11008
rect 13228 10996 13234 11008
rect 13228 10968 13273 10996
rect 13228 10956 13234 10968
rect 14550 10956 14556 11008
rect 14608 10996 14614 11008
rect 14829 10999 14887 11005
rect 14829 10996 14841 10999
rect 14608 10968 14841 10996
rect 14608 10956 14614 10968
rect 14829 10965 14841 10968
rect 14875 10965 14887 10999
rect 14829 10959 14887 10965
rect 15286 10956 15292 11008
rect 15344 10996 15350 11008
rect 16482 10996 16488 11008
rect 15344 10968 16488 10996
rect 15344 10956 15350 10968
rect 16482 10956 16488 10968
rect 16540 10956 16546 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 1489 10795 1547 10801
rect 1489 10761 1501 10795
rect 1535 10792 1547 10795
rect 1670 10792 1676 10804
rect 1535 10764 1676 10792
rect 1535 10761 1547 10764
rect 1489 10755 1547 10761
rect 1670 10752 1676 10764
rect 1728 10752 1734 10804
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 3142 10792 3148 10804
rect 3099 10764 3148 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 6730 10792 6736 10804
rect 4172 10764 6736 10792
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 4172 10656 4200 10764
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 7742 10792 7748 10804
rect 7703 10764 7748 10792
rect 7742 10752 7748 10764
rect 7800 10752 7806 10804
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11664 10764 11713 10792
rect 11664 10752 11670 10764
rect 11701 10761 11713 10764
rect 11747 10792 11759 10795
rect 12618 10792 12624 10804
rect 11747 10764 12624 10792
rect 11747 10761 11759 10764
rect 11701 10755 11759 10761
rect 12618 10752 12624 10764
rect 12676 10752 12682 10804
rect 14826 10752 14832 10804
rect 14884 10792 14890 10804
rect 15010 10792 15016 10804
rect 14884 10764 15016 10792
rect 14884 10752 14890 10764
rect 15010 10752 15016 10764
rect 15068 10752 15074 10804
rect 4338 10724 4344 10736
rect 4251 10696 4344 10724
rect 4338 10684 4344 10696
rect 4396 10724 4402 10736
rect 9677 10727 9735 10733
rect 4396 10696 7052 10724
rect 4396 10684 4402 10696
rect 7024 10668 7052 10696
rect 9677 10693 9689 10727
rect 9723 10724 9735 10727
rect 13262 10724 13268 10736
rect 9723 10696 13268 10724
rect 9723 10693 9735 10696
rect 9677 10687 9735 10693
rect 13262 10684 13268 10696
rect 13320 10684 13326 10736
rect 13832 10696 15148 10724
rect 13832 10668 13860 10696
rect 5534 10656 5540 10668
rect 5592 10665 5598 10668
rect 1719 10628 4200 10656
rect 5504 10628 5540 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 5534 10616 5540 10628
rect 5592 10619 5604 10665
rect 5810 10656 5816 10668
rect 5771 10628 5816 10656
rect 5592 10616 5598 10619
rect 5810 10616 5816 10628
rect 5868 10656 5874 10668
rect 6365 10659 6423 10665
rect 6365 10656 6377 10659
rect 5868 10628 6377 10656
rect 5868 10616 5874 10628
rect 6365 10625 6377 10628
rect 6411 10625 6423 10659
rect 6365 10619 6423 10625
rect 6632 10659 6690 10665
rect 6632 10625 6644 10659
rect 6678 10656 6690 10659
rect 6914 10656 6920 10668
rect 6678 10628 6920 10656
rect 6678 10625 6690 10628
rect 6632 10619 6690 10625
rect 6914 10616 6920 10628
rect 6972 10616 6978 10668
rect 7006 10616 7012 10668
rect 7064 10656 7070 10668
rect 7064 10628 8432 10656
rect 7064 10616 7070 10628
rect 5994 10548 6000 10600
rect 6052 10588 6058 10600
rect 6089 10591 6147 10597
rect 6089 10588 6101 10591
rect 6052 10560 6101 10588
rect 6052 10548 6058 10560
rect 6089 10557 6101 10560
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 2774 10480 2780 10532
rect 2832 10520 2838 10532
rect 4430 10520 4436 10532
rect 2832 10492 4436 10520
rect 2832 10480 2838 10492
rect 4430 10480 4436 10492
rect 4488 10480 4494 10532
rect 8404 10529 8432 10628
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 11066 10659 11124 10665
rect 11066 10656 11078 10659
rect 10836 10628 11078 10656
rect 10836 10616 10842 10628
rect 11066 10625 11078 10628
rect 11112 10625 11124 10659
rect 11066 10619 11124 10625
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11333 10659 11391 10665
rect 11333 10656 11345 10659
rect 11296 10628 11345 10656
rect 11296 10616 11302 10628
rect 11333 10625 11345 10628
rect 11379 10625 11391 10659
rect 11333 10619 11391 10625
rect 12825 10659 12883 10665
rect 12825 10625 12837 10659
rect 12871 10656 12883 10659
rect 12986 10656 12992 10668
rect 12871 10628 12992 10656
rect 12871 10625 12883 10628
rect 12825 10619 12883 10625
rect 12986 10616 12992 10628
rect 13044 10616 13050 10668
rect 13078 10616 13084 10668
rect 13136 10656 13142 10668
rect 13173 10659 13231 10665
rect 13173 10656 13185 10659
rect 13136 10628 13185 10656
rect 13136 10616 13142 10628
rect 13173 10625 13185 10628
rect 13219 10625 13231 10659
rect 13173 10619 13231 10625
rect 13440 10659 13498 10665
rect 13440 10625 13452 10659
rect 13486 10656 13498 10659
rect 13814 10656 13820 10668
rect 13486 10628 13820 10656
rect 13486 10625 13498 10628
rect 13440 10619 13498 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 15010 10656 15016 10668
rect 14971 10628 15016 10656
rect 15010 10616 15016 10628
rect 15068 10616 15074 10668
rect 15120 10656 15148 10696
rect 15120 10628 15240 10656
rect 14826 10548 14832 10600
rect 14884 10588 14890 10600
rect 15212 10597 15240 10628
rect 15105 10591 15163 10597
rect 15105 10588 15117 10591
rect 14884 10560 15117 10588
rect 14884 10548 14890 10560
rect 15105 10557 15117 10560
rect 15151 10557 15163 10591
rect 15105 10551 15163 10557
rect 15197 10591 15255 10597
rect 15197 10557 15209 10591
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 8389 10523 8447 10529
rect 8389 10489 8401 10523
rect 8435 10520 8447 10523
rect 10226 10520 10232 10532
rect 8435 10492 10232 10520
rect 8435 10489 8447 10492
rect 8389 10483 8447 10489
rect 10226 10480 10232 10492
rect 10284 10480 10290 10532
rect 14458 10480 14464 10532
rect 14516 10520 14522 10532
rect 14645 10523 14703 10529
rect 14645 10520 14657 10523
rect 14516 10492 14657 10520
rect 14516 10480 14522 10492
rect 14645 10489 14657 10492
rect 14691 10489 14703 10523
rect 15120 10520 15148 10551
rect 15473 10523 15531 10529
rect 15473 10520 15485 10523
rect 15120 10492 15485 10520
rect 14645 10483 14703 10489
rect 15473 10489 15485 10492
rect 15519 10489 15531 10523
rect 15473 10483 15531 10489
rect 5442 10412 5448 10464
rect 5500 10452 5506 10464
rect 5905 10455 5963 10461
rect 5905 10452 5917 10455
rect 5500 10424 5917 10452
rect 5500 10412 5506 10424
rect 5905 10421 5917 10424
rect 5951 10421 5963 10455
rect 9950 10452 9956 10464
rect 9911 10424 9956 10452
rect 5905 10415 5963 10421
rect 9950 10412 9956 10424
rect 10008 10412 10014 10464
rect 14553 10455 14611 10461
rect 14553 10421 14565 10455
rect 14599 10452 14611 10455
rect 14734 10452 14740 10464
rect 14599 10424 14740 10452
rect 14599 10421 14611 10424
rect 14553 10415 14611 10421
rect 14734 10412 14740 10424
rect 14792 10412 14798 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 3237 10251 3295 10257
rect 3237 10217 3249 10251
rect 3283 10248 3295 10251
rect 3326 10248 3332 10260
rect 3283 10220 3332 10248
rect 3283 10217 3295 10220
rect 3237 10211 3295 10217
rect 3326 10208 3332 10220
rect 3384 10208 3390 10260
rect 3605 10251 3663 10257
rect 3605 10217 3617 10251
rect 3651 10248 3663 10251
rect 3694 10248 3700 10260
rect 3651 10220 3700 10248
rect 3651 10217 3663 10220
rect 3605 10211 3663 10217
rect 3694 10208 3700 10220
rect 3752 10248 3758 10260
rect 4062 10248 4068 10260
rect 3752 10220 4068 10248
rect 3752 10208 3758 10220
rect 4062 10208 4068 10220
rect 4120 10208 4126 10260
rect 5534 10208 5540 10260
rect 5592 10248 5598 10260
rect 5629 10251 5687 10257
rect 5629 10248 5641 10251
rect 5592 10220 5641 10248
rect 5592 10208 5598 10220
rect 5629 10217 5641 10220
rect 5675 10217 5687 10251
rect 5629 10211 5687 10217
rect 7285 10251 7343 10257
rect 7285 10217 7297 10251
rect 7331 10248 7343 10251
rect 7331 10220 9352 10248
rect 7331 10217 7343 10220
rect 7285 10211 7343 10217
rect 7377 10183 7435 10189
rect 2884 10152 6132 10180
rect 2682 10112 2688 10124
rect 2643 10084 2688 10112
rect 2682 10072 2688 10084
rect 2740 10072 2746 10124
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10044 1731 10047
rect 1946 10044 1952 10056
rect 1719 10016 1808 10044
rect 1907 10016 1952 10044
rect 1719 10013 1731 10016
rect 1673 10007 1731 10013
rect 1486 9908 1492 9920
rect 1447 9880 1492 9908
rect 1486 9868 1492 9880
rect 1544 9868 1550 9920
rect 1780 9917 1808 10016
rect 1946 10004 1952 10016
rect 2004 10004 2010 10056
rect 2406 10044 2412 10056
rect 2367 10016 2412 10044
rect 2406 10004 2412 10016
rect 2464 10004 2470 10056
rect 2884 10053 2912 10152
rect 3694 10072 3700 10124
rect 3752 10112 3758 10124
rect 4246 10112 4252 10124
rect 3752 10084 4252 10112
rect 3752 10072 3758 10084
rect 4246 10072 4252 10084
rect 4304 10072 4310 10124
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10081 4491 10115
rect 4433 10075 4491 10081
rect 2869 10047 2927 10053
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 4154 10044 4160 10056
rect 4115 10016 4160 10044
rect 2869 10007 2927 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 4448 10044 4476 10075
rect 4522 10072 4528 10124
rect 4580 10112 4586 10124
rect 5258 10112 5264 10124
rect 4580 10084 5264 10112
rect 4580 10072 4586 10084
rect 5258 10072 5264 10084
rect 5316 10072 5322 10124
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4448 10016 4997 10044
rect 4985 10013 4997 10016
rect 5031 10044 5043 10047
rect 5031 10016 5764 10044
rect 5031 10013 5043 10016
rect 4985 10007 5043 10013
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 4249 9979 4307 9985
rect 2823 9948 3832 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 1765 9911 1823 9917
rect 1765 9877 1777 9911
rect 1811 9877 1823 9911
rect 1765 9871 1823 9877
rect 1854 9868 1860 9920
rect 1912 9908 1918 9920
rect 2041 9911 2099 9917
rect 2041 9908 2053 9911
rect 1912 9880 2053 9908
rect 1912 9868 1918 9880
rect 2041 9877 2053 9880
rect 2087 9877 2099 9911
rect 3326 9908 3332 9920
rect 3287 9880 3332 9908
rect 2041 9871 2099 9877
rect 3326 9868 3332 9880
rect 3384 9868 3390 9920
rect 3804 9917 3832 9948
rect 4249 9945 4261 9979
rect 4295 9976 4307 9979
rect 4522 9976 4528 9988
rect 4295 9948 4528 9976
rect 4295 9945 4307 9948
rect 4249 9939 4307 9945
rect 4522 9936 4528 9948
rect 4580 9936 4586 9988
rect 5442 9976 5448 9988
rect 4632 9948 5448 9976
rect 3789 9911 3847 9917
rect 3789 9877 3801 9911
rect 3835 9877 3847 9911
rect 3789 9871 3847 9877
rect 4430 9868 4436 9920
rect 4488 9908 4494 9920
rect 4632 9917 4660 9948
rect 5442 9936 5448 9948
rect 5500 9936 5506 9988
rect 4617 9911 4675 9917
rect 4617 9908 4629 9911
rect 4488 9880 4629 9908
rect 4488 9868 4494 9880
rect 4617 9877 4629 9880
rect 4663 9877 4675 9911
rect 4617 9871 4675 9877
rect 4893 9911 4951 9917
rect 4893 9877 4905 9911
rect 4939 9908 4951 9911
rect 5166 9908 5172 9920
rect 4939 9880 5172 9908
rect 4939 9877 4951 9880
rect 4893 9871 4951 9877
rect 5166 9868 5172 9880
rect 5224 9908 5230 9920
rect 5534 9908 5540 9920
rect 5224 9880 5540 9908
rect 5224 9868 5230 9880
rect 5534 9868 5540 9880
rect 5592 9868 5598 9920
rect 5736 9917 5764 10016
rect 5721 9911 5779 9917
rect 5721 9877 5733 9911
rect 5767 9877 5779 9911
rect 6104 9908 6132 10152
rect 7377 10149 7389 10183
rect 7423 10180 7435 10183
rect 7466 10180 7472 10192
rect 7423 10152 7472 10180
rect 7423 10149 7435 10152
rect 7377 10143 7435 10149
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 9324 10180 9352 10220
rect 9398 10208 9404 10260
rect 9456 10248 9462 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 9456 10220 9505 10248
rect 9456 10208 9462 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 11238 10208 11244 10260
rect 11296 10248 11302 10260
rect 11701 10251 11759 10257
rect 11701 10248 11713 10251
rect 11296 10220 11713 10248
rect 11296 10208 11302 10220
rect 11701 10217 11713 10220
rect 11747 10217 11759 10251
rect 12526 10248 12532 10260
rect 11701 10211 11759 10217
rect 12406 10220 12532 10248
rect 12406 10180 12434 10220
rect 12526 10208 12532 10220
rect 12584 10208 12590 10260
rect 14734 10180 14740 10192
rect 9324 10152 12434 10180
rect 13648 10152 14740 10180
rect 8757 10115 8815 10121
rect 8757 10081 8769 10115
rect 8803 10112 8815 10115
rect 8938 10112 8944 10124
rect 8803 10084 8944 10112
rect 8803 10081 8815 10084
rect 8757 10075 8815 10081
rect 8938 10072 8944 10084
rect 8996 10072 9002 10124
rect 9030 10072 9036 10124
rect 9088 10112 9094 10124
rect 9950 10112 9956 10124
rect 9088 10084 9956 10112
rect 9088 10072 9094 10084
rect 9950 10072 9956 10084
rect 10008 10112 10014 10124
rect 10137 10115 10195 10121
rect 10137 10112 10149 10115
rect 10008 10084 10149 10112
rect 10008 10072 10014 10084
rect 10137 10081 10149 10084
rect 10183 10112 10195 10115
rect 10870 10112 10876 10124
rect 10183 10084 10876 10112
rect 10183 10081 10195 10084
rect 10137 10075 10195 10081
rect 10870 10072 10876 10084
rect 10928 10072 10934 10124
rect 12066 10072 12072 10124
rect 12124 10112 12130 10124
rect 12805 10115 12863 10121
rect 12805 10112 12817 10115
rect 12124 10084 12817 10112
rect 12124 10072 12130 10084
rect 12805 10081 12817 10084
rect 12851 10112 12863 10115
rect 12894 10112 12900 10124
rect 12851 10084 12900 10112
rect 12851 10081 12863 10084
rect 12805 10075 12863 10081
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 12986 10072 12992 10124
rect 13044 10112 13050 10124
rect 13648 10121 13676 10152
rect 13633 10115 13691 10121
rect 13633 10112 13645 10115
rect 13044 10084 13645 10112
rect 13044 10072 13050 10084
rect 13633 10081 13645 10084
rect 13679 10081 13691 10115
rect 14550 10112 14556 10124
rect 14511 10084 14556 10112
rect 13633 10075 13691 10081
rect 14550 10072 14556 10084
rect 14608 10072 14614 10124
rect 14660 10121 14688 10152
rect 14734 10140 14740 10152
rect 14792 10140 14798 10192
rect 14645 10115 14703 10121
rect 14645 10081 14657 10115
rect 14691 10081 14703 10115
rect 14645 10075 14703 10081
rect 15010 10072 15016 10124
rect 15068 10112 15074 10124
rect 15105 10115 15163 10121
rect 15105 10112 15117 10115
rect 15068 10084 15117 10112
rect 15068 10072 15074 10084
rect 15105 10081 15117 10084
rect 15151 10081 15163 10115
rect 15105 10075 15163 10081
rect 6454 10004 6460 10056
rect 6512 10044 6518 10056
rect 7101 10047 7159 10053
rect 7101 10044 7113 10047
rect 6512 10016 7113 10044
rect 6512 10004 6518 10016
rect 7101 10013 7113 10016
rect 7147 10013 7159 10047
rect 7101 10007 7159 10013
rect 8501 10047 8559 10053
rect 8501 10013 8513 10047
rect 8547 10044 8559 10047
rect 9048 10044 9076 10072
rect 8547 10016 9076 10044
rect 9861 10047 9919 10053
rect 8547 10013 8559 10016
rect 8501 10007 8559 10013
rect 9861 10013 9873 10047
rect 9907 10044 9919 10047
rect 11514 10044 11520 10056
rect 9907 10016 11520 10044
rect 9907 10013 9919 10016
rect 9861 10007 9919 10013
rect 11514 10004 11520 10016
rect 11572 10004 11578 10056
rect 12621 10047 12679 10053
rect 12621 10044 12633 10047
rect 12406 10016 12633 10044
rect 6856 9979 6914 9985
rect 6856 9945 6868 9979
rect 6902 9976 6914 9979
rect 9122 9976 9128 9988
rect 6902 9948 9128 9976
rect 6902 9945 6914 9948
rect 6856 9939 6914 9945
rect 9122 9936 9128 9948
rect 9180 9936 9186 9988
rect 9398 9936 9404 9988
rect 9456 9976 9462 9988
rect 9456 9948 10180 9976
rect 9456 9936 9462 9948
rect 7190 9908 7196 9920
rect 6104 9880 7196 9908
rect 5721 9871 5779 9877
rect 7190 9868 7196 9880
rect 7248 9908 7254 9920
rect 8202 9908 8208 9920
rect 7248 9880 8208 9908
rect 7248 9868 7254 9880
rect 8202 9868 8208 9880
rect 8260 9868 8266 9920
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10152 9908 10180 9948
rect 10226 9936 10232 9988
rect 10284 9976 10290 9988
rect 10413 9979 10471 9985
rect 10413 9976 10425 9979
rect 10284 9948 10425 9976
rect 10284 9936 10290 9948
rect 10413 9945 10425 9948
rect 10459 9945 10471 9979
rect 12406 9976 12434 10016
rect 12621 10013 12633 10016
rect 12667 10044 12679 10047
rect 13446 10044 13452 10056
rect 12667 10016 13452 10044
rect 12667 10013 12679 10016
rect 12621 10007 12679 10013
rect 13446 10004 13452 10016
rect 13504 10004 13510 10056
rect 14458 10044 14464 10056
rect 14419 10016 14464 10044
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 15194 10004 15200 10056
rect 15252 10044 15258 10056
rect 15381 10047 15439 10053
rect 15381 10044 15393 10047
rect 15252 10016 15393 10044
rect 15252 10004 15258 10016
rect 15381 10013 15393 10016
rect 15427 10013 15439 10047
rect 15381 10007 15439 10013
rect 10413 9939 10471 9945
rect 10520 9948 12434 9976
rect 12713 9979 12771 9985
rect 10520 9908 10548 9948
rect 12713 9945 12725 9979
rect 12759 9976 12771 9979
rect 13262 9976 13268 9988
rect 12759 9948 13268 9976
rect 12759 9945 12771 9948
rect 12713 9939 12771 9945
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 10008 9880 10053 9908
rect 10152 9880 10548 9908
rect 10008 9868 10014 9880
rect 11054 9868 11060 9920
rect 11112 9908 11118 9920
rect 12253 9911 12311 9917
rect 12253 9908 12265 9911
rect 11112 9880 12265 9908
rect 11112 9868 11118 9880
rect 12253 9877 12265 9880
rect 12299 9877 12311 9911
rect 13078 9908 13084 9920
rect 13039 9880 13084 9908
rect 12253 9871 12311 9877
rect 13078 9868 13084 9880
rect 13136 9868 13142 9920
rect 13446 9908 13452 9920
rect 13407 9880 13452 9908
rect 13446 9868 13452 9880
rect 13504 9868 13510 9920
rect 13538 9868 13544 9920
rect 13596 9908 13602 9920
rect 14090 9908 14096 9920
rect 13596 9880 13641 9908
rect 14051 9880 14096 9908
rect 13596 9868 13602 9880
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 15562 9908 15568 9920
rect 15523 9880 15568 9908
rect 15562 9868 15568 9880
rect 15620 9868 15626 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 1394 9664 1400 9716
rect 1452 9704 1458 9716
rect 4154 9704 4160 9716
rect 1452 9676 4160 9704
rect 1452 9664 1458 9676
rect 4154 9664 4160 9676
rect 4212 9664 4218 9716
rect 4341 9707 4399 9713
rect 4341 9673 4353 9707
rect 4387 9704 4399 9707
rect 4387 9676 4568 9704
rect 4387 9673 4399 9676
rect 4341 9667 4399 9673
rect 2498 9596 2504 9648
rect 2556 9636 2562 9648
rect 2777 9639 2835 9645
rect 2777 9636 2789 9639
rect 2556 9608 2789 9636
rect 2556 9596 2562 9608
rect 2777 9605 2789 9608
rect 2823 9605 2835 9639
rect 4540 9636 4568 9676
rect 5258 9664 5264 9716
rect 5316 9704 5322 9716
rect 9398 9704 9404 9716
rect 5316 9676 5580 9704
rect 5316 9664 5322 9676
rect 5442 9636 5448 9648
rect 2777 9599 2835 9605
rect 3160 9608 4476 9636
rect 4540 9608 5448 9636
rect 3160 9580 3188 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 1762 9568 1768 9580
rect 1719 9540 1768 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 1762 9528 1768 9540
rect 1820 9528 1826 9580
rect 1949 9571 2007 9577
rect 1949 9537 1961 9571
rect 1995 9537 2007 9571
rect 1949 9531 2007 9537
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2406 9568 2412 9580
rect 2271 9540 2412 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 1964 9500 1992 9531
rect 2406 9528 2412 9540
rect 2464 9528 2470 9580
rect 3142 9568 3148 9580
rect 3055 9540 3148 9568
rect 3142 9528 3148 9540
rect 3200 9528 3206 9580
rect 4154 9528 4160 9580
rect 4212 9568 4218 9580
rect 4249 9571 4307 9577
rect 4249 9568 4261 9571
rect 4212 9540 4261 9568
rect 4212 9528 4218 9540
rect 4249 9537 4261 9540
rect 4295 9537 4307 9571
rect 4249 9531 4307 9537
rect 2498 9500 2504 9512
rect 1964 9472 2504 9500
rect 2498 9460 2504 9472
rect 2556 9460 2562 9512
rect 3053 9503 3111 9509
rect 3053 9469 3065 9503
rect 3099 9500 3111 9503
rect 3970 9500 3976 9512
rect 3099 9472 3976 9500
rect 3099 9469 3111 9472
rect 3053 9463 3111 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4448 9509 4476 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 5552 9636 5580 9676
rect 6012 9676 9404 9704
rect 5905 9639 5963 9645
rect 5905 9636 5917 9639
rect 5552 9608 5917 9636
rect 5905 9605 5917 9608
rect 5951 9605 5963 9639
rect 5905 9599 5963 9605
rect 4522 9528 4528 9580
rect 4580 9568 4586 9580
rect 4982 9568 4988 9580
rect 4580 9540 4988 9568
rect 4580 9528 4586 9540
rect 4982 9528 4988 9540
rect 5040 9568 5046 9580
rect 5169 9571 5227 9577
rect 5169 9568 5181 9571
rect 5040 9540 5181 9568
rect 5040 9528 5046 9540
rect 5169 9537 5181 9540
rect 5215 9537 5227 9571
rect 5169 9531 5227 9537
rect 5261 9571 5319 9577
rect 5261 9537 5273 9571
rect 5307 9568 5319 9571
rect 5534 9568 5540 9580
rect 5307 9540 5540 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5534 9528 5540 9540
rect 5592 9568 5598 9580
rect 6012 9568 6040 9676
rect 9398 9664 9404 9676
rect 9456 9664 9462 9716
rect 9858 9704 9864 9716
rect 9819 9676 9864 9704
rect 9858 9664 9864 9676
rect 9916 9664 9922 9716
rect 9950 9664 9956 9716
rect 10008 9704 10014 9716
rect 10229 9707 10287 9713
rect 10229 9704 10241 9707
rect 10008 9676 10241 9704
rect 10008 9664 10014 9676
rect 10229 9673 10241 9676
rect 10275 9673 10287 9707
rect 10229 9667 10287 9673
rect 10321 9707 10379 9713
rect 10321 9673 10333 9707
rect 10367 9673 10379 9707
rect 11514 9704 11520 9716
rect 11475 9676 11520 9704
rect 10321 9667 10379 9673
rect 6733 9639 6791 9645
rect 6733 9605 6745 9639
rect 6779 9636 6791 9639
rect 7926 9636 7932 9648
rect 6779 9608 7932 9636
rect 6779 9605 6791 9608
rect 6733 9599 6791 9605
rect 7926 9596 7932 9608
rect 7984 9596 7990 9648
rect 8389 9639 8447 9645
rect 8389 9605 8401 9639
rect 8435 9636 8447 9639
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8435 9608 8953 9636
rect 8435 9605 8447 9608
rect 8389 9599 8447 9605
rect 8941 9605 8953 9608
rect 8987 9636 8999 9639
rect 9122 9636 9128 9648
rect 8987 9608 9128 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 9769 9639 9827 9645
rect 9769 9605 9781 9639
rect 9815 9636 9827 9639
rect 10042 9636 10048 9648
rect 9815 9608 10048 9636
rect 9815 9605 9827 9608
rect 9769 9599 9827 9605
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10134 9596 10140 9648
rect 10192 9636 10198 9648
rect 10336 9636 10364 9667
rect 11514 9664 11520 9676
rect 11572 9664 11578 9716
rect 12805 9707 12863 9713
rect 12805 9673 12817 9707
rect 12851 9704 12863 9707
rect 13078 9704 13084 9716
rect 12851 9676 13084 9704
rect 12851 9673 12863 9676
rect 12805 9667 12863 9673
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13173 9707 13231 9713
rect 13173 9673 13185 9707
rect 13219 9704 13231 9707
rect 13446 9704 13452 9716
rect 13219 9676 13452 9704
rect 13219 9673 13231 9676
rect 13173 9667 13231 9673
rect 13446 9664 13452 9676
rect 13504 9664 13510 9716
rect 10192 9608 10364 9636
rect 10781 9639 10839 9645
rect 10192 9596 10198 9608
rect 10781 9605 10793 9639
rect 10827 9636 10839 9639
rect 11054 9636 11060 9648
rect 10827 9608 11060 9636
rect 10827 9605 10839 9608
rect 10781 9599 10839 9605
rect 11054 9596 11060 9608
rect 11112 9596 11118 9648
rect 11146 9596 11152 9648
rect 11204 9636 11210 9648
rect 11204 9608 11376 9636
rect 11204 9596 11210 9608
rect 5592 9540 6040 9568
rect 6089 9571 6147 9577
rect 5592 9528 5598 9540
rect 6089 9537 6101 9571
rect 6135 9568 6147 9571
rect 6822 9568 6828 9580
rect 6135 9540 6408 9568
rect 6135 9537 6147 9540
rect 6089 9531 6147 9537
rect 4433 9503 4491 9509
rect 4433 9469 4445 9503
rect 4479 9469 4491 9503
rect 5350 9500 5356 9512
rect 5311 9472 5356 9500
rect 4433 9463 4491 9469
rect 5350 9460 5356 9472
rect 5408 9460 5414 9512
rect 5626 9500 5632 9512
rect 5587 9472 5632 9500
rect 5626 9460 5632 9472
rect 5684 9460 5690 9512
rect 1670 9392 1676 9444
rect 1728 9432 1734 9444
rect 3881 9435 3939 9441
rect 3881 9432 3893 9435
rect 1728 9404 3893 9432
rect 1728 9392 1734 9404
rect 3881 9401 3893 9404
rect 3927 9401 3939 9435
rect 3881 9395 3939 9401
rect 4246 9392 4252 9444
rect 4304 9432 4310 9444
rect 6380 9432 6408 9540
rect 6564 9540 6828 9568
rect 6564 9509 6592 9540
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7558 9568 7564 9580
rect 7519 9540 7564 9568
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 8481 9571 8539 9577
rect 8481 9537 8493 9571
rect 8527 9568 8539 9571
rect 9398 9568 9404 9580
rect 8527 9540 9404 9568
rect 8527 9537 8539 9540
rect 8481 9531 8539 9537
rect 9398 9528 9404 9540
rect 9456 9528 9462 9580
rect 10689 9571 10747 9577
rect 9600 9540 10640 9568
rect 6549 9503 6607 9509
rect 6549 9469 6561 9503
rect 6595 9469 6607 9503
rect 6549 9463 6607 9469
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7650 9500 7656 9512
rect 6687 9472 7523 9500
rect 7611 9472 7656 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 6914 9432 6920 9444
rect 4304 9404 6123 9432
rect 6380 9404 6920 9432
rect 4304 9392 4310 9404
rect 1486 9364 1492 9376
rect 1447 9336 1492 9364
rect 1486 9324 1492 9336
rect 1544 9324 1550 9376
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 1765 9367 1823 9373
rect 1765 9364 1777 9367
rect 1636 9336 1777 9364
rect 1636 9324 1642 9336
rect 1765 9333 1777 9336
rect 1811 9333 1823 9367
rect 1765 9327 1823 9333
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2130 9364 2136 9376
rect 2087 9336 2136 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 2409 9367 2467 9373
rect 2409 9333 2421 9367
rect 2455 9364 2467 9367
rect 2498 9364 2504 9376
rect 2455 9336 2504 9364
rect 2455 9333 2467 9336
rect 2409 9327 2467 9333
rect 2498 9324 2504 9336
rect 2556 9324 2562 9376
rect 2590 9324 2596 9376
rect 2648 9364 2654 9376
rect 3789 9367 3847 9373
rect 2648 9336 2693 9364
rect 2648 9324 2654 9336
rect 3789 9333 3801 9367
rect 3835 9364 3847 9367
rect 4430 9364 4436 9376
rect 3835 9336 4436 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 4430 9324 4436 9336
rect 4488 9324 4494 9376
rect 4614 9324 4620 9376
rect 4672 9364 4678 9376
rect 4801 9367 4859 9373
rect 4801 9364 4813 9367
rect 4672 9336 4813 9364
rect 4672 9324 4678 9336
rect 4801 9333 4813 9336
rect 4847 9333 4859 9367
rect 6095 9364 6123 9404
rect 6914 9392 6920 9404
rect 6972 9392 6978 9444
rect 7098 9432 7104 9444
rect 7059 9404 7104 9432
rect 7098 9392 7104 9404
rect 7156 9392 7162 9444
rect 7495 9432 7523 9472
rect 7650 9460 7656 9472
rect 7708 9460 7714 9512
rect 7834 9500 7840 9512
rect 7795 9472 7840 9500
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9500 8723 9503
rect 9030 9500 9036 9512
rect 8711 9472 9036 9500
rect 8711 9469 8723 9472
rect 8665 9463 8723 9469
rect 9030 9460 9036 9472
rect 9088 9460 9094 9512
rect 9600 9509 9628 9540
rect 9585 9503 9643 9509
rect 9585 9469 9597 9503
rect 9631 9469 9643 9503
rect 9585 9463 9643 9469
rect 8021 9435 8079 9441
rect 8021 9432 8033 9435
rect 7495 9404 8033 9432
rect 8021 9401 8033 9404
rect 8067 9401 8079 9435
rect 8021 9395 8079 9401
rect 8938 9392 8944 9444
rect 8996 9432 9002 9444
rect 9217 9435 9275 9441
rect 9217 9432 9229 9435
rect 8996 9404 9229 9432
rect 8996 9392 9002 9404
rect 9217 9401 9229 9404
rect 9263 9401 9275 9435
rect 10612 9432 10640 9540
rect 10689 9537 10701 9571
rect 10735 9568 10747 9571
rect 11238 9568 11244 9580
rect 10735 9540 11244 9568
rect 10735 9537 10747 9540
rect 10689 9531 10747 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11348 9568 11376 9608
rect 11422 9596 11428 9648
rect 11480 9636 11486 9648
rect 11977 9639 12035 9645
rect 11977 9636 11989 9639
rect 11480 9608 11989 9636
rect 11480 9596 11486 9608
rect 11977 9605 11989 9608
rect 12023 9605 12035 9639
rect 11977 9599 12035 9605
rect 12713 9639 12771 9645
rect 12713 9605 12725 9639
rect 12759 9636 12771 9639
rect 14090 9636 14096 9648
rect 12759 9608 14096 9636
rect 12759 9605 12771 9608
rect 12713 9599 12771 9605
rect 14090 9596 14096 9608
rect 14148 9596 14154 9648
rect 14458 9636 14464 9648
rect 14200 9608 14464 9636
rect 11606 9568 11612 9580
rect 11348 9540 11612 9568
rect 11606 9528 11612 9540
rect 11664 9568 11670 9580
rect 11885 9571 11943 9577
rect 11885 9568 11897 9571
rect 11664 9540 11897 9568
rect 11664 9528 11670 9540
rect 11885 9537 11897 9540
rect 11931 9537 11943 9571
rect 11885 9531 11943 9537
rect 13446 9528 13452 9580
rect 13504 9568 13510 9580
rect 13541 9571 13599 9577
rect 13541 9568 13553 9571
rect 13504 9540 13553 9568
rect 13504 9528 13510 9540
rect 13541 9537 13553 9540
rect 13587 9568 13599 9571
rect 14200 9568 14228 9608
rect 14458 9596 14464 9608
rect 14516 9596 14522 9648
rect 13587 9540 14228 9568
rect 14369 9571 14427 9577
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 14369 9537 14381 9571
rect 14415 9568 14427 9571
rect 14826 9568 14832 9580
rect 14415 9540 14832 9568
rect 14415 9537 14427 9540
rect 14369 9531 14427 9537
rect 14826 9528 14832 9540
rect 14884 9528 14890 9580
rect 10870 9500 10876 9512
rect 10831 9472 10876 9500
rect 10870 9460 10876 9472
rect 10928 9460 10934 9512
rect 12066 9500 12072 9512
rect 11979 9472 12072 9500
rect 12066 9460 12072 9472
rect 12124 9460 12130 9512
rect 12618 9460 12624 9512
rect 12676 9500 12682 9512
rect 12897 9503 12955 9509
rect 12897 9500 12909 9503
rect 12676 9472 12909 9500
rect 12676 9460 12682 9472
rect 12897 9469 12909 9472
rect 12943 9469 12955 9503
rect 12897 9463 12955 9469
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9469 13691 9503
rect 13814 9500 13820 9512
rect 13775 9472 13820 9500
rect 13633 9463 13691 9469
rect 10778 9432 10784 9444
rect 10612 9404 10784 9432
rect 9217 9395 9275 9401
rect 10778 9392 10784 9404
rect 10836 9432 10842 9444
rect 12084 9432 12112 9460
rect 12342 9432 12348 9444
rect 10836 9404 12112 9432
rect 12303 9404 12348 9432
rect 10836 9392 10842 9404
rect 12342 9392 12348 9404
rect 12400 9392 12406 9444
rect 12526 9392 12532 9444
rect 12584 9432 12590 9444
rect 13648 9432 13676 9463
rect 13814 9460 13820 9472
rect 13872 9460 13878 9512
rect 14274 9460 14280 9512
rect 14332 9500 14338 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14332 9472 14473 9500
rect 14332 9460 14338 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 14550 9460 14556 9512
rect 14608 9500 14614 9512
rect 14608 9472 14653 9500
rect 14608 9460 14614 9472
rect 12584 9404 13676 9432
rect 12584 9392 12590 9404
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 15013 9435 15071 9441
rect 15013 9432 15025 9435
rect 13780 9404 15025 9432
rect 13780 9392 13786 9404
rect 15013 9401 15025 9404
rect 15059 9401 15071 9435
rect 15013 9395 15071 9401
rect 7193 9367 7251 9373
rect 7193 9364 7205 9367
rect 6095 9336 7205 9364
rect 4801 9327 4859 9333
rect 7193 9333 7205 9336
rect 7239 9333 7251 9367
rect 9030 9364 9036 9376
rect 8991 9336 9036 9364
rect 7193 9327 7251 9333
rect 9030 9324 9036 9336
rect 9088 9324 9094 9376
rect 9122 9324 9128 9376
rect 9180 9364 9186 9376
rect 9674 9364 9680 9376
rect 9180 9336 9680 9364
rect 9180 9324 9186 9336
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 11238 9364 11244 9376
rect 11199 9336 11244 9364
rect 11238 9324 11244 9336
rect 11296 9324 11302 9376
rect 12986 9324 12992 9376
rect 13044 9364 13050 9376
rect 14001 9367 14059 9373
rect 14001 9364 14013 9367
rect 13044 9336 14013 9364
rect 13044 9324 13050 9336
rect 14001 9333 14013 9336
rect 14047 9333 14059 9367
rect 14001 9327 14059 9333
rect 14458 9324 14464 9376
rect 14516 9364 14522 9376
rect 14918 9364 14924 9376
rect 14516 9336 14924 9364
rect 14516 9324 14522 9336
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 15289 9367 15347 9373
rect 15289 9333 15301 9367
rect 15335 9364 15347 9367
rect 15838 9364 15844 9376
rect 15335 9336 15844 9364
rect 15335 9333 15347 9336
rect 15289 9327 15347 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 3786 9160 3792 9172
rect 1780 9132 3556 9160
rect 3747 9132 3792 9160
rect 1670 8956 1676 8968
rect 1631 8928 1676 8956
rect 1670 8916 1676 8928
rect 1728 8916 1734 8968
rect 1780 8965 1808 9132
rect 3528 9024 3556 9132
rect 3786 9120 3792 9132
rect 3844 9120 3850 9172
rect 3970 9160 3976 9172
rect 3931 9132 3976 9160
rect 3970 9120 3976 9132
rect 4028 9120 4034 9172
rect 4154 9160 4160 9172
rect 4115 9132 4160 9160
rect 4154 9120 4160 9132
rect 4212 9120 4218 9172
rect 5902 9160 5908 9172
rect 4448 9132 5908 9160
rect 3605 9095 3663 9101
rect 3605 9061 3617 9095
rect 3651 9092 3663 9095
rect 3878 9092 3884 9104
rect 3651 9064 3884 9092
rect 3651 9061 3663 9064
rect 3605 9055 3663 9061
rect 3878 9052 3884 9064
rect 3936 9052 3942 9104
rect 4448 9024 4476 9132
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 7558 9120 7564 9172
rect 7616 9160 7622 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 7616 9132 8953 9160
rect 7616 9120 7622 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 9674 9120 9680 9172
rect 9732 9120 9738 9172
rect 8754 9092 8760 9104
rect 7576 9064 8760 9092
rect 7576 9036 7604 9064
rect 8754 9052 8760 9064
rect 8812 9052 8818 9104
rect 4614 9024 4620 9036
rect 3528 8996 4476 9024
rect 4575 8996 4620 9024
rect 4614 8984 4620 8996
rect 4672 8984 4678 9036
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 6454 9024 6460 9036
rect 4764 8996 4809 9024
rect 6415 8996 6460 9024
rect 4764 8984 4770 8996
rect 6454 8984 6460 8996
rect 6512 8984 6518 9036
rect 7558 8984 7564 9036
rect 7616 8984 7622 9036
rect 8202 9024 8208 9036
rect 8163 8996 8208 9024
rect 8202 8984 8208 8996
rect 8260 8984 8266 9036
rect 8846 8984 8852 9036
rect 8904 9024 8910 9036
rect 9493 9027 9551 9033
rect 9493 9024 9505 9027
rect 8904 8996 9505 9024
rect 8904 8984 8910 8996
rect 9493 8993 9505 8996
rect 9539 8993 9551 9027
rect 9692 9024 9720 9120
rect 14642 9052 14648 9104
rect 14700 9092 14706 9104
rect 14918 9092 14924 9104
rect 14700 9064 14924 9092
rect 14700 9052 14706 9064
rect 14918 9052 14924 9064
rect 14976 9052 14982 9104
rect 10778 9024 10784 9036
rect 9692 8996 10784 9024
rect 9493 8987 9551 8993
rect 10778 8984 10784 8996
rect 10836 8984 10842 9036
rect 12066 8984 12072 9036
rect 12124 9024 12130 9036
rect 12345 9027 12403 9033
rect 12345 9024 12357 9027
rect 12124 8996 12357 9024
rect 12124 8984 12130 8996
rect 12345 8993 12357 8996
rect 12391 8993 12403 9027
rect 12345 8987 12403 8993
rect 14553 9027 14611 9033
rect 14553 8993 14565 9027
rect 14599 9024 14611 9027
rect 15010 9024 15016 9036
rect 14599 8996 15016 9024
rect 14599 8993 14611 8996
rect 14553 8987 14611 8993
rect 15010 8984 15016 8996
rect 15068 8984 15074 9036
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8925 1823 8959
rect 1765 8919 1823 8925
rect 2225 8959 2283 8965
rect 2225 8925 2237 8959
rect 2271 8956 2283 8959
rect 3234 8956 3240 8968
rect 2271 8928 3240 8956
rect 2271 8925 2283 8928
rect 2225 8919 2283 8925
rect 3234 8916 3240 8928
rect 3292 8956 3298 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 3292 8928 4997 8956
rect 3292 8916 3298 8928
rect 4985 8925 4997 8928
rect 5031 8956 5043 8959
rect 5534 8956 5540 8968
rect 5031 8928 5540 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5534 8916 5540 8928
rect 5592 8956 5598 8968
rect 6472 8956 6500 8984
rect 7926 8956 7932 8968
rect 5592 8928 6500 8956
rect 7887 8928 7932 8956
rect 5592 8916 5598 8928
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 10134 8956 10140 8968
rect 10095 8928 10140 8956
rect 10134 8916 10140 8928
rect 10192 8916 10198 8968
rect 10873 8959 10931 8965
rect 10873 8925 10885 8959
rect 10919 8956 10931 8959
rect 10962 8956 10968 8968
rect 10919 8928 10968 8956
rect 10919 8925 10931 8928
rect 10873 8919 10931 8925
rect 10962 8916 10968 8928
rect 11020 8956 11026 8968
rect 12529 8959 12587 8965
rect 12529 8956 12541 8959
rect 11020 8928 11284 8956
rect 11020 8916 11026 8928
rect 2314 8888 2320 8900
rect 1964 8860 2320 8888
rect 1489 8823 1547 8829
rect 1489 8789 1501 8823
rect 1535 8820 1547 8823
rect 1670 8820 1676 8832
rect 1535 8792 1676 8820
rect 1535 8789 1547 8792
rect 1489 8783 1547 8789
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 1964 8829 1992 8860
rect 2314 8848 2320 8860
rect 2372 8848 2378 8900
rect 2492 8891 2550 8897
rect 2492 8857 2504 8891
rect 2538 8888 2550 8891
rect 3510 8888 3516 8900
rect 2538 8860 3516 8888
rect 2538 8857 2550 8860
rect 2492 8851 2550 8857
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 4430 8848 4436 8900
rect 4488 8888 4494 8900
rect 5230 8891 5288 8897
rect 5230 8888 5242 8891
rect 4488 8860 5242 8888
rect 4488 8848 4494 8860
rect 5230 8857 5242 8860
rect 5276 8857 5288 8891
rect 5230 8851 5288 8857
rect 5350 8848 5356 8900
rect 5408 8888 5414 8900
rect 6702 8891 6760 8897
rect 6702 8888 6714 8891
rect 5408 8860 6714 8888
rect 5408 8848 5414 8860
rect 6702 8857 6714 8860
rect 6748 8857 6760 8891
rect 6702 8851 6760 8857
rect 7190 8848 7196 8900
rect 7248 8888 7254 8900
rect 7248 8860 7705 8888
rect 7248 8848 7254 8860
rect 1949 8823 2007 8829
rect 1949 8789 1961 8823
rect 1995 8789 2007 8823
rect 1949 8783 2007 8789
rect 2133 8823 2191 8829
rect 2133 8789 2145 8823
rect 2179 8820 2191 8823
rect 4154 8820 4160 8832
rect 2179 8792 4160 8820
rect 2179 8789 2191 8792
rect 2133 8783 2191 8789
rect 4154 8780 4160 8792
rect 4212 8780 4218 8832
rect 4522 8820 4528 8832
rect 4483 8792 4528 8820
rect 4522 8780 4528 8792
rect 4580 8780 4586 8832
rect 6086 8780 6092 8832
rect 6144 8820 6150 8832
rect 6365 8823 6423 8829
rect 6365 8820 6377 8823
rect 6144 8792 6377 8820
rect 6144 8780 6150 8792
rect 6365 8789 6377 8792
rect 6411 8820 6423 8823
rect 7282 8820 7288 8832
rect 6411 8792 7288 8820
rect 6411 8789 6423 8792
rect 6365 8783 6423 8789
rect 7282 8780 7288 8792
rect 7340 8780 7346 8832
rect 7677 8820 7705 8860
rect 7742 8848 7748 8900
rect 7800 8888 7806 8900
rect 10594 8888 10600 8900
rect 7800 8860 10600 8888
rect 7800 8848 7806 8860
rect 10594 8848 10600 8860
rect 10652 8848 10658 8900
rect 10781 8891 10839 8897
rect 10781 8857 10793 8891
rect 10827 8888 10839 8891
rect 11118 8891 11176 8897
rect 11118 8888 11130 8891
rect 10827 8860 11130 8888
rect 10827 8857 10839 8860
rect 10781 8851 10839 8857
rect 11118 8857 11130 8860
rect 11164 8857 11176 8891
rect 11256 8888 11284 8928
rect 11992 8928 12541 8956
rect 11992 8888 12020 8928
rect 12529 8925 12541 8928
rect 12575 8956 12587 8959
rect 12575 8928 12940 8956
rect 12575 8925 12587 8928
rect 12529 8919 12587 8925
rect 12912 8900 12940 8928
rect 13354 8916 13360 8968
rect 13412 8956 13418 8968
rect 13722 8956 13728 8968
rect 13412 8928 13728 8956
rect 13412 8916 13418 8928
rect 13722 8916 13728 8928
rect 13780 8956 13786 8968
rect 14093 8959 14151 8965
rect 14093 8956 14105 8959
rect 13780 8928 14105 8956
rect 13780 8916 13786 8928
rect 14093 8925 14105 8928
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14642 8916 14648 8968
rect 14700 8956 14706 8968
rect 14829 8959 14887 8965
rect 14829 8956 14841 8959
rect 14700 8928 14841 8956
rect 14700 8916 14706 8928
rect 14829 8925 14841 8928
rect 14875 8925 14887 8959
rect 14829 8919 14887 8925
rect 15473 8959 15531 8965
rect 15473 8925 15485 8959
rect 15519 8956 15531 8959
rect 16022 8956 16028 8968
rect 15519 8928 16028 8956
rect 15519 8925 15531 8928
rect 15473 8919 15531 8925
rect 16022 8916 16028 8928
rect 16080 8916 16086 8968
rect 12796 8891 12854 8897
rect 12796 8888 12808 8891
rect 11256 8860 12020 8888
rect 12268 8860 12808 8888
rect 11118 8851 11176 8857
rect 7837 8823 7895 8829
rect 7837 8820 7849 8823
rect 7677 8792 7849 8820
rect 7837 8789 7849 8792
rect 7883 8789 7895 8823
rect 7837 8783 7895 8789
rect 9030 8780 9036 8832
rect 9088 8820 9094 8832
rect 9309 8823 9367 8829
rect 9309 8820 9321 8823
rect 9088 8792 9321 8820
rect 9088 8780 9094 8792
rect 9309 8789 9321 8792
rect 9355 8789 9367 8823
rect 9309 8783 9367 8789
rect 9398 8780 9404 8832
rect 9456 8820 9462 8832
rect 9766 8820 9772 8832
rect 9456 8792 9501 8820
rect 9727 8792 9772 8820
rect 9456 8780 9462 8792
rect 9766 8780 9772 8792
rect 9824 8780 9830 8832
rect 11974 8780 11980 8832
rect 12032 8820 12038 8832
rect 12268 8829 12296 8860
rect 12796 8857 12808 8860
rect 12842 8857 12854 8891
rect 12796 8851 12854 8857
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12032 8792 12265 8820
rect 12032 8780 12038 8792
rect 12253 8789 12265 8792
rect 12299 8789 12311 8823
rect 12820 8820 12848 8851
rect 12894 8848 12900 8900
rect 12952 8848 12958 8900
rect 14550 8888 14556 8900
rect 13004 8860 14556 8888
rect 13004 8820 13032 8860
rect 14550 8848 14556 8860
rect 14608 8848 14614 8900
rect 15289 8891 15347 8897
rect 15289 8857 15301 8891
rect 15335 8888 15347 8891
rect 15930 8888 15936 8900
rect 15335 8860 15936 8888
rect 15335 8857 15347 8860
rect 15289 8851 15347 8857
rect 15930 8848 15936 8860
rect 15988 8848 15994 8900
rect 12820 8792 13032 8820
rect 12253 8783 12311 8789
rect 13814 8780 13820 8832
rect 13872 8820 13878 8832
rect 13909 8823 13967 8829
rect 13909 8820 13921 8823
rect 13872 8792 13921 8820
rect 13872 8780 13878 8792
rect 13909 8789 13921 8792
rect 13955 8789 13967 8823
rect 14366 8820 14372 8832
rect 14327 8792 14372 8820
rect 13909 8783 13967 8789
rect 14366 8780 14372 8792
rect 14424 8780 14430 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 14645 8823 14703 8829
rect 14645 8820 14657 8823
rect 14516 8792 14657 8820
rect 14516 8780 14522 8792
rect 14645 8789 14657 8792
rect 14691 8789 14703 8823
rect 14645 8783 14703 8789
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 15013 8823 15071 8829
rect 15013 8820 15025 8823
rect 14792 8792 15025 8820
rect 14792 8780 14798 8792
rect 15013 8789 15025 8792
rect 15059 8789 15071 8823
rect 15013 8783 15071 8789
rect 15657 8823 15715 8829
rect 15657 8789 15669 8823
rect 15703 8820 15715 8823
rect 15746 8820 15752 8832
rect 15703 8792 15752 8820
rect 15703 8789 15715 8792
rect 15657 8783 15715 8789
rect 15746 8780 15752 8792
rect 15804 8780 15810 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 1762 8616 1768 8628
rect 1723 8588 1768 8616
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 3142 8576 3148 8628
rect 3200 8616 3206 8628
rect 3237 8619 3295 8625
rect 3237 8616 3249 8619
rect 3200 8588 3249 8616
rect 3200 8576 3206 8588
rect 3237 8585 3249 8588
rect 3283 8585 3295 8619
rect 3237 8579 3295 8585
rect 4154 8576 4160 8628
rect 4212 8616 4218 8628
rect 4709 8619 4767 8625
rect 4212 8588 4568 8616
rect 4212 8576 4218 8588
rect 4246 8548 4252 8560
rect 2240 8520 4252 8548
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1688 8412 1716 8443
rect 1854 8440 1860 8492
rect 1912 8480 1918 8492
rect 2240 8489 2268 8520
rect 4246 8508 4252 8520
rect 4304 8508 4310 8560
rect 1949 8483 2007 8489
rect 1949 8480 1961 8483
rect 1912 8452 1961 8480
rect 1912 8440 1918 8452
rect 1949 8449 1961 8452
rect 1995 8449 2007 8483
rect 1949 8443 2007 8449
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8449 2283 8483
rect 2498 8480 2504 8492
rect 2459 8452 2504 8480
rect 2225 8443 2283 8449
rect 2498 8440 2504 8452
rect 2556 8440 2562 8492
rect 2777 8483 2835 8489
rect 2777 8449 2789 8483
rect 2823 8449 2835 8483
rect 2777 8443 2835 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8480 3111 8483
rect 3142 8480 3148 8492
rect 3099 8452 3148 8480
rect 3099 8449 3111 8452
rect 3053 8443 3111 8449
rect 2792 8412 2820 8443
rect 3142 8440 3148 8452
rect 3200 8440 3206 8492
rect 3878 8440 3884 8492
rect 3936 8480 3942 8492
rect 4350 8483 4408 8489
rect 4350 8480 4362 8483
rect 3936 8452 4362 8480
rect 3936 8440 3942 8452
rect 4350 8449 4362 8452
rect 4396 8449 4408 8483
rect 4350 8443 4408 8449
rect 3602 8412 3608 8424
rect 1688 8384 2084 8412
rect 2792 8384 3608 8412
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 2056 8353 2084 8384
rect 3602 8372 3608 8384
rect 3660 8372 3666 8424
rect 4540 8412 4568 8588
rect 4709 8585 4721 8619
rect 4755 8616 4767 8619
rect 5350 8616 5356 8628
rect 4755 8588 5356 8616
rect 4755 8585 4767 8588
rect 4709 8579 4767 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5718 8616 5724 8628
rect 5679 8588 5724 8616
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5813 8619 5871 8625
rect 5813 8585 5825 8619
rect 5859 8616 5871 8619
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 5859 8588 8125 8616
rect 5859 8585 5871 8588
rect 5813 8579 5871 8585
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 8113 8579 8171 8585
rect 8941 8619 8999 8625
rect 8941 8585 8953 8619
rect 8987 8616 8999 8619
rect 9030 8616 9036 8628
rect 8987 8588 9036 8616
rect 8987 8585 8999 8588
rect 8941 8579 8999 8585
rect 9030 8576 9036 8588
rect 9088 8576 9094 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9858 8616 9864 8628
rect 9355 8588 9674 8616
rect 9819 8588 9864 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 5534 8548 5540 8560
rect 4816 8520 5540 8548
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8480 4675 8483
rect 4816 8480 4844 8520
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 6086 8548 6092 8560
rect 5920 8520 6092 8548
rect 4663 8452 4844 8480
rect 5353 8483 5411 8489
rect 4663 8449 4675 8452
rect 4617 8443 4675 8449
rect 5353 8449 5365 8483
rect 5399 8480 5411 8483
rect 5920 8480 5948 8520
rect 6086 8508 6092 8520
rect 6144 8508 6150 8560
rect 7101 8551 7159 8557
rect 6196 8520 7052 8548
rect 5399 8452 5948 8480
rect 5399 8449 5411 8452
rect 5353 8443 5411 8449
rect 5629 8415 5687 8421
rect 4540 8384 5589 8412
rect 2041 8347 2099 8353
rect 2041 8313 2053 8347
rect 2087 8313 2099 8347
rect 2041 8307 2099 8313
rect 2222 8304 2228 8356
rect 2280 8344 2286 8356
rect 2593 8347 2651 8353
rect 2593 8344 2605 8347
rect 2280 8316 2605 8344
rect 2280 8304 2286 8316
rect 2593 8313 2605 8316
rect 2639 8313 2651 8347
rect 2593 8307 2651 8313
rect 2869 8347 2927 8353
rect 2869 8313 2881 8347
rect 2915 8344 2927 8347
rect 3418 8344 3424 8356
rect 2915 8316 3424 8344
rect 2915 8313 2927 8316
rect 2869 8307 2927 8313
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 1762 8236 1768 8288
rect 1820 8276 1826 8288
rect 2317 8279 2375 8285
rect 2317 8276 2329 8279
rect 1820 8248 2329 8276
rect 1820 8236 1826 8248
rect 2317 8245 2329 8248
rect 2363 8245 2375 8279
rect 2317 8239 2375 8245
rect 3326 8236 3332 8288
rect 3384 8276 3390 8288
rect 3694 8276 3700 8288
rect 3384 8248 3700 8276
rect 3384 8236 3390 8248
rect 3694 8236 3700 8248
rect 3752 8236 3758 8288
rect 4246 8236 4252 8288
rect 4304 8276 4310 8288
rect 5166 8276 5172 8288
rect 4304 8248 5172 8276
rect 4304 8236 4310 8248
rect 5166 8236 5172 8248
rect 5224 8236 5230 8288
rect 5561 8276 5589 8384
rect 5629 8381 5641 8415
rect 5675 8412 5687 8415
rect 6196 8412 6224 8520
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 6365 8483 6423 8489
rect 6365 8480 6377 8483
rect 6328 8452 6377 8480
rect 6328 8440 6334 8452
rect 6365 8449 6377 8452
rect 6411 8449 6423 8483
rect 7024 8480 7052 8520
rect 7101 8517 7113 8551
rect 7147 8548 7159 8551
rect 8018 8548 8024 8560
rect 7147 8520 8024 8548
rect 7147 8517 7159 8520
rect 7101 8511 7159 8517
rect 8018 8508 8024 8520
rect 8076 8548 8082 8560
rect 9214 8548 9220 8560
rect 8076 8520 9220 8548
rect 8076 8508 8082 8520
rect 9214 8508 9220 8520
rect 9272 8508 9278 8560
rect 9646 8548 9674 8588
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8585 10011 8619
rect 9953 8579 10011 8585
rect 9766 8548 9772 8560
rect 9646 8520 9772 8548
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 8386 8480 8392 8492
rect 7024 8452 8392 8480
rect 6365 8443 6423 8449
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 8481 8483 8539 8489
rect 8481 8449 8493 8483
rect 8527 8480 8539 8483
rect 9122 8480 9128 8492
rect 8527 8452 9128 8480
rect 8527 8449 8539 8452
rect 8481 8443 8539 8449
rect 9122 8440 9128 8452
rect 9180 8440 9186 8492
rect 9876 8480 9904 8576
rect 9968 8548 9996 8579
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 10652 8588 12173 8616
rect 10652 8576 10658 8588
rect 12161 8585 12173 8588
rect 12207 8616 12219 8619
rect 12526 8616 12532 8628
rect 12207 8588 12434 8616
rect 12487 8588 12532 8616
rect 12207 8585 12219 8588
rect 12161 8579 12219 8585
rect 10134 8548 10140 8560
rect 9968 8520 10140 8548
rect 10134 8508 10140 8520
rect 10192 8548 10198 8560
rect 10870 8548 10876 8560
rect 10192 8520 10876 8548
rect 10192 8508 10198 8520
rect 10870 8508 10876 8520
rect 10928 8508 10934 8560
rect 10962 8508 10968 8560
rect 11020 8548 11026 8560
rect 12406 8548 12434 8588
rect 12526 8576 12532 8588
rect 12584 8576 12590 8628
rect 12897 8619 12955 8625
rect 12897 8585 12909 8619
rect 12943 8616 12955 8619
rect 12986 8616 12992 8628
rect 12943 8588 12992 8616
rect 12943 8585 12955 8588
rect 12897 8579 12955 8585
rect 12986 8576 12992 8588
rect 13044 8576 13050 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8616 13415 8619
rect 13538 8616 13544 8628
rect 13403 8588 13544 8616
rect 13403 8585 13415 8588
rect 13357 8579 13415 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 15286 8616 15292 8628
rect 14424 8588 15292 8616
rect 14424 8576 14430 8588
rect 15286 8576 15292 8588
rect 15344 8616 15350 8628
rect 16390 8616 16396 8628
rect 15344 8588 16396 8616
rect 15344 8576 15350 8588
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 12710 8548 12716 8560
rect 11020 8520 11376 8548
rect 12406 8520 12716 8548
rect 11020 8508 11026 8520
rect 11348 8489 11376 8520
rect 12710 8508 12716 8520
rect 12768 8508 12774 8560
rect 13814 8548 13820 8560
rect 12820 8520 13820 8548
rect 9416 8452 9904 8480
rect 11077 8483 11135 8489
rect 5675 8384 6224 8412
rect 6288 8384 6960 8412
rect 5675 8381 5687 8384
rect 5629 8375 5687 8381
rect 6181 8347 6239 8353
rect 6181 8313 6193 8347
rect 6227 8344 6239 8347
rect 6288 8344 6316 8384
rect 6227 8316 6316 8344
rect 6227 8313 6239 8316
rect 6181 8307 6239 8313
rect 6362 8304 6368 8356
rect 6420 8344 6426 8356
rect 6733 8347 6791 8353
rect 6733 8344 6745 8347
rect 6420 8316 6745 8344
rect 6420 8304 6426 8316
rect 6733 8313 6745 8316
rect 6779 8313 6791 8347
rect 6932 8344 6960 8384
rect 7098 8372 7104 8424
rect 7156 8412 7162 8424
rect 7193 8415 7251 8421
rect 7193 8412 7205 8415
rect 7156 8384 7205 8412
rect 7156 8372 7162 8384
rect 7193 8381 7205 8384
rect 7239 8381 7251 8415
rect 7193 8375 7251 8381
rect 7282 8372 7288 8424
rect 7340 8412 7346 8424
rect 7340 8384 7385 8412
rect 7340 8372 7346 8384
rect 7466 8372 7472 8424
rect 7524 8412 7530 8424
rect 7561 8415 7619 8421
rect 7561 8412 7573 8415
rect 7524 8384 7573 8412
rect 7524 8372 7530 8384
rect 7561 8381 7573 8384
rect 7607 8412 7619 8415
rect 7607 8384 8156 8412
rect 7607 8381 7619 8384
rect 7561 8375 7619 8381
rect 7650 8344 7656 8356
rect 6932 8316 7656 8344
rect 6733 8307 6791 8313
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 7742 8304 7748 8356
rect 7800 8344 7806 8356
rect 8128 8344 8156 8384
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8573 8415 8631 8421
rect 8573 8412 8585 8415
rect 8260 8384 8585 8412
rect 8260 8372 8266 8384
rect 8573 8381 8585 8384
rect 8619 8381 8631 8415
rect 8573 8375 8631 8381
rect 8662 8372 8668 8424
rect 8720 8412 8726 8424
rect 9416 8421 9444 8452
rect 11077 8449 11089 8483
rect 11123 8480 11135 8483
rect 11333 8483 11391 8489
rect 11123 8452 11284 8480
rect 11123 8449 11135 8452
rect 11077 8443 11135 8449
rect 9401 8415 9459 8421
rect 9401 8412 9413 8415
rect 8720 8384 8765 8412
rect 8864 8384 9413 8412
rect 8720 8372 8726 8384
rect 8864 8344 8892 8384
rect 9401 8381 9413 8384
rect 9447 8381 9459 8415
rect 9401 8375 9459 8381
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 11256 8412 11284 8452
rect 11333 8449 11345 8483
rect 11379 8449 11391 8483
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 11333 8443 11391 8449
rect 11808 8452 12081 8480
rect 11808 8424 11836 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 11514 8412 11520 8424
rect 11256 8384 11520 8412
rect 9493 8375 9551 8381
rect 7800 8316 7845 8344
rect 8128 8316 8892 8344
rect 7800 8304 7806 8316
rect 9214 8304 9220 8356
rect 9272 8344 9278 8356
rect 9508 8344 9536 8375
rect 11514 8372 11520 8384
rect 11572 8372 11578 8424
rect 11701 8415 11759 8421
rect 11701 8381 11713 8415
rect 11747 8412 11759 8415
rect 11790 8412 11796 8424
rect 11747 8384 11796 8412
rect 11747 8381 11759 8384
rect 11701 8375 11759 8381
rect 11790 8372 11796 8384
rect 11848 8372 11854 8424
rect 11974 8412 11980 8424
rect 11935 8384 11980 8412
rect 11974 8372 11980 8384
rect 12032 8372 12038 8424
rect 12820 8421 12848 8520
rect 13814 8508 13820 8520
rect 13872 8508 13878 8560
rect 12986 8480 12992 8492
rect 12947 8452 12992 8480
rect 12986 8440 12992 8452
rect 13044 8440 13050 8492
rect 13446 8480 13452 8492
rect 13407 8452 13452 8480
rect 13446 8440 13452 8452
rect 13504 8440 13510 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13832 8452 13921 8480
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 12805 8375 12863 8381
rect 9272 8316 9536 8344
rect 9272 8304 9278 8316
rect 11330 8304 11336 8356
rect 11388 8344 11394 8356
rect 13832 8353 13860 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 13817 8347 13875 8353
rect 13817 8344 13829 8347
rect 11388 8316 13829 8344
rect 11388 8304 11394 8316
rect 13817 8313 13829 8316
rect 13863 8313 13875 8347
rect 13817 8307 13875 8313
rect 5994 8276 6000 8288
rect 5561 8248 6000 8276
rect 5994 8236 6000 8248
rect 6052 8276 6058 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6052 8248 6561 8276
rect 6052 8236 6058 8248
rect 6549 8245 6561 8248
rect 6595 8245 6607 8279
rect 6549 8239 6607 8245
rect 7374 8236 7380 8288
rect 7432 8276 7438 8288
rect 7929 8279 7987 8285
rect 7929 8276 7941 8279
rect 7432 8248 7941 8276
rect 7432 8236 7438 8248
rect 7929 8245 7941 8248
rect 7975 8245 7987 8279
rect 7929 8239 7987 8245
rect 11698 8236 11704 8288
rect 11756 8276 11762 8288
rect 12710 8276 12716 8288
rect 11756 8248 12716 8276
rect 11756 8236 11762 8248
rect 12710 8236 12716 8248
rect 12768 8236 12774 8288
rect 15381 8279 15439 8285
rect 15381 8245 15393 8279
rect 15427 8276 15439 8279
rect 15654 8276 15660 8288
rect 15427 8248 15660 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 15654 8236 15660 8248
rect 15712 8236 15718 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 3694 8072 3700 8084
rect 2547 8044 3700 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 3694 8032 3700 8044
rect 3752 8032 3758 8084
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 5261 8075 5319 8081
rect 5261 8072 5273 8075
rect 4580 8044 5273 8072
rect 4580 8032 4586 8044
rect 5261 8041 5273 8044
rect 5307 8041 5319 8075
rect 5261 8035 5319 8041
rect 5718 8032 5724 8084
rect 5776 8072 5782 8084
rect 6089 8075 6147 8081
rect 6089 8072 6101 8075
rect 5776 8044 6101 8072
rect 5776 8032 5782 8044
rect 6089 8041 6101 8044
rect 6135 8041 6147 8075
rect 6089 8035 6147 8041
rect 8297 8075 8355 8081
rect 8297 8041 8309 8075
rect 8343 8072 8355 8075
rect 8386 8072 8392 8084
rect 8343 8044 8392 8072
rect 8343 8041 8355 8044
rect 8297 8035 8355 8041
rect 8386 8032 8392 8044
rect 8444 8072 8450 8084
rect 8846 8072 8852 8084
rect 8444 8044 8852 8072
rect 8444 8032 8450 8044
rect 8846 8032 8852 8044
rect 8904 8032 8910 8084
rect 8941 8075 8999 8081
rect 8941 8041 8953 8075
rect 8987 8072 8999 8075
rect 9398 8072 9404 8084
rect 8987 8044 9404 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9398 8032 9404 8044
rect 9456 8032 9462 8084
rect 9582 8032 9588 8084
rect 9640 8072 9646 8084
rect 9769 8075 9827 8081
rect 9769 8072 9781 8075
rect 9640 8044 9781 8072
rect 9640 8032 9646 8044
rect 9769 8041 9781 8044
rect 9815 8041 9827 8075
rect 9769 8035 9827 8041
rect 9858 8032 9864 8084
rect 9916 8072 9922 8084
rect 11241 8075 11299 8081
rect 11241 8072 11253 8075
rect 9916 8044 11253 8072
rect 9916 8032 9922 8044
rect 11241 8041 11253 8044
rect 11287 8072 11299 8075
rect 11698 8072 11704 8084
rect 11287 8044 11704 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 11698 8032 11704 8044
rect 11756 8072 11762 8084
rect 11882 8072 11888 8084
rect 11756 8044 11888 8072
rect 11756 8032 11762 8044
rect 11882 8032 11888 8044
rect 11940 8032 11946 8084
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 14093 8075 14151 8081
rect 14093 8072 14105 8075
rect 13044 8044 14105 8072
rect 13044 8032 13050 8044
rect 14093 8041 14105 8044
rect 14139 8041 14151 8075
rect 14918 8072 14924 8084
rect 14093 8035 14151 8041
rect 14292 8044 14924 8072
rect 14292 8016 14320 8044
rect 14918 8032 14924 8044
rect 14976 8072 14982 8084
rect 15105 8075 15163 8081
rect 15105 8072 15117 8075
rect 14976 8044 15117 8072
rect 14976 8032 14982 8044
rect 15105 8041 15117 8044
rect 15151 8041 15163 8075
rect 15105 8035 15163 8041
rect 1489 8007 1547 8013
rect 1489 7973 1501 8007
rect 1535 8004 1547 8007
rect 3050 8004 3056 8016
rect 1535 7976 3056 8004
rect 1535 7973 1547 7976
rect 1489 7967 1547 7973
rect 3050 7964 3056 7976
rect 3108 7964 3114 8016
rect 3510 7964 3516 8016
rect 3568 8004 3574 8016
rect 3789 8007 3847 8013
rect 3789 8004 3801 8007
rect 3568 7976 3801 8004
rect 3568 7964 3574 7976
rect 3789 7973 3801 7976
rect 3835 8004 3847 8007
rect 4154 8004 4160 8016
rect 3835 7976 4160 8004
rect 3835 7973 3847 7976
rect 3789 7967 3847 7973
rect 4154 7964 4160 7976
rect 4212 7964 4218 8016
rect 6454 8004 6460 8016
rect 5184 7976 6460 8004
rect 2590 7896 2596 7948
rect 2648 7896 2654 7948
rect 5184 7945 5212 7976
rect 6454 7964 6460 7976
rect 6512 8004 6518 8016
rect 6512 7976 6960 8004
rect 6512 7964 6518 7976
rect 5169 7939 5227 7945
rect 5169 7905 5181 7939
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5258 7896 5264 7948
rect 5316 7936 5322 7948
rect 5813 7939 5871 7945
rect 5813 7936 5825 7939
rect 5316 7908 5825 7936
rect 5316 7896 5322 7908
rect 5813 7905 5825 7908
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 6362 7896 6368 7948
rect 6420 7936 6426 7948
rect 6932 7945 6960 7976
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 9030 8004 9036 8016
rect 7984 7976 9036 8004
rect 7984 7964 7990 7976
rect 9030 7964 9036 7976
rect 9088 7964 9094 8016
rect 9953 8007 10011 8013
rect 9953 8004 9965 8007
rect 9416 7976 9965 8004
rect 9416 7948 9444 7976
rect 9953 7973 9965 7976
rect 9999 7973 10011 8007
rect 12618 8004 12624 8016
rect 9953 7967 10011 7973
rect 10152 7976 12624 8004
rect 6549 7939 6607 7945
rect 6549 7936 6561 7939
rect 6420 7908 6561 7936
rect 6420 7896 6426 7908
rect 6549 7905 6561 7908
rect 6595 7905 6607 7939
rect 6549 7899 6607 7905
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7905 6791 7939
rect 6733 7899 6791 7905
rect 6917 7939 6975 7945
rect 6917 7905 6929 7939
rect 6963 7905 6975 7939
rect 8478 7936 8484 7948
rect 8439 7908 8484 7936
rect 6917 7899 6975 7905
rect 1673 7871 1731 7877
rect 1673 7837 1685 7871
rect 1719 7868 1731 7871
rect 1762 7868 1768 7880
rect 1719 7840 1768 7868
rect 1719 7837 1731 7840
rect 1673 7831 1731 7837
rect 1762 7828 1768 7840
rect 1820 7828 1826 7880
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 2038 7868 2044 7880
rect 1995 7840 2044 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 2038 7828 2044 7840
rect 2096 7828 2102 7880
rect 2225 7871 2283 7877
rect 2225 7837 2237 7871
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 2317 7871 2375 7877
rect 2317 7837 2329 7871
rect 2363 7868 2375 7871
rect 2608 7868 2636 7896
rect 2363 7840 2636 7868
rect 3421 7871 3479 7877
rect 2363 7837 2375 7840
rect 2317 7831 2375 7837
rect 3421 7837 3433 7871
rect 3467 7868 3479 7871
rect 3510 7868 3516 7880
rect 3467 7840 3516 7868
rect 3467 7837 3479 7840
rect 3421 7831 3479 7837
rect 2240 7800 2268 7831
rect 3510 7828 3516 7840
rect 3568 7828 3574 7880
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5276 7868 5304 7896
rect 5626 7868 5632 7880
rect 4212 7840 5304 7868
rect 5587 7840 5632 7868
rect 4212 7828 4218 7840
rect 5626 7828 5632 7840
rect 5684 7828 5690 7880
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7868 5779 7871
rect 6178 7868 6184 7880
rect 5767 7840 6184 7868
rect 5767 7837 5779 7840
rect 5721 7831 5779 7837
rect 6178 7828 6184 7840
rect 6236 7828 6242 7880
rect 6748 7868 6776 7899
rect 8478 7896 8484 7908
rect 8536 7896 8542 7948
rect 9398 7936 9404 7948
rect 9359 7908 9404 7936
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 7190 7877 7196 7880
rect 7173 7871 7196 7877
rect 7173 7868 7185 7871
rect 6748 7840 7185 7868
rect 7173 7837 7185 7840
rect 7248 7868 7254 7880
rect 8662 7868 8668 7880
rect 7248 7840 8668 7868
rect 7173 7831 7196 7837
rect 7190 7828 7196 7831
rect 7248 7828 7254 7840
rect 8662 7828 8668 7840
rect 8720 7868 8726 7880
rect 9214 7868 9220 7880
rect 8720 7840 9220 7868
rect 8720 7828 8726 7840
rect 9214 7828 9220 7840
rect 9272 7868 9278 7880
rect 9508 7868 9536 7899
rect 9272 7840 9536 7868
rect 9272 7828 9278 7840
rect 2590 7800 2596 7812
rect 2240 7772 2596 7800
rect 2590 7760 2596 7772
rect 2648 7760 2654 7812
rect 2685 7803 2743 7809
rect 2685 7769 2697 7803
rect 2731 7800 2743 7803
rect 4246 7800 4252 7812
rect 2731 7772 4252 7800
rect 2731 7769 2743 7772
rect 2685 7763 2743 7769
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 4924 7803 4982 7809
rect 4924 7769 4936 7803
rect 4970 7800 4982 7803
rect 5166 7800 5172 7812
rect 4970 7772 5172 7800
rect 4970 7769 4982 7772
rect 4924 7763 4982 7769
rect 5166 7760 5172 7772
rect 5224 7760 5230 7812
rect 6457 7803 6515 7809
rect 6457 7769 6469 7803
rect 6503 7800 6515 7803
rect 7926 7800 7932 7812
rect 6503 7772 7932 7800
rect 6503 7769 6515 7772
rect 6457 7763 6515 7769
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 9309 7803 9367 7809
rect 9309 7769 9321 7803
rect 9355 7800 9367 7803
rect 9582 7800 9588 7812
rect 9355 7772 9588 7800
rect 9355 7769 9367 7772
rect 9309 7763 9367 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 1854 7732 1860 7744
rect 1811 7704 1860 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 1854 7692 1860 7704
rect 1912 7692 1918 7744
rect 2038 7732 2044 7744
rect 1999 7704 2044 7732
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 2832 7704 2877 7732
rect 2832 7692 2838 7704
rect 3326 7692 3332 7744
rect 3384 7732 3390 7744
rect 3513 7735 3571 7741
rect 3513 7732 3525 7735
rect 3384 7704 3525 7732
rect 3384 7692 3390 7704
rect 3513 7701 3525 7704
rect 3559 7701 3571 7735
rect 3513 7695 3571 7701
rect 3694 7692 3700 7744
rect 3752 7732 3758 7744
rect 5258 7732 5264 7744
rect 3752 7704 5264 7732
rect 3752 7692 3758 7704
rect 5258 7692 5264 7704
rect 5316 7692 5322 7744
rect 6362 7692 6368 7744
rect 6420 7732 6426 7744
rect 7466 7732 7472 7744
rect 6420 7704 7472 7732
rect 6420 7692 6426 7704
rect 7466 7692 7472 7704
rect 7524 7692 7530 7744
rect 8757 7735 8815 7741
rect 8757 7701 8769 7735
rect 8803 7732 8815 7735
rect 9122 7732 9128 7744
rect 8803 7704 9128 7732
rect 8803 7701 8815 7704
rect 8757 7695 8815 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 10152 7732 10180 7976
rect 12618 7964 12624 7976
rect 12676 8004 12682 8016
rect 13817 8007 13875 8013
rect 13817 8004 13829 8007
rect 12676 7976 13829 8004
rect 12676 7964 12682 7976
rect 10870 7936 10876 7948
rect 10831 7908 10876 7936
rect 10870 7896 10876 7908
rect 10928 7896 10934 7948
rect 11514 7896 11520 7948
rect 11572 7936 11578 7948
rect 11977 7939 12035 7945
rect 11977 7936 11989 7939
rect 11572 7908 11989 7936
rect 11572 7896 11578 7908
rect 11977 7905 11989 7908
rect 12023 7905 12035 7939
rect 11977 7899 12035 7905
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10778 7868 10784 7880
rect 10275 7840 10784 7868
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 11054 7828 11060 7880
rect 11112 7868 11118 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 11112 7840 12265 7868
rect 11112 7828 11118 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12710 7828 12716 7880
rect 12768 7868 12774 7880
rect 12989 7871 13047 7877
rect 12989 7868 13001 7871
rect 12768 7840 13001 7868
rect 12768 7828 12774 7840
rect 12989 7837 13001 7840
rect 13035 7837 13047 7871
rect 12989 7831 13047 7837
rect 10689 7803 10747 7809
rect 10689 7769 10701 7803
rect 10735 7800 10747 7803
rect 11793 7803 11851 7809
rect 10735 7772 11468 7800
rect 10735 7769 10747 7772
rect 10689 7763 10747 7769
rect 10318 7732 10324 7744
rect 9456 7704 10180 7732
rect 10279 7704 10324 7732
rect 9456 7692 9462 7704
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 10410 7692 10416 7744
rect 10468 7732 10474 7744
rect 11440 7741 11468 7772
rect 11793 7769 11805 7803
rect 11839 7800 11851 7803
rect 12802 7800 12808 7812
rect 11839 7772 12808 7800
rect 11839 7769 11851 7772
rect 11793 7763 11851 7769
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 10781 7735 10839 7741
rect 10781 7732 10793 7735
rect 10468 7704 10793 7732
rect 10468 7692 10474 7704
rect 10781 7701 10793 7704
rect 10827 7701 10839 7735
rect 10781 7695 10839 7701
rect 11425 7735 11483 7741
rect 11425 7701 11437 7735
rect 11471 7701 11483 7735
rect 11425 7695 11483 7701
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 11940 7704 11985 7732
rect 11940 7692 11946 7704
rect 12618 7692 12624 7744
rect 12676 7732 12682 7744
rect 12897 7735 12955 7741
rect 12897 7732 12909 7735
rect 12676 7704 12909 7732
rect 12676 7692 12682 7704
rect 12897 7701 12909 7704
rect 12943 7701 12955 7735
rect 12897 7695 12955 7701
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13096 7732 13124 7976
rect 13817 7973 13829 7976
rect 13863 7973 13875 8007
rect 13817 7967 13875 7973
rect 13170 7760 13176 7812
rect 13228 7800 13234 7812
rect 13541 7803 13599 7809
rect 13541 7800 13553 7803
rect 13228 7772 13553 7800
rect 13228 7760 13234 7772
rect 13541 7769 13553 7772
rect 13587 7800 13599 7803
rect 13722 7800 13728 7812
rect 13587 7772 13728 7800
rect 13587 7769 13599 7772
rect 13541 7763 13599 7769
rect 13722 7760 13728 7772
rect 13780 7760 13786 7812
rect 13832 7800 13860 7967
rect 14274 7964 14280 8016
rect 14332 7964 14338 8016
rect 14550 7896 14556 7948
rect 14608 7936 14614 7948
rect 14645 7939 14703 7945
rect 14645 7936 14657 7939
rect 14608 7908 14657 7936
rect 14608 7896 14614 7908
rect 14645 7905 14657 7908
rect 14691 7905 14703 7939
rect 14645 7899 14703 7905
rect 14366 7828 14372 7880
rect 14424 7868 14430 7880
rect 14461 7871 14519 7877
rect 14461 7868 14473 7871
rect 14424 7840 14473 7868
rect 14424 7828 14430 7840
rect 14461 7837 14473 7840
rect 14507 7837 14519 7871
rect 14461 7831 14519 7837
rect 14553 7803 14611 7809
rect 14553 7800 14565 7803
rect 13832 7772 14565 7800
rect 14553 7769 14565 7772
rect 14599 7800 14611 7803
rect 15286 7800 15292 7812
rect 14599 7772 15292 7800
rect 14599 7769 14611 7772
rect 14553 7763 14611 7769
rect 15286 7760 15292 7772
rect 15344 7760 15350 7812
rect 15381 7803 15439 7809
rect 15381 7769 15393 7803
rect 15427 7800 15439 7803
rect 16206 7800 16212 7812
rect 15427 7772 16212 7800
rect 15427 7769 15439 7772
rect 15381 7763 15439 7769
rect 16206 7760 16212 7772
rect 16264 7760 16270 7812
rect 13354 7732 13360 7744
rect 13044 7704 13124 7732
rect 13315 7704 13360 7732
rect 13044 7692 13050 7704
rect 13354 7692 13360 7704
rect 13412 7692 13418 7744
rect 13630 7732 13636 7744
rect 13591 7704 13636 7732
rect 13630 7692 13636 7704
rect 13688 7692 13694 7744
rect 14918 7732 14924 7744
rect 14879 7704 14924 7732
rect 14918 7692 14924 7704
rect 14976 7692 14982 7744
rect 15562 7732 15568 7744
rect 15523 7704 15568 7732
rect 15562 7692 15568 7704
rect 15620 7692 15626 7744
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 3053 7531 3111 7537
rect 3053 7497 3065 7531
rect 3099 7528 3111 7531
rect 3234 7528 3240 7540
rect 3099 7500 3240 7528
rect 3099 7497 3111 7500
rect 3053 7491 3111 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 3602 7488 3608 7540
rect 3660 7528 3666 7540
rect 4985 7531 5043 7537
rect 4985 7528 4997 7531
rect 3660 7500 4997 7528
rect 3660 7488 3666 7500
rect 4985 7497 4997 7500
rect 5031 7528 5043 7531
rect 5350 7528 5356 7540
rect 5031 7500 5356 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 5350 7488 5356 7500
rect 5408 7488 5414 7540
rect 5442 7488 5448 7540
rect 5500 7528 5506 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5500 7500 6377 7528
rect 5500 7488 5506 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7432 7500 7665 7528
rect 7432 7488 7438 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7834 7528 7840 7540
rect 7747 7500 7840 7528
rect 7653 7491 7711 7497
rect 7834 7488 7840 7500
rect 7892 7528 7898 7540
rect 10410 7528 10416 7540
rect 7892 7500 9352 7528
rect 10371 7500 10416 7528
rect 7892 7488 7898 7500
rect 2314 7420 2320 7472
rect 2372 7460 2378 7472
rect 3970 7460 3976 7472
rect 2372 7432 3976 7460
rect 2372 7420 2378 7432
rect 3970 7420 3976 7432
rect 4028 7420 4034 7472
rect 4338 7460 4344 7472
rect 4299 7432 4344 7460
rect 4338 7420 4344 7432
rect 4396 7420 4402 7472
rect 4525 7463 4583 7469
rect 4525 7429 4537 7463
rect 4571 7460 4583 7463
rect 5074 7460 5080 7472
rect 4571 7432 5080 7460
rect 4571 7429 4583 7432
rect 4525 7423 4583 7429
rect 5074 7420 5080 7432
rect 5132 7420 5138 7472
rect 5534 7420 5540 7472
rect 5592 7460 5598 7472
rect 6825 7463 6883 7469
rect 6825 7460 6837 7463
rect 5592 7432 6837 7460
rect 5592 7420 5598 7432
rect 6825 7429 6837 7432
rect 6871 7429 6883 7463
rect 6825 7423 6883 7429
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 8950 7463 9008 7469
rect 8950 7460 8962 7463
rect 8904 7432 8962 7460
rect 8904 7420 8910 7432
rect 8950 7429 8962 7432
rect 8996 7429 9008 7463
rect 9324 7460 9352 7500
rect 10410 7488 10416 7500
rect 10468 7488 10474 7540
rect 13449 7531 13507 7537
rect 13449 7497 13461 7531
rect 13495 7528 13507 7531
rect 13906 7528 13912 7540
rect 13495 7500 13912 7528
rect 13495 7497 13507 7500
rect 13449 7491 13507 7497
rect 13906 7488 13912 7500
rect 13964 7488 13970 7540
rect 14550 7488 14556 7540
rect 14608 7528 14614 7540
rect 15013 7531 15071 7537
rect 15013 7528 15025 7531
rect 14608 7500 15025 7528
rect 14608 7488 14614 7500
rect 15013 7497 15025 7500
rect 15059 7497 15071 7531
rect 15013 7491 15071 7497
rect 15657 7531 15715 7537
rect 15657 7497 15669 7531
rect 15703 7528 15715 7531
rect 16298 7528 16304 7540
rect 15703 7500 16304 7528
rect 15703 7497 15715 7500
rect 15657 7491 15715 7497
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 11054 7460 11060 7472
rect 9324 7432 11060 7460
rect 8950 7423 9008 7429
rect 11054 7420 11060 7432
rect 11112 7420 11118 7472
rect 11146 7420 11152 7472
rect 11204 7460 11210 7472
rect 11606 7460 11612 7472
rect 11204 7432 11612 7460
rect 11204 7420 11210 7432
rect 11606 7420 11612 7432
rect 11664 7460 11670 7472
rect 12342 7460 12348 7472
rect 11664 7432 12348 7460
rect 11664 7420 11670 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 12526 7420 12532 7472
rect 12584 7460 12590 7472
rect 12630 7463 12688 7469
rect 12630 7460 12642 7463
rect 12584 7432 12642 7460
rect 12584 7420 12590 7432
rect 12630 7429 12642 7432
rect 12676 7429 12688 7463
rect 12630 7423 12688 7429
rect 14366 7420 14372 7472
rect 14424 7460 14430 7472
rect 14829 7463 14887 7469
rect 14829 7460 14841 7463
rect 14424 7432 14841 7460
rect 14424 7420 14430 7432
rect 14829 7429 14841 7432
rect 14875 7429 14887 7463
rect 14829 7423 14887 7429
rect 1670 7392 1676 7404
rect 1631 7364 1676 7392
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 2041 7395 2099 7401
rect 2041 7361 2053 7395
rect 2087 7392 2099 7395
rect 2222 7392 2228 7404
rect 2087 7364 2228 7392
rect 2087 7361 2099 7364
rect 2041 7355 2099 7361
rect 2222 7352 2228 7364
rect 2280 7352 2286 7404
rect 2406 7352 2412 7404
rect 2464 7392 2470 7404
rect 2501 7395 2559 7401
rect 2501 7392 2513 7395
rect 2464 7364 2513 7392
rect 2464 7352 2470 7364
rect 2501 7361 2513 7364
rect 2547 7361 2559 7395
rect 2501 7355 2559 7361
rect 2682 7352 2688 7404
rect 2740 7392 2746 7404
rect 2740 7352 2774 7392
rect 3326 7352 3332 7404
rect 3384 7392 3390 7404
rect 4798 7392 4804 7404
rect 3384 7364 4804 7392
rect 3384 7352 3390 7364
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 5092 7392 5120 7420
rect 5626 7392 5632 7404
rect 5092 7364 5632 7392
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 5736 7364 5825 7392
rect 2746 7256 2774 7352
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3694 7324 3700 7336
rect 3108 7296 3700 7324
rect 3108 7284 3114 7296
rect 3694 7284 3700 7296
rect 3752 7284 3758 7336
rect 4614 7284 4620 7336
rect 4672 7324 4678 7336
rect 5074 7324 5080 7336
rect 4672 7296 5080 7324
rect 4672 7284 4678 7296
rect 5074 7284 5080 7296
rect 5132 7284 5138 7336
rect 5261 7327 5319 7333
rect 5261 7324 5273 7327
rect 5184 7296 5273 7324
rect 5184 7268 5212 7296
rect 5261 7293 5273 7296
rect 5307 7293 5319 7327
rect 5261 7287 5319 7293
rect 2746 7228 4752 7256
rect 1486 7188 1492 7200
rect 1447 7160 1492 7188
rect 1486 7148 1492 7160
rect 1544 7148 1550 7200
rect 1857 7191 1915 7197
rect 1857 7157 1869 7191
rect 1903 7188 1915 7191
rect 2222 7188 2228 7200
rect 1903 7160 2228 7188
rect 1903 7157 1915 7160
rect 1857 7151 1915 7157
rect 2222 7148 2228 7160
rect 2280 7148 2286 7200
rect 2317 7191 2375 7197
rect 2317 7157 2329 7191
rect 2363 7188 2375 7191
rect 2590 7188 2596 7200
rect 2363 7160 2596 7188
rect 2363 7157 2375 7160
rect 2317 7151 2375 7157
rect 2590 7148 2596 7160
rect 2648 7148 2654 7200
rect 4614 7188 4620 7200
rect 4575 7160 4620 7188
rect 4614 7148 4620 7160
rect 4672 7148 4678 7200
rect 4724 7188 4752 7228
rect 5166 7216 5172 7268
rect 5224 7216 5230 7268
rect 5736 7256 5764 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5905 7395 5963 7401
rect 5905 7361 5917 7395
rect 5951 7392 5963 7395
rect 5994 7392 6000 7404
rect 5951 7364 6000 7392
rect 5951 7361 5963 7364
rect 5905 7355 5963 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 6454 7352 6460 7404
rect 6512 7392 6518 7404
rect 6733 7395 6791 7401
rect 6733 7392 6745 7395
rect 6512 7364 6745 7392
rect 6512 7352 6518 7364
rect 6733 7361 6745 7364
rect 6779 7361 6791 7395
rect 7374 7392 7380 7404
rect 7335 7364 7380 7392
rect 6733 7355 6791 7361
rect 7374 7352 7380 7364
rect 7432 7352 7438 7404
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7392 7619 7395
rect 9217 7395 9275 7401
rect 7607 7364 9168 7392
rect 7607 7361 7619 7364
rect 7561 7355 7619 7361
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 6012 7296 6101 7324
rect 6012 7268 6040 7296
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6914 7324 6920 7336
rect 6875 7296 6920 7324
rect 6089 7287 6147 7293
rect 6914 7284 6920 7296
rect 6972 7284 6978 7336
rect 5276 7228 5764 7256
rect 5276 7188 5304 7228
rect 5442 7188 5448 7200
rect 4724 7160 5304 7188
rect 5403 7160 5448 7188
rect 5442 7148 5448 7160
rect 5500 7148 5506 7200
rect 5736 7188 5764 7228
rect 5994 7216 6000 7268
rect 6052 7216 6058 7268
rect 7576 7256 7604 7355
rect 9140 7324 9168 7364
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9858 7392 9864 7404
rect 9263 7364 9864 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 9858 7352 9864 7364
rect 9916 7352 9922 7404
rect 10045 7395 10103 7401
rect 10045 7361 10057 7395
rect 10091 7392 10103 7395
rect 12250 7392 12256 7404
rect 10091 7364 12256 7392
rect 10091 7361 10103 7364
rect 10045 7355 10103 7361
rect 12250 7352 12256 7364
rect 12308 7352 12314 7404
rect 12894 7392 12900 7404
rect 12855 7364 12900 7392
rect 12894 7352 12900 7364
rect 12952 7352 12958 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 15654 7392 15660 7404
rect 14783 7364 15660 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 15654 7352 15660 7364
rect 15712 7352 15718 7404
rect 9769 7327 9827 7333
rect 9140 7296 9628 7324
rect 9493 7259 9551 7265
rect 9493 7256 9505 7259
rect 6095 7228 7604 7256
rect 9232 7228 9505 7256
rect 6095 7188 6123 7228
rect 5736 7160 6123 7188
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7193 7191 7251 7197
rect 7193 7188 7205 7191
rect 6972 7160 7205 7188
rect 6972 7148 6978 7160
rect 7193 7157 7205 7160
rect 7239 7157 7251 7191
rect 7193 7151 7251 7157
rect 7650 7148 7656 7200
rect 7708 7188 7714 7200
rect 9232 7188 9260 7228
rect 9493 7225 9505 7228
rect 9539 7225 9551 7259
rect 9493 7219 9551 7225
rect 9398 7188 9404 7200
rect 7708 7160 9260 7188
rect 9359 7160 9404 7188
rect 7708 7148 7714 7160
rect 9398 7148 9404 7160
rect 9456 7148 9462 7200
rect 9600 7188 9628 7296
rect 9769 7293 9781 7327
rect 9815 7293 9827 7327
rect 9950 7324 9956 7336
rect 9911 7296 9956 7324
rect 9769 7287 9827 7293
rect 9784 7256 9812 7287
rect 9950 7284 9956 7296
rect 10008 7284 10014 7336
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 11146 7324 11152 7336
rect 10551 7296 11152 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 11146 7284 11152 7296
rect 11204 7284 11210 7336
rect 13906 7284 13912 7336
rect 13964 7324 13970 7336
rect 14826 7324 14832 7336
rect 13964 7296 14832 7324
rect 13964 7284 13970 7296
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15194 7284 15200 7336
rect 15252 7324 15258 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 15252 7296 15393 7324
rect 15252 7284 15258 7296
rect 15381 7293 15393 7296
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 11514 7256 11520 7268
rect 9784 7228 11520 7256
rect 11514 7216 11520 7228
rect 11572 7216 11578 7268
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 14550 7256 14556 7268
rect 14332 7228 14556 7256
rect 14332 7216 14338 7228
rect 14550 7216 14556 7228
rect 14608 7216 14614 7268
rect 9766 7188 9772 7200
rect 9600 7160 9772 7188
rect 9766 7148 9772 7160
rect 9824 7148 9830 7200
rect 10134 7148 10140 7200
rect 10192 7188 10198 7200
rect 10735 7191 10793 7197
rect 10735 7188 10747 7191
rect 10192 7160 10747 7188
rect 10192 7148 10198 7160
rect 10735 7157 10747 7160
rect 10781 7157 10793 7191
rect 10735 7151 10793 7157
rect 10870 7148 10876 7200
rect 10928 7188 10934 7200
rect 12618 7188 12624 7200
rect 10928 7160 12624 7188
rect 10928 7148 10934 7160
rect 12618 7148 12624 7160
rect 12676 7148 12682 7200
rect 15289 7191 15347 7197
rect 15289 7157 15301 7191
rect 15335 7188 15347 7191
rect 16114 7188 16120 7200
rect 15335 7160 16120 7188
rect 15335 7157 15347 7160
rect 15289 7151 15347 7157
rect 16114 7148 16120 7160
rect 16172 7188 16178 7200
rect 16574 7188 16580 7200
rect 16172 7160 16580 7188
rect 16172 7148 16178 7160
rect 16574 7148 16580 7160
rect 16632 7148 16638 7200
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 3605 6987 3663 6993
rect 3605 6953 3617 6987
rect 3651 6984 3663 6987
rect 5166 6984 5172 6996
rect 3651 6956 5172 6984
rect 3651 6953 3663 6956
rect 3605 6947 3663 6953
rect 5166 6944 5172 6956
rect 5224 6984 5230 6996
rect 5810 6984 5816 6996
rect 5224 6956 5816 6984
rect 5224 6944 5230 6956
rect 5810 6944 5816 6956
rect 5868 6944 5874 6996
rect 5997 6987 6055 6993
rect 5997 6953 6009 6987
rect 6043 6984 6055 6987
rect 6454 6984 6460 6996
rect 6043 6956 6460 6984
rect 6043 6953 6055 6956
rect 5997 6947 6055 6953
rect 6454 6944 6460 6956
rect 6512 6944 6518 6996
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 11241 6987 11299 6993
rect 11241 6984 11253 6987
rect 10008 6956 11253 6984
rect 10008 6944 10014 6956
rect 11241 6953 11253 6956
rect 11287 6953 11299 6987
rect 11241 6947 11299 6953
rect 11514 6944 11520 6996
rect 11572 6984 11578 6996
rect 12158 6984 12164 6996
rect 11572 6956 12164 6984
rect 11572 6944 11578 6956
rect 12158 6944 12164 6956
rect 12216 6944 12222 6996
rect 12526 6944 12532 6996
rect 12584 6944 12590 6996
rect 12618 6944 12624 6996
rect 12676 6984 12682 6996
rect 12676 6956 12756 6984
rect 12676 6944 12682 6956
rect 1394 6876 1400 6928
rect 1452 6916 1458 6928
rect 1946 6916 1952 6928
rect 1452 6888 1952 6916
rect 1452 6876 1458 6888
rect 1946 6876 1952 6888
rect 2004 6876 2010 6928
rect 4065 6919 4123 6925
rect 4065 6916 4077 6919
rect 3988 6888 4077 6916
rect 1581 6851 1639 6857
rect 1581 6817 1593 6851
rect 1627 6848 1639 6851
rect 1670 6848 1676 6860
rect 1627 6820 1676 6848
rect 1627 6817 1639 6820
rect 1581 6811 1639 6817
rect 1670 6808 1676 6820
rect 1728 6808 1734 6860
rect 2225 6783 2283 6789
rect 2225 6749 2237 6783
rect 2271 6780 2283 6783
rect 3234 6780 3240 6792
rect 2271 6752 3240 6780
rect 2271 6749 2283 6752
rect 2225 6743 2283 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 3384 6752 3464 6780
rect 3384 6740 3390 6752
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 1946 6712 1952 6724
rect 1719 6684 1952 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 1946 6672 1952 6684
rect 2004 6672 2010 6724
rect 2492 6715 2550 6721
rect 2492 6681 2504 6715
rect 2538 6712 2550 6715
rect 2774 6712 2780 6724
rect 2538 6684 2780 6712
rect 2538 6681 2550 6684
rect 2492 6675 2550 6681
rect 2774 6672 2780 6684
rect 2832 6672 2838 6724
rect 1762 6604 1768 6656
rect 1820 6644 1826 6656
rect 2133 6647 2191 6653
rect 1820 6616 1865 6644
rect 1820 6604 1826 6616
rect 2133 6613 2145 6647
rect 2179 6644 2191 6647
rect 3050 6644 3056 6656
rect 2179 6616 3056 6644
rect 2179 6613 2191 6616
rect 2133 6607 2191 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3436 6644 3464 6752
rect 3602 6740 3608 6792
rect 3660 6780 3666 6792
rect 3878 6780 3884 6792
rect 3660 6752 3884 6780
rect 3660 6740 3666 6752
rect 3878 6740 3884 6752
rect 3936 6740 3942 6792
rect 3988 6712 4016 6888
rect 4065 6885 4077 6888
rect 4111 6885 4123 6919
rect 4065 6879 4123 6885
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 11149 6919 11207 6925
rect 4212 6888 4844 6916
rect 4212 6876 4218 6888
rect 4246 6808 4252 6860
rect 4304 6808 4310 6860
rect 4540 6857 4568 6888
rect 4525 6851 4583 6857
rect 4525 6817 4537 6851
rect 4571 6817 4583 6851
rect 4525 6811 4583 6817
rect 4614 6808 4620 6860
rect 4672 6848 4678 6860
rect 4709 6851 4767 6857
rect 4709 6848 4721 6851
rect 4672 6820 4721 6848
rect 4672 6808 4678 6820
rect 4709 6817 4721 6820
rect 4755 6817 4767 6851
rect 4816 6848 4844 6888
rect 11149 6885 11161 6919
rect 11195 6885 11207 6919
rect 12544 6916 12572 6944
rect 12728 6916 12756 6956
rect 12802 6944 12808 6996
rect 12860 6984 12866 6996
rect 12897 6987 12955 6993
rect 12897 6984 12909 6987
rect 12860 6956 12909 6984
rect 12860 6944 12866 6956
rect 12897 6953 12909 6956
rect 12943 6953 12955 6987
rect 12897 6947 12955 6953
rect 14921 6987 14979 6993
rect 14921 6953 14933 6987
rect 14967 6984 14979 6987
rect 15286 6984 15292 6996
rect 14967 6956 15292 6984
rect 14967 6953 14979 6956
rect 14921 6947 14979 6953
rect 15286 6944 15292 6956
rect 15344 6944 15350 6996
rect 13722 6916 13728 6928
rect 11149 6879 11207 6885
rect 11808 6888 12664 6916
rect 12728 6888 13728 6916
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 4816 6820 5365 6848
rect 4709 6811 4767 6817
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5353 6811 5411 6817
rect 5442 6808 5448 6860
rect 5500 6848 5506 6860
rect 5537 6851 5595 6857
rect 5537 6848 5549 6851
rect 5500 6820 5549 6848
rect 5500 6808 5506 6820
rect 5537 6817 5549 6820
rect 5583 6817 5595 6851
rect 5537 6811 5595 6817
rect 5810 6808 5816 6860
rect 5868 6848 5874 6860
rect 5994 6848 6000 6860
rect 5868 6820 6000 6848
rect 5868 6808 5874 6820
rect 5994 6808 6000 6820
rect 6052 6848 6058 6860
rect 6641 6851 6699 6857
rect 6641 6848 6653 6851
rect 6052 6820 6653 6848
rect 6052 6808 6058 6820
rect 6641 6817 6653 6820
rect 6687 6817 6699 6851
rect 7466 6848 7472 6860
rect 7427 6820 7472 6848
rect 6641 6811 6699 6817
rect 7466 6808 7472 6820
rect 7524 6808 7530 6860
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6817 7711 6851
rect 8846 6848 8852 6860
rect 7653 6811 7711 6817
rect 8128 6820 8852 6848
rect 4264 6780 4292 6808
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 4264 6752 4353 6780
rect 4341 6749 4353 6752
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 5902 6740 5908 6792
rect 5960 6780 5966 6792
rect 6457 6783 6515 6789
rect 6457 6780 6469 6783
rect 5960 6752 6469 6780
rect 5960 6740 5966 6752
rect 6457 6749 6469 6752
rect 6503 6749 6515 6783
rect 6457 6743 6515 6749
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 7282 6780 7288 6792
rect 6595 6752 7288 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 7282 6740 7288 6752
rect 7340 6740 7346 6792
rect 4430 6712 4436 6724
rect 3988 6684 4436 6712
rect 4430 6672 4436 6684
rect 4488 6672 4494 6724
rect 4801 6715 4859 6721
rect 4801 6681 4813 6715
rect 4847 6712 4859 6715
rect 7377 6715 7435 6721
rect 4847 6684 6132 6712
rect 4847 6681 4859 6684
rect 4801 6675 4859 6681
rect 4157 6647 4215 6653
rect 4157 6644 4169 6647
rect 3436 6616 4169 6644
rect 4157 6613 4169 6616
rect 4203 6613 4215 6647
rect 4157 6607 4215 6613
rect 5169 6647 5227 6653
rect 5169 6613 5181 6647
rect 5215 6644 5227 6647
rect 5534 6644 5540 6656
rect 5215 6616 5540 6644
rect 5215 6613 5227 6616
rect 5169 6607 5227 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5626 6604 5632 6656
rect 5684 6644 5690 6656
rect 6104 6653 6132 6684
rect 7377 6681 7389 6715
rect 7423 6681 7435 6715
rect 7668 6712 7696 6811
rect 8128 6789 8156 6820
rect 8846 6808 8852 6820
rect 8904 6848 8910 6860
rect 9033 6851 9091 6857
rect 9033 6848 9045 6851
rect 8904 6820 9045 6848
rect 8904 6808 8910 6820
rect 9033 6817 9045 6820
rect 9079 6817 9091 6851
rect 11164 6848 11192 6879
rect 11808 6857 11836 6888
rect 11793 6851 11851 6857
rect 11793 6848 11805 6851
rect 11164 6820 11805 6848
rect 9033 6811 9091 6817
rect 11793 6817 11805 6820
rect 11839 6817 11851 6851
rect 11793 6811 11851 6817
rect 12342 6808 12348 6860
rect 12400 6848 12406 6860
rect 12636 6857 12664 6888
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 14553 6919 14611 6925
rect 14553 6885 14565 6919
rect 14599 6885 14611 6919
rect 15378 6916 15384 6928
rect 15339 6888 15384 6916
rect 14553 6879 14611 6885
rect 12529 6851 12587 6857
rect 12529 6848 12541 6851
rect 12400 6820 12541 6848
rect 12400 6808 12406 6820
rect 12529 6817 12541 6820
rect 12575 6817 12587 6851
rect 12529 6811 12587 6817
rect 12621 6851 12679 6857
rect 12621 6817 12633 6851
rect 12667 6848 12679 6851
rect 13449 6851 13507 6857
rect 13449 6848 13461 6851
rect 12667 6820 13461 6848
rect 12667 6817 12679 6820
rect 12621 6811 12679 6817
rect 13449 6817 13461 6820
rect 13495 6817 13507 6851
rect 13449 6811 13507 6817
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6749 8171 6783
rect 8113 6743 8171 6749
rect 9309 6783 9367 6789
rect 9309 6749 9321 6783
rect 9355 6780 9367 6783
rect 9674 6780 9680 6792
rect 9355 6752 9680 6780
rect 9355 6749 9367 6752
rect 9309 6743 9367 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9769 6783 9827 6789
rect 9769 6749 9781 6783
rect 9815 6780 9827 6783
rect 9858 6780 9864 6792
rect 9815 6752 9864 6780
rect 9815 6749 9827 6752
rect 9769 6743 9827 6749
rect 9858 6740 9864 6752
rect 9916 6740 9922 6792
rect 13265 6783 13323 6789
rect 13265 6749 13277 6783
rect 13311 6780 13323 6783
rect 13354 6780 13360 6792
rect 13311 6752 13360 6780
rect 13311 6749 13323 6752
rect 13265 6743 13323 6749
rect 13354 6740 13360 6752
rect 13412 6740 13418 6792
rect 14185 6783 14243 6789
rect 14185 6749 14197 6783
rect 14231 6780 14243 6783
rect 14274 6780 14280 6792
rect 14231 6752 14280 6780
rect 14231 6749 14243 6752
rect 14185 6743 14243 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 14568 6780 14596 6879
rect 15378 6876 15384 6888
rect 15436 6876 15442 6928
rect 14384 6752 14596 6780
rect 14737 6783 14795 6789
rect 8294 6712 8300 6724
rect 7668 6684 8300 6712
rect 7377 6675 7435 6681
rect 6089 6647 6147 6653
rect 5684 6616 5729 6644
rect 5684 6604 5690 6616
rect 6089 6613 6101 6647
rect 6135 6613 6147 6647
rect 7006 6644 7012 6656
rect 6967 6616 7012 6644
rect 6089 6607 6147 6613
rect 7006 6604 7012 6616
rect 7064 6604 7070 6656
rect 7392 6644 7420 6675
rect 8294 6672 8300 6684
rect 8352 6672 8358 6724
rect 8757 6715 8815 6721
rect 8757 6681 8769 6715
rect 8803 6712 8815 6715
rect 10014 6715 10072 6721
rect 10014 6712 10026 6715
rect 8803 6684 10026 6712
rect 8803 6681 8815 6684
rect 8757 6675 8815 6681
rect 10014 6681 10026 6684
rect 10060 6681 10072 6715
rect 12250 6712 12256 6724
rect 10014 6675 10072 6681
rect 10704 6684 11744 6712
rect 7926 6644 7932 6656
rect 7392 6616 7932 6644
rect 7926 6604 7932 6616
rect 7984 6604 7990 6656
rect 9217 6647 9275 6653
rect 9217 6613 9229 6647
rect 9263 6644 9275 6647
rect 9582 6644 9588 6656
rect 9263 6616 9588 6644
rect 9263 6613 9275 6616
rect 9217 6607 9275 6613
rect 9582 6604 9588 6616
rect 9640 6604 9646 6656
rect 9677 6647 9735 6653
rect 9677 6613 9689 6647
rect 9723 6644 9735 6647
rect 10704 6644 10732 6684
rect 11606 6644 11612 6656
rect 9723 6616 10732 6644
rect 11567 6616 11612 6644
rect 9723 6613 9735 6616
rect 9677 6607 9735 6613
rect 11606 6604 11612 6616
rect 11664 6604 11670 6656
rect 11716 6653 11744 6684
rect 12084 6684 12256 6712
rect 12084 6653 12112 6684
rect 12250 6672 12256 6684
rect 12308 6672 12314 6724
rect 13630 6672 13636 6724
rect 13688 6712 13694 6724
rect 14384 6712 14412 6752
rect 14737 6749 14749 6783
rect 14783 6780 14795 6783
rect 15470 6780 15476 6792
rect 14783 6752 15476 6780
rect 14783 6749 14795 6752
rect 14737 6743 14795 6749
rect 15470 6740 15476 6752
rect 15528 6740 15534 6792
rect 13688 6684 14412 6712
rect 13688 6672 13694 6684
rect 14550 6672 14556 6724
rect 14608 6712 14614 6724
rect 15013 6715 15071 6721
rect 15013 6712 15025 6715
rect 14608 6684 15025 6712
rect 14608 6672 14614 6684
rect 15013 6681 15025 6684
rect 15059 6681 15071 6715
rect 15194 6712 15200 6724
rect 15155 6684 15200 6712
rect 15013 6675 15071 6681
rect 15194 6672 15200 6684
rect 15252 6672 15258 6724
rect 15562 6712 15568 6724
rect 15475 6684 15568 6712
rect 15562 6672 15568 6684
rect 15620 6712 15626 6724
rect 16114 6712 16120 6724
rect 15620 6684 16120 6712
rect 15620 6672 15626 6684
rect 16114 6672 16120 6684
rect 16172 6672 16178 6724
rect 11701 6647 11759 6653
rect 11701 6613 11713 6647
rect 11747 6613 11759 6647
rect 11701 6607 11759 6613
rect 12069 6647 12127 6653
rect 12069 6613 12081 6647
rect 12115 6613 12127 6647
rect 12069 6607 12127 6613
rect 12437 6647 12495 6653
rect 12437 6613 12449 6647
rect 12483 6644 12495 6647
rect 12710 6644 12716 6656
rect 12483 6616 12716 6644
rect 12483 6613 12495 6616
rect 12437 6607 12495 6613
rect 12710 6604 12716 6616
rect 12768 6604 12774 6656
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13354 6644 13360 6656
rect 13228 6616 13360 6644
rect 13228 6604 13234 6616
rect 13354 6604 13360 6616
rect 13412 6644 13418 6656
rect 13725 6647 13783 6653
rect 13725 6644 13737 6647
rect 13412 6616 13737 6644
rect 13412 6604 13418 6616
rect 13725 6613 13737 6616
rect 13771 6613 13783 6647
rect 13725 6607 13783 6613
rect 14369 6647 14427 6653
rect 14369 6613 14381 6647
rect 14415 6644 14427 6647
rect 15378 6644 15384 6656
rect 14415 6616 15384 6644
rect 14415 6613 14427 6616
rect 14369 6607 14427 6613
rect 15378 6604 15384 6616
rect 15436 6604 15442 6656
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 1670 6400 1676 6452
rect 1728 6440 1734 6452
rect 2041 6443 2099 6449
rect 2041 6440 2053 6443
rect 1728 6412 2053 6440
rect 1728 6400 1734 6412
rect 2041 6409 2053 6412
rect 2087 6440 2099 6443
rect 4249 6443 4307 6449
rect 2087 6412 3556 6440
rect 2087 6409 2099 6412
rect 2041 6403 2099 6409
rect 3418 6372 3424 6384
rect 1688 6344 3424 6372
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1688 6313 1716 6344
rect 3418 6332 3424 6344
rect 3476 6332 3482 6384
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6304 1823 6307
rect 2406 6304 2412 6316
rect 1811 6276 2412 6304
rect 1811 6273 1823 6276
rect 1765 6267 1823 6273
rect 1504 6236 1532 6264
rect 1780 6236 1808 6267
rect 2406 6264 2412 6276
rect 2464 6264 2470 6316
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 3154 6307 3212 6313
rect 3154 6304 3166 6307
rect 2740 6276 3166 6304
rect 2740 6264 2746 6276
rect 3154 6273 3166 6276
rect 3200 6273 3212 6307
rect 3154 6267 3212 6273
rect 3418 6236 3424 6248
rect 1504 6208 1808 6236
rect 3379 6208 3424 6236
rect 3418 6196 3424 6208
rect 3476 6196 3482 6248
rect 3528 6236 3556 6412
rect 4249 6409 4261 6443
rect 4295 6440 4307 6443
rect 4617 6443 4675 6449
rect 4617 6440 4629 6443
rect 4295 6412 4629 6440
rect 4295 6409 4307 6412
rect 4249 6403 4307 6409
rect 4617 6409 4629 6412
rect 4663 6409 4675 6443
rect 4617 6403 4675 6409
rect 4985 6443 5043 6449
rect 4985 6409 4997 6443
rect 5031 6440 5043 6443
rect 5074 6440 5080 6452
rect 5031 6412 5080 6440
rect 5031 6409 5043 6412
rect 4985 6403 5043 6409
rect 5074 6400 5080 6412
rect 5132 6440 5138 6452
rect 7926 6440 7932 6452
rect 5132 6412 7932 6440
rect 5132 6400 5138 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8573 6443 8631 6449
rect 8573 6409 8585 6443
rect 8619 6440 8631 6443
rect 8846 6440 8852 6452
rect 8619 6412 8852 6440
rect 8619 6409 8631 6412
rect 8573 6403 8631 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 9582 6400 9588 6452
rect 9640 6440 9646 6452
rect 10042 6440 10048 6452
rect 9640 6412 10048 6440
rect 9640 6400 9646 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10870 6400 10876 6452
rect 10928 6400 10934 6452
rect 11054 6400 11060 6452
rect 11112 6440 11118 6452
rect 11149 6443 11207 6449
rect 11149 6440 11161 6443
rect 11112 6412 11161 6440
rect 11112 6400 11118 6412
rect 11149 6409 11161 6412
rect 11195 6409 11207 6443
rect 11149 6403 11207 6409
rect 11606 6400 11612 6452
rect 11664 6440 11670 6452
rect 11701 6443 11759 6449
rect 11701 6440 11713 6443
rect 11664 6412 11713 6440
rect 11664 6400 11670 6412
rect 11701 6409 11713 6412
rect 11747 6409 11759 6443
rect 11882 6440 11888 6452
rect 11843 6412 11888 6440
rect 11701 6403 11759 6409
rect 11882 6400 11888 6412
rect 11940 6400 11946 6452
rect 12253 6443 12311 6449
rect 12253 6409 12265 6443
rect 12299 6409 12311 6443
rect 12253 6403 12311 6409
rect 7742 6372 7748 6384
rect 5736 6344 7748 6372
rect 3697 6307 3755 6313
rect 3697 6273 3709 6307
rect 3743 6304 3755 6307
rect 3786 6304 3792 6316
rect 3743 6276 3792 6304
rect 3743 6273 3755 6276
rect 3697 6267 3755 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 4157 6307 4215 6313
rect 4157 6273 4169 6307
rect 4203 6304 4215 6307
rect 4203 6276 5304 6304
rect 4203 6273 4215 6276
rect 4157 6267 4215 6273
rect 4341 6239 4399 6245
rect 4341 6236 4353 6239
rect 3528 6208 4353 6236
rect 4341 6205 4353 6208
rect 4387 6205 4399 6239
rect 4341 6199 4399 6205
rect 4522 6196 4528 6248
rect 4580 6236 4586 6248
rect 5077 6239 5135 6245
rect 5077 6236 5089 6239
rect 4580 6208 5089 6236
rect 4580 6196 4586 6208
rect 5077 6205 5089 6208
rect 5123 6205 5135 6239
rect 5077 6199 5135 6205
rect 5169 6239 5227 6245
rect 5169 6205 5181 6239
rect 5215 6205 5227 6239
rect 5276 6236 5304 6276
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5736 6304 5764 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 8144 6375 8202 6381
rect 8144 6341 8156 6375
rect 8190 6372 8202 6375
rect 8294 6372 8300 6384
rect 8190 6344 8300 6372
rect 8190 6341 8202 6344
rect 8144 6335 8202 6341
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 9708 6375 9766 6381
rect 9708 6341 9720 6375
rect 9754 6372 9766 6375
rect 10888 6372 10916 6400
rect 9754 6344 10916 6372
rect 12268 6372 12296 6403
rect 12710 6400 12716 6452
rect 12768 6440 12774 6452
rect 13170 6440 13176 6452
rect 12768 6412 13176 6440
rect 12768 6400 12774 6412
rect 13170 6400 13176 6412
rect 13228 6400 13234 6452
rect 14274 6440 14280 6452
rect 14235 6412 14280 6440
rect 14274 6400 14280 6412
rect 14332 6400 14338 6452
rect 14461 6443 14519 6449
rect 14461 6409 14473 6443
rect 14507 6409 14519 6443
rect 14461 6403 14519 6409
rect 12434 6372 12440 6384
rect 12268 6344 12440 6372
rect 9754 6341 9766 6344
rect 9708 6335 9766 6341
rect 12434 6332 12440 6344
rect 12492 6372 12498 6384
rect 12618 6372 12624 6384
rect 12492 6344 12624 6372
rect 12492 6332 12498 6344
rect 12618 6332 12624 6344
rect 12676 6332 12682 6384
rect 12894 6332 12900 6384
rect 12952 6332 12958 6384
rect 12986 6332 12992 6384
rect 13044 6372 13050 6384
rect 13081 6375 13139 6381
rect 13081 6372 13093 6375
rect 13044 6344 13093 6372
rect 13044 6332 13050 6344
rect 13081 6341 13093 6344
rect 13127 6372 13139 6375
rect 13722 6372 13728 6384
rect 13127 6344 13728 6372
rect 13127 6341 13139 6344
rect 13081 6335 13139 6341
rect 13722 6332 13728 6344
rect 13780 6332 13786 6384
rect 13909 6375 13967 6381
rect 13909 6341 13921 6375
rect 13955 6372 13967 6375
rect 14476 6372 14504 6403
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 15286 6440 15292 6452
rect 14608 6412 15292 6440
rect 14608 6400 14614 6412
rect 15286 6400 15292 6412
rect 15344 6400 15350 6452
rect 15470 6372 15476 6384
rect 13955 6344 14504 6372
rect 14660 6344 15476 6372
rect 13955 6341 13967 6344
rect 13909 6335 13967 6341
rect 5408 6276 5764 6304
rect 5813 6307 5871 6313
rect 5408 6264 5414 6276
rect 5813 6273 5825 6307
rect 5859 6304 5871 6307
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 5859 6276 6377 6304
rect 5859 6273 5871 6276
rect 5813 6267 5871 6273
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 7760 6304 7788 6332
rect 7760 6276 9904 6304
rect 6365 6267 6423 6273
rect 5905 6239 5963 6245
rect 5276 6208 5488 6236
rect 5169 6199 5227 6205
rect 1486 6168 1492 6180
rect 1447 6140 1492 6168
rect 1486 6128 1492 6140
rect 1544 6128 1550 6180
rect 3970 6128 3976 6180
rect 4028 6168 4034 6180
rect 4982 6168 4988 6180
rect 4028 6140 4988 6168
rect 4028 6128 4034 6140
rect 4982 6128 4988 6140
rect 5040 6168 5046 6180
rect 5184 6168 5212 6199
rect 5460 6177 5488 6208
rect 5905 6205 5917 6239
rect 5951 6236 5963 6239
rect 5994 6236 6000 6248
rect 5951 6208 6000 6236
rect 5951 6205 5963 6208
rect 5905 6199 5963 6205
rect 5994 6196 6000 6208
rect 6052 6196 6058 6248
rect 6089 6239 6147 6245
rect 6089 6205 6101 6239
rect 6135 6236 6147 6239
rect 6178 6236 6184 6248
rect 6135 6208 6184 6236
rect 6135 6205 6147 6208
rect 6089 6199 6147 6205
rect 6178 6196 6184 6208
rect 6236 6196 6242 6248
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7374 6236 7380 6248
rect 6963 6208 7380 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7374 6196 7380 6208
rect 7432 6196 7438 6248
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6205 8447 6239
rect 9876 6236 9904 6276
rect 9950 6264 9956 6316
rect 10008 6304 10014 6316
rect 10962 6304 10968 6316
rect 10008 6276 10968 6304
rect 10008 6264 10014 6276
rect 10962 6264 10968 6276
rect 11020 6264 11026 6316
rect 11517 6307 11575 6313
rect 11517 6273 11529 6307
rect 11563 6273 11575 6307
rect 12342 6304 12348 6316
rect 12303 6276 12348 6304
rect 11517 6267 11575 6273
rect 9876 6208 9996 6236
rect 8389 6199 8447 6205
rect 5040 6140 5212 6168
rect 5445 6171 5503 6177
rect 5040 6128 5046 6140
rect 5445 6137 5457 6171
rect 5491 6137 5503 6171
rect 5445 6131 5503 6137
rect 1949 6103 2007 6109
rect 1949 6069 1961 6103
rect 1995 6100 2007 6103
rect 2222 6100 2228 6112
rect 1995 6072 2228 6100
rect 1995 6069 2007 6072
rect 1949 6063 2007 6069
rect 2222 6060 2228 6072
rect 2280 6060 2286 6112
rect 3513 6103 3571 6109
rect 3513 6069 3525 6103
rect 3559 6100 3571 6103
rect 3602 6100 3608 6112
rect 3559 6072 3608 6100
rect 3559 6069 3571 6072
rect 3513 6063 3571 6069
rect 3602 6060 3608 6072
rect 3660 6060 3666 6112
rect 3786 6100 3792 6112
rect 3747 6072 3792 6100
rect 3786 6060 3792 6072
rect 3844 6060 3850 6112
rect 6178 6060 6184 6112
rect 6236 6100 6242 6112
rect 7009 6103 7067 6109
rect 7009 6100 7021 6103
rect 6236 6072 7021 6100
rect 6236 6060 6242 6072
rect 7009 6069 7021 6072
rect 7055 6069 7067 6103
rect 8404 6100 8432 6199
rect 9968 6168 9996 6208
rect 10042 6196 10048 6248
rect 10100 6236 10106 6248
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 10100 6208 10241 6236
rect 10100 6196 10106 6208
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 10505 6239 10563 6245
rect 10505 6205 10517 6239
rect 10551 6205 10563 6239
rect 10505 6199 10563 6205
rect 10520 6168 10548 6199
rect 10778 6196 10784 6248
rect 10836 6236 10842 6248
rect 11532 6236 11560 6267
rect 12342 6264 12348 6276
rect 12400 6264 12406 6316
rect 12912 6304 12940 6332
rect 12912 6276 13032 6304
rect 12526 6236 12532 6248
rect 10836 6208 11560 6236
rect 12487 6208 12532 6236
rect 10836 6196 10842 6208
rect 12526 6196 12532 6208
rect 12584 6196 12590 6248
rect 12894 6236 12900 6248
rect 12855 6208 12900 6236
rect 12894 6196 12900 6208
rect 12952 6196 12958 6248
rect 13004 6245 13032 6276
rect 13464 6276 14044 6304
rect 12989 6239 13047 6245
rect 12989 6205 13001 6239
rect 13035 6205 13047 6239
rect 12989 6199 13047 6205
rect 12618 6168 12624 6180
rect 9968 6140 12624 6168
rect 12618 6128 12624 6140
rect 12676 6128 12682 6180
rect 13464 6177 13492 6276
rect 13725 6239 13783 6245
rect 13725 6205 13737 6239
rect 13771 6205 13783 6239
rect 13725 6199 13783 6205
rect 13449 6171 13507 6177
rect 13449 6137 13461 6171
rect 13495 6137 13507 6171
rect 13740 6168 13768 6199
rect 13814 6196 13820 6248
rect 13872 6236 13878 6248
rect 13872 6208 13917 6236
rect 13872 6196 13878 6208
rect 14016 6168 14044 6276
rect 14660 6168 14688 6344
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 14826 6304 14832 6316
rect 14787 6276 14832 6304
rect 14826 6264 14832 6276
rect 14884 6264 14890 6316
rect 15378 6304 15384 6316
rect 15339 6276 15384 6304
rect 15378 6264 15384 6276
rect 15436 6264 15442 6316
rect 14918 6236 14924 6248
rect 14879 6208 14924 6236
rect 14918 6196 14924 6208
rect 14976 6196 14982 6248
rect 15013 6239 15071 6245
rect 15013 6205 15025 6239
rect 15059 6205 15071 6239
rect 15013 6199 15071 6205
rect 13740 6140 13860 6168
rect 14016 6140 14688 6168
rect 13449 6131 13507 6137
rect 13832 6112 13860 6140
rect 9766 6100 9772 6112
rect 8404 6072 9772 6100
rect 7009 6063 7067 6069
rect 9766 6060 9772 6072
rect 9824 6060 9830 6112
rect 10042 6100 10048 6112
rect 10003 6072 10048 6100
rect 10042 6060 10048 6072
rect 10100 6060 10106 6112
rect 13814 6060 13820 6112
rect 13872 6060 13878 6112
rect 14458 6060 14464 6112
rect 14516 6100 14522 6112
rect 15028 6100 15056 6199
rect 15562 6100 15568 6112
rect 14516 6072 15056 6100
rect 15523 6072 15568 6100
rect 14516 6060 14522 6072
rect 15562 6060 15568 6072
rect 15620 6060 15626 6112
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 3881 5899 3939 5905
rect 3881 5865 3893 5899
rect 3927 5896 3939 5899
rect 4154 5896 4160 5908
rect 3927 5868 4160 5896
rect 3927 5865 3939 5868
rect 3881 5859 3939 5865
rect 4154 5856 4160 5868
rect 4212 5896 4218 5908
rect 4212 5868 5856 5896
rect 4212 5856 4218 5868
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5797 2835 5831
rect 2777 5791 2835 5797
rect 2869 5831 2927 5837
rect 2869 5797 2881 5831
rect 2915 5828 2927 5831
rect 3142 5828 3148 5840
rect 2915 5800 3148 5828
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 2792 5760 2820 5791
rect 3142 5788 3148 5800
rect 3200 5788 3206 5840
rect 5828 5828 5856 5868
rect 5902 5856 5908 5908
rect 5960 5896 5966 5908
rect 5960 5868 8892 5896
rect 5960 5856 5966 5868
rect 5994 5828 6000 5840
rect 5828 5800 6000 5828
rect 5994 5788 6000 5800
rect 6052 5828 6058 5840
rect 6052 5800 6408 5828
rect 6052 5788 6058 5800
rect 3510 5760 3516 5772
rect 2792 5732 3516 5760
rect 3510 5720 3516 5732
rect 3568 5720 3574 5772
rect 6178 5720 6184 5772
rect 6236 5760 6242 5772
rect 6273 5763 6331 5769
rect 6273 5760 6285 5763
rect 6236 5732 6285 5760
rect 6236 5720 6242 5732
rect 6273 5729 6285 5732
rect 6319 5729 6331 5763
rect 6380 5760 6408 5800
rect 6454 5788 6460 5840
rect 6512 5828 6518 5840
rect 6917 5831 6975 5837
rect 6917 5828 6929 5831
rect 6512 5800 6929 5828
rect 6512 5788 6518 5800
rect 6917 5797 6929 5800
rect 6963 5797 6975 5831
rect 6917 5791 6975 5797
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8864 5828 8892 5868
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 9214 5896 9220 5908
rect 8996 5868 9041 5896
rect 9175 5868 9220 5896
rect 8996 5856 9002 5868
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 9306 5856 9312 5908
rect 9364 5896 9370 5908
rect 9582 5896 9588 5908
rect 9364 5868 9588 5896
rect 9364 5856 9370 5868
rect 9582 5856 9588 5868
rect 9640 5856 9646 5908
rect 10134 5896 10140 5908
rect 9876 5868 10140 5896
rect 9876 5840 9904 5868
rect 10134 5856 10140 5868
rect 10192 5856 10198 5908
rect 10962 5856 10968 5908
rect 11020 5896 11026 5908
rect 11330 5896 11336 5908
rect 11020 5868 11336 5896
rect 11020 5856 11026 5868
rect 11330 5856 11336 5868
rect 11388 5896 11394 5908
rect 11701 5899 11759 5905
rect 11701 5896 11713 5899
rect 11388 5868 11713 5896
rect 11388 5856 11394 5868
rect 11701 5865 11713 5868
rect 11747 5865 11759 5899
rect 13538 5896 13544 5908
rect 11701 5859 11759 5865
rect 13096 5868 13544 5896
rect 9858 5828 9864 5840
rect 7524 5800 8800 5828
rect 8864 5800 9864 5828
rect 7524 5788 7530 5800
rect 7653 5763 7711 5769
rect 6380 5732 7512 5760
rect 6273 5723 6331 5729
rect 1397 5695 1455 5701
rect 1397 5661 1409 5695
rect 1443 5692 1455 5695
rect 3050 5692 3056 5704
rect 1443 5664 3056 5692
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3237 5695 3295 5701
rect 3237 5661 3249 5695
rect 3283 5692 3295 5695
rect 3786 5692 3792 5704
rect 3283 5664 3792 5692
rect 3283 5661 3295 5664
rect 3237 5655 3295 5661
rect 3786 5652 3792 5664
rect 3844 5652 3850 5704
rect 5353 5695 5411 5701
rect 5353 5661 5365 5695
rect 5399 5692 5411 5695
rect 5626 5692 5632 5704
rect 5399 5664 5632 5692
rect 5399 5661 5411 5664
rect 5353 5655 5411 5661
rect 5626 5652 5632 5664
rect 5684 5652 5690 5704
rect 6089 5695 6147 5701
rect 6089 5661 6101 5695
rect 6135 5692 6147 5695
rect 6457 5695 6515 5701
rect 6135 5664 6316 5692
rect 6135 5661 6147 5664
rect 6089 5655 6147 5661
rect 6288 5636 6316 5664
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 7006 5692 7012 5704
rect 6503 5664 7012 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 7006 5652 7012 5664
rect 7064 5652 7070 5704
rect 7374 5692 7380 5704
rect 7335 5664 7380 5692
rect 7374 5652 7380 5664
rect 7432 5652 7438 5704
rect 7484 5701 7512 5732
rect 7653 5729 7665 5763
rect 7699 5760 7711 5763
rect 8294 5760 8300 5772
rect 7699 5732 8300 5760
rect 7699 5729 7711 5732
rect 7653 5723 7711 5729
rect 8294 5720 8300 5732
rect 8352 5760 8358 5772
rect 8389 5763 8447 5769
rect 8389 5760 8401 5763
rect 8352 5732 8401 5760
rect 8352 5720 8358 5732
rect 8389 5729 8401 5732
rect 8435 5729 8447 5763
rect 8662 5760 8668 5772
rect 8623 5732 8668 5760
rect 8389 5723 8447 5729
rect 8662 5720 8668 5732
rect 8720 5720 8726 5772
rect 8772 5760 8800 5800
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 10134 5760 10140 5772
rect 8772 5732 9444 5760
rect 10095 5732 10140 5760
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5692 7527 5695
rect 7558 5692 7564 5704
rect 7515 5664 7564 5692
rect 7515 5661 7527 5664
rect 7469 5655 7527 5661
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8202 5652 8208 5704
rect 8260 5652 8266 5704
rect 8680 5692 8708 5720
rect 9416 5701 9444 5732
rect 10134 5720 10140 5732
rect 10192 5720 10198 5772
rect 12802 5760 12808 5772
rect 12763 5732 12808 5760
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 9401 5695 9459 5701
rect 8680 5688 8993 5692
rect 8680 5668 9076 5688
rect 9125 5671 9183 5677
rect 9125 5668 9137 5671
rect 8680 5664 9137 5668
rect 8965 5660 9137 5664
rect 1670 5633 1676 5636
rect 1664 5624 1676 5633
rect 1631 5596 1676 5624
rect 1664 5587 1676 5596
rect 1670 5584 1676 5587
rect 1728 5584 1734 5636
rect 3326 5624 3332 5636
rect 3287 5596 3332 5624
rect 3326 5584 3332 5596
rect 3384 5584 3390 5636
rect 5074 5624 5080 5636
rect 5132 5633 5138 5636
rect 5044 5596 5080 5624
rect 5074 5584 5080 5596
rect 5132 5587 5144 5633
rect 5132 5584 5138 5587
rect 6270 5584 6276 5636
rect 6328 5584 6334 5636
rect 6549 5627 6607 5633
rect 6549 5593 6561 5627
rect 6595 5624 6607 5627
rect 8220 5624 8248 5652
rect 9048 5640 9137 5660
rect 9125 5637 9137 5640
rect 9171 5637 9183 5671
rect 9401 5661 9413 5695
rect 9447 5661 9459 5695
rect 10042 5692 10048 5704
rect 9401 5655 9459 5661
rect 9968 5664 10048 5692
rect 8297 5627 8355 5633
rect 9125 5631 9183 5637
rect 8297 5624 8309 5627
rect 6595 5596 7052 5624
rect 8220 5596 8309 5624
rect 6595 5593 6607 5596
rect 6549 5587 6607 5593
rect 2682 5516 2688 5568
rect 2740 5556 2746 5568
rect 3970 5556 3976 5568
rect 2740 5528 3976 5556
rect 2740 5516 2746 5528
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 5445 5559 5503 5565
rect 5445 5525 5457 5559
rect 5491 5556 5503 5559
rect 5994 5556 6000 5568
rect 5491 5528 6000 5556
rect 5491 5525 5503 5528
rect 5445 5519 5503 5525
rect 5994 5516 6000 5528
rect 6052 5516 6058 5568
rect 7024 5565 7052 5596
rect 8297 5593 8309 5596
rect 8343 5593 8355 5627
rect 9968 5624 9996 5664
rect 10042 5652 10048 5664
rect 10100 5692 10106 5704
rect 11698 5692 11704 5704
rect 10100 5664 11704 5692
rect 10100 5652 10106 5664
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 12618 5692 12624 5704
rect 12579 5664 12624 5692
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 8297 5587 8355 5593
rect 8680 5596 8993 5624
rect 7009 5559 7067 5565
rect 7009 5525 7021 5559
rect 7055 5525 7067 5559
rect 7834 5556 7840 5568
rect 7795 5528 7840 5556
rect 7009 5519 7067 5525
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 8110 5516 8116 5568
rect 8168 5556 8174 5568
rect 8205 5559 8263 5565
rect 8205 5556 8217 5559
rect 8168 5528 8217 5556
rect 8168 5516 8174 5528
rect 8205 5525 8217 5528
rect 8251 5556 8263 5559
rect 8680 5556 8708 5596
rect 8251 5528 8708 5556
rect 8965 5556 8993 5596
rect 9232 5596 9996 5624
rect 9232 5556 9260 5596
rect 10226 5584 10232 5636
rect 10284 5624 10290 5636
rect 10413 5627 10471 5633
rect 10413 5624 10425 5627
rect 10284 5596 10425 5624
rect 10284 5584 10290 5596
rect 10413 5593 10425 5596
rect 10459 5593 10471 5627
rect 10413 5587 10471 5593
rect 8965 5528 9260 5556
rect 8251 5525 8263 5528
rect 8205 5519 8263 5525
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 9585 5559 9643 5565
rect 9585 5556 9597 5559
rect 9364 5528 9597 5556
rect 9364 5516 9370 5528
rect 9585 5525 9597 5528
rect 9631 5525 9643 5559
rect 9950 5556 9956 5568
rect 9911 5528 9956 5556
rect 9585 5519 9643 5525
rect 9950 5516 9956 5528
rect 10008 5516 10014 5568
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 12253 5559 12311 5565
rect 12253 5556 12265 5559
rect 10091 5528 12265 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 12253 5525 12265 5528
rect 12299 5525 12311 5559
rect 12710 5556 12716 5568
rect 12671 5528 12716 5556
rect 12253 5519 12311 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 12986 5516 12992 5568
rect 13044 5556 13050 5568
rect 13096 5556 13124 5868
rect 13538 5856 13544 5868
rect 13596 5856 13602 5908
rect 14829 5899 14887 5905
rect 14829 5865 14841 5899
rect 14875 5896 14887 5899
rect 14918 5896 14924 5908
rect 14875 5868 14924 5896
rect 14875 5865 14887 5868
rect 14829 5859 14887 5865
rect 14918 5856 14924 5868
rect 14976 5856 14982 5908
rect 13817 5831 13875 5837
rect 13817 5797 13829 5831
rect 13863 5828 13875 5831
rect 15378 5828 15384 5840
rect 13863 5800 15384 5828
rect 13863 5797 13875 5800
rect 13817 5791 13875 5797
rect 15378 5788 15384 5800
rect 15436 5788 15442 5840
rect 13265 5763 13323 5769
rect 13265 5729 13277 5763
rect 13311 5760 13323 5763
rect 13538 5760 13544 5772
rect 13311 5732 13544 5760
rect 13311 5729 13323 5732
rect 13265 5723 13323 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 14277 5763 14335 5769
rect 14277 5729 14289 5763
rect 14323 5760 14335 5763
rect 15473 5763 15531 5769
rect 15473 5760 15485 5763
rect 14323 5732 15485 5760
rect 14323 5729 14335 5732
rect 14277 5723 14335 5729
rect 15473 5729 15485 5732
rect 15519 5760 15531 5763
rect 15562 5760 15568 5772
rect 15519 5732 15568 5760
rect 15519 5729 15531 5732
rect 15473 5723 15531 5729
rect 15562 5720 15568 5732
rect 15620 5720 15626 5772
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 15286 5692 15292 5704
rect 14507 5664 15292 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 15286 5652 15292 5664
rect 15344 5652 15350 5704
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5692 15439 5695
rect 16482 5692 16488 5704
rect 15427 5664 16488 5692
rect 15427 5661 15439 5664
rect 15381 5655 15439 5661
rect 16482 5652 16488 5664
rect 16540 5652 16546 5704
rect 13449 5627 13507 5633
rect 13449 5593 13461 5627
rect 13495 5624 13507 5627
rect 13906 5624 13912 5636
rect 13495 5596 13912 5624
rect 13495 5593 13507 5596
rect 13449 5587 13507 5593
rect 13906 5584 13912 5596
rect 13964 5584 13970 5636
rect 13357 5559 13415 5565
rect 13357 5556 13369 5559
rect 13044 5528 13369 5556
rect 13044 5516 13050 5528
rect 13357 5525 13369 5528
rect 13403 5525 13415 5559
rect 13357 5519 13415 5525
rect 14274 5516 14280 5568
rect 14332 5556 14338 5568
rect 14369 5559 14427 5565
rect 14369 5556 14381 5559
rect 14332 5528 14381 5556
rect 14332 5516 14338 5528
rect 14369 5525 14381 5528
rect 14415 5525 14427 5559
rect 14369 5519 14427 5525
rect 14826 5516 14832 5568
rect 14884 5556 14890 5568
rect 14921 5559 14979 5565
rect 14921 5556 14933 5559
rect 14884 5528 14933 5556
rect 14884 5516 14890 5528
rect 14921 5525 14933 5528
rect 14967 5525 14979 5559
rect 15286 5556 15292 5568
rect 15247 5528 15292 5556
rect 14921 5519 14979 5525
rect 15286 5516 15292 5528
rect 15344 5516 15350 5568
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 1486 5352 1492 5364
rect 1447 5324 1492 5352
rect 1486 5312 1492 5324
rect 1544 5312 1550 5364
rect 1762 5352 1768 5364
rect 1723 5324 1768 5352
rect 1762 5312 1768 5324
rect 1820 5312 1826 5364
rect 2130 5312 2136 5364
rect 2188 5312 2194 5364
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 2866 5352 2872 5364
rect 2280 5324 2872 5352
rect 2280 5312 2286 5324
rect 2866 5312 2872 5324
rect 2924 5312 2930 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3418 5352 3424 5364
rect 3108 5324 3424 5352
rect 3108 5312 3114 5324
rect 3418 5312 3424 5324
rect 3476 5352 3482 5364
rect 3476 5324 3832 5352
rect 3476 5312 3482 5324
rect 2148 5284 2176 5312
rect 3804 5296 3832 5324
rect 5810 5312 5816 5364
rect 5868 5352 5874 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5868 5324 6469 5352
rect 5868 5312 5874 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7101 5355 7159 5361
rect 7101 5321 7113 5355
rect 7147 5352 7159 5355
rect 7834 5352 7840 5364
rect 7147 5324 7840 5352
rect 7147 5321 7159 5324
rect 7101 5315 7159 5321
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 7929 5355 7987 5361
rect 7929 5321 7941 5355
rect 7975 5352 7987 5355
rect 8018 5352 8024 5364
rect 7975 5324 8024 5352
rect 7975 5321 7987 5324
rect 7929 5315 7987 5321
rect 8018 5312 8024 5324
rect 8076 5312 8082 5364
rect 8294 5312 8300 5364
rect 8352 5352 8358 5364
rect 8389 5355 8447 5361
rect 8389 5352 8401 5355
rect 8352 5324 8401 5352
rect 8352 5312 8358 5324
rect 8389 5321 8401 5324
rect 8435 5321 8447 5355
rect 8389 5315 8447 5321
rect 9953 5355 10011 5361
rect 9953 5321 9965 5355
rect 9999 5352 10011 5355
rect 10134 5352 10140 5364
rect 9999 5324 10140 5352
rect 9999 5321 10011 5324
rect 9953 5315 10011 5321
rect 10134 5312 10140 5324
rect 10192 5352 10198 5364
rect 10962 5352 10968 5364
rect 10192 5324 10968 5352
rect 10192 5312 10198 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11517 5355 11575 5361
rect 11517 5321 11529 5355
rect 11563 5321 11575 5355
rect 11517 5315 11575 5321
rect 1688 5256 2176 5284
rect 1688 5225 1716 5256
rect 2498 5244 2504 5296
rect 2556 5284 2562 5296
rect 3142 5284 3148 5296
rect 2556 5256 3148 5284
rect 2556 5244 2562 5256
rect 3142 5244 3148 5256
rect 3200 5244 3206 5296
rect 3786 5244 3792 5296
rect 3844 5284 3850 5296
rect 5626 5284 5632 5296
rect 3844 5256 5632 5284
rect 3844 5244 3850 5256
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5185 1731 5219
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 1673 5179 1731 5185
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 2774 5176 2780 5228
rect 2832 5216 2838 5228
rect 3878 5216 3884 5228
rect 2832 5188 3884 5216
rect 2832 5176 2838 5188
rect 3878 5176 3884 5188
rect 3936 5176 3942 5228
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4154 5216 4160 5228
rect 4028 5188 4160 5216
rect 4028 5176 4034 5188
rect 4154 5176 4160 5188
rect 4212 5176 4218 5228
rect 4338 5216 4344 5228
rect 4299 5188 4344 5216
rect 4338 5176 4344 5188
rect 4396 5176 4402 5228
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4816 5225 4844 5256
rect 5626 5244 5632 5256
rect 5684 5244 5690 5296
rect 6196 5256 7328 5284
rect 6196 5228 6224 5256
rect 4801 5219 4859 5225
rect 4488 5188 4533 5216
rect 4488 5176 4494 5188
rect 4801 5185 4813 5219
rect 4847 5185 4859 5219
rect 4801 5179 4859 5185
rect 5068 5219 5126 5225
rect 5068 5185 5080 5219
rect 5114 5216 5126 5219
rect 6178 5216 6184 5228
rect 5114 5188 6184 5216
rect 5114 5185 5126 5188
rect 5068 5179 5126 5185
rect 6178 5176 6184 5188
rect 6236 5176 6242 5228
rect 6362 5176 6368 5228
rect 6420 5216 6426 5228
rect 6641 5219 6699 5225
rect 6641 5216 6653 5219
rect 6420 5188 6653 5216
rect 6420 5176 6426 5188
rect 6641 5185 6653 5188
rect 6687 5185 6699 5219
rect 6641 5179 6699 5185
rect 2222 5148 2228 5160
rect 2183 5120 2228 5148
rect 2222 5108 2228 5120
rect 2280 5108 2286 5160
rect 2409 5151 2467 5157
rect 2409 5117 2421 5151
rect 2455 5148 2467 5151
rect 2498 5148 2504 5160
rect 2455 5120 2504 5148
rect 2455 5117 2467 5120
rect 2409 5111 2467 5117
rect 2498 5108 2504 5120
rect 2556 5148 2562 5160
rect 2682 5148 2688 5160
rect 2556 5120 2688 5148
rect 2556 5108 2562 5120
rect 2682 5108 2688 5120
rect 2740 5108 2746 5160
rect 2866 5108 2872 5160
rect 2924 5148 2930 5160
rect 4522 5148 4528 5160
rect 2924 5120 4528 5148
rect 2924 5108 2930 5120
rect 4522 5108 4528 5120
rect 4580 5108 4586 5160
rect 7190 5148 7196 5160
rect 7151 5120 7196 5148
rect 7190 5108 7196 5120
rect 7248 5108 7254 5160
rect 7300 5157 7328 5256
rect 10686 5244 10692 5296
rect 10744 5284 10750 5296
rect 11088 5287 11146 5293
rect 11088 5284 11100 5287
rect 10744 5256 11100 5284
rect 10744 5244 10750 5256
rect 11088 5253 11100 5256
rect 11134 5284 11146 5287
rect 11532 5284 11560 5315
rect 11974 5312 11980 5364
rect 12032 5352 12038 5364
rect 12989 5355 13047 5361
rect 12989 5352 13001 5355
rect 12032 5324 13001 5352
rect 12032 5312 12038 5324
rect 12989 5321 13001 5324
rect 13035 5321 13047 5355
rect 12989 5315 13047 5321
rect 13170 5312 13176 5364
rect 13228 5352 13234 5364
rect 13449 5355 13507 5361
rect 13449 5352 13461 5355
rect 13228 5324 13461 5352
rect 13228 5312 13234 5324
rect 13449 5321 13461 5324
rect 13495 5321 13507 5355
rect 13449 5315 13507 5321
rect 13906 5312 13912 5364
rect 13964 5352 13970 5364
rect 14369 5355 14427 5361
rect 14369 5352 14381 5355
rect 13964 5324 14381 5352
rect 13964 5312 13970 5324
rect 14369 5321 14381 5324
rect 14415 5352 14427 5355
rect 15102 5352 15108 5364
rect 14415 5324 15108 5352
rect 14415 5321 14427 5324
rect 14369 5315 14427 5321
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 12802 5284 12808 5296
rect 11134 5256 12808 5284
rect 11134 5253 11146 5256
rect 11088 5247 11146 5253
rect 12802 5244 12808 5256
rect 12860 5244 12866 5296
rect 15654 5284 15660 5296
rect 15615 5256 15660 5284
rect 15654 5244 15660 5256
rect 15712 5244 15718 5296
rect 9122 5176 9128 5228
rect 9180 5216 9186 5228
rect 9502 5219 9560 5225
rect 9502 5216 9514 5219
rect 9180 5188 9514 5216
rect 9180 5176 9186 5188
rect 9502 5185 9514 5188
rect 9548 5185 9560 5219
rect 9766 5216 9772 5228
rect 9727 5188 9772 5216
rect 9502 5179 9560 5185
rect 9766 5176 9772 5188
rect 9824 5176 9830 5228
rect 11330 5216 11336 5228
rect 11291 5188 11336 5216
rect 11330 5176 11336 5188
rect 11388 5176 11394 5228
rect 12641 5219 12699 5225
rect 12641 5185 12653 5219
rect 12687 5216 12699 5219
rect 13357 5219 13415 5225
rect 12687 5188 13308 5216
rect 12687 5185 12699 5188
rect 12641 5179 12699 5185
rect 7285 5151 7343 5157
rect 7285 5117 7297 5151
rect 7331 5117 7343 5151
rect 7285 5111 7343 5117
rect 7374 5108 7380 5160
rect 7432 5148 7438 5160
rect 7653 5151 7711 5157
rect 7653 5148 7665 5151
rect 7432 5120 7665 5148
rect 7432 5108 7438 5120
rect 7653 5117 7665 5120
rect 7699 5117 7711 5151
rect 7653 5111 7711 5117
rect 7837 5151 7895 5157
rect 7837 5117 7849 5151
rect 7883 5117 7895 5151
rect 7837 5111 7895 5117
rect 12897 5151 12955 5157
rect 12897 5117 12909 5151
rect 12943 5117 12955 5151
rect 12897 5111 12955 5117
rect 4246 5040 4252 5092
rect 4304 5080 4310 5092
rect 4304 5052 4844 5080
rect 4304 5040 4310 5052
rect 4154 4972 4160 5024
rect 4212 5012 4218 5024
rect 4617 5015 4675 5021
rect 4617 5012 4629 5015
rect 4212 4984 4629 5012
rect 4212 4972 4218 4984
rect 4617 4981 4629 4984
rect 4663 4981 4675 5015
rect 4816 5012 4844 5052
rect 6362 5040 6368 5092
rect 6420 5080 6426 5092
rect 6733 5083 6791 5089
rect 6733 5080 6745 5083
rect 6420 5052 6745 5080
rect 6420 5040 6426 5052
rect 6733 5049 6745 5052
rect 6779 5049 6791 5083
rect 6733 5043 6791 5049
rect 7098 5040 7104 5092
rect 7156 5080 7162 5092
rect 7852 5080 7880 5111
rect 8018 5080 8024 5092
rect 7156 5052 8024 5080
rect 7156 5040 7162 5052
rect 8018 5040 8024 5052
rect 8076 5040 8082 5092
rect 6086 5012 6092 5024
rect 4816 4984 6092 5012
rect 4617 4975 4675 4981
rect 6086 4972 6092 4984
rect 6144 4972 6150 5024
rect 6181 5015 6239 5021
rect 6181 4981 6193 5015
rect 6227 5012 6239 5015
rect 6270 5012 6276 5024
rect 6227 4984 6276 5012
rect 6227 4981 6239 4984
rect 6181 4975 6239 4981
rect 6270 4972 6276 4984
rect 6328 4972 6334 5024
rect 8294 5012 8300 5024
rect 8255 4984 8300 5012
rect 8294 4972 8300 4984
rect 8352 4972 8358 5024
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 11054 5012 11060 5024
rect 10100 4984 11060 5012
rect 10100 4972 10106 4984
rect 11054 4972 11060 4984
rect 11112 4972 11118 5024
rect 12526 4972 12532 5024
rect 12584 5012 12590 5024
rect 12912 5012 12940 5111
rect 13280 5080 13308 5188
rect 13357 5185 13369 5219
rect 13403 5216 13415 5219
rect 16298 5216 16304 5228
rect 13403 5188 16304 5216
rect 13403 5185 13415 5188
rect 13357 5179 13415 5185
rect 16298 5176 16304 5188
rect 16356 5176 16362 5228
rect 13538 5148 13544 5160
rect 13499 5120 13544 5148
rect 13538 5108 13544 5120
rect 13596 5108 13602 5160
rect 14734 5080 14740 5092
rect 13280 5052 14740 5080
rect 14734 5040 14740 5052
rect 14792 5040 14798 5092
rect 12584 4984 12940 5012
rect 12584 4972 12590 4984
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 2222 4768 2228 4820
rect 2280 4808 2286 4820
rect 2869 4811 2927 4817
rect 2869 4808 2881 4811
rect 2280 4780 2881 4808
rect 2280 4768 2286 4780
rect 2869 4777 2881 4780
rect 2915 4777 2927 4811
rect 7098 4808 7104 4820
rect 2869 4771 2927 4777
rect 3804 4780 7104 4808
rect 2406 4700 2412 4752
rect 2464 4700 2470 4752
rect 3804 4740 3832 4780
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7190 4768 7196 4820
rect 7248 4808 7254 4820
rect 7929 4811 7987 4817
rect 7929 4808 7941 4811
rect 7248 4780 7941 4808
rect 7248 4768 7254 4780
rect 7929 4777 7941 4780
rect 7975 4777 7987 4811
rect 7929 4771 7987 4777
rect 9214 4768 9220 4820
rect 9272 4808 9278 4820
rect 11422 4808 11428 4820
rect 9272 4780 11428 4808
rect 9272 4768 9278 4780
rect 11422 4768 11428 4780
rect 11480 4768 11486 4820
rect 12437 4811 12495 4817
rect 12437 4777 12449 4811
rect 12483 4808 12495 4811
rect 13722 4808 13728 4820
rect 12483 4780 13728 4808
rect 12483 4777 12495 4780
rect 12437 4771 12495 4777
rect 13722 4768 13728 4780
rect 13780 4768 13786 4820
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 13909 4811 13967 4817
rect 13909 4808 13921 4811
rect 13872 4780 13921 4808
rect 13872 4768 13878 4780
rect 13909 4777 13921 4780
rect 13955 4777 13967 4811
rect 14734 4808 14740 4820
rect 14695 4780 14740 4808
rect 13909 4771 13967 4777
rect 2516 4712 3832 4740
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 2038 4604 2044 4616
rect 1719 4576 2044 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 2038 4564 2044 4576
rect 2096 4564 2102 4616
rect 2424 4613 2452 4700
rect 2516 4681 2544 4712
rect 5074 4700 5080 4752
rect 5132 4740 5138 4752
rect 5169 4743 5227 4749
rect 5169 4740 5181 4743
rect 5132 4712 5181 4740
rect 5132 4700 5138 4712
rect 5169 4709 5181 4712
rect 5215 4709 5227 4743
rect 5169 4703 5227 4709
rect 5626 4700 5632 4752
rect 5684 4740 5690 4752
rect 5684 4712 5948 4740
rect 5684 4700 5690 4712
rect 2501 4675 2559 4681
rect 2501 4641 2513 4675
rect 2547 4641 2559 4675
rect 2682 4672 2688 4684
rect 2643 4644 2688 4672
rect 2501 4635 2559 4641
rect 2682 4632 2688 4644
rect 2740 4672 2746 4684
rect 3513 4675 3571 4681
rect 3513 4672 3525 4675
rect 2740 4644 3525 4672
rect 2740 4632 2746 4644
rect 3513 4641 3525 4644
rect 3559 4641 3571 4675
rect 3786 4672 3792 4684
rect 3747 4644 3792 4672
rect 3513 4635 3571 4641
rect 2409 4607 2467 4613
rect 2409 4573 2421 4607
rect 2455 4573 2467 4607
rect 2409 4567 2467 4573
rect 3234 4564 3240 4616
rect 3292 4604 3298 4616
rect 3329 4607 3387 4613
rect 3329 4604 3341 4607
rect 3292 4576 3341 4604
rect 3292 4564 3298 4576
rect 3329 4573 3341 4576
rect 3375 4573 3387 4607
rect 3528 4604 3556 4635
rect 3786 4632 3792 4644
rect 3844 4632 3850 4684
rect 5092 4604 5120 4700
rect 5920 4684 5948 4712
rect 7558 4700 7564 4752
rect 7616 4740 7622 4752
rect 7745 4743 7803 4749
rect 7745 4740 7757 4743
rect 7616 4712 7757 4740
rect 7616 4700 7622 4712
rect 7745 4709 7757 4712
rect 7791 4740 7803 4743
rect 7791 4712 9444 4740
rect 7791 4709 7803 4712
rect 7745 4703 7803 4709
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 5960 4644 6005 4672
rect 5960 4632 5966 4644
rect 8294 4632 8300 4684
rect 8352 4672 8358 4684
rect 8389 4675 8447 4681
rect 8389 4672 8401 4675
rect 8352 4644 8401 4672
rect 8352 4632 8358 4644
rect 8389 4641 8401 4644
rect 8435 4641 8447 4675
rect 8389 4635 8447 4641
rect 8478 4632 8484 4684
rect 8536 4672 8542 4684
rect 9125 4675 9183 4681
rect 8536 4644 8581 4672
rect 8536 4632 8542 4644
rect 9125 4641 9137 4675
rect 9171 4672 9183 4675
rect 9214 4672 9220 4684
rect 9171 4644 9220 4672
rect 9171 4641 9183 4644
rect 9125 4635 9183 4641
rect 9214 4632 9220 4644
rect 9272 4632 9278 4684
rect 5258 4604 5264 4616
rect 3528 4576 5120 4604
rect 5219 4576 5264 4604
rect 3329 4567 3387 4573
rect 5258 4564 5264 4576
rect 5316 4564 5322 4616
rect 5813 4607 5871 4613
rect 5813 4573 5825 4607
rect 5859 4600 5871 4607
rect 5859 4573 5948 4600
rect 5813 4572 5948 4573
rect 5813 4567 5871 4572
rect 1949 4539 2007 4545
rect 1949 4505 1961 4539
rect 1995 4536 2007 4539
rect 4056 4539 4114 4545
rect 1995 4508 4016 4536
rect 1995 4505 2007 4508
rect 1949 4499 2007 4505
rect 3988 4480 4016 4508
rect 4056 4505 4068 4539
rect 4102 4536 4114 4539
rect 4338 4536 4344 4548
rect 4102 4508 4344 4536
rect 4102 4505 4114 4508
rect 4056 4499 4114 4505
rect 4338 4496 4344 4508
rect 4396 4496 4402 4548
rect 5166 4496 5172 4548
rect 5224 4536 5230 4548
rect 5920 4536 5948 4572
rect 5994 4564 6000 4616
rect 6052 4604 6058 4616
rect 6161 4607 6219 4613
rect 6161 4604 6173 4607
rect 6052 4576 6173 4604
rect 6052 4564 6058 4576
rect 6161 4573 6173 4576
rect 6207 4573 6219 4607
rect 6161 4567 6219 4573
rect 7653 4607 7711 4613
rect 7653 4573 7665 4607
rect 7699 4604 7711 4607
rect 8938 4604 8944 4616
rect 7699 4576 8944 4604
rect 7699 4573 7711 4576
rect 7653 4567 7711 4573
rect 8938 4564 8944 4576
rect 8996 4564 9002 4616
rect 9416 4613 9444 4712
rect 9674 4700 9680 4752
rect 9732 4740 9738 4752
rect 11330 4740 11336 4752
rect 9732 4712 10732 4740
rect 11291 4712 11336 4740
rect 9732 4700 9738 4712
rect 9769 4675 9827 4681
rect 9769 4641 9781 4675
rect 9815 4672 9827 4675
rect 10594 4672 10600 4684
rect 9815 4644 10600 4672
rect 9815 4641 9827 4644
rect 9769 4635 9827 4641
rect 10594 4632 10600 4644
rect 10652 4632 10658 4684
rect 10704 4681 10732 4712
rect 11330 4700 11336 4712
rect 11388 4700 11394 4752
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4641 10747 4675
rect 11606 4672 11612 4684
rect 10689 4635 10747 4641
rect 10796 4644 11612 4672
rect 9401 4607 9459 4613
rect 9401 4573 9413 4607
rect 9447 4573 9459 4607
rect 9401 4567 9459 4573
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4604 9919 4607
rect 10042 4604 10048 4616
rect 9907 4576 10048 4604
rect 9907 4573 9919 4576
rect 9861 4567 9919 4573
rect 10042 4564 10048 4576
rect 10100 4564 10106 4616
rect 10134 4564 10140 4616
rect 10192 4604 10198 4616
rect 10413 4607 10471 4613
rect 10413 4604 10425 4607
rect 10192 4576 10425 4604
rect 10192 4564 10198 4576
rect 10413 4573 10425 4576
rect 10459 4573 10471 4607
rect 10796 4604 10824 4644
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 11885 4675 11943 4681
rect 11885 4641 11897 4675
rect 11931 4641 11943 4675
rect 11885 4635 11943 4641
rect 11977 4675 12035 4681
rect 11977 4641 11989 4675
rect 12023 4672 12035 4675
rect 12023 4644 12664 4672
rect 12023 4641 12035 4644
rect 11977 4635 12035 4641
rect 10413 4567 10471 4573
rect 10520 4576 10824 4604
rect 7558 4536 7564 4548
rect 5224 4508 5856 4536
rect 5920 4508 7564 4536
rect 5224 4496 5230 4508
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 2041 4471 2099 4477
rect 2041 4437 2053 4471
rect 2087 4468 2099 4471
rect 2222 4468 2228 4480
rect 2087 4440 2228 4468
rect 2087 4437 2099 4440
rect 2041 4431 2099 4437
rect 2222 4428 2228 4440
rect 2280 4428 2286 4480
rect 3237 4471 3295 4477
rect 3237 4437 3249 4471
rect 3283 4468 3295 4471
rect 3510 4468 3516 4480
rect 3283 4440 3516 4468
rect 3283 4437 3295 4440
rect 3237 4431 3295 4437
rect 3510 4428 3516 4440
rect 3568 4428 3574 4480
rect 3970 4428 3976 4480
rect 4028 4428 4034 4480
rect 5442 4468 5448 4480
rect 5403 4440 5448 4468
rect 5442 4428 5448 4440
rect 5500 4428 5506 4480
rect 5626 4468 5632 4480
rect 5587 4440 5632 4468
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 5828 4468 5856 4508
rect 7558 4496 7564 4508
rect 7616 4496 7622 4548
rect 10520 4536 10548 4576
rect 10870 4564 10876 4616
rect 10928 4604 10934 4616
rect 11517 4607 11575 4613
rect 11517 4604 11529 4607
rect 10928 4576 11529 4604
rect 10928 4564 10934 4576
rect 11517 4573 11529 4576
rect 11563 4604 11575 4607
rect 11790 4604 11796 4616
rect 11563 4576 11796 4604
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 11790 4564 11796 4576
rect 11848 4564 11854 4616
rect 10244 4508 10548 4536
rect 7006 4468 7012 4480
rect 5828 4440 7012 4468
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7282 4468 7288 4480
rect 7243 4440 7288 4468
rect 7282 4428 7288 4440
rect 7340 4428 7346 4480
rect 7466 4468 7472 4480
rect 7427 4440 7472 4468
rect 7466 4428 7472 4440
rect 7524 4428 7530 4480
rect 8294 4468 8300 4480
rect 8255 4440 8300 4468
rect 8294 4428 8300 4440
rect 8352 4468 8358 4480
rect 9030 4468 9036 4480
rect 8352 4440 9036 4468
rect 8352 4428 8358 4440
rect 9030 4428 9036 4440
rect 9088 4428 9094 4480
rect 9214 4468 9220 4480
rect 9175 4440 9220 4468
rect 9214 4428 9220 4440
rect 9272 4428 9278 4480
rect 9398 4428 9404 4480
rect 9456 4468 9462 4480
rect 9674 4468 9680 4480
rect 9456 4440 9680 4468
rect 9456 4428 9462 4440
rect 9674 4428 9680 4440
rect 9732 4428 9738 4480
rect 9953 4471 10011 4477
rect 9953 4437 9965 4471
rect 9999 4468 10011 4471
rect 10244 4468 10272 4508
rect 9999 4440 10272 4468
rect 9999 4437 10011 4440
rect 9953 4431 10011 4437
rect 10318 4428 10324 4480
rect 10376 4468 10382 4480
rect 11900 4468 11928 4635
rect 12526 4604 12532 4616
rect 12487 4576 12532 4604
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 12636 4604 12664 4644
rect 13814 4604 13820 4616
rect 12636 4576 13820 4604
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 13924 4604 13952 4771
rect 14734 4768 14740 4780
rect 14792 4768 14798 4820
rect 15657 4675 15715 4681
rect 15657 4641 15669 4675
rect 15703 4672 15715 4675
rect 15746 4672 15752 4684
rect 15703 4644 15752 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 15746 4632 15752 4644
rect 15804 4632 15810 4684
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13924 4576 14105 4604
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4573 15439 4607
rect 15381 4567 15439 4573
rect 12069 4539 12127 4545
rect 12069 4505 12081 4539
rect 12115 4536 12127 4539
rect 12618 4536 12624 4548
rect 12115 4508 12624 4536
rect 12115 4505 12127 4508
rect 12069 4499 12127 4505
rect 12618 4496 12624 4508
rect 12676 4496 12682 4548
rect 12796 4539 12854 4545
rect 12796 4536 12808 4539
rect 12728 4508 12808 4536
rect 12728 4468 12756 4508
rect 12796 4505 12808 4508
rect 12842 4536 12854 4539
rect 14458 4536 14464 4548
rect 12842 4508 14464 4536
rect 12842 4505 12854 4508
rect 12796 4499 12854 4505
rect 14458 4496 14464 4508
rect 14516 4496 14522 4548
rect 15396 4536 15424 4567
rect 15654 4536 15660 4548
rect 15396 4508 15660 4536
rect 15654 4496 15660 4508
rect 15712 4536 15718 4548
rect 16390 4536 16396 4548
rect 15712 4508 16396 4536
rect 15712 4496 15718 4508
rect 16390 4496 16396 4508
rect 16448 4496 16454 4548
rect 10376 4440 10421 4468
rect 11900 4440 12756 4468
rect 10376 4428 10382 4440
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1394 4224 1400 4276
rect 1452 4264 1458 4276
rect 1765 4267 1823 4273
rect 1765 4264 1777 4267
rect 1452 4236 1777 4264
rect 1452 4224 1458 4236
rect 1765 4233 1777 4236
rect 1811 4233 1823 4267
rect 2682 4264 2688 4276
rect 1765 4227 1823 4233
rect 2332 4236 2688 4264
rect 2332 4196 2360 4236
rect 2682 4224 2688 4236
rect 2740 4224 2746 4276
rect 3510 4224 3516 4276
rect 3568 4264 3574 4276
rect 4430 4264 4436 4276
rect 3568 4236 4436 4264
rect 3568 4224 3574 4236
rect 4430 4224 4436 4236
rect 4488 4224 4494 4276
rect 4614 4224 4620 4276
rect 4672 4264 4678 4276
rect 5626 4264 5632 4276
rect 4672 4236 5632 4264
rect 4672 4224 4678 4236
rect 5626 4224 5632 4236
rect 5684 4224 5690 4276
rect 6362 4224 6368 4276
rect 6420 4264 6426 4276
rect 6825 4267 6883 4273
rect 6825 4264 6837 4267
rect 6420 4236 6837 4264
rect 6420 4224 6426 4236
rect 6825 4233 6837 4236
rect 6871 4233 6883 4267
rect 9582 4264 9588 4276
rect 6825 4227 6883 4233
rect 8864 4236 9588 4264
rect 3786 4196 3792 4208
rect 1596 4168 2360 4196
rect 2424 4168 3792 4196
rect 1596 4069 1624 4168
rect 2424 4128 2452 4168
rect 3786 4156 3792 4168
rect 3844 4156 3850 4208
rect 4522 4156 4528 4208
rect 4580 4196 4586 4208
rect 4580 4168 6408 4196
rect 4580 4156 4586 4168
rect 2240 4100 2452 4128
rect 2492 4131 2550 4137
rect 1581 4063 1639 4069
rect 1581 4029 1593 4063
rect 1627 4029 1639 4063
rect 1581 4023 1639 4029
rect 1670 4020 1676 4072
rect 1728 4060 1734 4072
rect 1728 4032 1773 4060
rect 1728 4020 1734 4032
rect 2038 4020 2044 4072
rect 2096 4060 2102 4072
rect 2240 4069 2268 4100
rect 2492 4097 2504 4131
rect 2538 4128 2550 4131
rect 3510 4128 3516 4140
rect 2538 4100 3516 4128
rect 2538 4097 2550 4100
rect 2492 4091 2550 4097
rect 3510 4088 3516 4100
rect 3568 4088 3574 4140
rect 3697 4132 3755 4137
rect 3620 4131 3755 4132
rect 3620 4104 3709 4131
rect 2225 4063 2283 4069
rect 2225 4060 2237 4063
rect 2096 4032 2237 4060
rect 2096 4020 2102 4032
rect 2225 4029 2237 4032
rect 2271 4029 2283 4063
rect 2225 4023 2283 4029
rect 198 3952 204 4004
rect 256 3992 262 4004
rect 256 3964 2268 3992
rect 256 3952 262 3964
rect 2130 3924 2136 3936
rect 2091 3896 2136 3924
rect 2130 3884 2136 3896
rect 2188 3884 2194 3936
rect 2240 3924 2268 3964
rect 3620 3936 3648 4104
rect 3697 4097 3709 4104
rect 3743 4097 3755 4131
rect 4338 4128 4344 4140
rect 4299 4100 4344 4128
rect 3697 4091 3755 4097
rect 4338 4088 4344 4100
rect 4396 4088 4402 4140
rect 5258 4088 5264 4140
rect 5316 4128 5322 4140
rect 5546 4131 5604 4137
rect 5546 4128 5558 4131
rect 5316 4100 5558 4128
rect 5316 4088 5322 4100
rect 5546 4097 5558 4100
rect 5592 4097 5604 4131
rect 5546 4091 5604 4097
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4128 5871 4131
rect 5902 4128 5908 4140
rect 5859 4100 5908 4128
rect 5859 4097 5871 4100
rect 5813 4091 5871 4097
rect 5902 4088 5908 4100
rect 5960 4088 5966 4140
rect 6181 4131 6239 4137
rect 6181 4097 6193 4131
rect 6227 4097 6239 4131
rect 6380 4128 6408 4168
rect 6454 4156 6460 4208
rect 6512 4196 6518 4208
rect 6733 4199 6791 4205
rect 6733 4196 6745 4199
rect 6512 4168 6745 4196
rect 6512 4156 6518 4168
rect 6733 4165 6745 4168
rect 6779 4165 6791 4199
rect 8662 4196 8668 4208
rect 6733 4159 6791 4165
rect 6840 4168 8668 4196
rect 6840 4128 6868 4168
rect 8662 4156 8668 4168
rect 8720 4156 8726 4208
rect 7282 4128 7288 4140
rect 6380 4100 6868 4128
rect 7243 4100 7288 4128
rect 6181 4091 6239 4097
rect 6196 3992 6224 4091
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 8205 4131 8263 4137
rect 8205 4097 8217 4131
rect 8251 4128 8263 4131
rect 8864 4128 8892 4236
rect 9582 4224 9588 4236
rect 9640 4224 9646 4276
rect 9858 4224 9864 4276
rect 9916 4224 9922 4276
rect 10045 4267 10103 4273
rect 10045 4233 10057 4267
rect 10091 4264 10103 4267
rect 10134 4264 10140 4276
rect 10091 4236 10140 4264
rect 10091 4233 10103 4236
rect 10045 4227 10103 4233
rect 10134 4224 10140 4236
rect 10192 4224 10198 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 12069 4267 12127 4273
rect 12069 4264 12081 4267
rect 11480 4236 12081 4264
rect 11480 4224 11486 4236
rect 12069 4233 12081 4236
rect 12115 4233 12127 4267
rect 12069 4227 12127 4233
rect 12437 4267 12495 4273
rect 12437 4233 12449 4267
rect 12483 4264 12495 4267
rect 12618 4264 12624 4276
rect 12483 4236 12624 4264
rect 12483 4233 12495 4236
rect 12437 4227 12495 4233
rect 12618 4224 12624 4236
rect 12676 4224 12682 4276
rect 12710 4224 12716 4276
rect 12768 4224 12774 4276
rect 13814 4224 13820 4276
rect 13872 4264 13878 4276
rect 14921 4267 14979 4273
rect 14921 4264 14933 4267
rect 13872 4236 14933 4264
rect 13872 4224 13878 4236
rect 14921 4233 14933 4236
rect 14967 4233 14979 4267
rect 14921 4227 14979 4233
rect 15289 4267 15347 4273
rect 15289 4233 15301 4267
rect 15335 4264 15347 4267
rect 15470 4264 15476 4276
rect 15335 4236 15476 4264
rect 15335 4233 15347 4236
rect 15289 4227 15347 4233
rect 15470 4224 15476 4236
rect 15528 4224 15534 4276
rect 9876 4196 9904 4224
rect 10152 4196 10180 4224
rect 12728 4196 12756 4224
rect 9140 4168 9536 4196
rect 9876 4168 10088 4196
rect 10152 4168 12756 4196
rect 8251 4100 8892 4128
rect 8941 4131 8999 4137
rect 8251 4097 8263 4100
rect 8205 4091 8263 4097
rect 8941 4097 8953 4131
rect 8987 4128 8999 4131
rect 9030 4128 9036 4140
rect 8987 4100 9036 4128
rect 8987 4097 8999 4100
rect 8941 4091 8999 4097
rect 9030 4088 9036 4100
rect 9088 4088 9094 4140
rect 6270 4020 6276 4072
rect 6328 4060 6334 4072
rect 9140 4069 9168 4168
rect 9398 4128 9404 4140
rect 9359 4100 9404 4128
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 6917 4063 6975 4069
rect 6917 4060 6929 4063
rect 6328 4032 6929 4060
rect 6328 4020 6334 4032
rect 6917 4029 6929 4032
rect 6963 4029 6975 4063
rect 6917 4023 6975 4029
rect 9125 4063 9183 4069
rect 9125 4029 9137 4063
rect 9171 4029 9183 4063
rect 9306 4060 9312 4072
rect 9267 4032 9312 4060
rect 9125 4023 9183 4029
rect 9306 4020 9312 4032
rect 9364 4020 9370 4072
rect 9508 4060 9536 4168
rect 9582 4088 9588 4140
rect 9640 4128 9646 4140
rect 9861 4131 9919 4137
rect 9861 4128 9873 4131
rect 9640 4100 9873 4128
rect 9640 4088 9646 4100
rect 9861 4097 9873 4100
rect 9907 4097 9919 4131
rect 10060 4128 10088 4168
rect 14550 4156 14556 4208
rect 14608 4156 14614 4208
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10060 4100 10517 4128
rect 9861 4091 9919 4097
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10597 4131 10655 4137
rect 10597 4097 10609 4131
rect 10643 4128 10655 4131
rect 10778 4128 10784 4140
rect 10643 4100 10784 4128
rect 10643 4097 10655 4100
rect 10597 4091 10655 4097
rect 9876 4060 9904 4091
rect 10778 4088 10784 4100
rect 10836 4088 10842 4140
rect 11054 4128 11060 4140
rect 11015 4100 11060 4128
rect 11054 4088 11060 4100
rect 11112 4088 11118 4140
rect 11974 4128 11980 4140
rect 11935 4100 11980 4128
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12796 4131 12854 4137
rect 12796 4128 12808 4131
rect 12406 4100 12808 4128
rect 10686 4060 10692 4072
rect 9508 4032 9674 4060
rect 9876 4032 10364 4060
rect 10647 4032 10692 4060
rect 8021 3995 8079 4001
rect 8021 3992 8033 3995
rect 6196 3964 8033 3992
rect 8021 3961 8033 3964
rect 8067 3961 8079 3995
rect 8021 3955 8079 3961
rect 8110 3952 8116 4004
rect 8168 3992 8174 4004
rect 9490 3992 9496 4004
rect 8168 3964 9496 3992
rect 8168 3952 8174 3964
rect 9490 3952 9496 3964
rect 9548 3952 9554 4004
rect 9646 3992 9674 4032
rect 9858 3992 9864 4004
rect 9646 3964 9864 3992
rect 9858 3952 9864 3964
rect 9916 3952 9922 4004
rect 9950 3952 9956 4004
rect 10008 3992 10014 4004
rect 10137 3995 10195 4001
rect 10137 3992 10149 3995
rect 10008 3964 10149 3992
rect 10008 3952 10014 3964
rect 10137 3961 10149 3964
rect 10183 3961 10195 3995
rect 10336 3992 10364 4032
rect 10686 4020 10692 4032
rect 10744 4020 10750 4072
rect 11241 4063 11299 4069
rect 11241 4029 11253 4063
rect 11287 4060 11299 4063
rect 11330 4060 11336 4072
rect 11287 4032 11336 4060
rect 11287 4029 11299 4032
rect 11241 4023 11299 4029
rect 11330 4020 11336 4032
rect 11388 4020 11394 4072
rect 11885 4063 11943 4069
rect 11885 4029 11897 4063
rect 11931 4029 11943 4063
rect 11885 4023 11943 4029
rect 11517 3995 11575 4001
rect 11517 3992 11529 3995
rect 10336 3964 11529 3992
rect 10137 3955 10195 3961
rect 11517 3961 11529 3964
rect 11563 3961 11575 3995
rect 11900 3992 11928 4023
rect 12406 3992 12434 4100
rect 12796 4097 12808 4100
rect 12842 4128 12854 4131
rect 13722 4128 13728 4140
rect 12842 4100 13728 4128
rect 12842 4097 12854 4100
rect 12796 4091 12854 4097
rect 13722 4088 13728 4100
rect 13780 4088 13786 4140
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 14568 4128 14596 4156
rect 14826 4128 14832 4140
rect 13872 4100 14596 4128
rect 14787 4100 14832 4128
rect 13872 4088 13878 4100
rect 14826 4088 14832 4100
rect 14884 4088 14890 4140
rect 15378 4088 15384 4140
rect 15436 4128 15442 4140
rect 15436 4100 15481 4128
rect 15436 4088 15442 4100
rect 12526 4020 12532 4072
rect 12584 4060 12590 4072
rect 14553 4063 14611 4069
rect 14553 4060 14565 4063
rect 12584 4032 12677 4060
rect 13556 4032 14565 4060
rect 12584 4020 12590 4032
rect 11900 3964 12434 3992
rect 11517 3955 11575 3961
rect 3234 3924 3240 3936
rect 2240 3896 3240 3924
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3602 3924 3608 3936
rect 3563 3896 3608 3924
rect 3602 3884 3608 3896
rect 3660 3884 3666 3936
rect 5626 3884 5632 3936
rect 5684 3924 5690 3936
rect 5997 3927 6055 3933
rect 5997 3924 6009 3927
rect 5684 3896 6009 3924
rect 5684 3884 5690 3896
rect 5997 3893 6009 3896
rect 6043 3893 6055 3927
rect 5997 3887 6055 3893
rect 6086 3884 6092 3936
rect 6144 3924 6150 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 6144 3896 6377 3924
rect 6144 3884 6150 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 7650 3884 7656 3936
rect 7708 3924 7714 3936
rect 7929 3927 7987 3933
rect 7929 3924 7941 3927
rect 7708 3896 7941 3924
rect 7708 3884 7714 3896
rect 7929 3893 7941 3896
rect 7975 3893 7987 3927
rect 7929 3887 7987 3893
rect 8297 3927 8355 3933
rect 8297 3893 8309 3927
rect 8343 3924 8355 3927
rect 8478 3924 8484 3936
rect 8343 3896 8484 3924
rect 8343 3893 8355 3896
rect 8297 3887 8355 3893
rect 8478 3884 8484 3896
rect 8536 3884 8542 3936
rect 9674 3884 9680 3936
rect 9732 3924 9738 3936
rect 9769 3927 9827 3933
rect 9769 3924 9781 3927
rect 9732 3896 9781 3924
rect 9732 3884 9738 3896
rect 9769 3893 9781 3896
rect 9815 3893 9827 3927
rect 9769 3887 9827 3893
rect 11606 3884 11612 3936
rect 11664 3924 11670 3936
rect 12544 3924 12572 4020
rect 11664 3896 12572 3924
rect 11664 3884 11670 3896
rect 12802 3884 12808 3936
rect 12860 3924 12866 3936
rect 13556 3924 13584 4032
rect 14553 4029 14565 4032
rect 14599 4029 14611 4063
rect 14553 4023 14611 4029
rect 13909 3995 13967 4001
rect 13909 3961 13921 3995
rect 13955 3992 13967 3995
rect 14458 3992 14464 4004
rect 13955 3964 14464 3992
rect 13955 3961 13967 3964
rect 13909 3955 13967 3961
rect 14458 3952 14464 3964
rect 14516 3952 14522 4004
rect 14844 3992 14872 4088
rect 15562 4060 15568 4072
rect 15523 4032 15568 4060
rect 15562 4020 15568 4032
rect 15620 4020 15626 4072
rect 16482 3992 16488 4004
rect 14844 3964 16488 3992
rect 16482 3952 16488 3964
rect 16540 3952 16546 4004
rect 12860 3896 13584 3924
rect 12860 3884 12866 3896
rect 14550 3884 14556 3936
rect 14608 3924 14614 3936
rect 15838 3924 15844 3936
rect 14608 3896 15844 3924
rect 14608 3884 14614 3896
rect 15838 3884 15844 3896
rect 15896 3884 15902 3936
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 1946 3720 1952 3732
rect 1907 3692 1952 3720
rect 1946 3680 1952 3692
rect 2004 3680 2010 3732
rect 3234 3680 3240 3732
rect 3292 3720 3298 3732
rect 7374 3720 7380 3732
rect 3292 3692 5948 3720
rect 7335 3692 7380 3720
rect 3292 3680 3298 3692
rect 1026 3612 1032 3664
rect 1084 3652 1090 3664
rect 1673 3655 1731 3661
rect 1673 3652 1685 3655
rect 1084 3624 1685 3652
rect 1084 3612 1090 3624
rect 1673 3621 1685 3624
rect 1719 3621 1731 3655
rect 2314 3652 2320 3664
rect 1673 3615 1731 3621
rect 1780 3624 2320 3652
rect 566 3544 572 3596
rect 624 3584 630 3596
rect 1780 3584 1808 3624
rect 2314 3612 2320 3624
rect 2372 3612 2378 3664
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 3142 3652 3148 3664
rect 2915 3624 3148 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 3142 3612 3148 3624
rect 3200 3612 3206 3664
rect 5442 3652 5448 3664
rect 3436 3624 5448 3652
rect 624 3556 1808 3584
rect 624 3544 630 3556
rect 2222 3544 2228 3596
rect 2280 3584 2286 3596
rect 2409 3587 2467 3593
rect 2409 3584 2421 3587
rect 2280 3556 2421 3584
rect 2280 3544 2286 3556
rect 2409 3553 2421 3556
rect 2455 3553 2467 3587
rect 2409 3547 2467 3553
rect 2498 3544 2504 3596
rect 2556 3584 2562 3596
rect 3436 3584 3464 3624
rect 5442 3612 5448 3624
rect 5500 3612 5506 3664
rect 5920 3652 5948 3692
rect 7374 3680 7380 3692
rect 7432 3680 7438 3732
rect 9125 3723 9183 3729
rect 9125 3720 9137 3723
rect 7484 3692 9137 3720
rect 7484 3652 7512 3692
rect 9125 3689 9137 3692
rect 9171 3689 9183 3723
rect 9125 3683 9183 3689
rect 9398 3680 9404 3732
rect 9456 3720 9462 3732
rect 9585 3723 9643 3729
rect 9585 3720 9597 3723
rect 9456 3692 9597 3720
rect 9456 3680 9462 3692
rect 9585 3689 9597 3692
rect 9631 3689 9643 3723
rect 12986 3720 12992 3732
rect 9585 3683 9643 3689
rect 10060 3692 12992 3720
rect 9766 3652 9772 3664
rect 5920 3624 7512 3652
rect 8772 3624 9772 3652
rect 2556 3556 2601 3584
rect 2700 3556 3464 3584
rect 3513 3587 3571 3593
rect 2556 3544 2562 3556
rect 1854 3516 1860 3528
rect 1815 3488 1860 3516
rect 1854 3476 1860 3488
rect 1912 3476 1918 3528
rect 2130 3476 2136 3528
rect 2188 3516 2194 3528
rect 2317 3519 2375 3525
rect 2317 3516 2329 3519
rect 2188 3488 2329 3516
rect 2188 3476 2194 3488
rect 2317 3485 2329 3488
rect 2363 3485 2375 3519
rect 2317 3479 2375 3485
rect 2222 3408 2228 3460
rect 2280 3448 2286 3460
rect 2700 3448 2728 3556
rect 3513 3553 3525 3587
rect 3559 3584 3571 3587
rect 3602 3584 3608 3596
rect 3559 3556 3608 3584
rect 3559 3553 3571 3556
rect 3513 3547 3571 3553
rect 3602 3544 3608 3556
rect 3660 3544 3666 3596
rect 4430 3544 4436 3596
rect 4488 3584 4494 3596
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4488 3556 4537 3584
rect 4488 3544 4494 3556
rect 4525 3553 4537 3556
rect 4571 3553 4583 3587
rect 4525 3547 4583 3553
rect 5077 3587 5135 3593
rect 5077 3553 5089 3587
rect 5123 3584 5135 3587
rect 5258 3584 5264 3596
rect 5123 3556 5264 3584
rect 5123 3553 5135 3556
rect 5077 3547 5135 3553
rect 5258 3544 5264 3556
rect 5316 3584 5322 3596
rect 6362 3584 6368 3596
rect 5316 3556 6368 3584
rect 5316 3544 5322 3556
rect 6362 3544 6368 3556
rect 6420 3544 6426 3596
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7193 3587 7251 3593
rect 7193 3553 7205 3587
rect 7239 3584 7251 3587
rect 7282 3584 7288 3596
rect 7239 3556 7288 3584
rect 7239 3553 7251 3556
rect 7193 3547 7251 3553
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 8772 3593 8800 3624
rect 9766 3612 9772 3624
rect 9824 3612 9830 3664
rect 8757 3587 8815 3593
rect 8757 3553 8769 3587
rect 8803 3553 8815 3587
rect 10060 3584 10088 3692
rect 12986 3680 12992 3692
rect 13044 3720 13050 3732
rect 13538 3720 13544 3732
rect 13044 3692 13544 3720
rect 13044 3680 13050 3692
rect 13538 3680 13544 3692
rect 13596 3680 13602 3732
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 10376 3624 14872 3652
rect 10376 3612 10382 3624
rect 8757 3547 8815 3553
rect 9324 3556 10088 3584
rect 10137 3587 10195 3593
rect 3329 3519 3387 3525
rect 3329 3485 3341 3519
rect 3375 3516 3387 3519
rect 5169 3519 5227 3525
rect 3375 3488 5129 3516
rect 3375 3485 3387 3488
rect 3329 3479 3387 3485
rect 2280 3420 2728 3448
rect 3237 3451 3295 3457
rect 2280 3408 2286 3420
rect 3237 3417 3249 3451
rect 3283 3448 3295 3451
rect 3283 3420 4016 3448
rect 3283 3417 3295 3420
rect 3237 3411 3295 3417
rect 1489 3383 1547 3389
rect 1489 3349 1501 3383
rect 1535 3380 1547 3383
rect 3602 3380 3608 3392
rect 1535 3352 3608 3380
rect 1535 3349 1547 3352
rect 1489 3343 1547 3349
rect 3602 3340 3608 3352
rect 3660 3340 3666 3392
rect 3878 3380 3884 3392
rect 3839 3352 3884 3380
rect 3878 3340 3884 3352
rect 3936 3340 3942 3392
rect 3988 3389 4016 3420
rect 3973 3383 4031 3389
rect 3973 3349 3985 3383
rect 4019 3349 4031 3383
rect 4338 3380 4344 3392
rect 4299 3352 4344 3380
rect 3973 3343 4031 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 5101 3380 5129 3488
rect 5169 3485 5181 3519
rect 5215 3516 5227 3519
rect 5718 3516 5724 3528
rect 5215 3488 5724 3516
rect 5215 3485 5227 3488
rect 5169 3479 5227 3485
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 6089 3519 6147 3525
rect 6089 3485 6101 3519
rect 6135 3516 6147 3519
rect 7098 3516 7104 3528
rect 6135 3488 7104 3516
rect 6135 3485 6147 3488
rect 6089 3479 6147 3485
rect 7098 3476 7104 3488
rect 7156 3516 7162 3528
rect 7558 3516 7564 3528
rect 7156 3488 7564 3516
rect 7156 3476 7162 3488
rect 7558 3476 7564 3488
rect 7616 3476 7622 3528
rect 8478 3476 8484 3528
rect 8536 3525 8542 3528
rect 8536 3516 8548 3525
rect 8536 3488 8581 3516
rect 8536 3479 8548 3488
rect 8536 3476 8542 3479
rect 8662 3476 8668 3528
rect 8720 3516 8726 3528
rect 8941 3519 8999 3525
rect 8941 3516 8953 3519
rect 8720 3488 8953 3516
rect 8720 3476 8726 3488
rect 8941 3485 8953 3488
rect 8987 3485 8999 3519
rect 9324 3516 9352 3556
rect 10137 3553 10149 3587
rect 10183 3584 10195 3587
rect 10962 3584 10968 3596
rect 10183 3556 10968 3584
rect 10183 3553 10195 3556
rect 10137 3547 10195 3553
rect 10962 3544 10968 3556
rect 11020 3584 11026 3596
rect 12805 3587 12863 3593
rect 12805 3584 12817 3587
rect 11020 3556 12817 3584
rect 11020 3544 11026 3556
rect 12805 3553 12817 3556
rect 12851 3553 12863 3587
rect 12805 3547 12863 3553
rect 13078 3544 13084 3596
rect 13136 3544 13142 3596
rect 13170 3544 13176 3596
rect 13228 3584 13234 3596
rect 13814 3584 13820 3596
rect 13228 3556 13820 3584
rect 13228 3544 13234 3556
rect 13814 3544 13820 3556
rect 13872 3584 13878 3596
rect 13909 3587 13967 3593
rect 13909 3584 13921 3587
rect 13872 3556 13921 3584
rect 13872 3544 13878 3556
rect 13909 3553 13921 3556
rect 13955 3553 13967 3587
rect 13909 3547 13967 3553
rect 14458 3544 14464 3596
rect 14516 3584 14522 3596
rect 14553 3587 14611 3593
rect 14553 3584 14565 3587
rect 14516 3556 14565 3584
rect 14516 3544 14522 3556
rect 14553 3553 14565 3556
rect 14599 3584 14611 3587
rect 14642 3584 14648 3596
rect 14599 3556 14648 3584
rect 14599 3553 14611 3556
rect 14553 3547 14611 3553
rect 14642 3544 14648 3556
rect 14700 3544 14706 3596
rect 14844 3593 14872 3624
rect 14829 3587 14887 3593
rect 14829 3553 14841 3587
rect 14875 3553 14887 3587
rect 14829 3547 14887 3553
rect 15286 3544 15292 3596
rect 15344 3584 15350 3596
rect 15473 3587 15531 3593
rect 15473 3584 15485 3587
rect 15344 3556 15485 3584
rect 15344 3544 15350 3556
rect 15473 3553 15485 3556
rect 15519 3553 15531 3587
rect 15473 3547 15531 3553
rect 9490 3516 9496 3528
rect 8941 3479 8999 3485
rect 9048 3488 9352 3516
rect 9451 3488 9496 3516
rect 5442 3408 5448 3460
rect 5500 3448 5506 3460
rect 9048 3448 9076 3488
rect 9490 3476 9496 3488
rect 9548 3476 9554 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10100 3488 10145 3516
rect 10100 3476 10106 3488
rect 10226 3476 10232 3528
rect 10284 3516 10290 3528
rect 10413 3519 10471 3525
rect 10413 3516 10425 3519
rect 10284 3488 10425 3516
rect 10284 3476 10290 3488
rect 10413 3485 10425 3488
rect 10459 3485 10471 3519
rect 10413 3479 10471 3485
rect 11882 3476 11888 3528
rect 11940 3516 11946 3528
rect 12713 3519 12771 3525
rect 12713 3516 12725 3519
rect 11940 3488 12725 3516
rect 11940 3476 11946 3488
rect 12713 3485 12725 3488
rect 12759 3485 12771 3519
rect 13096 3516 13124 3544
rect 13538 3516 13544 3528
rect 13096 3488 13544 3516
rect 12713 3479 12771 3485
rect 13538 3476 13544 3488
rect 13596 3516 13602 3528
rect 13633 3519 13691 3525
rect 13633 3516 13645 3519
rect 13596 3488 13645 3516
rect 13596 3476 13602 3488
rect 13633 3485 13645 3488
rect 13679 3485 13691 3519
rect 14090 3516 14096 3528
rect 14051 3488 14096 3516
rect 13633 3479 13691 3485
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 14277 3519 14335 3525
rect 14277 3485 14289 3519
rect 14323 3516 14335 3519
rect 14918 3516 14924 3528
rect 14323 3488 14924 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 14918 3476 14924 3488
rect 14976 3516 14982 3528
rect 15930 3516 15936 3528
rect 14976 3488 15936 3516
rect 14976 3476 14982 3488
rect 15930 3476 15936 3488
rect 15988 3476 15994 3528
rect 12158 3448 12164 3460
rect 5500 3420 9076 3448
rect 9140 3420 9628 3448
rect 5500 3408 5506 3420
rect 5166 3380 5172 3392
rect 4488 3352 4533 3380
rect 5101 3352 5172 3380
rect 4488 3340 4494 3352
rect 5166 3340 5172 3352
rect 5224 3340 5230 3392
rect 5258 3340 5264 3392
rect 5316 3380 5322 3392
rect 5316 3352 5361 3380
rect 5316 3340 5322 3352
rect 5534 3340 5540 3392
rect 5592 3380 5598 3392
rect 5629 3383 5687 3389
rect 5629 3380 5641 3383
rect 5592 3352 5641 3380
rect 5592 3340 5598 3352
rect 5629 3349 5641 3352
rect 5675 3349 5687 3383
rect 5629 3343 5687 3349
rect 5718 3340 5724 3392
rect 5776 3380 5782 3392
rect 6181 3383 6239 3389
rect 5776 3352 5821 3380
rect 5776 3340 5782 3352
rect 6181 3349 6193 3383
rect 6227 3380 6239 3383
rect 6549 3383 6607 3389
rect 6549 3380 6561 3383
rect 6227 3352 6561 3380
rect 6227 3349 6239 3352
rect 6181 3343 6239 3349
rect 6549 3349 6561 3352
rect 6595 3349 6607 3383
rect 6549 3343 6607 3349
rect 6917 3383 6975 3389
rect 6917 3349 6929 3383
rect 6963 3380 6975 3383
rect 7742 3380 7748 3392
rect 6963 3352 7748 3380
rect 6963 3349 6975 3352
rect 6917 3343 6975 3349
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 7834 3340 7840 3392
rect 7892 3380 7898 3392
rect 9140 3380 9168 3420
rect 9306 3380 9312 3392
rect 7892 3352 9168 3380
rect 9267 3352 9312 3380
rect 7892 3340 7898 3352
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9600 3380 9628 3420
rect 9876 3420 12164 3448
rect 9876 3380 9904 3420
rect 12158 3408 12164 3420
rect 12216 3408 12222 3460
rect 9600 3352 9904 3380
rect 9953 3383 10011 3389
rect 9953 3349 9965 3383
rect 9999 3380 10011 3383
rect 10042 3380 10048 3392
rect 9999 3352 10048 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 10042 3340 10048 3352
rect 10100 3340 10106 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 11701 3383 11759 3389
rect 11701 3380 11713 3383
rect 11664 3352 11713 3380
rect 11664 3340 11670 3352
rect 11701 3349 11713 3352
rect 11747 3349 11759 3383
rect 11701 3343 11759 3349
rect 11882 3340 11888 3392
rect 11940 3380 11946 3392
rect 12253 3383 12311 3389
rect 12253 3380 12265 3383
rect 11940 3352 12265 3380
rect 11940 3340 11946 3352
rect 12253 3349 12265 3352
rect 12299 3349 12311 3383
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 12253 3343 12311 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 3881 3179 3939 3185
rect 3881 3176 3893 3179
rect 1504 3148 3893 3176
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 1394 2796 1400 2848
rect 1452 2836 1458 2848
rect 1504 2836 1532 3148
rect 3881 3145 3893 3148
rect 3927 3145 3939 3179
rect 3881 3139 3939 3145
rect 4341 3179 4399 3185
rect 4341 3145 4353 3179
rect 4387 3176 4399 3179
rect 4430 3176 4436 3188
rect 4387 3148 4436 3176
rect 4387 3145 4399 3148
rect 4341 3139 4399 3145
rect 4430 3136 4436 3148
rect 4488 3136 4494 3188
rect 4709 3179 4767 3185
rect 4709 3145 4721 3179
rect 4755 3145 4767 3179
rect 5166 3176 5172 3188
rect 5127 3148 5172 3176
rect 4709 3139 4767 3145
rect 1762 3068 1768 3120
rect 1820 3108 1826 3120
rect 2308 3111 2366 3117
rect 1820 3080 2268 3108
rect 1820 3068 1826 3080
rect 1946 3040 1952 3052
rect 1907 3012 1952 3040
rect 1946 3000 1952 3012
rect 2004 3000 2010 3052
rect 2038 3000 2044 3052
rect 2096 3040 2102 3052
rect 2240 3040 2268 3080
rect 2308 3077 2320 3111
rect 2354 3108 2366 3111
rect 3510 3108 3516 3120
rect 2354 3080 3516 3108
rect 2354 3077 2366 3080
rect 2308 3071 2366 3077
rect 3510 3068 3516 3080
rect 3568 3068 3574 3120
rect 4154 3108 4160 3120
rect 3620 3080 4160 3108
rect 3620 3040 3648 3080
rect 4154 3068 4160 3080
rect 4212 3068 4218 3120
rect 4724 3108 4752 3139
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5534 3176 5540 3188
rect 5495 3148 5540 3176
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 5629 3179 5687 3185
rect 5629 3145 5641 3179
rect 5675 3176 5687 3179
rect 5718 3176 5724 3188
rect 5675 3148 5724 3176
rect 5675 3145 5687 3148
rect 5629 3139 5687 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 7466 3176 7472 3188
rect 6512 3148 7472 3176
rect 6512 3136 6518 3148
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 10134 3176 10140 3188
rect 7576 3148 10140 3176
rect 5074 3108 5080 3120
rect 4724 3080 5080 3108
rect 5074 3068 5080 3080
rect 5132 3108 5138 3120
rect 6365 3111 6423 3117
rect 5132 3080 6316 3108
rect 5132 3068 5138 3080
rect 2096 3012 2141 3040
rect 2240 3012 3648 3040
rect 3697 3043 3755 3049
rect 2096 3000 2102 3012
rect 3697 3009 3709 3043
rect 3743 3040 3755 3043
rect 4062 3040 4068 3052
rect 3743 3012 4068 3040
rect 3743 3009 3755 3012
rect 3697 3003 3755 3009
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 6178 3040 6184 3052
rect 6139 3012 6184 3040
rect 4249 3003 4307 3009
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3292 2944 3648 2972
rect 3292 2932 3298 2944
rect 1581 2907 1639 2913
rect 1581 2873 1593 2907
rect 1627 2904 1639 2907
rect 1854 2904 1860 2916
rect 1627 2876 1860 2904
rect 1627 2873 1639 2876
rect 1581 2867 1639 2873
rect 1854 2864 1860 2876
rect 1912 2864 1918 2916
rect 3142 2864 3148 2916
rect 3200 2864 3206 2916
rect 3510 2904 3516 2916
rect 3471 2876 3516 2904
rect 3510 2864 3516 2876
rect 3568 2864 3574 2916
rect 3620 2904 3648 2944
rect 3786 2932 3792 2984
rect 3844 2972 3850 2984
rect 4264 2972 4292 3003
rect 6178 3000 6184 3012
rect 6236 3000 6242 3052
rect 6288 3040 6316 3080
rect 6365 3077 6377 3111
rect 6411 3108 6423 3111
rect 7576 3108 7604 3148
rect 10134 3136 10140 3148
rect 10192 3176 10198 3188
rect 11054 3176 11060 3188
rect 10192 3148 11060 3176
rect 10192 3136 10198 3148
rect 11054 3136 11060 3148
rect 11112 3136 11118 3188
rect 11238 3136 11244 3188
rect 11296 3176 11302 3188
rect 11885 3179 11943 3185
rect 11885 3176 11897 3179
rect 11296 3148 11897 3176
rect 11296 3136 11302 3148
rect 11885 3145 11897 3148
rect 11931 3145 11943 3179
rect 11885 3139 11943 3145
rect 11977 3179 12035 3185
rect 11977 3145 11989 3179
rect 12023 3176 12035 3179
rect 12066 3176 12072 3188
rect 12023 3148 12072 3176
rect 12023 3145 12035 3148
rect 11977 3139 12035 3145
rect 12066 3136 12072 3148
rect 12124 3136 12130 3188
rect 13078 3176 13084 3188
rect 12544 3148 13084 3176
rect 6411 3080 7604 3108
rect 6411 3077 6423 3080
rect 6365 3071 6423 3077
rect 7650 3068 7656 3120
rect 7708 3117 7714 3120
rect 7708 3108 7720 3117
rect 11606 3108 11612 3120
rect 7708 3080 7753 3108
rect 7944 3080 11612 3108
rect 7708 3071 7720 3080
rect 7708 3068 7714 3071
rect 7834 3040 7840 3052
rect 6288 3012 7840 3040
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 7944 3049 7972 3080
rect 9784 3052 9812 3080
rect 7929 3043 7987 3049
rect 7929 3009 7941 3043
rect 7975 3009 7987 3043
rect 7929 3003 7987 3009
rect 8018 3000 8024 3052
rect 8076 3040 8082 3052
rect 8202 3040 8208 3052
rect 8076 3012 8121 3040
rect 8163 3012 8208 3040
rect 8076 3000 8082 3012
rect 8202 3000 8208 3012
rect 8260 3000 8266 3052
rect 9513 3043 9571 3049
rect 9513 3009 9525 3043
rect 9559 3040 9571 3043
rect 9559 3012 9720 3040
rect 9559 3009 9571 3012
rect 9513 3003 9571 3009
rect 3844 2944 4292 2972
rect 4801 2975 4859 2981
rect 3844 2932 3850 2944
rect 4801 2941 4813 2975
rect 4847 2941 4859 2975
rect 4801 2935 4859 2941
rect 4893 2975 4951 2981
rect 4893 2941 4905 2975
rect 4939 2972 4951 2975
rect 5442 2972 5448 2984
rect 4939 2944 5028 2972
rect 4939 2941 4951 2944
rect 4893 2935 4951 2941
rect 4065 2907 4123 2913
rect 4065 2904 4077 2907
rect 3620 2876 4077 2904
rect 4065 2873 4077 2876
rect 4111 2873 4123 2907
rect 4065 2867 4123 2873
rect 4246 2864 4252 2916
rect 4304 2904 4310 2916
rect 4816 2904 4844 2935
rect 5000 2916 5028 2944
rect 5101 2944 5448 2972
rect 4304 2876 4844 2904
rect 4304 2864 4310 2876
rect 4982 2864 4988 2916
rect 5040 2864 5046 2916
rect 1452 2808 1532 2836
rect 1765 2839 1823 2845
rect 1452 2796 1458 2808
rect 1765 2805 1777 2839
rect 1811 2836 1823 2839
rect 3160 2836 3188 2864
rect 1811 2808 3188 2836
rect 3421 2839 3479 2845
rect 1811 2805 1823 2808
rect 1765 2799 1823 2805
rect 3421 2805 3433 2839
rect 3467 2836 3479 2839
rect 5101 2836 5129 2944
rect 5442 2932 5448 2944
rect 5500 2932 5506 2984
rect 5718 2972 5724 2984
rect 5679 2944 5724 2972
rect 5718 2932 5724 2944
rect 5776 2932 5782 2984
rect 9692 2972 9720 3012
rect 9766 3000 9772 3052
rect 9824 3040 9830 3052
rect 9824 3012 9869 3040
rect 9824 3000 9830 3012
rect 10962 3000 10968 3052
rect 11020 3049 11026 3052
rect 11256 3049 11284 3080
rect 11606 3068 11612 3080
rect 11664 3108 11670 3120
rect 12544 3108 12572 3148
rect 13078 3136 13084 3148
rect 13136 3136 13142 3188
rect 14461 3179 14519 3185
rect 14461 3145 14473 3179
rect 14507 3176 14519 3179
rect 15562 3176 15568 3188
rect 14507 3148 15568 3176
rect 14507 3145 14519 3148
rect 14461 3139 14519 3145
rect 12710 3108 12716 3120
rect 11664 3080 12572 3108
rect 12671 3080 12716 3108
rect 11664 3068 11670 3080
rect 12710 3068 12716 3080
rect 12768 3068 12774 3120
rect 12986 3068 12992 3120
rect 13044 3108 13050 3120
rect 13326 3111 13384 3117
rect 13326 3108 13338 3111
rect 13044 3080 13338 3108
rect 13044 3068 13050 3080
rect 13326 3077 13338 3080
rect 13372 3077 13384 3111
rect 13326 3071 13384 3077
rect 13722 3068 13728 3120
rect 13780 3108 13786 3120
rect 14476 3108 14504 3139
rect 15562 3136 15568 3148
rect 15620 3136 15626 3188
rect 13780 3080 14504 3108
rect 13780 3068 13786 3080
rect 11020 3040 11032 3049
rect 11241 3043 11299 3049
rect 11020 3012 11192 3040
rect 11020 3003 11032 3012
rect 11020 3000 11026 3003
rect 11164 2972 11192 3012
rect 11241 3009 11253 3043
rect 11287 3009 11299 3043
rect 11241 3003 11299 3009
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 12529 3043 12587 3049
rect 11756 3012 12204 3040
rect 11756 3000 11762 3012
rect 12069 2975 12127 2981
rect 9692 2944 9904 2972
rect 11164 2944 11652 2972
rect 9876 2916 9904 2944
rect 5166 2864 5172 2916
rect 5224 2904 5230 2916
rect 6362 2904 6368 2916
rect 5224 2876 6368 2904
rect 5224 2864 5230 2876
rect 6362 2864 6368 2876
rect 6420 2904 6426 2916
rect 6549 2907 6607 2913
rect 6549 2904 6561 2907
rect 6420 2876 6561 2904
rect 6420 2864 6426 2876
rect 6549 2873 6561 2876
rect 6595 2873 6607 2907
rect 9858 2904 9864 2916
rect 9819 2876 9864 2904
rect 6549 2867 6607 2873
rect 9858 2864 9864 2876
rect 9916 2864 9922 2916
rect 11624 2904 11652 2944
rect 12069 2941 12081 2975
rect 12115 2941 12127 2975
rect 12176 2972 12204 3012
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 12897 3043 12955 3049
rect 12897 3009 12909 3043
rect 12943 3009 12955 3043
rect 13078 3040 13084 3052
rect 13039 3012 13084 3040
rect 12897 3003 12955 3009
rect 12345 2975 12403 2981
rect 12345 2972 12357 2975
rect 12176 2944 12357 2972
rect 12069 2935 12127 2941
rect 12345 2941 12357 2944
rect 12391 2941 12403 2975
rect 12544 2972 12572 3003
rect 12710 2972 12716 2984
rect 12544 2944 12716 2972
rect 12345 2935 12403 2941
rect 12084 2904 12112 2935
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 11624 2876 12112 2904
rect 3467 2808 5129 2836
rect 3467 2805 3479 2808
rect 3421 2799 3479 2805
rect 5258 2796 5264 2848
rect 5316 2836 5322 2848
rect 5997 2839 6055 2845
rect 5997 2836 6009 2839
rect 5316 2808 6009 2836
rect 5316 2796 5322 2808
rect 5997 2805 6009 2808
rect 6043 2805 6055 2839
rect 5997 2799 6055 2805
rect 8389 2839 8447 2845
rect 8389 2805 8401 2839
rect 8435 2836 8447 2839
rect 9030 2836 9036 2848
rect 8435 2808 9036 2836
rect 8435 2805 8447 2808
rect 8389 2799 8447 2805
rect 9030 2796 9036 2808
rect 9088 2836 9094 2848
rect 9582 2836 9588 2848
rect 9088 2808 9588 2836
rect 9088 2796 9094 2808
rect 9582 2796 9588 2808
rect 9640 2796 9646 2848
rect 11238 2796 11244 2848
rect 11296 2836 11302 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11296 2808 11529 2836
rect 11296 2796 11302 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 11517 2799 11575 2805
rect 11606 2796 11612 2848
rect 11664 2836 11670 2848
rect 12912 2836 12940 3003
rect 13078 3000 13084 3012
rect 13136 3000 13142 3052
rect 13814 3000 13820 3052
rect 13872 3040 13878 3052
rect 13872 3012 14596 3040
rect 13872 3000 13878 3012
rect 14568 2981 14596 3012
rect 14734 3000 14740 3052
rect 14792 3040 14798 3052
rect 14829 3043 14887 3049
rect 14829 3040 14841 3043
rect 14792 3012 14841 3040
rect 14792 3000 14798 3012
rect 14829 3009 14841 3012
rect 14875 3009 14887 3043
rect 15470 3040 15476 3052
rect 15431 3012 15476 3040
rect 14829 3003 14887 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 14553 2975 14611 2981
rect 14553 2941 14565 2975
rect 14599 2972 14611 2975
rect 16022 2972 16028 2984
rect 14599 2944 16028 2972
rect 14599 2941 14611 2944
rect 14553 2935 14611 2941
rect 16022 2932 16028 2944
rect 16080 2932 16086 2984
rect 16206 2904 16212 2916
rect 14016 2876 16212 2904
rect 14016 2836 14044 2876
rect 16206 2864 16212 2876
rect 16264 2864 16270 2916
rect 11664 2808 14044 2836
rect 15657 2839 15715 2845
rect 11664 2796 11670 2808
rect 15657 2805 15669 2839
rect 15703 2836 15715 2839
rect 16942 2836 16948 2848
rect 15703 2808 16948 2836
rect 15703 2805 15715 2808
rect 15657 2799 15715 2805
rect 16942 2796 16948 2808
rect 17000 2796 17006 2848
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 3510 2632 3516 2644
rect 1627 2604 3516 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 3510 2592 3516 2604
rect 3568 2592 3574 2644
rect 4338 2592 4344 2644
rect 4396 2632 4402 2644
rect 4525 2635 4583 2641
rect 4525 2632 4537 2635
rect 4396 2604 4537 2632
rect 4396 2592 4402 2604
rect 4525 2601 4537 2604
rect 4571 2601 4583 2635
rect 4525 2595 4583 2601
rect 5629 2635 5687 2641
rect 5629 2601 5641 2635
rect 5675 2632 5687 2635
rect 7742 2632 7748 2644
rect 5675 2604 7748 2632
rect 5675 2601 5687 2604
rect 5629 2595 5687 2601
rect 7742 2592 7748 2604
rect 7800 2592 7806 2644
rect 8113 2635 8171 2641
rect 8113 2601 8125 2635
rect 8159 2632 8171 2635
rect 9030 2632 9036 2644
rect 8159 2604 8892 2632
rect 8991 2604 9036 2632
rect 8159 2601 8171 2604
rect 8113 2595 8171 2601
rect 2041 2567 2099 2573
rect 2041 2533 2053 2567
rect 2087 2533 2099 2567
rect 2041 2527 2099 2533
rect 2685 2567 2743 2573
rect 2685 2533 2697 2567
rect 2731 2564 2743 2567
rect 3970 2564 3976 2576
rect 2731 2536 3976 2564
rect 2731 2533 2743 2536
rect 2685 2527 2743 2533
rect 2056 2496 2084 2527
rect 3970 2524 3976 2536
rect 4028 2524 4034 2576
rect 4249 2567 4307 2573
rect 4249 2533 4261 2567
rect 4295 2564 4307 2567
rect 5534 2564 5540 2576
rect 4295 2536 5540 2564
rect 4295 2533 4307 2536
rect 4249 2527 4307 2533
rect 5534 2524 5540 2536
rect 5592 2524 5598 2576
rect 8205 2567 8263 2573
rect 8205 2564 8217 2567
rect 6196 2536 8217 2564
rect 4338 2496 4344 2508
rect 2056 2468 4344 2496
rect 4338 2456 4344 2468
rect 4396 2456 4402 2508
rect 5166 2496 5172 2508
rect 5127 2468 5172 2496
rect 5166 2456 5172 2468
rect 5224 2456 5230 2508
rect 1578 2388 1584 2440
rect 1636 2428 1642 2440
rect 1765 2431 1823 2437
rect 1765 2428 1777 2431
rect 1636 2400 1777 2428
rect 1636 2388 1642 2400
rect 1765 2397 1777 2400
rect 1811 2397 1823 2431
rect 1765 2391 1823 2397
rect 1854 2388 1860 2440
rect 1912 2428 1918 2440
rect 2498 2428 2504 2440
rect 1912 2400 1957 2428
rect 2459 2400 2504 2428
rect 1912 2388 1918 2400
rect 2498 2388 2504 2400
rect 2556 2388 2562 2440
rect 2869 2431 2927 2437
rect 2869 2397 2881 2431
rect 2915 2397 2927 2431
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 2869 2391 2927 2397
rect 2884 2360 2912 2391
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3602 2428 3608 2440
rect 3563 2400 3608 2428
rect 3602 2388 3608 2400
rect 3660 2388 3666 2440
rect 4062 2428 4068 2440
rect 4023 2400 4068 2428
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 5258 2428 5264 2440
rect 4479 2400 5264 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5810 2428 5816 2440
rect 5771 2400 5816 2428
rect 5810 2388 5816 2400
rect 5868 2388 5874 2440
rect 6196 2437 6224 2536
rect 8205 2533 8217 2536
rect 8251 2533 8263 2567
rect 8205 2527 8263 2533
rect 8294 2524 8300 2576
rect 8352 2564 8358 2576
rect 8481 2567 8539 2573
rect 8481 2564 8493 2567
rect 8352 2536 8493 2564
rect 8352 2524 8358 2536
rect 8481 2533 8493 2536
rect 8527 2533 8539 2567
rect 8864 2564 8892 2604
rect 9030 2592 9036 2604
rect 9088 2592 9094 2644
rect 10042 2592 10048 2644
rect 10100 2632 10106 2644
rect 10413 2635 10471 2641
rect 10413 2632 10425 2635
rect 10100 2604 10425 2632
rect 10100 2592 10106 2604
rect 10413 2601 10425 2604
rect 10459 2632 10471 2635
rect 10778 2632 10784 2644
rect 10459 2604 10784 2632
rect 10459 2601 10471 2604
rect 10413 2595 10471 2601
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 10962 2592 10968 2644
rect 11020 2632 11026 2644
rect 11020 2604 11836 2632
rect 11020 2592 11026 2604
rect 9122 2564 9128 2576
rect 8864 2536 9128 2564
rect 8481 2527 8539 2533
rect 9122 2524 9128 2536
rect 9180 2524 9186 2576
rect 10505 2567 10563 2573
rect 10505 2564 10517 2567
rect 9416 2536 10517 2564
rect 8110 2496 8116 2508
rect 6886 2468 8116 2496
rect 6181 2431 6239 2437
rect 6181 2397 6193 2431
rect 6227 2397 6239 2431
rect 6181 2391 6239 2397
rect 6472 2400 6776 2428
rect 3326 2360 3332 2372
rect 2884 2332 3332 2360
rect 3326 2320 3332 2332
rect 3384 2320 3390 2372
rect 4614 2360 4620 2372
rect 3436 2332 4620 2360
rect 2314 2292 2320 2304
rect 2275 2264 2320 2292
rect 2314 2252 2320 2264
rect 2372 2252 2378 2304
rect 3050 2292 3056 2304
rect 3011 2264 3056 2292
rect 3050 2252 3056 2264
rect 3108 2252 3114 2304
rect 3436 2301 3464 2332
rect 4614 2320 4620 2332
rect 4672 2320 4678 2372
rect 4985 2363 5043 2369
rect 4985 2329 4997 2363
rect 5031 2360 5043 2363
rect 5350 2360 5356 2372
rect 5031 2332 5356 2360
rect 5031 2329 5043 2332
rect 4985 2323 5043 2329
rect 5350 2320 5356 2332
rect 5408 2320 5414 2372
rect 6472 2360 6500 2400
rect 6012 2332 6500 2360
rect 3421 2295 3479 2301
rect 3421 2261 3433 2295
rect 3467 2261 3479 2295
rect 3878 2292 3884 2304
rect 3839 2264 3884 2292
rect 3421 2255 3479 2261
rect 3878 2252 3884 2264
rect 3936 2252 3942 2304
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4893 2295 4951 2301
rect 4893 2292 4905 2295
rect 4212 2264 4905 2292
rect 4212 2252 4218 2264
rect 4893 2261 4905 2264
rect 4939 2261 4951 2295
rect 5442 2292 5448 2304
rect 5403 2264 5448 2292
rect 4893 2255 4951 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 6012 2301 6040 2332
rect 6546 2320 6552 2372
rect 6604 2360 6610 2372
rect 6748 2360 6776 2400
rect 6886 2360 6914 2468
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 6953 2431 7011 2437
rect 6953 2397 6965 2431
rect 6999 2428 7011 2431
rect 7374 2428 7380 2440
rect 6999 2400 7380 2428
rect 6999 2397 7011 2400
rect 6953 2391 7011 2397
rect 7374 2388 7380 2400
rect 7432 2388 7438 2440
rect 7466 2388 7472 2440
rect 7524 2437 7530 2440
rect 7524 2431 7538 2437
rect 7526 2428 7538 2431
rect 7526 2400 7569 2428
rect 7526 2397 7538 2400
rect 7524 2391 7538 2397
rect 7524 2388 7530 2391
rect 8386 2388 8392 2440
rect 8444 2428 8450 2440
rect 9214 2428 9220 2440
rect 8444 2400 9220 2428
rect 8444 2388 8450 2400
rect 9214 2388 9220 2400
rect 9272 2388 9278 2440
rect 9416 2437 9444 2536
rect 10505 2533 10517 2536
rect 10551 2533 10563 2567
rect 10505 2527 10563 2533
rect 10686 2524 10692 2576
rect 10744 2564 10750 2576
rect 10744 2536 11560 2564
rect 10744 2524 10750 2536
rect 9582 2496 9588 2508
rect 9543 2468 9588 2496
rect 9582 2456 9588 2468
rect 9640 2456 9646 2508
rect 9858 2456 9864 2508
rect 9916 2496 9922 2508
rect 11532 2505 11560 2536
rect 11057 2499 11115 2505
rect 11057 2496 11069 2499
rect 9916 2468 11069 2496
rect 9916 2456 9922 2468
rect 11057 2465 11069 2468
rect 11103 2465 11115 2499
rect 11057 2459 11115 2465
rect 11517 2499 11575 2505
rect 11517 2465 11529 2499
rect 11563 2496 11575 2499
rect 11698 2496 11704 2508
rect 11563 2468 11704 2496
rect 11563 2465 11575 2468
rect 11517 2459 11575 2465
rect 11698 2456 11704 2468
rect 11756 2456 11762 2508
rect 11808 2505 11836 2604
rect 13722 2592 13728 2644
rect 13780 2632 13786 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 13780 2604 15485 2632
rect 13780 2592 13786 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 15473 2595 15531 2601
rect 15010 2564 15016 2576
rect 13280 2536 15016 2564
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2465 11851 2499
rect 11793 2459 11851 2465
rect 12526 2456 12532 2508
rect 12584 2496 12590 2508
rect 13280 2505 13308 2536
rect 15010 2524 15016 2536
rect 15068 2524 15074 2576
rect 13265 2499 13323 2505
rect 13265 2496 13277 2499
rect 12584 2468 13277 2496
rect 12584 2456 12590 2468
rect 13265 2465 13277 2468
rect 13311 2465 13323 2499
rect 13265 2459 13323 2465
rect 13725 2499 13783 2505
rect 13725 2465 13737 2499
rect 13771 2496 13783 2499
rect 15470 2496 15476 2508
rect 13771 2468 15476 2496
rect 13771 2465 13783 2468
rect 13725 2459 13783 2465
rect 15470 2456 15476 2468
rect 15528 2456 15534 2508
rect 9401 2431 9459 2437
rect 9401 2397 9413 2431
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 9493 2431 9551 2437
rect 9493 2397 9505 2431
rect 9539 2428 9551 2431
rect 9674 2428 9680 2440
rect 9539 2400 9680 2428
rect 9539 2397 9551 2400
rect 9493 2391 9551 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10042 2428 10048 2440
rect 10003 2400 10048 2428
rect 10042 2388 10048 2400
rect 10100 2388 10106 2440
rect 10226 2428 10232 2440
rect 10187 2400 10232 2428
rect 10226 2388 10232 2400
rect 10284 2388 10290 2440
rect 10873 2431 10931 2437
rect 10873 2397 10885 2431
rect 10919 2428 10931 2431
rect 11238 2428 11244 2440
rect 10919 2400 11244 2428
rect 10919 2397 10931 2400
rect 10873 2391 10931 2397
rect 11238 2388 11244 2400
rect 11296 2388 11302 2440
rect 12986 2428 12992 2440
rect 12947 2400 12992 2428
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13906 2428 13912 2440
rect 13867 2400 13912 2428
rect 13906 2388 13912 2400
rect 13964 2388 13970 2440
rect 14550 2428 14556 2440
rect 14511 2400 14556 2428
rect 14550 2388 14556 2400
rect 14608 2388 14614 2440
rect 14826 2428 14832 2440
rect 14787 2400 14832 2428
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 7190 2360 7196 2372
rect 6604 2332 6649 2360
rect 6748 2332 6914 2360
rect 7151 2332 7196 2360
rect 6604 2320 6610 2332
rect 7190 2320 7196 2332
rect 7248 2320 7254 2372
rect 8018 2360 8024 2372
rect 7300 2332 8024 2360
rect 5997 2295 6055 2301
rect 5997 2261 6009 2295
rect 6043 2261 6055 2295
rect 5997 2255 6055 2261
rect 6362 2252 6368 2304
rect 6420 2292 6426 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 6420 2264 6469 2292
rect 6420 2252 6426 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 6825 2295 6883 2301
rect 6825 2261 6837 2295
rect 6871 2292 6883 2295
rect 7006 2292 7012 2304
rect 6871 2264 7012 2292
rect 6871 2261 6883 2264
rect 6825 2255 6883 2261
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7300 2301 7328 2332
rect 8018 2320 8024 2332
rect 8076 2360 8082 2372
rect 8665 2363 8723 2369
rect 8665 2360 8677 2363
rect 8076 2332 8677 2360
rect 8076 2320 8082 2332
rect 8665 2329 8677 2332
rect 8711 2329 8723 2363
rect 8665 2323 8723 2329
rect 10965 2363 11023 2369
rect 10965 2329 10977 2363
rect 11011 2360 11023 2363
rect 11882 2360 11888 2372
rect 11011 2332 11888 2360
rect 11011 2329 11023 2332
rect 10965 2323 11023 2329
rect 11882 2320 11888 2332
rect 11940 2320 11946 2372
rect 12710 2320 12716 2372
rect 12768 2360 12774 2372
rect 13538 2360 13544 2372
rect 12768 2332 13544 2360
rect 12768 2320 12774 2332
rect 13538 2320 13544 2332
rect 13596 2360 13602 2372
rect 14277 2363 14335 2369
rect 14277 2360 14289 2363
rect 13596 2332 14289 2360
rect 13596 2320 13602 2332
rect 14277 2329 14289 2332
rect 14323 2329 14335 2363
rect 14277 2323 14335 2329
rect 7285 2295 7343 2301
rect 7285 2261 7297 2295
rect 7331 2261 7343 2295
rect 7285 2255 7343 2261
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 9953 2295 10011 2301
rect 9953 2292 9965 2295
rect 7708 2264 9965 2292
rect 7708 2252 7714 2264
rect 9953 2261 9965 2264
rect 9999 2261 10011 2295
rect 9953 2255 10011 2261
rect 10042 2252 10048 2304
rect 10100 2292 10106 2304
rect 13722 2292 13728 2304
rect 10100 2264 13728 2292
rect 10100 2252 10106 2264
rect 13722 2252 13728 2264
rect 13780 2252 13786 2304
rect 14182 2292 14188 2304
rect 14143 2264 14188 2292
rect 14182 2252 14188 2264
rect 14240 2292 14246 2304
rect 16390 2292 16396 2304
rect 14240 2264 16396 2292
rect 14240 2252 14246 2264
rect 16390 2252 16396 2264
rect 16448 2252 16454 2304
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 2314 2048 2320 2100
rect 2372 2088 2378 2100
rect 5166 2088 5172 2100
rect 2372 2060 5172 2088
rect 2372 2048 2378 2060
rect 5166 2048 5172 2060
rect 5224 2048 5230 2100
rect 5442 2048 5448 2100
rect 5500 2088 5506 2100
rect 9766 2088 9772 2100
rect 5500 2060 9772 2088
rect 5500 2048 5506 2060
rect 9766 2048 9772 2060
rect 9824 2088 9830 2100
rect 10226 2088 10232 2100
rect 9824 2060 10232 2088
rect 9824 2048 9830 2060
rect 10226 2048 10232 2060
rect 10284 2048 10290 2100
rect 13538 2048 13544 2100
rect 13596 2088 13602 2100
rect 14550 2088 14556 2100
rect 13596 2060 14556 2088
rect 13596 2048 13602 2060
rect 14550 2048 14556 2060
rect 14608 2048 14614 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 5994 2020 6000 2032
rect 3108 1992 6000 2020
rect 3108 1980 3114 1992
rect 5994 1980 6000 1992
rect 6052 1980 6058 2032
rect 11422 1980 11428 2032
rect 11480 2020 11486 2032
rect 14182 2020 14188 2032
rect 11480 1992 14188 2020
rect 11480 1980 11486 1992
rect 14182 1980 14188 1992
rect 14240 1980 14246 2032
rect 3602 1912 3608 1964
rect 3660 1952 3666 1964
rect 9306 1952 9312 1964
rect 3660 1924 9312 1952
rect 3660 1912 3666 1924
rect 9306 1912 9312 1924
rect 9364 1912 9370 1964
rect 2498 1844 2504 1896
rect 2556 1884 2562 1896
rect 4522 1884 4528 1896
rect 2556 1856 4528 1884
rect 2556 1844 2562 1856
rect 4522 1844 4528 1856
rect 4580 1844 4586 1896
rect 6546 1844 6552 1896
rect 6604 1884 6610 1896
rect 8846 1884 8852 1896
rect 6604 1856 8852 1884
rect 6604 1844 6610 1856
rect 8846 1844 8852 1856
rect 8904 1844 8910 1896
rect 9214 1844 9220 1896
rect 9272 1884 9278 1896
rect 13354 1884 13360 1896
rect 9272 1856 13360 1884
rect 9272 1844 9278 1856
rect 13354 1844 13360 1856
rect 13412 1844 13418 1896
rect 3694 1776 3700 1828
rect 3752 1816 3758 1828
rect 6362 1816 6368 1828
rect 3752 1788 6368 1816
rect 3752 1776 3758 1788
rect 6362 1776 6368 1788
rect 6420 1816 6426 1828
rect 8202 1816 8208 1828
rect 6420 1788 8208 1816
rect 6420 1776 6426 1788
rect 8202 1776 8208 1788
rect 8260 1776 8266 1828
rect 5534 1708 5540 1760
rect 5592 1748 5598 1760
rect 7282 1748 7288 1760
rect 5592 1720 7288 1748
rect 5592 1708 5598 1720
rect 7282 1708 7288 1720
rect 7340 1708 7346 1760
rect 7374 1708 7380 1760
rect 7432 1748 7438 1760
rect 10318 1748 10324 1760
rect 7432 1720 10324 1748
rect 7432 1708 7438 1720
rect 10318 1708 10324 1720
rect 10376 1708 10382 1760
rect 1670 1640 1676 1692
rect 1728 1680 1734 1692
rect 8294 1680 8300 1692
rect 1728 1652 8300 1680
rect 1728 1640 1734 1652
rect 8294 1640 8300 1652
rect 8352 1640 8358 1692
rect 3878 1572 3884 1624
rect 3936 1612 3942 1624
rect 6822 1612 6828 1624
rect 3936 1584 6828 1612
rect 3936 1572 3942 1584
rect 6822 1572 6828 1584
rect 6880 1572 6886 1624
<< via1 >>
rect 6460 17620 6512 17672
rect 8392 17620 8444 17672
rect 5540 17552 5592 17604
rect 6736 17552 6788 17604
rect 7288 17552 7340 17604
rect 12532 17552 12584 17604
rect 204 17484 256 17536
rect 3792 17484 3844 17536
rect 9036 17484 9088 17536
rect 11428 17484 11480 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 1768 17280 1820 17332
rect 2228 17280 2280 17332
rect 2596 17280 2648 17332
rect 3056 17280 3108 17332
rect 3424 17280 3476 17332
rect 4620 17280 4672 17332
rect 5908 17280 5960 17332
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 3700 17212 3752 17264
rect 5632 17212 5684 17264
rect 3148 17144 3200 17196
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 3792 17187 3844 17196
rect 3792 17153 3793 17187
rect 3793 17153 3827 17187
rect 3827 17153 3844 17187
rect 4344 17187 4396 17196
rect 3792 17144 3844 17153
rect 3240 17076 3292 17128
rect 4344 17153 4353 17187
rect 4353 17153 4387 17187
rect 4387 17153 4396 17187
rect 4344 17144 4396 17153
rect 4436 17187 4488 17196
rect 4436 17153 4445 17187
rect 4445 17153 4479 17187
rect 4479 17153 4488 17187
rect 4436 17144 4488 17153
rect 4620 17144 4672 17196
rect 5172 17187 5224 17196
rect 5172 17153 5181 17187
rect 5181 17153 5215 17187
rect 5215 17153 5224 17187
rect 5172 17144 5224 17153
rect 5632 17076 5684 17128
rect 3332 17008 3384 17060
rect 4252 17008 4304 17060
rect 5448 17008 5500 17060
rect 3976 16983 4028 16992
rect 3976 16949 3985 16983
rect 3985 16949 4019 16983
rect 4019 16949 4028 16983
rect 3976 16940 4028 16949
rect 5540 16940 5592 16992
rect 7104 17212 7156 17264
rect 8852 17280 8904 17332
rect 7564 17212 7616 17264
rect 11520 17212 11572 17264
rect 11704 17255 11756 17264
rect 11704 17221 11713 17255
rect 11713 17221 11747 17255
rect 11747 17221 11756 17255
rect 11704 17212 11756 17221
rect 5908 17187 5960 17196
rect 5908 17153 5917 17187
rect 5917 17153 5951 17187
rect 5951 17153 5960 17187
rect 5908 17144 5960 17153
rect 6000 17144 6052 17196
rect 7196 17144 7248 17196
rect 7380 17187 7432 17196
rect 7380 17153 7389 17187
rect 7389 17153 7423 17187
rect 7423 17153 7432 17187
rect 7380 17144 7432 17153
rect 6828 17008 6880 17060
rect 7472 17076 7524 17128
rect 9312 17144 9364 17196
rect 9588 17187 9640 17196
rect 9588 17153 9597 17187
rect 9597 17153 9631 17187
rect 9631 17153 9640 17187
rect 9588 17144 9640 17153
rect 10048 17187 10100 17196
rect 10048 17153 10057 17187
rect 10057 17153 10091 17187
rect 10091 17153 10100 17187
rect 10048 17144 10100 17153
rect 11888 17187 11940 17196
rect 11888 17153 11897 17187
rect 11897 17153 11931 17187
rect 11931 17153 11940 17187
rect 11888 17144 11940 17153
rect 12624 17144 12676 17196
rect 8116 17076 8168 17128
rect 8208 17008 8260 17060
rect 6460 16940 6512 16992
rect 7104 16940 7156 16992
rect 8024 16940 8076 16992
rect 9220 17008 9272 17060
rect 8944 16983 8996 16992
rect 8944 16949 8953 16983
rect 8953 16949 8987 16983
rect 8987 16949 8996 16983
rect 8944 16940 8996 16949
rect 11060 17119 11112 17128
rect 11060 17085 11069 17119
rect 11069 17085 11103 17119
rect 11103 17085 11112 17119
rect 11060 17076 11112 17085
rect 10692 17008 10744 17060
rect 11152 17008 11204 17060
rect 11428 17076 11480 17128
rect 11704 17076 11756 17128
rect 12072 17076 12124 17128
rect 12440 17119 12492 17128
rect 12440 17085 12449 17119
rect 12449 17085 12483 17119
rect 12483 17085 12492 17119
rect 12440 17076 12492 17085
rect 15752 17212 15804 17264
rect 14832 17144 14884 17196
rect 13452 17076 13504 17128
rect 13820 17076 13872 17128
rect 15844 17008 15896 17060
rect 10140 16940 10192 16992
rect 10232 16940 10284 16992
rect 10784 16940 10836 16992
rect 11888 16940 11940 16992
rect 12532 16940 12584 16992
rect 13084 16940 13136 16992
rect 15384 16940 15436 16992
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 1860 16779 1912 16788
rect 1860 16745 1869 16779
rect 1869 16745 1903 16779
rect 1903 16745 1912 16779
rect 1860 16736 1912 16745
rect 2688 16736 2740 16788
rect 3792 16736 3844 16788
rect 4436 16779 4488 16788
rect 4436 16745 4445 16779
rect 4445 16745 4479 16779
rect 4479 16745 4488 16779
rect 4436 16736 4488 16745
rect 5172 16736 5224 16788
rect 5816 16736 5868 16788
rect 7104 16736 7156 16788
rect 8852 16736 8904 16788
rect 9588 16736 9640 16788
rect 10692 16779 10744 16788
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 11060 16736 11112 16788
rect 1492 16711 1544 16720
rect 1492 16677 1501 16711
rect 1501 16677 1535 16711
rect 1535 16677 1544 16711
rect 1492 16668 1544 16677
rect 3148 16668 3200 16720
rect 6000 16668 6052 16720
rect 1952 16532 2004 16584
rect 2412 16575 2464 16584
rect 2412 16541 2421 16575
rect 2421 16541 2455 16575
rect 2455 16541 2464 16575
rect 2412 16532 2464 16541
rect 2504 16575 2556 16584
rect 2504 16541 2513 16575
rect 2513 16541 2547 16575
rect 2547 16541 2556 16575
rect 2504 16532 2556 16541
rect 2964 16532 3016 16584
rect 2596 16464 2648 16516
rect 3516 16532 3568 16584
rect 3792 16464 3844 16516
rect 940 16396 992 16448
rect 4528 16532 4580 16584
rect 6184 16600 6236 16652
rect 6920 16668 6972 16720
rect 11336 16668 11388 16720
rect 5172 16532 5224 16584
rect 6368 16532 6420 16584
rect 8116 16600 8168 16652
rect 7748 16532 7800 16584
rect 8300 16532 8352 16584
rect 11796 16600 11848 16652
rect 11060 16532 11112 16584
rect 13820 16600 13872 16652
rect 7840 16464 7892 16516
rect 5080 16396 5132 16448
rect 6092 16439 6144 16448
rect 6092 16405 6101 16439
rect 6101 16405 6135 16439
rect 6135 16405 6144 16439
rect 6092 16396 6144 16405
rect 6460 16439 6512 16448
rect 6460 16405 6469 16439
rect 6469 16405 6503 16439
rect 6503 16405 6512 16439
rect 6460 16396 6512 16405
rect 8024 16396 8076 16448
rect 9220 16464 9272 16516
rect 9588 16507 9640 16516
rect 9588 16473 9622 16507
rect 9622 16473 9640 16507
rect 9588 16464 9640 16473
rect 10140 16464 10192 16516
rect 11888 16464 11940 16516
rect 13176 16507 13228 16516
rect 13176 16473 13194 16507
rect 13194 16473 13228 16507
rect 13176 16464 13228 16473
rect 13544 16464 13596 16516
rect 16028 16464 16080 16516
rect 9956 16396 10008 16448
rect 10784 16439 10836 16448
rect 10784 16405 10793 16439
rect 10793 16405 10827 16439
rect 10827 16405 10836 16439
rect 10784 16396 10836 16405
rect 11060 16396 11112 16448
rect 11428 16396 11480 16448
rect 12532 16396 12584 16448
rect 13360 16396 13412 16448
rect 15476 16439 15528 16448
rect 15476 16405 15485 16439
rect 15485 16405 15519 16439
rect 15519 16405 15528 16439
rect 15476 16396 15528 16405
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 572 16192 624 16244
rect 2136 16192 2188 16244
rect 3240 16192 3292 16244
rect 3608 16192 3660 16244
rect 4344 16235 4396 16244
rect 4344 16201 4353 16235
rect 4353 16201 4387 16235
rect 4387 16201 4396 16235
rect 4344 16192 4396 16201
rect 4620 16192 4672 16244
rect 5540 16192 5592 16244
rect 5908 16192 5960 16244
rect 6368 16235 6420 16244
rect 6368 16201 6377 16235
rect 6377 16201 6411 16235
rect 6411 16201 6420 16235
rect 6368 16192 6420 16201
rect 7012 16192 7064 16244
rect 7840 16235 7892 16244
rect 2228 16124 2280 16176
rect 1584 16056 1636 16108
rect 1768 16099 1820 16108
rect 1768 16065 1777 16099
rect 1777 16065 1811 16099
rect 1811 16065 1820 16099
rect 1768 16056 1820 16065
rect 2596 16056 2648 16108
rect 2320 15988 2372 16040
rect 3240 16056 3292 16108
rect 4436 16124 4488 16176
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 3792 16056 3844 16108
rect 3976 16056 4028 16108
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 2964 15988 3016 16040
rect 4988 16056 5040 16108
rect 4712 15988 4764 16040
rect 5356 16056 5408 16108
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 7932 16192 7984 16244
rect 9128 16192 9180 16244
rect 10784 16192 10836 16244
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 12532 16192 12584 16244
rect 14556 16192 14608 16244
rect 5540 15988 5592 16040
rect 1400 15920 1452 15972
rect 2412 15920 2464 15972
rect 3700 15963 3752 15972
rect 3700 15929 3709 15963
rect 3709 15929 3743 15963
rect 3743 15929 3752 15963
rect 3700 15920 3752 15929
rect 3884 15920 3936 15972
rect 6184 16056 6236 16108
rect 7472 16099 7524 16108
rect 7472 16065 7490 16099
rect 7490 16065 7524 16099
rect 7472 16056 7524 16065
rect 7748 16099 7800 16108
rect 7748 16065 7757 16099
rect 7757 16065 7791 16099
rect 7791 16065 7800 16099
rect 7748 16056 7800 16065
rect 8944 16124 8996 16176
rect 9220 16124 9272 16176
rect 11244 16167 11296 16176
rect 8300 16056 8352 16108
rect 10140 15988 10192 16040
rect 10692 16056 10744 16108
rect 11244 16133 11253 16167
rect 11253 16133 11287 16167
rect 11287 16133 11296 16167
rect 11244 16124 11296 16133
rect 12900 16124 12952 16176
rect 16580 16192 16632 16244
rect 15660 16167 15712 16176
rect 15660 16133 15669 16167
rect 15669 16133 15703 16167
rect 15703 16133 15712 16167
rect 15660 16124 15712 16133
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 6276 15920 6328 15972
rect 9956 15920 10008 15972
rect 11520 15988 11572 16040
rect 11980 16031 12032 16040
rect 11980 15997 11989 16031
rect 11989 15997 12023 16031
rect 12023 15997 12032 16031
rect 11980 15988 12032 15997
rect 13176 16056 13228 16108
rect 13268 16056 13320 16108
rect 13544 16056 13596 16108
rect 11060 15963 11112 15972
rect 11060 15929 11069 15963
rect 11069 15929 11103 15963
rect 11103 15929 11112 15963
rect 11060 15920 11112 15929
rect 11336 15920 11388 15972
rect 15568 15988 15620 16040
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 3608 15895 3660 15904
rect 3608 15861 3617 15895
rect 3617 15861 3651 15895
rect 3651 15861 3660 15895
rect 3608 15852 3660 15861
rect 5724 15852 5776 15904
rect 6000 15852 6052 15904
rect 8116 15852 8168 15904
rect 9588 15852 9640 15904
rect 9772 15895 9824 15904
rect 9772 15861 9781 15895
rect 9781 15861 9815 15895
rect 9815 15861 9824 15895
rect 9772 15852 9824 15861
rect 10784 15895 10836 15904
rect 10784 15861 10793 15895
rect 10793 15861 10827 15895
rect 10827 15861 10836 15895
rect 10784 15852 10836 15861
rect 11520 15852 11572 15904
rect 13912 15920 13964 15972
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 1584 15648 1636 15700
rect 1768 15691 1820 15700
rect 1768 15657 1777 15691
rect 1777 15657 1811 15691
rect 1811 15657 1820 15691
rect 1768 15648 1820 15657
rect 1952 15648 2004 15700
rect 2504 15648 2556 15700
rect 2688 15691 2740 15700
rect 2688 15657 2697 15691
rect 2697 15657 2731 15691
rect 2731 15657 2740 15691
rect 2688 15648 2740 15657
rect 3332 15648 3384 15700
rect 3608 15691 3660 15700
rect 3608 15657 3617 15691
rect 3617 15657 3651 15691
rect 3651 15657 3660 15691
rect 3608 15648 3660 15657
rect 4436 15648 4488 15700
rect 4528 15648 4580 15700
rect 5264 15648 5316 15700
rect 6184 15648 6236 15700
rect 7380 15648 7432 15700
rect 9956 15691 10008 15700
rect 9956 15657 9965 15691
rect 9965 15657 9999 15691
rect 9999 15657 10008 15691
rect 9956 15648 10008 15657
rect 10048 15648 10100 15700
rect 13268 15648 13320 15700
rect 15384 15648 15436 15700
rect 2596 15580 2648 15632
rect 4068 15623 4120 15632
rect 4068 15589 4077 15623
rect 4077 15589 4111 15623
rect 4111 15589 4120 15623
rect 4068 15580 4120 15589
rect 4528 15512 4580 15564
rect 7012 15580 7064 15632
rect 1952 15487 2004 15496
rect 1952 15453 1961 15487
rect 1961 15453 1995 15487
rect 1995 15453 2004 15487
rect 1952 15444 2004 15453
rect 2320 15487 2372 15496
rect 2320 15453 2329 15487
rect 2329 15453 2363 15487
rect 2363 15453 2372 15487
rect 2320 15444 2372 15453
rect 2504 15444 2556 15496
rect 3148 15487 3200 15496
rect 3148 15453 3157 15487
rect 3157 15453 3191 15487
rect 3191 15453 3200 15487
rect 3148 15444 3200 15453
rect 4436 15444 4488 15496
rect 5724 15444 5776 15496
rect 3424 15308 3476 15360
rect 4344 15308 4396 15360
rect 9772 15512 9824 15564
rect 9956 15512 10008 15564
rect 10784 15580 10836 15632
rect 7104 15444 7156 15496
rect 7288 15487 7340 15496
rect 7288 15453 7297 15487
rect 7297 15453 7331 15487
rect 7331 15453 7340 15487
rect 7288 15444 7340 15453
rect 7564 15487 7616 15496
rect 7564 15453 7573 15487
rect 7573 15453 7607 15487
rect 7607 15453 7616 15487
rect 7564 15444 7616 15453
rect 9128 15487 9180 15496
rect 9128 15453 9137 15487
rect 9137 15453 9171 15487
rect 9171 15453 9180 15487
rect 9128 15444 9180 15453
rect 10968 15512 11020 15564
rect 11336 15512 11388 15564
rect 11704 15512 11756 15564
rect 13728 15580 13780 15632
rect 13636 15512 13688 15564
rect 14924 15512 14976 15564
rect 12992 15444 13044 15496
rect 14188 15444 14240 15496
rect 14464 15444 14516 15496
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 8116 15376 8168 15428
rect 9036 15376 9088 15428
rect 5448 15308 5500 15360
rect 7380 15308 7432 15360
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 9496 15351 9548 15360
rect 9496 15317 9505 15351
rect 9505 15317 9539 15351
rect 9539 15317 9548 15351
rect 9496 15308 9548 15317
rect 10048 15351 10100 15360
rect 10048 15317 10057 15351
rect 10057 15317 10091 15351
rect 10091 15317 10100 15351
rect 10048 15308 10100 15317
rect 10232 15308 10284 15360
rect 10692 15376 10744 15428
rect 10784 15308 10836 15360
rect 11336 15351 11388 15360
rect 11336 15317 11345 15351
rect 11345 15317 11379 15351
rect 11379 15317 11388 15351
rect 11336 15308 11388 15317
rect 11520 15308 11572 15360
rect 15936 15444 15988 15496
rect 16120 15444 16172 15496
rect 15660 15419 15712 15428
rect 15660 15385 15669 15419
rect 15669 15385 15703 15419
rect 15703 15385 15712 15419
rect 15660 15376 15712 15385
rect 12900 15308 12952 15360
rect 13084 15351 13136 15360
rect 13084 15317 13093 15351
rect 13093 15317 13127 15351
rect 13127 15317 13136 15351
rect 13084 15308 13136 15317
rect 13268 15308 13320 15360
rect 13636 15351 13688 15360
rect 13636 15317 13645 15351
rect 13645 15317 13679 15351
rect 13679 15317 13688 15351
rect 13636 15308 13688 15317
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 4528 15104 4580 15156
rect 5816 15147 5868 15156
rect 5816 15113 5825 15147
rect 5825 15113 5859 15147
rect 5859 15113 5868 15147
rect 5816 15104 5868 15113
rect 6092 15104 6144 15156
rect 6460 15104 6512 15156
rect 6920 15104 6972 15156
rect 7288 15104 7340 15156
rect 9496 15147 9548 15156
rect 9496 15113 9505 15147
rect 9505 15113 9539 15147
rect 9539 15113 9548 15147
rect 9496 15104 9548 15113
rect 10048 15104 10100 15156
rect 10876 15104 10928 15156
rect 10968 15104 11020 15156
rect 11980 15104 12032 15156
rect 2688 15011 2740 15020
rect 5724 15036 5776 15088
rect 2688 14977 2706 15011
rect 2706 14977 2740 15011
rect 2688 14968 2740 14977
rect 3332 15011 3384 15020
rect 3332 14977 3366 15011
rect 3366 14977 3384 15011
rect 3332 14968 3384 14977
rect 4252 14968 4304 15020
rect 5172 14968 5224 15020
rect 5356 14968 5408 15020
rect 5448 14968 5500 15020
rect 9036 15036 9088 15088
rect 10232 15079 10284 15088
rect 10232 15045 10266 15079
rect 10266 15045 10284 15079
rect 10232 15036 10284 15045
rect 12164 15036 12216 15088
rect 12808 15104 12860 15156
rect 12900 15104 12952 15156
rect 15200 15104 15252 15156
rect 15568 15147 15620 15156
rect 15568 15113 15577 15147
rect 15577 15113 15611 15147
rect 15611 15113 15620 15147
rect 15568 15104 15620 15113
rect 15016 15036 15068 15088
rect 15292 15036 15344 15088
rect 6736 15011 6788 15020
rect 6736 14977 6745 15011
rect 6745 14977 6779 15011
rect 6779 14977 6788 15011
rect 6736 14968 6788 14977
rect 7104 14968 7156 15020
rect 7196 14968 7248 15020
rect 8760 14968 8812 15020
rect 8944 14968 8996 15020
rect 12256 14968 12308 15020
rect 12624 14968 12676 15020
rect 13912 14968 13964 15020
rect 14372 14968 14424 15020
rect 14648 14968 14700 15020
rect 15108 15011 15160 15020
rect 15108 14977 15117 15011
rect 15117 14977 15151 15011
rect 15151 14977 15160 15011
rect 15108 14968 15160 14977
rect 4068 14900 4120 14952
rect 1584 14807 1636 14816
rect 1584 14773 1593 14807
rect 1593 14773 1627 14807
rect 1627 14773 1636 14807
rect 1584 14764 1636 14773
rect 4620 14832 4672 14884
rect 6368 14900 6420 14952
rect 6920 14900 6972 14952
rect 7012 14943 7064 14952
rect 7012 14909 7021 14943
rect 7021 14909 7055 14943
rect 7055 14909 7064 14943
rect 7656 14943 7708 14952
rect 7012 14900 7064 14909
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 7288 14832 7340 14884
rect 8208 14900 8260 14952
rect 8852 14943 8904 14952
rect 8852 14909 8861 14943
rect 8861 14909 8895 14943
rect 8895 14909 8904 14943
rect 8852 14900 8904 14909
rect 9772 14900 9824 14952
rect 4252 14764 4304 14816
rect 4436 14807 4488 14816
rect 4436 14773 4445 14807
rect 4445 14773 4479 14807
rect 4479 14773 4488 14807
rect 4436 14764 4488 14773
rect 4528 14807 4580 14816
rect 4528 14773 4537 14807
rect 4537 14773 4571 14807
rect 4571 14773 4580 14807
rect 4528 14764 4580 14773
rect 5172 14764 5224 14816
rect 8852 14764 8904 14816
rect 9312 14764 9364 14816
rect 9864 14764 9916 14816
rect 10968 14900 11020 14952
rect 12440 14943 12492 14952
rect 11520 14875 11572 14884
rect 11520 14841 11529 14875
rect 11529 14841 11563 14875
rect 11563 14841 11572 14875
rect 11520 14832 11572 14841
rect 12440 14909 12449 14943
rect 12449 14909 12483 14943
rect 12483 14909 12492 14943
rect 12440 14900 12492 14909
rect 13084 14900 13136 14952
rect 13728 14900 13780 14952
rect 14556 14900 14608 14952
rect 14740 14900 14792 14952
rect 10968 14764 11020 14816
rect 11888 14807 11940 14816
rect 11888 14773 11897 14807
rect 11897 14773 11931 14807
rect 11931 14773 11940 14807
rect 11888 14764 11940 14773
rect 12900 14832 12952 14884
rect 15108 14832 15160 14884
rect 14740 14764 14792 14816
rect 15844 14832 15896 14884
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 1492 14603 1544 14612
rect 1492 14569 1501 14603
rect 1501 14569 1535 14603
rect 1535 14569 1544 14603
rect 1492 14560 1544 14569
rect 2872 14535 2924 14544
rect 2872 14501 2881 14535
rect 2881 14501 2915 14535
rect 2915 14501 2924 14535
rect 2872 14492 2924 14501
rect 1584 14424 1636 14476
rect 3332 14424 3384 14476
rect 3700 14424 3752 14476
rect 4068 14424 4120 14476
rect 5632 14492 5684 14544
rect 6092 14492 6144 14544
rect 7656 14560 7708 14612
rect 10508 14492 10560 14544
rect 2964 14288 3016 14340
rect 4528 14288 4580 14340
rect 2320 14263 2372 14272
rect 2320 14229 2329 14263
rect 2329 14229 2363 14263
rect 2363 14229 2372 14263
rect 2320 14220 2372 14229
rect 2780 14263 2832 14272
rect 2780 14229 2789 14263
rect 2789 14229 2823 14263
rect 2823 14229 2832 14263
rect 2780 14220 2832 14229
rect 3608 14220 3660 14272
rect 3884 14263 3936 14272
rect 3884 14229 3893 14263
rect 3893 14229 3927 14263
rect 3927 14229 3936 14263
rect 3884 14220 3936 14229
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4712 14331 4764 14340
rect 4712 14297 4746 14331
rect 4746 14297 4764 14331
rect 4712 14288 4764 14297
rect 5356 14288 5408 14340
rect 9220 14424 9272 14476
rect 10324 14467 10376 14476
rect 10324 14433 10333 14467
rect 10333 14433 10367 14467
rect 10367 14433 10376 14467
rect 10324 14424 10376 14433
rect 5724 14356 5776 14408
rect 7748 14356 7800 14408
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 6460 14331 6512 14340
rect 5632 14220 5684 14272
rect 6460 14297 6494 14331
rect 6494 14297 6512 14331
rect 6460 14288 6512 14297
rect 6828 14288 6880 14340
rect 7012 14220 7064 14272
rect 8116 14220 8168 14272
rect 8760 14288 8812 14340
rect 8852 14220 8904 14272
rect 9128 14288 9180 14340
rect 11888 14560 11940 14612
rect 16948 14560 17000 14612
rect 13728 14492 13780 14544
rect 15108 14492 15160 14544
rect 12532 14424 12584 14476
rect 12716 14424 12768 14476
rect 12992 14424 13044 14476
rect 10968 14399 11020 14408
rect 10968 14365 10977 14399
rect 10977 14365 11011 14399
rect 11011 14365 11020 14399
rect 10968 14356 11020 14365
rect 11704 14356 11756 14408
rect 12716 14331 12768 14340
rect 9496 14220 9548 14272
rect 9680 14220 9732 14272
rect 10324 14220 10376 14272
rect 10692 14220 10744 14272
rect 10876 14263 10928 14272
rect 10876 14229 10885 14263
rect 10885 14229 10919 14263
rect 10919 14229 10928 14263
rect 10876 14220 10928 14229
rect 12716 14297 12725 14331
rect 12725 14297 12759 14331
rect 12759 14297 12768 14331
rect 12716 14288 12768 14297
rect 12900 14331 12952 14340
rect 12900 14297 12909 14331
rect 12909 14297 12943 14331
rect 12943 14297 12952 14331
rect 12900 14288 12952 14297
rect 11980 14220 12032 14272
rect 13176 14356 13228 14408
rect 13820 14356 13872 14408
rect 13728 14288 13780 14340
rect 15292 14288 15344 14340
rect 15384 14220 15436 14272
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 2872 14016 2924 14068
rect 2964 14059 3016 14068
rect 2964 14025 2973 14059
rect 2973 14025 3007 14059
rect 3007 14025 3016 14059
rect 2964 14016 3016 14025
rect 3608 14016 3660 14068
rect 4160 14059 4212 14068
rect 4160 14025 4169 14059
rect 4169 14025 4203 14059
rect 4203 14025 4212 14059
rect 4160 14016 4212 14025
rect 4252 14016 4304 14068
rect 5172 14016 5224 14068
rect 2780 13948 2832 14000
rect 3240 13948 3292 14000
rect 4528 13948 4580 14000
rect 5448 14016 5500 14068
rect 7380 14059 7432 14068
rect 7380 14025 7389 14059
rect 7389 14025 7423 14059
rect 7423 14025 7432 14059
rect 7380 14016 7432 14025
rect 7656 14016 7708 14068
rect 2596 13880 2648 13932
rect 4344 13880 4396 13932
rect 6920 13948 6972 14000
rect 10140 14016 10192 14068
rect 10324 14016 10376 14068
rect 11980 14059 12032 14068
rect 11980 14025 11989 14059
rect 11989 14025 12023 14059
rect 12023 14025 12032 14059
rect 11980 14016 12032 14025
rect 12808 14059 12860 14068
rect 9579 13948 9631 14000
rect 10968 13948 11020 14000
rect 11244 13948 11296 14000
rect 12808 14025 12817 14059
rect 12817 14025 12851 14059
rect 12851 14025 12860 14059
rect 12808 14016 12860 14025
rect 12900 14016 12952 14068
rect 13268 14016 13320 14068
rect 13360 14016 13412 14068
rect 13728 14016 13780 14068
rect 12624 13948 12676 14000
rect 1492 13787 1544 13796
rect 1492 13753 1501 13787
rect 1501 13753 1535 13787
rect 1535 13753 1544 13787
rect 1492 13744 1544 13753
rect 2688 13812 2740 13864
rect 3884 13812 3936 13864
rect 3976 13744 4028 13796
rect 4160 13812 4212 13864
rect 4620 13812 4672 13864
rect 5908 13880 5960 13932
rect 7564 13880 7616 13932
rect 7748 13923 7800 13932
rect 7748 13889 7757 13923
rect 7757 13889 7791 13923
rect 7791 13889 7800 13923
rect 7748 13880 7800 13889
rect 8024 13923 8076 13932
rect 8024 13889 8058 13923
rect 8058 13889 8076 13923
rect 8024 13880 8076 13889
rect 8300 13880 8352 13932
rect 8760 13880 8812 13932
rect 9312 13880 9364 13932
rect 10508 13880 10560 13932
rect 14004 13948 14056 14000
rect 6828 13812 6880 13864
rect 7012 13855 7064 13864
rect 7012 13821 7021 13855
rect 7021 13821 7055 13855
rect 7055 13821 7064 13855
rect 7012 13812 7064 13821
rect 5632 13744 5684 13796
rect 6184 13744 6236 13796
rect 9220 13744 9272 13796
rect 10508 13744 10560 13796
rect 11704 13744 11756 13796
rect 12164 13744 12216 13796
rect 4436 13676 4488 13728
rect 6368 13719 6420 13728
rect 6368 13685 6377 13719
rect 6377 13685 6411 13719
rect 6411 13685 6420 13719
rect 6368 13676 6420 13685
rect 8024 13676 8076 13728
rect 10140 13676 10192 13728
rect 11244 13676 11296 13728
rect 11888 13676 11940 13728
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 12992 13812 13044 13864
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13360 13855 13412 13864
rect 13360 13821 13369 13855
rect 13369 13821 13403 13855
rect 13403 13821 13412 13855
rect 13360 13812 13412 13821
rect 13912 13855 13964 13864
rect 13912 13821 13921 13855
rect 13921 13821 13955 13855
rect 13955 13821 13964 13855
rect 13912 13812 13964 13821
rect 15476 13855 15528 13864
rect 15476 13821 15485 13855
rect 15485 13821 15519 13855
rect 15519 13821 15528 13855
rect 15476 13812 15528 13821
rect 15752 13812 15804 13864
rect 15016 13676 15068 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 2320 13472 2372 13524
rect 5172 13515 5224 13524
rect 5172 13481 5181 13515
rect 5181 13481 5215 13515
rect 5215 13481 5224 13515
rect 5172 13472 5224 13481
rect 5724 13515 5776 13524
rect 5724 13481 5733 13515
rect 5733 13481 5767 13515
rect 5767 13481 5776 13515
rect 5724 13472 5776 13481
rect 7288 13472 7340 13524
rect 7472 13472 7524 13524
rect 8852 13472 8904 13524
rect 9588 13515 9640 13524
rect 9588 13481 9597 13515
rect 9597 13481 9631 13515
rect 9631 13481 9640 13515
rect 9588 13472 9640 13481
rect 10968 13472 11020 13524
rect 13820 13472 13872 13524
rect 13912 13472 13964 13524
rect 4160 13404 4212 13456
rect 5816 13404 5868 13456
rect 9956 13404 10008 13456
rect 10876 13404 10928 13456
rect 12072 13404 12124 13456
rect 12256 13447 12308 13456
rect 12256 13413 12265 13447
rect 12265 13413 12299 13447
rect 12299 13413 12308 13447
rect 12256 13404 12308 13413
rect 14280 13404 14332 13456
rect 15292 13404 15344 13456
rect 2872 13336 2924 13388
rect 3240 13336 3292 13388
rect 3884 13336 3936 13388
rect 1308 13200 1360 13252
rect 2228 13200 2280 13252
rect 3148 13268 3200 13320
rect 3516 13311 3568 13320
rect 3516 13277 3525 13311
rect 3525 13277 3559 13311
rect 3559 13277 3568 13311
rect 3516 13268 3568 13277
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 6368 13336 6420 13388
rect 8760 13379 8812 13388
rect 8760 13345 8769 13379
rect 8769 13345 8803 13379
rect 8803 13345 8812 13379
rect 8760 13336 8812 13345
rect 10140 13379 10192 13388
rect 10140 13345 10149 13379
rect 10149 13345 10183 13379
rect 10183 13345 10192 13379
rect 10140 13336 10192 13345
rect 14372 13336 14424 13388
rect 15568 13379 15620 13388
rect 15568 13345 15577 13379
rect 15577 13345 15611 13379
rect 15611 13345 15620 13379
rect 15568 13336 15620 13345
rect 6276 13268 6328 13320
rect 9128 13268 9180 13320
rect 3240 13200 3292 13252
rect 5356 13200 5408 13252
rect 7012 13243 7064 13252
rect 7012 13209 7021 13243
rect 7021 13209 7055 13243
rect 7055 13209 7064 13243
rect 7012 13200 7064 13209
rect 8668 13200 8720 13252
rect 9588 13200 9640 13252
rect 9680 13200 9732 13252
rect 10232 13200 10284 13252
rect 11336 13200 11388 13252
rect 12808 13268 12860 13320
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 1952 13175 2004 13184
rect 1952 13141 1961 13175
rect 1961 13141 1995 13175
rect 1995 13141 2004 13175
rect 1952 13132 2004 13141
rect 3424 13132 3476 13184
rect 6828 13132 6880 13184
rect 6920 13132 6972 13184
rect 8024 13132 8076 13184
rect 11520 13132 11572 13184
rect 12440 13200 12492 13252
rect 12624 13200 12676 13252
rect 13268 13200 13320 13252
rect 14096 13268 14148 13320
rect 13912 13200 13964 13252
rect 14188 13132 14240 13184
rect 14556 13175 14608 13184
rect 14556 13141 14565 13175
rect 14565 13141 14599 13175
rect 14599 13141 14608 13175
rect 15660 13200 15712 13252
rect 14556 13132 14608 13141
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 1952 12928 2004 12980
rect 3240 12971 3292 12980
rect 3240 12937 3249 12971
rect 3249 12937 3283 12971
rect 3283 12937 3292 12971
rect 3240 12928 3292 12937
rect 4620 12928 4672 12980
rect 5080 12928 5132 12980
rect 5356 12971 5408 12980
rect 5356 12937 5365 12971
rect 5365 12937 5399 12971
rect 5399 12937 5408 12971
rect 5356 12928 5408 12937
rect 6736 12971 6788 12980
rect 6736 12937 6745 12971
rect 6745 12937 6779 12971
rect 6779 12937 6788 12971
rect 6736 12928 6788 12937
rect 7472 12928 7524 12980
rect 8116 12928 8168 12980
rect 2136 12835 2188 12844
rect 2136 12801 2170 12835
rect 2170 12801 2188 12835
rect 5264 12903 5316 12912
rect 5264 12869 5273 12903
rect 5273 12869 5307 12903
rect 5307 12869 5316 12903
rect 5264 12860 5316 12869
rect 6184 12860 6236 12912
rect 9312 12928 9364 12980
rect 9864 12928 9916 12980
rect 10968 12971 11020 12980
rect 10968 12937 10977 12971
rect 10977 12937 11011 12971
rect 11011 12937 11020 12971
rect 10968 12928 11020 12937
rect 11244 12928 11296 12980
rect 11520 12971 11572 12980
rect 11520 12937 11529 12971
rect 11529 12937 11563 12971
rect 11563 12937 11572 12971
rect 11520 12928 11572 12937
rect 12072 12928 12124 12980
rect 14096 12928 14148 12980
rect 14740 12928 14792 12980
rect 14832 12928 14884 12980
rect 12992 12903 13044 12912
rect 2136 12792 2188 12801
rect 3148 12792 3200 12844
rect 4068 12792 4120 12844
rect 6460 12792 6512 12844
rect 8116 12835 8168 12844
rect 6828 12767 6880 12776
rect 2872 12656 2924 12708
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 8116 12801 8125 12835
rect 8125 12801 8159 12835
rect 8159 12801 8168 12835
rect 8116 12792 8168 12801
rect 7104 12724 7156 12776
rect 7840 12767 7892 12776
rect 7840 12733 7849 12767
rect 7849 12733 7883 12767
rect 7883 12733 7892 12767
rect 7840 12724 7892 12733
rect 12992 12869 13001 12903
rect 13001 12869 13035 12903
rect 13035 12869 13044 12903
rect 12992 12860 13044 12869
rect 9220 12792 9272 12844
rect 9772 12792 9824 12844
rect 9956 12792 10008 12844
rect 10508 12792 10560 12844
rect 11520 12792 11572 12844
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 1584 12631 1636 12640
rect 1584 12597 1593 12631
rect 1593 12597 1627 12631
rect 1627 12597 1636 12631
rect 1584 12588 1636 12597
rect 2228 12588 2280 12640
rect 9036 12656 9088 12708
rect 10784 12724 10836 12776
rect 11704 12724 11756 12776
rect 11980 12767 12032 12776
rect 11980 12733 11989 12767
rect 11989 12733 12023 12767
rect 12023 12733 12032 12767
rect 11980 12724 12032 12733
rect 12808 12767 12860 12776
rect 9772 12656 9824 12708
rect 10048 12656 10100 12708
rect 12808 12733 12817 12767
rect 12817 12733 12851 12767
rect 12851 12733 12860 12767
rect 12808 12724 12860 12733
rect 13268 12767 13320 12776
rect 13268 12733 13277 12767
rect 13277 12733 13311 12767
rect 13311 12733 13320 12767
rect 13268 12724 13320 12733
rect 13820 12724 13872 12776
rect 14280 12767 14332 12776
rect 14280 12733 14289 12767
rect 14289 12733 14323 12767
rect 14323 12733 14332 12767
rect 14280 12724 14332 12733
rect 15016 12792 15068 12844
rect 15108 12792 15160 12844
rect 15568 12792 15620 12844
rect 16304 12724 16356 12776
rect 12532 12656 12584 12708
rect 15292 12656 15344 12708
rect 6092 12588 6144 12640
rect 6460 12588 6512 12640
rect 9128 12588 9180 12640
rect 10140 12588 10192 12640
rect 10968 12588 11020 12640
rect 11152 12588 11204 12640
rect 13636 12588 13688 12640
rect 15016 12588 15068 12640
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 2136 12427 2188 12436
rect 2136 12393 2145 12427
rect 2145 12393 2179 12427
rect 2179 12393 2188 12427
rect 2136 12384 2188 12393
rect 3332 12384 3384 12436
rect 3424 12384 3476 12436
rect 5080 12384 5132 12436
rect 5264 12384 5316 12436
rect 2504 12316 2556 12368
rect 2596 12316 2648 12368
rect 1400 12180 1452 12232
rect 2320 12087 2372 12096
rect 2320 12053 2329 12087
rect 2329 12053 2363 12087
rect 2363 12053 2372 12087
rect 2320 12044 2372 12053
rect 3608 12316 3660 12368
rect 3240 12248 3292 12300
rect 5172 12248 5224 12300
rect 8300 12384 8352 12436
rect 10692 12427 10744 12436
rect 10692 12393 10701 12427
rect 10701 12393 10735 12427
rect 10735 12393 10744 12427
rect 10692 12384 10744 12393
rect 10968 12427 11020 12436
rect 10968 12393 10977 12427
rect 10977 12393 11011 12427
rect 11011 12393 11020 12427
rect 10968 12384 11020 12393
rect 12440 12384 12492 12436
rect 15660 12427 15712 12436
rect 15660 12393 15669 12427
rect 15669 12393 15703 12427
rect 15703 12393 15712 12427
rect 15660 12384 15712 12393
rect 10784 12316 10836 12368
rect 11060 12316 11112 12368
rect 12532 12248 12584 12300
rect 13452 12248 13504 12300
rect 13636 12248 13688 12300
rect 14096 12248 14148 12300
rect 16028 12248 16080 12300
rect 5540 12180 5592 12232
rect 5816 12223 5868 12232
rect 5816 12189 5825 12223
rect 5825 12189 5859 12223
rect 5859 12189 5868 12223
rect 5816 12180 5868 12189
rect 2872 12112 2924 12164
rect 3516 12112 3568 12164
rect 4068 12112 4120 12164
rect 4988 12112 5040 12164
rect 6092 12155 6144 12164
rect 6092 12121 6126 12155
rect 6126 12121 6144 12155
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 11244 12180 11296 12232
rect 12808 12180 12860 12232
rect 6092 12112 6144 12121
rect 4620 12044 4672 12096
rect 5080 12044 5132 12096
rect 5448 12044 5500 12096
rect 6368 12044 6420 12096
rect 6828 12044 6880 12096
rect 9312 12112 9364 12164
rect 10784 12112 10836 12164
rect 11428 12155 11480 12164
rect 11428 12121 11462 12155
rect 11462 12121 11480 12155
rect 11428 12112 11480 12121
rect 14740 12180 14792 12232
rect 15292 12223 15344 12232
rect 15292 12189 15301 12223
rect 15301 12189 15335 12223
rect 15335 12189 15344 12223
rect 15292 12180 15344 12189
rect 8852 12044 8904 12096
rect 13452 12112 13504 12164
rect 15108 12112 15160 12164
rect 12532 12087 12584 12096
rect 12532 12053 12541 12087
rect 12541 12053 12575 12087
rect 12575 12053 12584 12087
rect 12532 12044 12584 12053
rect 12624 12044 12676 12096
rect 13176 12044 13228 12096
rect 14096 12044 14148 12096
rect 15292 12044 15344 12096
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 3240 11840 3292 11892
rect 4068 11840 4120 11892
rect 5172 11883 5224 11892
rect 5172 11849 5181 11883
rect 5181 11849 5215 11883
rect 5215 11849 5224 11883
rect 5172 11840 5224 11849
rect 6000 11883 6052 11892
rect 6000 11849 6009 11883
rect 6009 11849 6043 11883
rect 6043 11849 6052 11883
rect 6000 11840 6052 11849
rect 6460 11840 6512 11892
rect 7748 11883 7800 11892
rect 3424 11772 3476 11824
rect 5908 11772 5960 11824
rect 7748 11849 7757 11883
rect 7757 11849 7791 11883
rect 7791 11849 7800 11883
rect 7748 11840 7800 11849
rect 9312 11883 9364 11892
rect 9312 11849 9321 11883
rect 9321 11849 9355 11883
rect 9355 11849 9364 11883
rect 9312 11840 9364 11849
rect 9680 11840 9732 11892
rect 10140 11840 10192 11892
rect 11888 11840 11940 11892
rect 3148 11704 3200 11756
rect 3608 11704 3660 11756
rect 4252 11747 4304 11756
rect 4252 11713 4261 11747
rect 4261 11713 4295 11747
rect 4295 11713 4304 11747
rect 4252 11704 4304 11713
rect 4988 11704 5040 11756
rect 5632 11704 5684 11756
rect 6000 11704 6052 11756
rect 6460 11704 6512 11756
rect 3332 11679 3384 11688
rect 3332 11645 3341 11679
rect 3341 11645 3375 11679
rect 3375 11645 3384 11679
rect 3332 11636 3384 11645
rect 3792 11636 3844 11688
rect 4896 11636 4948 11688
rect 3516 11568 3568 11620
rect 5448 11568 5500 11620
rect 6828 11636 6880 11688
rect 7840 11679 7892 11688
rect 7840 11645 7849 11679
rect 7849 11645 7883 11679
rect 7883 11645 7892 11679
rect 7840 11636 7892 11645
rect 7380 11568 7432 11620
rect 11336 11772 11388 11824
rect 13176 11840 13228 11892
rect 13360 11840 13412 11892
rect 14096 11840 14148 11892
rect 14464 11840 14516 11892
rect 14740 11883 14792 11892
rect 14740 11849 14749 11883
rect 14749 11849 14783 11883
rect 14783 11849 14792 11883
rect 14740 11840 14792 11849
rect 14832 11840 14884 11892
rect 15752 11840 15804 11892
rect 8300 11704 8352 11756
rect 10140 11704 10192 11756
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 12808 11772 12860 11824
rect 13452 11815 13504 11824
rect 11980 11704 12032 11713
rect 8300 11568 8352 11620
rect 11428 11636 11480 11688
rect 12348 11636 12400 11688
rect 13452 11781 13461 11815
rect 13461 11781 13495 11815
rect 13495 11781 13504 11815
rect 13452 11772 13504 11781
rect 15384 11815 15436 11824
rect 15384 11781 15393 11815
rect 15393 11781 15427 11815
rect 15427 11781 15436 11815
rect 15384 11772 15436 11781
rect 14648 11704 14700 11756
rect 15108 11747 15160 11756
rect 13728 11636 13780 11688
rect 14464 11679 14516 11688
rect 14464 11645 14473 11679
rect 14473 11645 14507 11679
rect 14507 11645 14516 11679
rect 14464 11636 14516 11645
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 15384 11636 15436 11688
rect 16120 11636 16172 11688
rect 12532 11568 12584 11620
rect 12992 11611 13044 11620
rect 12992 11577 13001 11611
rect 13001 11577 13035 11611
rect 13035 11577 13044 11611
rect 12992 11568 13044 11577
rect 1400 11543 1452 11552
rect 1400 11509 1409 11543
rect 1409 11509 1443 11543
rect 1443 11509 1452 11543
rect 1400 11500 1452 11509
rect 2412 11500 2464 11552
rect 3884 11543 3936 11552
rect 3884 11509 3893 11543
rect 3893 11509 3927 11543
rect 3927 11509 3936 11543
rect 3884 11500 3936 11509
rect 4344 11500 4396 11552
rect 4988 11500 5040 11552
rect 5264 11500 5316 11552
rect 8392 11500 8444 11552
rect 10968 11500 11020 11552
rect 11612 11500 11664 11552
rect 12348 11500 12400 11552
rect 12440 11543 12492 11552
rect 12440 11509 12449 11543
rect 12449 11509 12483 11543
rect 12483 11509 12492 11543
rect 12440 11500 12492 11509
rect 12808 11500 12860 11552
rect 13084 11500 13136 11552
rect 13360 11500 13412 11552
rect 16120 11500 16172 11552
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 3608 11339 3660 11348
rect 3608 11305 3617 11339
rect 3617 11305 3651 11339
rect 3651 11305 3660 11339
rect 3608 11296 3660 11305
rect 3792 11339 3844 11348
rect 3792 11305 3801 11339
rect 3801 11305 3835 11339
rect 3835 11305 3844 11339
rect 3792 11296 3844 11305
rect 4252 11296 4304 11348
rect 6460 11339 6512 11348
rect 6460 11305 6469 11339
rect 6469 11305 6503 11339
rect 6503 11305 6512 11339
rect 6460 11296 6512 11305
rect 8852 11296 8904 11348
rect 10140 11339 10192 11348
rect 2872 11228 2924 11280
rect 1400 11160 1452 11212
rect 2412 11160 2464 11212
rect 2780 11160 2832 11212
rect 3424 11160 3476 11212
rect 1676 11135 1728 11144
rect 1676 11101 1685 11135
rect 1685 11101 1719 11135
rect 1719 11101 1728 11135
rect 1676 11092 1728 11101
rect 2044 11024 2096 11076
rect 2872 11024 2924 11076
rect 3056 11092 3108 11144
rect 5724 11160 5776 11212
rect 10140 11305 10149 11339
rect 10149 11305 10183 11339
rect 10183 11305 10192 11339
rect 10140 11296 10192 11305
rect 7748 11160 7800 11212
rect 8116 11160 8168 11212
rect 8392 11203 8444 11212
rect 8392 11169 8401 11203
rect 8401 11169 8435 11203
rect 8435 11169 8444 11203
rect 8392 11160 8444 11169
rect 9036 11160 9088 11212
rect 3884 11024 3936 11076
rect 4436 11024 4488 11076
rect 4896 11067 4948 11076
rect 4896 11033 4914 11067
rect 4914 11033 4948 11067
rect 6920 11092 6972 11144
rect 7472 11092 7524 11144
rect 9772 11160 9824 11212
rect 11152 11228 11204 11280
rect 10784 11203 10836 11212
rect 10140 11092 10192 11144
rect 10784 11169 10793 11203
rect 10793 11169 10827 11203
rect 10827 11169 10836 11203
rect 10784 11160 10836 11169
rect 11244 11160 11296 11212
rect 10876 11092 10928 11144
rect 11428 11092 11480 11144
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 12900 11092 12952 11144
rect 13544 11296 13596 11348
rect 15384 11296 15436 11348
rect 15476 11296 15528 11348
rect 15936 11228 15988 11280
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 13636 11160 13688 11212
rect 13820 11160 13872 11212
rect 14556 11160 14608 11212
rect 15200 11092 15252 11144
rect 4896 11024 4948 11033
rect 1492 10999 1544 11008
rect 1492 10965 1501 10999
rect 1501 10965 1535 10999
rect 1535 10965 1544 10999
rect 1492 10956 1544 10965
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 5724 10999 5776 11008
rect 3240 10956 3292 10965
rect 5724 10965 5733 10999
rect 5733 10965 5767 10999
rect 5767 10965 5776 10999
rect 6460 11024 6512 11076
rect 7104 11067 7156 11076
rect 7104 11033 7113 11067
rect 7113 11033 7147 11067
rect 7147 11033 7156 11067
rect 7104 11024 7156 11033
rect 6736 10999 6788 11008
rect 5724 10956 5776 10965
rect 6736 10965 6745 10999
rect 6745 10965 6779 10999
rect 6779 10965 6788 10999
rect 6736 10956 6788 10965
rect 7932 10999 7984 11008
rect 7932 10965 7941 10999
rect 7941 10965 7975 10999
rect 7975 10965 7984 10999
rect 7932 10956 7984 10965
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 9588 10956 9640 11008
rect 15384 11024 15436 11076
rect 12900 10956 12952 11008
rect 13176 10999 13228 11008
rect 13176 10965 13185 10999
rect 13185 10965 13219 10999
rect 13219 10965 13228 10999
rect 13176 10956 13228 10965
rect 14556 10956 14608 11008
rect 15292 10956 15344 11008
rect 16488 10956 16540 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 1676 10752 1728 10804
rect 3148 10752 3200 10804
rect 6736 10752 6788 10804
rect 7748 10795 7800 10804
rect 7748 10761 7757 10795
rect 7757 10761 7791 10795
rect 7791 10761 7800 10795
rect 7748 10752 7800 10761
rect 11612 10752 11664 10804
rect 12624 10752 12676 10804
rect 14832 10752 14884 10804
rect 15016 10752 15068 10804
rect 4344 10727 4396 10736
rect 4344 10693 4353 10727
rect 4353 10693 4387 10727
rect 4387 10693 4396 10727
rect 4344 10684 4396 10693
rect 13268 10684 13320 10736
rect 5540 10659 5592 10668
rect 5540 10625 5558 10659
rect 5558 10625 5592 10659
rect 5540 10616 5592 10625
rect 5816 10659 5868 10668
rect 5816 10625 5825 10659
rect 5825 10625 5859 10659
rect 5859 10625 5868 10659
rect 5816 10616 5868 10625
rect 6920 10616 6972 10668
rect 7012 10616 7064 10668
rect 6000 10548 6052 10600
rect 2780 10480 2832 10532
rect 4436 10523 4488 10532
rect 4436 10489 4445 10523
rect 4445 10489 4479 10523
rect 4479 10489 4488 10523
rect 4436 10480 4488 10489
rect 10784 10616 10836 10668
rect 11244 10616 11296 10668
rect 12992 10616 13044 10668
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 13820 10616 13872 10668
rect 15016 10659 15068 10668
rect 15016 10625 15025 10659
rect 15025 10625 15059 10659
rect 15059 10625 15068 10659
rect 15016 10616 15068 10625
rect 14832 10548 14884 10600
rect 10232 10480 10284 10532
rect 14464 10480 14516 10532
rect 5448 10412 5500 10464
rect 9956 10455 10008 10464
rect 9956 10421 9965 10455
rect 9965 10421 9999 10455
rect 9999 10421 10008 10455
rect 9956 10412 10008 10421
rect 14740 10412 14792 10464
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 3332 10208 3384 10260
rect 3700 10208 3752 10260
rect 4068 10208 4120 10260
rect 5540 10208 5592 10260
rect 2688 10115 2740 10124
rect 2688 10081 2697 10115
rect 2697 10081 2731 10115
rect 2731 10081 2740 10115
rect 2688 10072 2740 10081
rect 1952 10047 2004 10056
rect 1492 9911 1544 9920
rect 1492 9877 1501 9911
rect 1501 9877 1535 9911
rect 1535 9877 1544 9911
rect 1492 9868 1544 9877
rect 1952 10013 1961 10047
rect 1961 10013 1995 10047
rect 1995 10013 2004 10047
rect 1952 10004 2004 10013
rect 2412 10047 2464 10056
rect 2412 10013 2421 10047
rect 2421 10013 2455 10047
rect 2455 10013 2464 10047
rect 2412 10004 2464 10013
rect 3700 10072 3752 10124
rect 4252 10072 4304 10124
rect 4160 10047 4212 10056
rect 4160 10013 4169 10047
rect 4169 10013 4203 10047
rect 4203 10013 4212 10047
rect 4160 10004 4212 10013
rect 4528 10072 4580 10124
rect 5264 10072 5316 10124
rect 1860 9868 1912 9920
rect 3332 9911 3384 9920
rect 3332 9877 3341 9911
rect 3341 9877 3375 9911
rect 3375 9877 3384 9911
rect 3332 9868 3384 9877
rect 4528 9936 4580 9988
rect 4436 9868 4488 9920
rect 5448 9936 5500 9988
rect 5172 9868 5224 9920
rect 5540 9868 5592 9920
rect 7472 10140 7524 10192
rect 9404 10208 9456 10260
rect 11244 10208 11296 10260
rect 12532 10208 12584 10260
rect 8944 10072 8996 10124
rect 9036 10072 9088 10124
rect 9956 10072 10008 10124
rect 10876 10072 10928 10124
rect 12072 10072 12124 10124
rect 12900 10072 12952 10124
rect 12992 10072 13044 10124
rect 14556 10115 14608 10124
rect 14556 10081 14565 10115
rect 14565 10081 14599 10115
rect 14599 10081 14608 10115
rect 14556 10072 14608 10081
rect 14740 10140 14792 10192
rect 15016 10072 15068 10124
rect 6460 10004 6512 10056
rect 11520 10004 11572 10056
rect 9128 9936 9180 9988
rect 9404 9936 9456 9988
rect 7196 9868 7248 9920
rect 8208 9868 8260 9920
rect 9956 9911 10008 9920
rect 9956 9877 9965 9911
rect 9965 9877 9999 9911
rect 9999 9877 10008 9911
rect 10232 9936 10284 9988
rect 13452 10004 13504 10056
rect 14464 10047 14516 10056
rect 14464 10013 14473 10047
rect 14473 10013 14507 10047
rect 14507 10013 14516 10047
rect 14464 10004 14516 10013
rect 15200 10004 15252 10056
rect 13268 9936 13320 9988
rect 9956 9868 10008 9877
rect 11060 9868 11112 9920
rect 13084 9911 13136 9920
rect 13084 9877 13093 9911
rect 13093 9877 13127 9911
rect 13127 9877 13136 9911
rect 13084 9868 13136 9877
rect 13452 9911 13504 9920
rect 13452 9877 13461 9911
rect 13461 9877 13495 9911
rect 13495 9877 13504 9911
rect 13452 9868 13504 9877
rect 13544 9911 13596 9920
rect 13544 9877 13553 9911
rect 13553 9877 13587 9911
rect 13587 9877 13596 9911
rect 14096 9911 14148 9920
rect 13544 9868 13596 9877
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 15568 9911 15620 9920
rect 15568 9877 15577 9911
rect 15577 9877 15611 9911
rect 15611 9877 15620 9911
rect 15568 9868 15620 9877
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 1400 9664 1452 9716
rect 4160 9664 4212 9716
rect 2504 9596 2556 9648
rect 5264 9664 5316 9716
rect 1768 9528 1820 9580
rect 2412 9528 2464 9580
rect 3148 9571 3200 9580
rect 3148 9537 3157 9571
rect 3157 9537 3191 9571
rect 3191 9537 3200 9571
rect 3148 9528 3200 9537
rect 4160 9528 4212 9580
rect 2504 9460 2556 9512
rect 3976 9460 4028 9512
rect 5448 9596 5500 9648
rect 4528 9528 4580 9580
rect 4988 9528 5040 9580
rect 5540 9528 5592 9580
rect 9404 9664 9456 9716
rect 9864 9707 9916 9716
rect 9864 9673 9873 9707
rect 9873 9673 9907 9707
rect 9907 9673 9916 9707
rect 9864 9664 9916 9673
rect 9956 9664 10008 9716
rect 11520 9707 11572 9716
rect 7932 9596 7984 9648
rect 9128 9596 9180 9648
rect 10048 9596 10100 9648
rect 10140 9596 10192 9648
rect 11520 9673 11529 9707
rect 11529 9673 11563 9707
rect 11563 9673 11572 9707
rect 11520 9664 11572 9673
rect 13084 9664 13136 9716
rect 13452 9664 13504 9716
rect 11060 9596 11112 9648
rect 11152 9596 11204 9648
rect 5356 9503 5408 9512
rect 5356 9469 5365 9503
rect 5365 9469 5399 9503
rect 5399 9469 5408 9503
rect 5356 9460 5408 9469
rect 5632 9503 5684 9512
rect 5632 9469 5641 9503
rect 5641 9469 5675 9503
rect 5675 9469 5684 9503
rect 5632 9460 5684 9469
rect 1676 9392 1728 9444
rect 4252 9392 4304 9444
rect 6828 9528 6880 9580
rect 7564 9571 7616 9580
rect 7564 9537 7573 9571
rect 7573 9537 7607 9571
rect 7607 9537 7616 9571
rect 7564 9528 7616 9537
rect 9404 9528 9456 9580
rect 7656 9503 7708 9512
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 1584 9324 1636 9376
rect 2136 9324 2188 9376
rect 2504 9324 2556 9376
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 4436 9324 4488 9376
rect 4620 9324 4672 9376
rect 6920 9392 6972 9444
rect 7104 9435 7156 9444
rect 7104 9401 7113 9435
rect 7113 9401 7147 9435
rect 7147 9401 7156 9435
rect 7104 9392 7156 9401
rect 7656 9469 7665 9503
rect 7665 9469 7699 9503
rect 7699 9469 7708 9503
rect 7656 9460 7708 9469
rect 7840 9503 7892 9512
rect 7840 9469 7849 9503
rect 7849 9469 7883 9503
rect 7883 9469 7892 9503
rect 7840 9460 7892 9469
rect 9036 9460 9088 9512
rect 8944 9392 8996 9444
rect 11244 9528 11296 9580
rect 11428 9596 11480 9648
rect 14096 9596 14148 9648
rect 11612 9528 11664 9580
rect 13452 9528 13504 9580
rect 14464 9596 14516 9648
rect 14832 9528 14884 9580
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 12072 9503 12124 9512
rect 12072 9469 12081 9503
rect 12081 9469 12115 9503
rect 12115 9469 12124 9503
rect 12072 9460 12124 9469
rect 12624 9460 12676 9512
rect 13820 9503 13872 9512
rect 10784 9392 10836 9444
rect 12348 9435 12400 9444
rect 12348 9401 12357 9435
rect 12357 9401 12391 9435
rect 12391 9401 12400 9435
rect 12348 9392 12400 9401
rect 12532 9392 12584 9444
rect 13820 9469 13829 9503
rect 13829 9469 13863 9503
rect 13863 9469 13872 9503
rect 13820 9460 13872 9469
rect 14280 9460 14332 9512
rect 14556 9503 14608 9512
rect 14556 9469 14565 9503
rect 14565 9469 14599 9503
rect 14599 9469 14608 9503
rect 14556 9460 14608 9469
rect 13728 9392 13780 9444
rect 9036 9367 9088 9376
rect 9036 9333 9045 9367
rect 9045 9333 9079 9367
rect 9079 9333 9088 9367
rect 9036 9324 9088 9333
rect 9128 9324 9180 9376
rect 9680 9324 9732 9376
rect 11244 9367 11296 9376
rect 11244 9333 11253 9367
rect 11253 9333 11287 9367
rect 11287 9333 11296 9367
rect 11244 9324 11296 9333
rect 12992 9324 13044 9376
rect 14464 9324 14516 9376
rect 14924 9367 14976 9376
rect 14924 9333 14933 9367
rect 14933 9333 14967 9367
rect 14967 9333 14976 9367
rect 14924 9324 14976 9333
rect 15844 9324 15896 9376
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 3792 9163 3844 9172
rect 1676 8959 1728 8968
rect 1676 8925 1685 8959
rect 1685 8925 1719 8959
rect 1719 8925 1728 8959
rect 1676 8916 1728 8925
rect 3792 9129 3801 9163
rect 3801 9129 3835 9163
rect 3835 9129 3844 9163
rect 3792 9120 3844 9129
rect 3976 9163 4028 9172
rect 3976 9129 3985 9163
rect 3985 9129 4019 9163
rect 4019 9129 4028 9163
rect 3976 9120 4028 9129
rect 4160 9163 4212 9172
rect 4160 9129 4169 9163
rect 4169 9129 4203 9163
rect 4203 9129 4212 9163
rect 4160 9120 4212 9129
rect 3884 9052 3936 9104
rect 5908 9120 5960 9172
rect 7564 9120 7616 9172
rect 9680 9120 9732 9172
rect 8760 9052 8812 9104
rect 4620 9027 4672 9036
rect 4620 8993 4629 9027
rect 4629 8993 4663 9027
rect 4663 8993 4672 9027
rect 4620 8984 4672 8993
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 6460 9027 6512 9036
rect 4712 8984 4764 8993
rect 6460 8993 6469 9027
rect 6469 8993 6503 9027
rect 6503 8993 6512 9027
rect 6460 8984 6512 8993
rect 7564 8984 7616 9036
rect 8208 9027 8260 9036
rect 8208 8993 8217 9027
rect 8217 8993 8251 9027
rect 8251 8993 8260 9027
rect 8208 8984 8260 8993
rect 8852 8984 8904 9036
rect 14648 9052 14700 9104
rect 14924 9052 14976 9104
rect 10784 8984 10836 9036
rect 12072 8984 12124 9036
rect 15016 8984 15068 9036
rect 3240 8916 3292 8968
rect 5540 8916 5592 8968
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 10140 8959 10192 8968
rect 10140 8925 10149 8959
rect 10149 8925 10183 8959
rect 10183 8925 10192 8959
rect 10140 8916 10192 8925
rect 10968 8916 11020 8968
rect 1676 8780 1728 8832
rect 2320 8848 2372 8900
rect 3516 8848 3568 8900
rect 4436 8848 4488 8900
rect 5356 8848 5408 8900
rect 7196 8848 7248 8900
rect 4160 8780 4212 8832
rect 4528 8823 4580 8832
rect 4528 8789 4537 8823
rect 4537 8789 4571 8823
rect 4571 8789 4580 8823
rect 4528 8780 4580 8789
rect 6092 8780 6144 8832
rect 7288 8780 7340 8832
rect 7748 8848 7800 8900
rect 10600 8848 10652 8900
rect 13360 8916 13412 8968
rect 13728 8916 13780 8968
rect 14648 8916 14700 8968
rect 16028 8916 16080 8968
rect 9036 8780 9088 8832
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 9772 8823 9824 8832
rect 9404 8780 9456 8789
rect 9772 8789 9781 8823
rect 9781 8789 9815 8823
rect 9815 8789 9824 8823
rect 9772 8780 9824 8789
rect 11980 8780 12032 8832
rect 12900 8848 12952 8900
rect 14556 8848 14608 8900
rect 15936 8848 15988 8900
rect 13820 8780 13872 8832
rect 14372 8823 14424 8832
rect 14372 8789 14381 8823
rect 14381 8789 14415 8823
rect 14415 8789 14424 8823
rect 14372 8780 14424 8789
rect 14464 8780 14516 8832
rect 14740 8780 14792 8832
rect 15752 8780 15804 8832
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 1768 8619 1820 8628
rect 1768 8585 1777 8619
rect 1777 8585 1811 8619
rect 1811 8585 1820 8619
rect 1768 8576 1820 8585
rect 3148 8576 3200 8628
rect 4160 8576 4212 8628
rect 1860 8440 1912 8492
rect 4252 8508 4304 8560
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 3148 8440 3200 8492
rect 3884 8440 3936 8492
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 3608 8372 3660 8424
rect 5356 8576 5408 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 9036 8576 9088 8628
rect 9864 8619 9916 8628
rect 5540 8508 5592 8560
rect 6092 8508 6144 8560
rect 2228 8304 2280 8356
rect 3424 8304 3476 8356
rect 1768 8236 1820 8288
rect 3332 8236 3384 8288
rect 3700 8236 3752 8288
rect 4252 8236 4304 8288
rect 5172 8236 5224 8288
rect 6276 8440 6328 8492
rect 8024 8508 8076 8560
rect 9220 8508 9272 8560
rect 9864 8585 9873 8619
rect 9873 8585 9907 8619
rect 9907 8585 9916 8619
rect 9864 8576 9916 8585
rect 9772 8508 9824 8560
rect 8392 8440 8444 8492
rect 9128 8440 9180 8492
rect 10600 8576 10652 8628
rect 12532 8619 12584 8628
rect 10140 8508 10192 8560
rect 10876 8508 10928 8560
rect 10968 8508 11020 8560
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 12992 8576 13044 8628
rect 13544 8576 13596 8628
rect 14372 8576 14424 8628
rect 15292 8576 15344 8628
rect 16396 8576 16448 8628
rect 12716 8508 12768 8560
rect 6368 8304 6420 8356
rect 7104 8372 7156 8424
rect 7288 8415 7340 8424
rect 7288 8381 7297 8415
rect 7297 8381 7331 8415
rect 7331 8381 7340 8415
rect 7288 8372 7340 8381
rect 7472 8372 7524 8424
rect 7656 8304 7708 8356
rect 7748 8347 7800 8356
rect 7748 8313 7757 8347
rect 7757 8313 7791 8347
rect 7791 8313 7800 8347
rect 8208 8372 8260 8424
rect 8668 8415 8720 8424
rect 8668 8381 8677 8415
rect 8677 8381 8711 8415
rect 8711 8381 8720 8415
rect 8668 8372 8720 8381
rect 7748 8304 7800 8313
rect 9220 8304 9272 8356
rect 11520 8372 11572 8424
rect 11796 8372 11848 8424
rect 11980 8415 12032 8424
rect 11980 8381 11989 8415
rect 11989 8381 12023 8415
rect 12023 8381 12032 8415
rect 11980 8372 12032 8381
rect 13820 8508 13872 8560
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13452 8483 13504 8492
rect 13452 8449 13461 8483
rect 13461 8449 13495 8483
rect 13495 8449 13504 8483
rect 13452 8440 13504 8449
rect 11336 8304 11388 8356
rect 6000 8236 6052 8288
rect 7380 8236 7432 8288
rect 11704 8236 11756 8288
rect 12716 8236 12768 8288
rect 15660 8236 15712 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 3700 8032 3752 8084
rect 4528 8032 4580 8084
rect 5724 8032 5776 8084
rect 8392 8032 8444 8084
rect 8852 8032 8904 8084
rect 9404 8032 9456 8084
rect 9588 8032 9640 8084
rect 9864 8032 9916 8084
rect 11704 8032 11756 8084
rect 11888 8032 11940 8084
rect 12992 8032 13044 8084
rect 14924 8032 14976 8084
rect 3056 7964 3108 8016
rect 3516 7964 3568 8016
rect 4160 7964 4212 8016
rect 2596 7896 2648 7948
rect 6460 7964 6512 8016
rect 5264 7896 5316 7948
rect 6368 7896 6420 7948
rect 7932 7964 7984 8016
rect 9036 7964 9088 8016
rect 8484 7939 8536 7948
rect 1768 7828 1820 7880
rect 2044 7828 2096 7880
rect 3516 7828 3568 7880
rect 4160 7828 4212 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 6184 7828 6236 7880
rect 8484 7905 8493 7939
rect 8493 7905 8527 7939
rect 8527 7905 8536 7939
rect 8484 7896 8536 7905
rect 9404 7939 9456 7948
rect 9404 7905 9413 7939
rect 9413 7905 9447 7939
rect 9447 7905 9456 7939
rect 9404 7896 9456 7905
rect 7196 7871 7248 7880
rect 7196 7837 7219 7871
rect 7219 7837 7248 7871
rect 7196 7828 7248 7837
rect 8668 7828 8720 7880
rect 9220 7828 9272 7880
rect 2596 7760 2648 7812
rect 4252 7760 4304 7812
rect 5172 7760 5224 7812
rect 7932 7760 7984 7812
rect 9588 7760 9640 7812
rect 1860 7692 1912 7744
rect 2044 7735 2096 7744
rect 2044 7701 2053 7735
rect 2053 7701 2087 7735
rect 2087 7701 2096 7735
rect 2044 7692 2096 7701
rect 2780 7735 2832 7744
rect 2780 7701 2789 7735
rect 2789 7701 2823 7735
rect 2823 7701 2832 7735
rect 2780 7692 2832 7701
rect 3332 7692 3384 7744
rect 3700 7692 3752 7744
rect 5264 7692 5316 7744
rect 6368 7692 6420 7744
rect 7472 7692 7524 7744
rect 9128 7692 9180 7744
rect 9404 7692 9456 7744
rect 12624 7964 12676 8016
rect 10876 7939 10928 7948
rect 10876 7905 10885 7939
rect 10885 7905 10919 7939
rect 10919 7905 10928 7939
rect 10876 7896 10928 7905
rect 11520 7896 11572 7948
rect 10784 7828 10836 7880
rect 11060 7828 11112 7880
rect 12716 7828 12768 7880
rect 10324 7735 10376 7744
rect 10324 7701 10333 7735
rect 10333 7701 10367 7735
rect 10367 7701 10376 7735
rect 10324 7692 10376 7701
rect 10416 7692 10468 7744
rect 12808 7760 12860 7812
rect 11888 7735 11940 7744
rect 11888 7701 11897 7735
rect 11897 7701 11931 7735
rect 11931 7701 11940 7735
rect 11888 7692 11940 7701
rect 12624 7692 12676 7744
rect 12992 7692 13044 7744
rect 13176 7760 13228 7812
rect 13728 7760 13780 7812
rect 14280 7964 14332 8016
rect 14556 7896 14608 7948
rect 14372 7828 14424 7880
rect 15292 7760 15344 7812
rect 16212 7760 16264 7812
rect 13360 7735 13412 7744
rect 13360 7701 13369 7735
rect 13369 7701 13403 7735
rect 13403 7701 13412 7735
rect 13360 7692 13412 7701
rect 13636 7735 13688 7744
rect 13636 7701 13645 7735
rect 13645 7701 13679 7735
rect 13679 7701 13688 7735
rect 13636 7692 13688 7701
rect 14924 7735 14976 7744
rect 14924 7701 14933 7735
rect 14933 7701 14967 7735
rect 14967 7701 14976 7735
rect 14924 7692 14976 7701
rect 15568 7735 15620 7744
rect 15568 7701 15577 7735
rect 15577 7701 15611 7735
rect 15611 7701 15620 7735
rect 15568 7692 15620 7701
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 3240 7488 3292 7540
rect 3608 7488 3660 7540
rect 5356 7488 5408 7540
rect 5448 7488 5500 7540
rect 7380 7488 7432 7540
rect 7840 7531 7892 7540
rect 7840 7497 7849 7531
rect 7849 7497 7883 7531
rect 7883 7497 7892 7531
rect 10416 7531 10468 7540
rect 7840 7488 7892 7497
rect 2320 7420 2372 7472
rect 3976 7420 4028 7472
rect 4344 7463 4396 7472
rect 4344 7429 4353 7463
rect 4353 7429 4387 7463
rect 4387 7429 4396 7463
rect 4344 7420 4396 7429
rect 5080 7420 5132 7472
rect 5540 7420 5592 7472
rect 8852 7420 8904 7472
rect 10416 7497 10425 7531
rect 10425 7497 10459 7531
rect 10459 7497 10468 7531
rect 10416 7488 10468 7497
rect 13912 7488 13964 7540
rect 14556 7488 14608 7540
rect 16304 7488 16356 7540
rect 11060 7420 11112 7472
rect 11152 7420 11204 7472
rect 11612 7420 11664 7472
rect 12348 7420 12400 7472
rect 12532 7420 12584 7472
rect 14372 7420 14424 7472
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 2228 7352 2280 7404
rect 2412 7352 2464 7404
rect 2688 7352 2740 7404
rect 3332 7352 3384 7404
rect 4804 7352 4856 7404
rect 5632 7352 5684 7404
rect 3056 7284 3108 7336
rect 3700 7284 3752 7336
rect 4620 7284 4672 7336
rect 5080 7327 5132 7336
rect 5080 7293 5089 7327
rect 5089 7293 5123 7327
rect 5123 7293 5132 7327
rect 5080 7284 5132 7293
rect 1492 7191 1544 7200
rect 1492 7157 1501 7191
rect 1501 7157 1535 7191
rect 1535 7157 1544 7191
rect 1492 7148 1544 7157
rect 2228 7148 2280 7200
rect 2596 7148 2648 7200
rect 4620 7191 4672 7200
rect 4620 7157 4629 7191
rect 4629 7157 4663 7191
rect 4663 7157 4672 7191
rect 4620 7148 4672 7157
rect 5172 7216 5224 7268
rect 6000 7352 6052 7404
rect 6460 7352 6512 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 6920 7327 6972 7336
rect 6920 7293 6929 7327
rect 6929 7293 6963 7327
rect 6963 7293 6972 7327
rect 6920 7284 6972 7293
rect 5448 7191 5500 7200
rect 5448 7157 5457 7191
rect 5457 7157 5491 7191
rect 5491 7157 5500 7191
rect 5448 7148 5500 7157
rect 6000 7216 6052 7268
rect 9864 7352 9916 7404
rect 12256 7352 12308 7404
rect 12900 7395 12952 7404
rect 12900 7361 12909 7395
rect 12909 7361 12943 7395
rect 12943 7361 12952 7395
rect 12900 7352 12952 7361
rect 15660 7352 15712 7404
rect 6920 7148 6972 7200
rect 7656 7148 7708 7200
rect 9404 7191 9456 7200
rect 9404 7157 9413 7191
rect 9413 7157 9447 7191
rect 9447 7157 9456 7191
rect 9404 7148 9456 7157
rect 9956 7327 10008 7336
rect 9956 7293 9965 7327
rect 9965 7293 9999 7327
rect 9999 7293 10008 7327
rect 9956 7284 10008 7293
rect 11152 7284 11204 7336
rect 13912 7284 13964 7336
rect 14832 7284 14884 7336
rect 15200 7284 15252 7336
rect 11520 7259 11572 7268
rect 11520 7225 11529 7259
rect 11529 7225 11563 7259
rect 11563 7225 11572 7259
rect 11520 7216 11572 7225
rect 14280 7216 14332 7268
rect 14556 7216 14608 7268
rect 9772 7148 9824 7200
rect 10140 7148 10192 7200
rect 10876 7148 10928 7200
rect 12624 7148 12676 7200
rect 16120 7148 16172 7200
rect 16580 7148 16632 7200
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 5172 6944 5224 6996
rect 5816 6944 5868 6996
rect 6460 6944 6512 6996
rect 9956 6944 10008 6996
rect 11520 6944 11572 6996
rect 12164 6944 12216 6996
rect 12532 6944 12584 6996
rect 12624 6944 12676 6996
rect 1400 6876 1452 6928
rect 1952 6876 2004 6928
rect 1676 6808 1728 6860
rect 3240 6740 3292 6792
rect 3332 6740 3384 6792
rect 1952 6672 2004 6724
rect 2780 6672 2832 6724
rect 1768 6647 1820 6656
rect 1768 6613 1777 6647
rect 1777 6613 1811 6647
rect 1811 6613 1820 6647
rect 1768 6604 1820 6613
rect 3056 6604 3108 6656
rect 3608 6740 3660 6792
rect 3884 6783 3936 6792
rect 3884 6749 3893 6783
rect 3893 6749 3927 6783
rect 3927 6749 3936 6783
rect 3884 6740 3936 6749
rect 4160 6876 4212 6928
rect 4252 6808 4304 6860
rect 4620 6808 4672 6860
rect 12808 6944 12860 6996
rect 15292 6944 15344 6996
rect 5448 6808 5500 6860
rect 5816 6808 5868 6860
rect 6000 6808 6052 6860
rect 7472 6851 7524 6860
rect 7472 6817 7481 6851
rect 7481 6817 7515 6851
rect 7515 6817 7524 6851
rect 7472 6808 7524 6817
rect 5908 6740 5960 6792
rect 7288 6740 7340 6792
rect 4436 6672 4488 6724
rect 5540 6604 5592 6656
rect 5632 6647 5684 6656
rect 5632 6613 5641 6647
rect 5641 6613 5675 6647
rect 5675 6613 5684 6647
rect 8852 6808 8904 6860
rect 12348 6808 12400 6860
rect 13728 6876 13780 6928
rect 15384 6919 15436 6928
rect 9680 6740 9732 6792
rect 9864 6740 9916 6792
rect 13360 6740 13412 6792
rect 14280 6740 14332 6792
rect 15384 6885 15393 6919
rect 15393 6885 15427 6919
rect 15427 6885 15436 6919
rect 15384 6876 15436 6885
rect 5632 6604 5684 6613
rect 7012 6647 7064 6656
rect 7012 6613 7021 6647
rect 7021 6613 7055 6647
rect 7055 6613 7064 6647
rect 7012 6604 7064 6613
rect 8300 6672 8352 6724
rect 7932 6647 7984 6656
rect 7932 6613 7941 6647
rect 7941 6613 7975 6647
rect 7975 6613 7984 6647
rect 7932 6604 7984 6613
rect 9588 6604 9640 6656
rect 11612 6647 11664 6656
rect 11612 6613 11621 6647
rect 11621 6613 11655 6647
rect 11655 6613 11664 6647
rect 11612 6604 11664 6613
rect 12256 6672 12308 6724
rect 13636 6672 13688 6724
rect 15476 6740 15528 6792
rect 14556 6672 14608 6724
rect 15200 6715 15252 6724
rect 15200 6681 15209 6715
rect 15209 6681 15243 6715
rect 15243 6681 15252 6715
rect 15200 6672 15252 6681
rect 15568 6715 15620 6724
rect 15568 6681 15577 6715
rect 15577 6681 15611 6715
rect 15611 6681 15620 6715
rect 15568 6672 15620 6681
rect 16120 6672 16172 6724
rect 12716 6604 12768 6656
rect 13176 6604 13228 6656
rect 13360 6647 13412 6656
rect 13360 6613 13369 6647
rect 13369 6613 13403 6647
rect 13403 6613 13412 6647
rect 13360 6604 13412 6613
rect 15384 6604 15436 6656
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 1676 6400 1728 6452
rect 1492 6264 1544 6316
rect 3424 6332 3476 6384
rect 2412 6264 2464 6316
rect 2688 6264 2740 6316
rect 3424 6239 3476 6248
rect 3424 6205 3433 6239
rect 3433 6205 3467 6239
rect 3467 6205 3476 6239
rect 3424 6196 3476 6205
rect 5080 6400 5132 6452
rect 7932 6400 7984 6452
rect 8852 6400 8904 6452
rect 9588 6400 9640 6452
rect 10048 6400 10100 6452
rect 10876 6400 10928 6452
rect 11060 6400 11112 6452
rect 11612 6400 11664 6452
rect 11888 6443 11940 6452
rect 11888 6409 11897 6443
rect 11897 6409 11931 6443
rect 11931 6409 11940 6443
rect 11888 6400 11940 6409
rect 3792 6264 3844 6316
rect 4528 6196 4580 6248
rect 5356 6264 5408 6316
rect 7748 6332 7800 6384
rect 8300 6332 8352 6384
rect 12716 6400 12768 6452
rect 13176 6400 13228 6452
rect 14280 6443 14332 6452
rect 14280 6409 14289 6443
rect 14289 6409 14323 6443
rect 14323 6409 14332 6443
rect 14280 6400 14332 6409
rect 12440 6332 12492 6384
rect 12624 6332 12676 6384
rect 12900 6332 12952 6384
rect 12992 6332 13044 6384
rect 13728 6332 13780 6384
rect 14556 6400 14608 6452
rect 15292 6400 15344 6452
rect 1492 6171 1544 6180
rect 1492 6137 1501 6171
rect 1501 6137 1535 6171
rect 1535 6137 1544 6171
rect 1492 6128 1544 6137
rect 3976 6128 4028 6180
rect 4988 6128 5040 6180
rect 6000 6196 6052 6248
rect 6184 6196 6236 6248
rect 7380 6196 7432 6248
rect 9956 6307 10008 6316
rect 9956 6273 9965 6307
rect 9965 6273 9999 6307
rect 9999 6273 10008 6307
rect 9956 6264 10008 6273
rect 10968 6264 11020 6316
rect 12348 6307 12400 6316
rect 2228 6060 2280 6112
rect 3608 6060 3660 6112
rect 3792 6103 3844 6112
rect 3792 6069 3801 6103
rect 3801 6069 3835 6103
rect 3835 6069 3844 6103
rect 3792 6060 3844 6069
rect 6184 6060 6236 6112
rect 10048 6196 10100 6248
rect 10784 6196 10836 6248
rect 12348 6273 12357 6307
rect 12357 6273 12391 6307
rect 12391 6273 12400 6307
rect 12348 6264 12400 6273
rect 12532 6239 12584 6248
rect 12532 6205 12541 6239
rect 12541 6205 12575 6239
rect 12575 6205 12584 6239
rect 12532 6196 12584 6205
rect 12900 6239 12952 6248
rect 12900 6205 12909 6239
rect 12909 6205 12943 6239
rect 12943 6205 12952 6239
rect 12900 6196 12952 6205
rect 12624 6128 12676 6180
rect 13820 6239 13872 6248
rect 13820 6205 13829 6239
rect 13829 6205 13863 6239
rect 13863 6205 13872 6239
rect 13820 6196 13872 6205
rect 15476 6332 15528 6384
rect 14832 6307 14884 6316
rect 14832 6273 14841 6307
rect 14841 6273 14875 6307
rect 14875 6273 14884 6307
rect 14832 6264 14884 6273
rect 15384 6307 15436 6316
rect 15384 6273 15393 6307
rect 15393 6273 15427 6307
rect 15427 6273 15436 6307
rect 15384 6264 15436 6273
rect 14924 6239 14976 6248
rect 14924 6205 14933 6239
rect 14933 6205 14967 6239
rect 14967 6205 14976 6239
rect 14924 6196 14976 6205
rect 9772 6060 9824 6112
rect 10048 6103 10100 6112
rect 10048 6069 10057 6103
rect 10057 6069 10091 6103
rect 10091 6069 10100 6103
rect 10048 6060 10100 6069
rect 13820 6060 13872 6112
rect 14464 6060 14516 6112
rect 15568 6103 15620 6112
rect 15568 6069 15577 6103
rect 15577 6069 15611 6103
rect 15611 6069 15620 6103
rect 15568 6060 15620 6069
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 4160 5856 4212 5908
rect 3148 5788 3200 5840
rect 5908 5856 5960 5908
rect 6000 5788 6052 5840
rect 3516 5763 3568 5772
rect 3516 5729 3525 5763
rect 3525 5729 3559 5763
rect 3559 5729 3568 5763
rect 3516 5720 3568 5729
rect 6184 5720 6236 5772
rect 6460 5788 6512 5840
rect 7472 5788 7524 5840
rect 8944 5899 8996 5908
rect 8944 5865 8953 5899
rect 8953 5865 8987 5899
rect 8987 5865 8996 5899
rect 9220 5899 9272 5908
rect 8944 5856 8996 5865
rect 9220 5865 9229 5899
rect 9229 5865 9263 5899
rect 9263 5865 9272 5899
rect 9220 5856 9272 5865
rect 9312 5856 9364 5908
rect 9588 5856 9640 5908
rect 10140 5856 10192 5908
rect 10968 5856 11020 5908
rect 11336 5856 11388 5908
rect 3056 5652 3108 5704
rect 3792 5652 3844 5704
rect 5632 5652 5684 5704
rect 7012 5652 7064 5704
rect 7380 5695 7432 5704
rect 7380 5661 7389 5695
rect 7389 5661 7423 5695
rect 7423 5661 7432 5695
rect 7380 5652 7432 5661
rect 8300 5720 8352 5772
rect 8668 5763 8720 5772
rect 8668 5729 8677 5763
rect 8677 5729 8711 5763
rect 8711 5729 8720 5763
rect 8668 5720 8720 5729
rect 9864 5788 9916 5840
rect 10140 5763 10192 5772
rect 7564 5652 7616 5704
rect 8208 5652 8260 5704
rect 10140 5729 10149 5763
rect 10149 5729 10183 5763
rect 10183 5729 10192 5763
rect 10140 5720 10192 5729
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 1676 5627 1728 5636
rect 1676 5593 1710 5627
rect 1710 5593 1728 5627
rect 1676 5584 1728 5593
rect 3332 5627 3384 5636
rect 3332 5593 3341 5627
rect 3341 5593 3375 5627
rect 3375 5593 3384 5627
rect 3332 5584 3384 5593
rect 5080 5627 5132 5636
rect 5080 5593 5098 5627
rect 5098 5593 5132 5627
rect 5080 5584 5132 5593
rect 6276 5584 6328 5636
rect 2688 5516 2740 5568
rect 3976 5559 4028 5568
rect 3976 5525 3985 5559
rect 3985 5525 4019 5559
rect 4019 5525 4028 5559
rect 3976 5516 4028 5525
rect 6000 5516 6052 5568
rect 10048 5652 10100 5704
rect 11704 5652 11756 5704
rect 12624 5695 12676 5704
rect 12624 5661 12633 5695
rect 12633 5661 12667 5695
rect 12667 5661 12676 5695
rect 12624 5652 12676 5661
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 8116 5516 8168 5568
rect 10232 5584 10284 5636
rect 9312 5516 9364 5568
rect 9956 5559 10008 5568
rect 9956 5525 9965 5559
rect 9965 5525 9999 5559
rect 9999 5525 10008 5559
rect 9956 5516 10008 5525
rect 12716 5559 12768 5568
rect 12716 5525 12725 5559
rect 12725 5525 12759 5559
rect 12759 5525 12768 5559
rect 12716 5516 12768 5525
rect 12992 5516 13044 5568
rect 13544 5856 13596 5908
rect 14924 5856 14976 5908
rect 15384 5788 15436 5840
rect 13544 5720 13596 5772
rect 15568 5720 15620 5772
rect 15292 5652 15344 5704
rect 16488 5652 16540 5704
rect 13912 5584 13964 5636
rect 14280 5516 14332 5568
rect 14832 5516 14884 5568
rect 15292 5559 15344 5568
rect 15292 5525 15301 5559
rect 15301 5525 15335 5559
rect 15335 5525 15344 5559
rect 15292 5516 15344 5525
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 1492 5355 1544 5364
rect 1492 5321 1501 5355
rect 1501 5321 1535 5355
rect 1535 5321 1544 5355
rect 1492 5312 1544 5321
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 2136 5312 2188 5364
rect 2228 5312 2280 5364
rect 2872 5312 2924 5364
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 3424 5312 3476 5364
rect 5816 5312 5868 5364
rect 7840 5312 7892 5364
rect 8024 5312 8076 5364
rect 8300 5312 8352 5364
rect 10140 5312 10192 5364
rect 10968 5312 11020 5364
rect 2504 5244 2556 5296
rect 3148 5244 3200 5296
rect 3792 5244 3844 5296
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 2780 5176 2832 5228
rect 3884 5176 3936 5228
rect 3976 5176 4028 5228
rect 4160 5176 4212 5228
rect 4344 5219 4396 5228
rect 4344 5185 4353 5219
rect 4353 5185 4387 5219
rect 4387 5185 4396 5219
rect 4344 5176 4396 5185
rect 4436 5219 4488 5228
rect 4436 5185 4445 5219
rect 4445 5185 4479 5219
rect 4479 5185 4488 5219
rect 5632 5244 5684 5296
rect 4436 5176 4488 5185
rect 6184 5176 6236 5228
rect 6368 5176 6420 5228
rect 2228 5151 2280 5160
rect 2228 5117 2237 5151
rect 2237 5117 2271 5151
rect 2271 5117 2280 5151
rect 2228 5108 2280 5117
rect 2504 5108 2556 5160
rect 2688 5108 2740 5160
rect 2872 5108 2924 5160
rect 4528 5108 4580 5160
rect 7196 5151 7248 5160
rect 7196 5117 7205 5151
rect 7205 5117 7239 5151
rect 7239 5117 7248 5151
rect 7196 5108 7248 5117
rect 10692 5244 10744 5296
rect 11980 5312 12032 5364
rect 13176 5312 13228 5364
rect 13912 5312 13964 5364
rect 15108 5312 15160 5364
rect 12808 5244 12860 5296
rect 15660 5287 15712 5296
rect 15660 5253 15669 5287
rect 15669 5253 15703 5287
rect 15703 5253 15712 5287
rect 15660 5244 15712 5253
rect 9128 5176 9180 5228
rect 9772 5219 9824 5228
rect 9772 5185 9781 5219
rect 9781 5185 9815 5219
rect 9815 5185 9824 5219
rect 9772 5176 9824 5185
rect 11336 5219 11388 5228
rect 11336 5185 11345 5219
rect 11345 5185 11379 5219
rect 11379 5185 11388 5219
rect 11336 5176 11388 5185
rect 7380 5108 7432 5160
rect 4252 5040 4304 5092
rect 4160 4972 4212 5024
rect 6368 5040 6420 5092
rect 7104 5040 7156 5092
rect 8024 5040 8076 5092
rect 6092 4972 6144 5024
rect 6276 4972 6328 5024
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 10048 4972 10100 5024
rect 11060 4972 11112 5024
rect 12532 4972 12584 5024
rect 16304 5176 16356 5228
rect 13544 5151 13596 5160
rect 13544 5117 13553 5151
rect 13553 5117 13587 5151
rect 13587 5117 13596 5151
rect 13544 5108 13596 5117
rect 14740 5040 14792 5092
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 2228 4768 2280 4820
rect 2412 4700 2464 4752
rect 7104 4768 7156 4820
rect 7196 4768 7248 4820
rect 9220 4768 9272 4820
rect 11428 4768 11480 4820
rect 13728 4768 13780 4820
rect 13820 4768 13872 4820
rect 14740 4811 14792 4820
rect 2044 4564 2096 4616
rect 5080 4700 5132 4752
rect 5632 4700 5684 4752
rect 2688 4675 2740 4684
rect 2688 4641 2697 4675
rect 2697 4641 2731 4675
rect 2731 4641 2740 4675
rect 2688 4632 2740 4641
rect 3792 4675 3844 4684
rect 3240 4564 3292 4616
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 7564 4700 7616 4752
rect 5908 4675 5960 4684
rect 5908 4641 5917 4675
rect 5917 4641 5951 4675
rect 5951 4641 5960 4675
rect 5908 4632 5960 4641
rect 8300 4632 8352 4684
rect 8484 4675 8536 4684
rect 8484 4641 8493 4675
rect 8493 4641 8527 4675
rect 8527 4641 8536 4675
rect 8484 4632 8536 4641
rect 9220 4632 9272 4684
rect 5264 4607 5316 4616
rect 5264 4573 5273 4607
rect 5273 4573 5307 4607
rect 5307 4573 5316 4607
rect 5264 4564 5316 4573
rect 4344 4496 4396 4548
rect 5172 4496 5224 4548
rect 6000 4564 6052 4616
rect 8944 4564 8996 4616
rect 9680 4700 9732 4752
rect 11336 4743 11388 4752
rect 10600 4632 10652 4684
rect 11336 4709 11345 4743
rect 11345 4709 11379 4743
rect 11379 4709 11388 4743
rect 11336 4700 11388 4709
rect 10048 4564 10100 4616
rect 10140 4564 10192 4616
rect 11612 4632 11664 4684
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2228 4428 2280 4480
rect 3516 4428 3568 4480
rect 3976 4428 4028 4480
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 5632 4471 5684 4480
rect 5632 4437 5641 4471
rect 5641 4437 5675 4471
rect 5675 4437 5684 4471
rect 5632 4428 5684 4437
rect 7564 4496 7616 4548
rect 10876 4564 10928 4616
rect 11796 4564 11848 4616
rect 7012 4428 7064 4480
rect 7288 4471 7340 4480
rect 7288 4437 7297 4471
rect 7297 4437 7331 4471
rect 7331 4437 7340 4471
rect 7288 4428 7340 4437
rect 7472 4471 7524 4480
rect 7472 4437 7481 4471
rect 7481 4437 7515 4471
rect 7515 4437 7524 4471
rect 7472 4428 7524 4437
rect 8300 4471 8352 4480
rect 8300 4437 8309 4471
rect 8309 4437 8343 4471
rect 8343 4437 8352 4471
rect 8300 4428 8352 4437
rect 9036 4428 9088 4480
rect 9220 4471 9272 4480
rect 9220 4437 9229 4471
rect 9229 4437 9263 4471
rect 9263 4437 9272 4471
rect 9220 4428 9272 4437
rect 9404 4428 9456 4480
rect 9680 4428 9732 4480
rect 10324 4471 10376 4480
rect 10324 4437 10333 4471
rect 10333 4437 10367 4471
rect 10367 4437 10376 4471
rect 12532 4607 12584 4616
rect 12532 4573 12541 4607
rect 12541 4573 12575 4607
rect 12575 4573 12584 4607
rect 12532 4564 12584 4573
rect 13820 4564 13872 4616
rect 14740 4777 14749 4811
rect 14749 4777 14783 4811
rect 14783 4777 14792 4811
rect 14740 4768 14792 4777
rect 15752 4632 15804 4684
rect 12624 4496 12676 4548
rect 14464 4496 14516 4548
rect 15660 4496 15712 4548
rect 16396 4496 16448 4548
rect 10324 4428 10376 4437
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 1400 4224 1452 4276
rect 2688 4224 2740 4276
rect 3516 4224 3568 4276
rect 4436 4267 4488 4276
rect 4436 4233 4445 4267
rect 4445 4233 4479 4267
rect 4479 4233 4488 4267
rect 4436 4224 4488 4233
rect 4620 4224 4672 4276
rect 5632 4224 5684 4276
rect 6368 4224 6420 4276
rect 3792 4156 3844 4208
rect 4528 4156 4580 4208
rect 1676 4063 1728 4072
rect 1676 4029 1685 4063
rect 1685 4029 1719 4063
rect 1719 4029 1728 4063
rect 1676 4020 1728 4029
rect 2044 4020 2096 4072
rect 3516 4088 3568 4140
rect 204 3952 256 4004
rect 2136 3927 2188 3936
rect 2136 3893 2145 3927
rect 2145 3893 2179 3927
rect 2179 3893 2188 3927
rect 2136 3884 2188 3893
rect 4344 4131 4396 4140
rect 4344 4097 4353 4131
rect 4353 4097 4387 4131
rect 4387 4097 4396 4131
rect 4344 4088 4396 4097
rect 5264 4088 5316 4140
rect 5908 4088 5960 4140
rect 6460 4156 6512 4208
rect 8668 4156 8720 4208
rect 7288 4131 7340 4140
rect 7288 4097 7297 4131
rect 7297 4097 7331 4131
rect 7331 4097 7340 4131
rect 7288 4088 7340 4097
rect 9588 4224 9640 4276
rect 9864 4224 9916 4276
rect 10140 4224 10192 4276
rect 11428 4224 11480 4276
rect 12624 4224 12676 4276
rect 12716 4224 12768 4276
rect 13820 4224 13872 4276
rect 15476 4224 15528 4276
rect 9036 4088 9088 4140
rect 6276 4020 6328 4072
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 9312 4063 9364 4072
rect 9312 4029 9321 4063
rect 9321 4029 9355 4063
rect 9355 4029 9364 4063
rect 9312 4020 9364 4029
rect 9588 4088 9640 4140
rect 14556 4156 14608 4208
rect 10784 4088 10836 4140
rect 11060 4131 11112 4140
rect 11060 4097 11069 4131
rect 11069 4097 11103 4131
rect 11103 4097 11112 4131
rect 11060 4088 11112 4097
rect 11980 4131 12032 4140
rect 11980 4097 11989 4131
rect 11989 4097 12023 4131
rect 12023 4097 12032 4131
rect 11980 4088 12032 4097
rect 10692 4063 10744 4072
rect 8116 3952 8168 4004
rect 9496 3952 9548 4004
rect 9864 3952 9916 4004
rect 9956 3952 10008 4004
rect 10692 4029 10701 4063
rect 10701 4029 10735 4063
rect 10735 4029 10744 4063
rect 10692 4020 10744 4029
rect 11336 4020 11388 4072
rect 13728 4088 13780 4140
rect 13820 4088 13872 4140
rect 14832 4131 14884 4140
rect 14832 4097 14841 4131
rect 14841 4097 14875 4131
rect 14875 4097 14884 4131
rect 14832 4088 14884 4097
rect 15384 4131 15436 4140
rect 15384 4097 15393 4131
rect 15393 4097 15427 4131
rect 15427 4097 15436 4131
rect 15384 4088 15436 4097
rect 12532 4063 12584 4072
rect 12532 4029 12541 4063
rect 12541 4029 12575 4063
rect 12575 4029 12584 4063
rect 12532 4020 12584 4029
rect 3240 3884 3292 3936
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 5632 3884 5684 3936
rect 6092 3884 6144 3936
rect 7656 3884 7708 3936
rect 8484 3884 8536 3936
rect 9680 3884 9732 3936
rect 11612 3884 11664 3936
rect 12808 3884 12860 3936
rect 14464 3952 14516 4004
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 16488 3952 16540 4004
rect 14556 3884 14608 3936
rect 15844 3884 15896 3936
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 1952 3723 2004 3732
rect 1952 3689 1961 3723
rect 1961 3689 1995 3723
rect 1995 3689 2004 3723
rect 1952 3680 2004 3689
rect 3240 3680 3292 3732
rect 7380 3723 7432 3732
rect 1032 3612 1084 3664
rect 572 3544 624 3596
rect 2320 3612 2372 3664
rect 3148 3612 3200 3664
rect 2228 3544 2280 3596
rect 2504 3587 2556 3596
rect 2504 3553 2513 3587
rect 2513 3553 2547 3587
rect 2547 3553 2556 3587
rect 5448 3612 5500 3664
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 9404 3680 9456 3732
rect 2504 3544 2556 3553
rect 1860 3519 1912 3528
rect 1860 3485 1869 3519
rect 1869 3485 1903 3519
rect 1903 3485 1912 3519
rect 1860 3476 1912 3485
rect 2136 3476 2188 3528
rect 2228 3408 2280 3460
rect 3608 3544 3660 3596
rect 4436 3544 4488 3596
rect 5264 3544 5316 3596
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 7288 3544 7340 3596
rect 9772 3612 9824 3664
rect 12992 3680 13044 3732
rect 13544 3680 13596 3732
rect 10324 3612 10376 3664
rect 3608 3340 3660 3392
rect 3884 3383 3936 3392
rect 3884 3349 3893 3383
rect 3893 3349 3927 3383
rect 3927 3349 3936 3383
rect 3884 3340 3936 3349
rect 4344 3383 4396 3392
rect 4344 3349 4353 3383
rect 4353 3349 4387 3383
rect 4387 3349 4396 3383
rect 4344 3340 4396 3349
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 5724 3476 5776 3528
rect 7104 3476 7156 3528
rect 7564 3476 7616 3528
rect 8484 3519 8536 3528
rect 8484 3485 8502 3519
rect 8502 3485 8536 3519
rect 8484 3476 8536 3485
rect 8668 3476 8720 3528
rect 10968 3544 11020 3596
rect 13084 3544 13136 3596
rect 13176 3544 13228 3596
rect 13820 3544 13872 3596
rect 14464 3544 14516 3596
rect 14648 3544 14700 3596
rect 15292 3544 15344 3596
rect 9496 3519 9548 3528
rect 5448 3408 5500 3460
rect 9496 3485 9505 3519
rect 9505 3485 9539 3519
rect 9539 3485 9548 3519
rect 9496 3476 9548 3485
rect 10048 3519 10100 3528
rect 10048 3485 10057 3519
rect 10057 3485 10091 3519
rect 10091 3485 10100 3519
rect 10048 3476 10100 3485
rect 10232 3476 10284 3528
rect 11888 3476 11940 3528
rect 13544 3476 13596 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 14924 3476 14976 3528
rect 15936 3476 15988 3528
rect 4436 3340 4488 3349
rect 5172 3340 5224 3392
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 5540 3340 5592 3392
rect 5724 3383 5776 3392
rect 5724 3349 5733 3383
rect 5733 3349 5767 3383
rect 5767 3349 5776 3383
rect 5724 3340 5776 3349
rect 7748 3340 7800 3392
rect 7840 3340 7892 3392
rect 9312 3383 9364 3392
rect 9312 3349 9321 3383
rect 9321 3349 9355 3383
rect 9355 3349 9364 3383
rect 9312 3340 9364 3349
rect 12164 3408 12216 3460
rect 10048 3340 10100 3392
rect 11612 3340 11664 3392
rect 11888 3340 11940 3392
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 1400 2796 1452 2848
rect 4436 3136 4488 3188
rect 5172 3179 5224 3188
rect 1768 3068 1820 3120
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 3516 3068 3568 3120
rect 4160 3068 4212 3120
rect 5172 3145 5181 3179
rect 5181 3145 5215 3179
rect 5215 3145 5224 3179
rect 5172 3136 5224 3145
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 5724 3136 5776 3188
rect 6460 3136 6512 3188
rect 7472 3136 7524 3188
rect 5080 3068 5132 3120
rect 2044 3000 2096 3009
rect 4068 3000 4120 3052
rect 6184 3043 6236 3052
rect 3240 2932 3292 2984
rect 1860 2864 1912 2916
rect 3148 2864 3200 2916
rect 3516 2907 3568 2916
rect 3516 2873 3525 2907
rect 3525 2873 3559 2907
rect 3559 2873 3568 2907
rect 3516 2864 3568 2873
rect 3792 2932 3844 2984
rect 6184 3009 6193 3043
rect 6193 3009 6227 3043
rect 6227 3009 6236 3043
rect 6184 3000 6236 3009
rect 10140 3136 10192 3188
rect 11060 3136 11112 3188
rect 11244 3136 11296 3188
rect 12072 3136 12124 3188
rect 7656 3111 7708 3120
rect 7656 3077 7674 3111
rect 7674 3077 7708 3111
rect 7656 3068 7708 3077
rect 7840 3000 7892 3052
rect 8024 3043 8076 3052
rect 8024 3009 8033 3043
rect 8033 3009 8067 3043
rect 8067 3009 8076 3043
rect 8208 3043 8260 3052
rect 8024 3000 8076 3009
rect 8208 3009 8217 3043
rect 8217 3009 8251 3043
rect 8251 3009 8260 3043
rect 8208 3000 8260 3009
rect 4252 2864 4304 2916
rect 4988 2864 5040 2916
rect 5448 2932 5500 2984
rect 5724 2975 5776 2984
rect 5724 2941 5733 2975
rect 5733 2941 5767 2975
rect 5767 2941 5776 2975
rect 5724 2932 5776 2941
rect 9772 3043 9824 3052
rect 9772 3009 9781 3043
rect 9781 3009 9815 3043
rect 9815 3009 9824 3043
rect 9772 3000 9824 3009
rect 10968 3043 11020 3052
rect 11612 3068 11664 3120
rect 13084 3136 13136 3188
rect 12716 3111 12768 3120
rect 12716 3077 12725 3111
rect 12725 3077 12759 3111
rect 12759 3077 12768 3111
rect 12716 3068 12768 3077
rect 12992 3068 13044 3120
rect 13728 3068 13780 3120
rect 15568 3136 15620 3188
rect 10968 3009 10986 3043
rect 10986 3009 11020 3043
rect 10968 3000 11020 3009
rect 11704 3000 11756 3052
rect 5172 2864 5224 2916
rect 6368 2864 6420 2916
rect 9864 2907 9916 2916
rect 9864 2873 9873 2907
rect 9873 2873 9907 2907
rect 9907 2873 9916 2907
rect 9864 2864 9916 2873
rect 13084 3043 13136 3052
rect 12716 2932 12768 2984
rect 5264 2796 5316 2848
rect 9036 2796 9088 2848
rect 9588 2796 9640 2848
rect 11244 2796 11296 2848
rect 11612 2796 11664 2848
rect 13084 3009 13093 3043
rect 13093 3009 13127 3043
rect 13127 3009 13136 3043
rect 13084 3000 13136 3009
rect 13820 3000 13872 3052
rect 14740 3000 14792 3052
rect 15476 3043 15528 3052
rect 15476 3009 15485 3043
rect 15485 3009 15519 3043
rect 15519 3009 15528 3043
rect 15476 3000 15528 3009
rect 16028 2932 16080 2984
rect 16212 2864 16264 2916
rect 16948 2796 17000 2848
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 3516 2592 3568 2644
rect 4344 2592 4396 2644
rect 7748 2592 7800 2644
rect 9036 2635 9088 2644
rect 3976 2524 4028 2576
rect 5540 2524 5592 2576
rect 4344 2456 4396 2508
rect 5172 2499 5224 2508
rect 5172 2465 5181 2499
rect 5181 2465 5215 2499
rect 5215 2465 5224 2499
rect 5172 2456 5224 2465
rect 1584 2388 1636 2440
rect 1860 2431 1912 2440
rect 1860 2397 1869 2431
rect 1869 2397 1903 2431
rect 1903 2397 1912 2431
rect 2504 2431 2556 2440
rect 1860 2388 1912 2397
rect 2504 2397 2513 2431
rect 2513 2397 2547 2431
rect 2547 2397 2556 2431
rect 2504 2388 2556 2397
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 3608 2431 3660 2440
rect 3608 2397 3617 2431
rect 3617 2397 3651 2431
rect 3651 2397 3660 2431
rect 3608 2388 3660 2397
rect 4068 2431 4120 2440
rect 4068 2397 4077 2431
rect 4077 2397 4111 2431
rect 4111 2397 4120 2431
rect 4068 2388 4120 2397
rect 5264 2388 5316 2440
rect 5816 2431 5868 2440
rect 5816 2397 5825 2431
rect 5825 2397 5859 2431
rect 5859 2397 5868 2431
rect 5816 2388 5868 2397
rect 8300 2524 8352 2576
rect 9036 2601 9045 2635
rect 9045 2601 9079 2635
rect 9079 2601 9088 2635
rect 9036 2592 9088 2601
rect 10048 2592 10100 2644
rect 10784 2592 10836 2644
rect 10968 2592 11020 2644
rect 9128 2524 9180 2576
rect 3332 2320 3384 2372
rect 2320 2295 2372 2304
rect 2320 2261 2329 2295
rect 2329 2261 2363 2295
rect 2363 2261 2372 2295
rect 2320 2252 2372 2261
rect 3056 2295 3108 2304
rect 3056 2261 3065 2295
rect 3065 2261 3099 2295
rect 3099 2261 3108 2295
rect 3056 2252 3108 2261
rect 4620 2320 4672 2372
rect 5356 2320 5408 2372
rect 3884 2295 3936 2304
rect 3884 2261 3893 2295
rect 3893 2261 3927 2295
rect 3927 2261 3936 2295
rect 3884 2252 3936 2261
rect 4160 2252 4212 2304
rect 5448 2295 5500 2304
rect 5448 2261 5457 2295
rect 5457 2261 5491 2295
rect 5491 2261 5500 2295
rect 5448 2252 5500 2261
rect 6552 2363 6604 2372
rect 6552 2329 6561 2363
rect 6561 2329 6595 2363
rect 6595 2329 6604 2363
rect 8116 2456 8168 2508
rect 7380 2388 7432 2440
rect 7472 2431 7524 2440
rect 7472 2397 7492 2431
rect 7492 2397 7524 2431
rect 7472 2388 7524 2397
rect 8392 2431 8444 2440
rect 8392 2397 8401 2431
rect 8401 2397 8435 2431
rect 8435 2397 8444 2431
rect 8392 2388 8444 2397
rect 9220 2388 9272 2440
rect 10692 2524 10744 2576
rect 9588 2499 9640 2508
rect 9588 2465 9597 2499
rect 9597 2465 9631 2499
rect 9631 2465 9640 2499
rect 9588 2456 9640 2465
rect 9864 2456 9916 2508
rect 11704 2456 11756 2508
rect 13728 2592 13780 2644
rect 12532 2456 12584 2508
rect 15016 2524 15068 2576
rect 15476 2456 15528 2508
rect 9680 2388 9732 2440
rect 10048 2431 10100 2440
rect 10048 2397 10057 2431
rect 10057 2397 10091 2431
rect 10091 2397 10100 2431
rect 10048 2388 10100 2397
rect 10232 2431 10284 2440
rect 10232 2397 10241 2431
rect 10241 2397 10275 2431
rect 10275 2397 10284 2431
rect 10232 2388 10284 2397
rect 11244 2388 11296 2440
rect 12992 2431 13044 2440
rect 12992 2397 13001 2431
rect 13001 2397 13035 2431
rect 13035 2397 13044 2431
rect 12992 2388 13044 2397
rect 13912 2431 13964 2440
rect 13912 2397 13921 2431
rect 13921 2397 13955 2431
rect 13955 2397 13964 2431
rect 13912 2388 13964 2397
rect 14556 2431 14608 2440
rect 14556 2397 14565 2431
rect 14565 2397 14599 2431
rect 14599 2397 14608 2431
rect 14556 2388 14608 2397
rect 14832 2431 14884 2440
rect 14832 2397 14841 2431
rect 14841 2397 14875 2431
rect 14875 2397 14884 2431
rect 14832 2388 14884 2397
rect 7196 2363 7248 2372
rect 6552 2320 6604 2329
rect 7196 2329 7205 2363
rect 7205 2329 7239 2363
rect 7239 2329 7248 2363
rect 7196 2320 7248 2329
rect 6368 2252 6420 2304
rect 7012 2252 7064 2304
rect 8024 2320 8076 2372
rect 11888 2320 11940 2372
rect 12716 2320 12768 2372
rect 13544 2320 13596 2372
rect 7656 2252 7708 2304
rect 10048 2252 10100 2304
rect 13728 2252 13780 2304
rect 14188 2295 14240 2304
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 16396 2252 16448 2304
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 2320 2048 2372 2100
rect 5172 2048 5224 2100
rect 5448 2048 5500 2100
rect 9772 2048 9824 2100
rect 10232 2048 10284 2100
rect 13544 2048 13596 2100
rect 14556 2048 14608 2100
rect 3056 1980 3108 2032
rect 6000 1980 6052 2032
rect 11428 1980 11480 2032
rect 14188 1980 14240 2032
rect 3608 1912 3660 1964
rect 9312 1912 9364 1964
rect 2504 1844 2556 1896
rect 4528 1844 4580 1896
rect 6552 1844 6604 1896
rect 8852 1844 8904 1896
rect 9220 1844 9272 1896
rect 13360 1844 13412 1896
rect 3700 1776 3752 1828
rect 6368 1776 6420 1828
rect 8208 1776 8260 1828
rect 5540 1708 5592 1760
rect 7288 1708 7340 1760
rect 7380 1708 7432 1760
rect 10324 1708 10376 1760
rect 1676 1640 1728 1692
rect 8300 1640 8352 1692
rect 3884 1572 3936 1624
rect 6828 1572 6880 1624
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 938 19200 994 20000
rect 1398 19200 1454 20000
rect 1766 19200 1822 20000
rect 2226 19200 2282 20000
rect 2594 19200 2650 20000
rect 3054 19200 3110 20000
rect 3422 19200 3478 20000
rect 3882 19200 3938 20000
rect 4250 19200 4306 20000
rect 4618 19200 4674 20000
rect 5078 19200 5134 20000
rect 5446 19200 5502 20000
rect 5906 19200 5962 20000
rect 6274 19200 6330 20000
rect 6734 19200 6790 20000
rect 7102 19200 7158 20000
rect 7562 19200 7618 20000
rect 7930 19200 7986 20000
rect 8390 19200 8446 20000
rect 8758 19200 8814 20000
rect 9126 19200 9182 20000
rect 9586 19200 9642 20000
rect 9954 19200 10010 20000
rect 10414 19200 10470 20000
rect 10520 19230 10732 19258
rect 216 17542 244 19200
rect 204 17536 256 17542
rect 204 17478 256 17484
rect 584 16250 612 19200
rect 952 16454 980 19200
rect 940 16448 992 16454
rect 940 16390 992 16396
rect 572 16244 624 16250
rect 572 16186 624 16192
rect 1412 15978 1440 19200
rect 1780 17338 1808 19200
rect 1858 17640 1914 17649
rect 1858 17575 1914 17584
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1872 16794 1900 17575
rect 2240 17338 2268 19200
rect 2608 17338 2636 19200
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 1860 16788 1912 16794
rect 1860 16730 1912 16736
rect 1492 16720 1544 16726
rect 1490 16688 1492 16697
rect 1544 16688 1546 16697
rect 1490 16623 1546 16632
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1400 15972 1452 15978
rect 1400 15914 1452 15920
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15745 1532 15846
rect 1490 15736 1546 15745
rect 1596 15706 1624 16050
rect 1780 15706 1808 16050
rect 1964 15706 1992 16526
rect 2148 16250 2176 17138
rect 2792 16980 2820 19071
rect 3068 17338 3096 19200
rect 3330 18592 3386 18601
rect 3330 18527 3386 18536
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3148 17196 3200 17202
rect 3344 17184 3372 18527
rect 3436 17338 3464 19200
rect 3792 17536 3844 17542
rect 3792 17478 3844 17484
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3608 17196 3660 17202
rect 3344 17156 3464 17184
rect 3148 17138 3200 17144
rect 2700 16952 2820 16980
rect 2700 16794 2728 16952
rect 2824 16892 3132 16912
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16816 3132 16836
rect 2688 16788 2740 16794
rect 2688 16730 2740 16736
rect 3160 16726 3188 17138
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3148 16720 3200 16726
rect 3148 16662 3200 16668
rect 2412 16584 2464 16590
rect 2412 16526 2464 16532
rect 2504 16584 2556 16590
rect 2504 16526 2556 16532
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2228 16176 2280 16182
rect 2228 16118 2280 16124
rect 1490 15671 1546 15680
rect 1584 15700 1636 15706
rect 1584 15642 1636 15648
rect 1768 15700 1820 15706
rect 1768 15642 1820 15648
rect 1952 15700 2004 15706
rect 1952 15642 2004 15648
rect 1952 15496 2004 15502
rect 1952 15438 2004 15444
rect 1584 14816 1636 14822
rect 1490 14784 1546 14793
rect 1584 14758 1636 14764
rect 1490 14719 1546 14728
rect 1504 14618 1532 14719
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1596 14482 1624 14758
rect 1584 14476 1636 14482
rect 1584 14418 1636 14424
rect 1964 14113 1992 15438
rect 1950 14104 2006 14113
rect 1950 14039 2006 14048
rect 1490 13832 1546 13841
rect 1490 13767 1492 13776
rect 1544 13767 1546 13776
rect 1492 13738 1544 13744
rect 2240 13705 2268 16118
rect 2320 16040 2372 16046
rect 2320 15982 2372 15988
rect 2332 15722 2360 15982
rect 2424 15978 2452 16526
rect 2412 15972 2464 15978
rect 2412 15914 2464 15920
rect 2332 15694 2452 15722
rect 2516 15706 2544 16526
rect 2596 16516 2648 16522
rect 2596 16458 2648 16464
rect 2608 16402 2636 16458
rect 2608 16374 2728 16402
rect 2596 16108 2648 16114
rect 2596 16050 2648 16056
rect 2318 15600 2374 15609
rect 2318 15535 2374 15544
rect 2332 15502 2360 15535
rect 2320 15496 2372 15502
rect 2320 15438 2372 15444
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2226 13696 2282 13705
rect 2226 13631 2282 13640
rect 2240 13258 2268 13631
rect 2332 13530 2360 14214
rect 2320 13524 2372 13530
rect 2320 13466 2372 13472
rect 1308 13252 1360 13258
rect 1308 13194 1360 13200
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 204 4004 256 4010
rect 204 3946 256 3952
rect 216 800 244 3946
rect 1032 3664 1084 3670
rect 1032 3606 1084 3612
rect 572 3596 624 3602
rect 572 3538 624 3544
rect 584 800 612 3538
rect 1044 800 1072 3606
rect 1320 2938 1348 13194
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1952 13184 2004 13190
rect 1952 13126 2004 13132
rect 1504 12889 1532 13126
rect 1964 12986 1992 13126
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1490 12880 1546 12889
rect 1490 12815 1546 12824
rect 2136 12844 2188 12850
rect 2136 12786 2188 12792
rect 1584 12640 1636 12646
rect 1584 12582 1636 12588
rect 1596 12481 1624 12582
rect 1582 12472 1638 12481
rect 2148 12442 2176 12786
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 1582 12407 1638 12416
rect 2136 12436 2188 12442
rect 2136 12378 2188 12384
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11558 1440 12174
rect 1400 11552 1452 11558
rect 1400 11494 1452 11500
rect 1412 11218 1440 11494
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1492 11008 1544 11014
rect 1490 10976 1492 10985
rect 1544 10976 1546 10985
rect 1490 10911 1546 10920
rect 1688 10810 1716 11086
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1858 10704 1914 10713
rect 1858 10639 1914 10648
rect 1490 10024 1546 10033
rect 1490 9959 1546 9968
rect 1504 9926 1532 9959
rect 1872 9926 1900 10639
rect 1952 10056 2004 10062
rect 1952 9998 2004 10004
rect 1492 9920 1544 9926
rect 1860 9920 1912 9926
rect 1492 9862 1544 9868
rect 1858 9888 1860 9897
rect 1912 9888 1914 9897
rect 1858 9823 1914 9832
rect 1400 9716 1452 9722
rect 1400 9658 1452 9664
rect 1412 7018 1440 9658
rect 1768 9580 1820 9586
rect 1768 9522 1820 9528
rect 1676 9444 1728 9450
rect 1676 9386 1728 9392
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1504 9081 1532 9318
rect 1490 9072 1546 9081
rect 1490 9007 1546 9016
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 1504 8129 1532 8298
rect 1490 8120 1546 8129
rect 1490 8055 1546 8064
rect 1492 7200 1544 7206
rect 1490 7168 1492 7177
rect 1544 7168 1546 7177
rect 1490 7103 1546 7112
rect 1412 6990 1532 7018
rect 1400 6928 1452 6934
rect 1400 6870 1452 6876
rect 1412 4282 1440 6870
rect 1504 6322 1532 6990
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1490 6216 1546 6225
rect 1490 6151 1492 6160
rect 1544 6151 1546 6160
rect 1492 6122 1544 6128
rect 1492 5364 1544 5370
rect 1492 5306 1544 5312
rect 1504 5273 1532 5306
rect 1490 5264 1546 5273
rect 1490 5199 1546 5208
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4321 1532 4422
rect 1490 4312 1546 4321
rect 1400 4276 1452 4282
rect 1490 4247 1546 4256
rect 1400 4218 1452 4224
rect 1398 4040 1454 4049
rect 1398 3975 1454 3984
rect 1412 3058 1440 3975
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1320 2910 1532 2938
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 1412 800 1440 2790
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1398 0 1454 800
rect 1504 513 1532 2910
rect 1596 2446 1624 9318
rect 1688 8974 1716 9386
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 7410 1716 8774
rect 1780 8634 1808 9522
rect 1964 9489 1992 9998
rect 1950 9480 2006 9489
rect 1950 9415 2006 9424
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1768 8288 1820 8294
rect 1768 8230 1820 8236
rect 1780 7886 1808 8230
rect 1768 7880 1820 7886
rect 1872 7857 1900 8434
rect 2056 7886 2084 11018
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2044 7880 2096 7886
rect 1768 7822 1820 7828
rect 1858 7848 1914 7857
rect 1858 7783 1914 7792
rect 1964 7828 2044 7834
rect 1964 7822 2096 7828
rect 1964 7806 2084 7822
rect 1860 7744 1912 7750
rect 1860 7686 1912 7692
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1676 6860 1728 6866
rect 1676 6802 1728 6808
rect 1688 6458 1716 6802
rect 1768 6656 1820 6662
rect 1768 6598 1820 6604
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1688 5642 1716 6394
rect 1676 5636 1728 5642
rect 1676 5578 1728 5584
rect 1780 5370 1808 6598
rect 1768 5364 1820 5370
rect 1768 5306 1820 5312
rect 1676 4072 1728 4078
rect 1676 4014 1728 4020
rect 1584 2440 1636 2446
rect 1584 2382 1636 2388
rect 1688 1698 1716 4014
rect 1872 3534 1900 7686
rect 1964 6934 1992 7806
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1952 6928 2004 6934
rect 1952 6870 2004 6876
rect 1952 6724 2004 6730
rect 1952 6666 2004 6672
rect 1964 3738 1992 6666
rect 2056 4622 2084 7686
rect 2148 5370 2176 9318
rect 2240 8673 2268 12582
rect 2424 12209 2452 15694
rect 2504 15700 2556 15706
rect 2504 15642 2556 15648
rect 2608 15638 2636 16050
rect 2700 15706 2728 16374
rect 2976 16046 3004 16526
rect 3252 16250 3280 17070
rect 3332 17060 3384 17066
rect 3332 17002 3384 17008
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3240 16108 3292 16114
rect 3240 16050 3292 16056
rect 2964 16040 3016 16046
rect 2964 15982 3016 15988
rect 2824 15804 3132 15824
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15728 3132 15748
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2596 15632 2648 15638
rect 2596 15574 2648 15580
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 3148 15496 3200 15502
rect 3148 15438 3200 15444
rect 2516 12374 2544 15438
rect 2688 15020 2740 15026
rect 2688 14962 2740 14968
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2608 12374 2636 13874
rect 2700 13870 2728 14962
rect 2824 14716 3132 14736
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14640 3132 14660
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2780 14272 2832 14278
rect 2780 14214 2832 14220
rect 2792 14006 2820 14214
rect 2884 14074 2912 14486
rect 2964 14340 3016 14346
rect 2964 14282 3016 14288
rect 2976 14074 3004 14282
rect 2872 14068 2924 14074
rect 2872 14010 2924 14016
rect 2964 14068 3016 14074
rect 2964 14010 3016 14016
rect 2780 14000 2832 14006
rect 2780 13942 2832 13948
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2824 13628 3132 13648
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13552 3132 13572
rect 2872 13388 2924 13394
rect 2872 13330 2924 13336
rect 2884 12714 2912 13330
rect 3160 13326 3188 15438
rect 3252 14362 3280 16050
rect 3344 15706 3372 17002
rect 3436 16114 3464 17156
rect 3608 17138 3660 17144
rect 3516 16584 3568 16590
rect 3516 16526 3568 16532
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3424 15360 3476 15366
rect 3424 15302 3476 15308
rect 3332 15020 3384 15026
rect 3332 14962 3384 14968
rect 3344 14482 3372 14962
rect 3332 14476 3384 14482
rect 3332 14418 3384 14424
rect 3252 14334 3372 14362
rect 3240 14000 3292 14006
rect 3238 13968 3240 13977
rect 3292 13968 3294 13977
rect 3238 13903 3294 13912
rect 3344 13410 3372 14334
rect 3436 13433 3464 15302
rect 3252 13394 3372 13410
rect 3240 13388 3372 13394
rect 3292 13382 3372 13388
rect 3422 13424 3478 13433
rect 3528 13410 3556 16526
rect 3620 16250 3648 17138
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3606 16008 3662 16017
rect 3712 15978 3740 17206
rect 3804 17202 3832 17478
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3792 16788 3844 16794
rect 3896 16776 3924 19200
rect 4264 17066 4292 19200
rect 4632 17338 4660 19200
rect 4698 17436 5006 17456
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17360 5006 17380
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4344 17196 4396 17202
rect 4344 17138 4396 17144
rect 4436 17196 4488 17202
rect 4436 17138 4488 17144
rect 4620 17196 4672 17202
rect 4620 17138 4672 17144
rect 4252 17060 4304 17066
rect 4252 17002 4304 17008
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 3844 16748 3924 16776
rect 3792 16730 3844 16736
rect 3988 16697 4016 16934
rect 3974 16688 4030 16697
rect 3974 16623 4030 16632
rect 3790 16552 3846 16561
rect 3790 16487 3792 16496
rect 3844 16487 3846 16496
rect 3792 16458 3844 16464
rect 4356 16250 4384 17138
rect 4448 16794 4476 17138
rect 4436 16788 4488 16794
rect 4436 16730 4488 16736
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4344 16244 4396 16250
rect 4344 16186 4396 16192
rect 4436 16176 4488 16182
rect 4066 16144 4122 16153
rect 3792 16108 3844 16114
rect 3792 16050 3844 16056
rect 3976 16108 4028 16114
rect 4436 16118 4488 16124
rect 4066 16079 4122 16088
rect 4252 16108 4304 16114
rect 3976 16050 4028 16056
rect 3606 15943 3662 15952
rect 3700 15972 3752 15978
rect 3620 15910 3648 15943
rect 3700 15914 3752 15920
rect 3608 15904 3660 15910
rect 3608 15846 3660 15852
rect 3606 15736 3662 15745
rect 3606 15671 3608 15680
rect 3660 15671 3662 15680
rect 3608 15642 3660 15648
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3608 14272 3660 14278
rect 3608 14214 3660 14220
rect 3620 14074 3648 14214
rect 3608 14068 3660 14074
rect 3608 14010 3660 14016
rect 3528 13382 3648 13410
rect 3422 13359 3478 13368
rect 3240 13330 3292 13336
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3240 13252 3292 13258
rect 3240 13194 3292 13200
rect 3252 12986 3280 13194
rect 3424 13184 3476 13190
rect 3424 13126 3476 13132
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3148 12844 3200 12850
rect 3148 12786 3200 12792
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2824 12540 3132 12560
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12464 3132 12484
rect 2504 12368 2556 12374
rect 2504 12310 2556 12316
rect 2596 12368 2648 12374
rect 2596 12310 2648 12316
rect 2410 12200 2466 12209
rect 2872 12164 2924 12170
rect 2410 12135 2466 12144
rect 2320 12096 2372 12102
rect 2320 12038 2372 12044
rect 2332 11937 2360 12038
rect 2318 11928 2374 11937
rect 2318 11863 2374 11872
rect 2424 11642 2452 12135
rect 2700 12124 2872 12152
rect 2424 11614 2544 11642
rect 2412 11552 2464 11558
rect 2412 11494 2464 11500
rect 2424 11218 2452 11494
rect 2412 11212 2464 11218
rect 2412 11154 2464 11160
rect 2412 10056 2464 10062
rect 2410 10024 2412 10033
rect 2464 10024 2466 10033
rect 2410 9959 2466 9968
rect 2516 9654 2544 11614
rect 2700 11354 2728 12124
rect 2872 12106 2924 12112
rect 3160 11762 3188 12786
rect 3252 12306 3280 12922
rect 3330 12472 3386 12481
rect 3436 12442 3464 13126
rect 3330 12407 3332 12416
rect 3384 12407 3386 12416
rect 3424 12436 3476 12442
rect 3332 12378 3384 12384
rect 3424 12378 3476 12384
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3528 12170 3556 13262
rect 3620 12753 3648 13382
rect 3606 12744 3662 12753
rect 3606 12679 3662 12688
rect 3606 12608 3662 12617
rect 3606 12543 3662 12552
rect 3620 12374 3648 12543
rect 3608 12368 3660 12374
rect 3608 12310 3660 12316
rect 3516 12164 3568 12170
rect 3516 12106 3568 12112
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3148 11756 3200 11762
rect 3148 11698 3200 11704
rect 2824 11452 3132 11472
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11376 3132 11396
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2872 11280 2924 11286
rect 2872 11222 2924 11228
rect 2780 11212 2832 11218
rect 2780 11154 2832 11160
rect 2792 11098 2820 11154
rect 2700 11070 2820 11098
rect 2884 11082 2912 11222
rect 3056 11144 3108 11150
rect 3160 11132 3188 11698
rect 3108 11104 3188 11132
rect 3056 11086 3108 11092
rect 2872 11076 2924 11082
rect 2700 10554 2728 11070
rect 2872 11018 2924 11024
rect 3160 10810 3188 11104
rect 3252 11014 3280 11834
rect 3424 11824 3476 11830
rect 3424 11766 3476 11772
rect 3332 11688 3384 11694
rect 3332 11630 3384 11636
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 2700 10538 2820 10554
rect 2700 10532 2832 10538
rect 2700 10526 2780 10532
rect 2700 10130 2728 10526
rect 2780 10474 2832 10480
rect 2824 10364 3132 10384
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10288 3132 10308
rect 3344 10266 3372 11630
rect 3436 11218 3464 11766
rect 3528 11626 3556 12106
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3516 11620 3568 11626
rect 3516 11562 3568 11568
rect 3620 11354 3648 11698
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3712 10266 3740 14418
rect 3804 12481 3832 16050
rect 3884 15972 3936 15978
rect 3884 15914 3936 15920
rect 3896 14278 3924 15914
rect 3884 14272 3936 14278
rect 3884 14214 3936 14220
rect 3896 13977 3924 14214
rect 3882 13968 3938 13977
rect 3882 13903 3938 13912
rect 3988 13920 4016 16050
rect 4080 15638 4108 16079
rect 4252 16050 4304 16056
rect 4068 15632 4120 15638
rect 4068 15574 4120 15580
rect 4264 15337 4292 16050
rect 4448 15706 4476 16118
rect 4540 15706 4568 16526
rect 4632 16250 4660 17138
rect 5092 16454 5120 19200
rect 5172 17196 5224 17202
rect 5172 17138 5224 17144
rect 5184 16794 5212 17138
rect 5460 17066 5488 19200
rect 5540 17604 5592 17610
rect 5540 17546 5592 17552
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5552 16998 5580 17546
rect 5920 17338 5948 19200
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5632 17264 5684 17270
rect 5684 17224 5764 17252
rect 5632 17206 5684 17212
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5172 16584 5224 16590
rect 5172 16526 5224 16532
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 4698 16348 5006 16368
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16272 5006 16292
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4988 16108 5040 16114
rect 5040 16068 5120 16096
rect 4988 16050 5040 16056
rect 4712 16040 4764 16046
rect 4712 15982 4764 15988
rect 4436 15700 4488 15706
rect 4436 15642 4488 15648
rect 4528 15700 4580 15706
rect 4528 15642 4580 15648
rect 4528 15564 4580 15570
rect 4528 15506 4580 15512
rect 4436 15496 4488 15502
rect 4436 15438 4488 15444
rect 4344 15360 4396 15366
rect 4250 15328 4306 15337
rect 4344 15302 4396 15308
rect 4250 15263 4306 15272
rect 4356 15144 4384 15302
rect 4172 15116 4384 15144
rect 4068 14952 4120 14958
rect 4068 14894 4120 14900
rect 4080 14482 4108 14894
rect 4068 14476 4120 14482
rect 4068 14418 4120 14424
rect 4172 14385 4200 15116
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4264 14822 4292 14962
rect 4342 14920 4398 14929
rect 4342 14855 4398 14864
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14074 4200 14214
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4252 14068 4304 14074
rect 4252 14010 4304 14016
rect 3988 13892 4108 13920
rect 3884 13864 3936 13870
rect 3884 13806 3936 13812
rect 3896 13394 3924 13806
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3988 13326 4016 13738
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4080 12850 4108 13892
rect 4160 13864 4212 13870
rect 4160 13806 4212 13812
rect 4172 13462 4200 13806
rect 4160 13456 4212 13462
rect 4160 13398 4212 13404
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 3790 12472 3846 12481
rect 3790 12407 3846 12416
rect 4080 12170 4108 12786
rect 4264 12434 4292 14010
rect 4356 13938 4384 14855
rect 4448 14822 4476 15438
rect 4540 15162 4568 15506
rect 4724 15473 4752 15982
rect 4710 15464 4766 15473
rect 4710 15399 4766 15408
rect 4698 15260 5006 15280
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15184 5006 15204
rect 4528 15156 4580 15162
rect 4528 15098 4580 15104
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4436 14816 4488 14822
rect 4436 14758 4488 14764
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4344 13932 4396 13938
rect 4344 13874 4396 13880
rect 4448 13734 4476 14758
rect 4540 14346 4568 14758
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4526 14104 4582 14113
rect 4526 14039 4582 14048
rect 4540 14006 4568 14039
rect 4528 14000 4580 14006
rect 4528 13942 4580 13948
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4172 12406 4292 12434
rect 4068 12164 4120 12170
rect 4068 12106 4120 12112
rect 4080 11898 4108 12106
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 3974 11792 4030 11801
rect 3974 11727 4030 11736
rect 3792 11688 3844 11694
rect 3792 11630 3844 11636
rect 3804 11354 3832 11630
rect 3884 11552 3936 11558
rect 3884 11494 3936 11500
rect 3792 11348 3844 11354
rect 3792 11290 3844 11296
rect 3896 11082 3924 11494
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3700 10260 3752 10266
rect 3700 10202 3752 10208
rect 2688 10124 2740 10130
rect 2688 10066 2740 10072
rect 3700 10124 3752 10130
rect 3700 10066 3752 10072
rect 3332 9920 3384 9926
rect 3330 9888 3332 9897
rect 3384 9888 3386 9897
rect 3330 9823 3386 9832
rect 2504 9648 2556 9654
rect 2502 9616 2504 9625
rect 2556 9616 2558 9625
rect 2412 9580 2464 9586
rect 2502 9551 2558 9560
rect 3148 9580 3200 9586
rect 2412 9522 2464 9528
rect 3148 9522 3200 9528
rect 2320 8900 2372 8906
rect 2320 8842 2372 8848
rect 2226 8664 2282 8673
rect 2226 8599 2282 8608
rect 2228 8356 2280 8362
rect 2228 8298 2280 8304
rect 2240 7410 2268 8298
rect 2332 7478 2360 8842
rect 2424 8242 2452 9522
rect 2504 9512 2556 9518
rect 2504 9454 2556 9460
rect 2516 9382 2544 9454
rect 2504 9376 2556 9382
rect 2504 9318 2556 9324
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2516 9081 2544 9318
rect 2502 9072 2558 9081
rect 2502 9007 2558 9016
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2516 8401 2544 8434
rect 2502 8392 2558 8401
rect 2502 8327 2558 8336
rect 2424 8214 2544 8242
rect 2320 7472 2372 7478
rect 2320 7414 2372 7420
rect 2228 7404 2280 7410
rect 2228 7346 2280 7352
rect 2412 7404 2464 7410
rect 2412 7346 2464 7352
rect 2228 7200 2280 7206
rect 2228 7142 2280 7148
rect 2240 6914 2268 7142
rect 2240 6886 2360 6914
rect 2228 6112 2280 6118
rect 2228 6054 2280 6060
rect 2240 5370 2268 6054
rect 2136 5364 2188 5370
rect 2136 5306 2188 5312
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2134 5264 2190 5273
rect 2134 5199 2136 5208
rect 2188 5199 2190 5208
rect 2136 5170 2188 5176
rect 2228 5160 2280 5166
rect 2228 5102 2280 5108
rect 2240 4826 2268 5102
rect 2228 4820 2280 4826
rect 2228 4762 2280 4768
rect 2044 4616 2096 4622
rect 2044 4558 2096 4564
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2044 4072 2096 4078
rect 2044 4014 2096 4020
rect 1952 3732 2004 3738
rect 1952 3674 2004 3680
rect 1860 3528 1912 3534
rect 1860 3470 1912 3476
rect 1768 3120 1820 3126
rect 1768 3062 1820 3068
rect 1950 3088 2006 3097
rect 1780 2292 1808 3062
rect 2056 3058 2084 4014
rect 2136 3936 2188 3942
rect 2136 3878 2188 3884
rect 2148 3534 2176 3878
rect 2240 3602 2268 4422
rect 2332 3670 2360 6886
rect 2424 6497 2452 7346
rect 2410 6488 2466 6497
rect 2410 6423 2466 6432
rect 2412 6316 2464 6322
rect 2412 6258 2464 6264
rect 2424 4758 2452 6258
rect 2516 5302 2544 8214
rect 2608 7970 2636 9318
rect 2824 9276 3132 9296
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9200 3132 9220
rect 3160 8634 3188 9522
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3148 8492 3200 8498
rect 3148 8434 3200 8440
rect 2824 8188 3132 8208
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8112 3132 8132
rect 3056 8016 3108 8022
rect 2608 7954 2728 7970
rect 3056 7958 3108 7964
rect 2596 7948 2728 7954
rect 2648 7942 2728 7948
rect 2596 7890 2648 7896
rect 2596 7812 2648 7818
rect 2596 7754 2648 7760
rect 2608 7449 2636 7754
rect 2594 7440 2650 7449
rect 2700 7410 2728 7942
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 2594 7375 2650 7384
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2596 7200 2648 7206
rect 2792 7188 2820 7686
rect 3068 7342 3096 7958
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2596 7142 2648 7148
rect 2700 7160 2820 7188
rect 2504 5296 2556 5302
rect 2504 5238 2556 5244
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2412 4752 2464 4758
rect 2412 4694 2464 4700
rect 2320 3664 2372 3670
rect 2320 3606 2372 3612
rect 2516 3602 2544 5102
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2504 3596 2556 3602
rect 2504 3538 2556 3544
rect 2136 3528 2188 3534
rect 2136 3470 2188 3476
rect 2228 3460 2280 3466
rect 2228 3402 2280 3408
rect 1950 3023 1952 3032
rect 2004 3023 2006 3032
rect 2044 3052 2096 3058
rect 1952 2994 2004 3000
rect 2044 2994 2096 3000
rect 1860 2916 1912 2922
rect 1860 2858 1912 2864
rect 1872 2446 1900 2858
rect 1860 2440 1912 2446
rect 1860 2382 1912 2388
rect 1780 2264 1900 2292
rect 1676 1692 1728 1698
rect 1676 1634 1728 1640
rect 1872 800 1900 2264
rect 2240 800 2268 3402
rect 2504 2440 2556 2446
rect 2504 2382 2556 2388
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2332 2106 2360 2246
rect 2320 2100 2372 2106
rect 2320 2042 2372 2048
rect 2516 1902 2544 2382
rect 2504 1896 2556 1902
rect 2504 1838 2556 1844
rect 2608 1748 2636 7142
rect 2700 6914 2728 7160
rect 2824 7100 3132 7120
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7024 3132 7044
rect 2700 6886 2820 6914
rect 2792 6730 2820 6886
rect 2780 6724 2832 6730
rect 2780 6666 2832 6672
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 2700 5574 2728 6258
rect 3068 6225 3096 6598
rect 3054 6216 3110 6225
rect 3054 6151 3110 6160
rect 2824 6012 3132 6032
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5936 3132 5956
rect 3160 5846 3188 8434
rect 3252 7546 3280 8910
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 7750 3372 8230
rect 3332 7744 3384 7750
rect 3332 7686 3384 7692
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3252 6798 3280 7482
rect 3344 7410 3372 7686
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3344 6644 3372 6734
rect 3252 6616 3372 6644
rect 3148 5840 3200 5846
rect 3148 5782 3200 5788
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2688 5568 2740 5574
rect 2688 5510 2740 5516
rect 2700 5166 2728 5510
rect 3068 5370 3096 5646
rect 2872 5364 2924 5370
rect 2872 5306 2924 5312
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2688 5160 2740 5166
rect 2688 5102 2740 5108
rect 2792 5012 2820 5170
rect 2884 5166 2912 5306
rect 3148 5296 3200 5302
rect 3148 5238 3200 5244
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2700 4984 2820 5012
rect 2700 4808 2728 4984
rect 2824 4924 3132 4944
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4848 3132 4868
rect 2700 4780 2820 4808
rect 2688 4684 2740 4690
rect 2688 4626 2740 4632
rect 2700 4282 2728 4626
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2792 4026 2820 4780
rect 2700 3998 2820 4026
rect 2700 3720 2728 3998
rect 2824 3836 3132 3856
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3760 3132 3780
rect 2700 3692 2820 3720
rect 2792 2836 2820 3692
rect 3160 3670 3188 5238
rect 3252 4706 3280 6616
rect 3436 6390 3464 8298
rect 3528 8022 3556 8842
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3516 8016 3568 8022
rect 3516 7958 3568 7964
rect 3516 7880 3568 7886
rect 3516 7822 3568 7828
rect 3424 6384 3476 6390
rect 3424 6326 3476 6332
rect 3424 6248 3476 6254
rect 3330 6216 3386 6225
rect 3424 6190 3476 6196
rect 3330 6151 3386 6160
rect 3344 5642 3372 6151
rect 3332 5636 3384 5642
rect 3332 5578 3384 5584
rect 3436 5370 3464 6190
rect 3528 5778 3556 7822
rect 3620 7546 3648 8366
rect 3712 8294 3740 10066
rect 3988 9518 4016 11727
rect 4066 10568 4122 10577
rect 4066 10503 4122 10512
rect 4080 10266 4108 10503
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 9178 4016 9454
rect 3792 9172 3844 9178
rect 3792 9114 3844 9120
rect 3976 9172 4028 9178
rect 3976 9114 4028 9120
rect 3700 8288 3752 8294
rect 3700 8230 3752 8236
rect 3700 8084 3752 8090
rect 3700 8026 3752 8032
rect 3712 7750 3740 8026
rect 3700 7744 3752 7750
rect 3700 7686 3752 7692
rect 3608 7540 3660 7546
rect 3608 7482 3660 7488
rect 3700 7336 3752 7342
rect 3700 7278 3752 7284
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3620 6225 3648 6734
rect 3606 6216 3662 6225
rect 3606 6151 3662 6160
rect 3608 6112 3660 6118
rect 3608 6054 3660 6060
rect 3516 5772 3568 5778
rect 3516 5714 3568 5720
rect 3514 5536 3570 5545
rect 3514 5471 3570 5480
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3422 5264 3478 5273
rect 3422 5199 3478 5208
rect 3252 4678 3372 4706
rect 3240 4616 3292 4622
rect 3238 4584 3240 4593
rect 3292 4584 3294 4593
rect 3238 4519 3294 4528
rect 3252 4049 3280 4519
rect 3238 4040 3294 4049
rect 3238 3975 3294 3984
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3738 3280 3878
rect 3240 3732 3292 3738
rect 3240 3674 3292 3680
rect 3148 3664 3200 3670
rect 3148 3606 3200 3612
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 3148 2916 3200 2922
rect 3148 2858 3200 2864
rect 2700 2808 2820 2836
rect 2700 2530 2728 2808
rect 2824 2748 3132 2768
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2672 3132 2692
rect 2700 2502 2820 2530
rect 2608 1720 2728 1748
rect 2700 800 2728 1720
rect 2792 1465 2820 2502
rect 3056 2304 3108 2310
rect 3056 2246 3108 2252
rect 3068 2038 3096 2246
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 2778 1456 2834 1465
rect 3160 1442 3188 2858
rect 3252 2446 3280 2926
rect 3240 2440 3292 2446
rect 3240 2382 3292 2388
rect 3344 2378 3372 4678
rect 3436 2417 3464 5199
rect 3528 4486 3556 5471
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3516 4276 3568 4282
rect 3516 4218 3568 4224
rect 3528 4146 3556 4218
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3620 4026 3648 6054
rect 3528 3998 3648 4026
rect 3528 3126 3556 3998
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3620 3602 3648 3878
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 3608 3392 3660 3398
rect 3712 3369 3740 7278
rect 3804 6322 3832 9114
rect 3884 9104 3936 9110
rect 3884 9046 3936 9052
rect 3896 8945 3924 9046
rect 3882 8936 3938 8945
rect 3882 8871 3938 8880
rect 3896 8498 3924 8871
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 3988 8378 4016 9114
rect 3896 8350 4016 8378
rect 3896 6798 3924 8350
rect 4080 7585 4108 10202
rect 4172 10062 4200 12406
rect 4252 11756 4304 11762
rect 4252 11698 4304 11704
rect 4264 11354 4292 11698
rect 4344 11552 4396 11558
rect 4344 11494 4396 11500
rect 4252 11348 4304 11354
rect 4252 11290 4304 11296
rect 4356 11234 4384 11494
rect 4264 11206 4384 11234
rect 4264 10130 4292 11206
rect 4436 11076 4488 11082
rect 4436 11018 4488 11024
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 4252 10124 4304 10130
rect 4252 10066 4304 10072
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 4172 9722 4200 9998
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4160 9580 4212 9586
rect 4160 9522 4212 9528
rect 4172 9178 4200 9522
rect 4252 9444 4304 9450
rect 4252 9386 4304 9392
rect 4160 9172 4212 9178
rect 4160 9114 4212 9120
rect 4158 9072 4214 9081
rect 4158 9007 4214 9016
rect 4172 8838 4200 9007
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 4158 8664 4214 8673
rect 4158 8599 4160 8608
rect 4212 8599 4214 8608
rect 4160 8570 4212 8576
rect 4264 8566 4292 9386
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4252 8288 4304 8294
rect 4252 8230 4304 8236
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4172 7886 4200 7958
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4066 7576 4122 7585
rect 4066 7511 4122 7520
rect 3976 7472 4028 7478
rect 3976 7414 4028 7420
rect 4066 7440 4122 7449
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3988 6644 4016 7414
rect 4066 7375 4122 7384
rect 4080 6746 4108 7375
rect 4172 6934 4200 7822
rect 4264 7818 4292 8230
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4264 6866 4292 7754
rect 4356 7478 4384 10678
rect 4448 10538 4476 11018
rect 4436 10532 4488 10538
rect 4436 10474 4488 10480
rect 4540 10130 4568 13942
rect 4632 13870 4660 14826
rect 4710 14376 4766 14385
rect 4710 14311 4712 14320
rect 4764 14311 4766 14320
rect 4712 14282 4764 14288
rect 4698 14172 5006 14192
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14096 5006 14116
rect 4620 13864 4672 13870
rect 4620 13806 4672 13812
rect 4632 12986 4660 13806
rect 4698 13084 5006 13104
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13008 5006 13028
rect 5092 12986 5120 16068
rect 5184 15026 5212 16526
rect 5540 16244 5592 16250
rect 5540 16186 5592 16192
rect 5552 16153 5580 16186
rect 5538 16144 5594 16153
rect 5356 16108 5408 16114
rect 5538 16079 5594 16088
rect 5356 16050 5408 16056
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5184 14074 5212 14758
rect 5172 14068 5224 14074
rect 5172 14010 5224 14016
rect 5172 13524 5224 13530
rect 5172 13466 5224 13472
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 5080 12980 5132 12986
rect 5080 12922 5132 12928
rect 4986 12744 5042 12753
rect 4986 12679 5042 12688
rect 5000 12170 5028 12679
rect 5092 12442 5120 12922
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5078 12336 5134 12345
rect 5184 12306 5212 13466
rect 5276 12918 5304 15642
rect 5368 15201 5396 16050
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5552 15745 5580 15982
rect 5538 15736 5594 15745
rect 5538 15671 5594 15680
rect 5448 15360 5500 15366
rect 5448 15302 5500 15308
rect 5354 15192 5410 15201
rect 5354 15127 5410 15136
rect 5460 15026 5488 15302
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5368 14346 5396 14962
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5368 13954 5396 14282
rect 5460 14074 5488 14962
rect 5552 14521 5580 15671
rect 5644 14550 5672 17070
rect 5736 15910 5764 17224
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5724 15904 5776 15910
rect 5724 15846 5776 15852
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 15094 5764 15438
rect 5828 15162 5856 16730
rect 5920 16250 5948 17138
rect 6012 16726 6040 17138
rect 6000 16720 6052 16726
rect 6000 16662 6052 16668
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 6000 15904 6052 15910
rect 6000 15846 6052 15852
rect 5816 15156 5868 15162
rect 5816 15098 5868 15104
rect 5724 15088 5776 15094
rect 5724 15030 5776 15036
rect 5632 14544 5684 14550
rect 5538 14512 5594 14521
rect 5632 14486 5684 14492
rect 5538 14447 5594 14456
rect 5736 14414 5764 15030
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5814 14376 5870 14385
rect 5632 14272 5684 14278
rect 5632 14214 5684 14220
rect 5448 14068 5500 14074
rect 5448 14010 5500 14016
rect 5538 13968 5594 13977
rect 5368 13926 5488 13954
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5368 12986 5396 13194
rect 5356 12980 5408 12986
rect 5356 12922 5408 12928
rect 5264 12912 5316 12918
rect 5264 12854 5316 12860
rect 5264 12436 5316 12442
rect 5460 12434 5488 13926
rect 5538 13903 5594 13912
rect 5552 13682 5580 13903
rect 5644 13802 5672 14214
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5552 13654 5672 13682
rect 5264 12378 5316 12384
rect 5368 12406 5488 12434
rect 5078 12271 5134 12280
rect 5172 12300 5224 12306
rect 4988 12164 5040 12170
rect 4988 12106 5040 12112
rect 5092 12102 5120 12271
rect 5172 12242 5224 12248
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 5080 12096 5132 12102
rect 5080 12038 5132 12044
rect 4528 10124 4580 10130
rect 4528 10066 4580 10072
rect 4540 9994 4568 10066
rect 4528 9988 4580 9994
rect 4528 9930 4580 9936
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9674 4476 9862
rect 4632 9704 4660 12038
rect 4698 11996 5006 12016
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11920 5006 11940
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 4896 11688 4948 11694
rect 4896 11630 4948 11636
rect 4908 11082 4936 11630
rect 5000 11558 5028 11698
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4698 10908 5006 10928
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10832 5006 10852
rect 4698 9820 5006 9840
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9744 5006 9764
rect 4632 9676 4844 9704
rect 4448 9646 4568 9674
rect 4540 9586 4568 9646
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4436 9376 4488 9382
rect 4436 9318 4488 9324
rect 4620 9376 4672 9382
rect 4620 9318 4672 9324
rect 4448 8906 4476 9318
rect 4632 9042 4660 9318
rect 4620 9036 4672 9042
rect 4620 8978 4672 8984
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4724 8945 4752 8978
rect 4710 8936 4766 8945
rect 4436 8900 4488 8906
rect 4710 8871 4766 8880
rect 4436 8842 4488 8848
rect 4528 8832 4580 8838
rect 4434 8800 4490 8809
rect 4816 8820 4844 9676
rect 4988 9580 5040 9586
rect 4988 9522 5040 9528
rect 5000 9353 5028 9522
rect 4986 9344 5042 9353
rect 4986 9279 5042 9288
rect 4528 8774 4580 8780
rect 4632 8792 4844 8820
rect 4434 8735 4490 8744
rect 4448 8401 4476 8735
rect 4434 8392 4490 8401
rect 4434 8327 4490 8336
rect 4344 7472 4396 7478
rect 4344 7414 4396 7420
rect 4252 6860 4304 6866
rect 4252 6802 4304 6808
rect 4080 6718 4292 6746
rect 3988 6616 4108 6644
rect 3792 6316 3844 6322
rect 3844 6276 3924 6304
rect 3792 6258 3844 6264
rect 3792 6112 3844 6118
rect 3792 6054 3844 6060
rect 3804 5710 3832 6054
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3792 5296 3844 5302
rect 3792 5238 3844 5244
rect 3804 4690 3832 5238
rect 3896 5234 3924 6276
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5574 4016 6122
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3804 4214 3832 4626
rect 3988 4570 4016 5170
rect 3896 4542 4016 4570
rect 3792 4208 3844 4214
rect 3792 4150 3844 4156
rect 3896 3482 3924 4542
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3804 3454 3924 3482
rect 3608 3334 3660 3340
rect 3698 3360 3754 3369
rect 3516 3120 3568 3126
rect 3516 3062 3568 3068
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3528 2825 3556 2858
rect 3514 2816 3570 2825
rect 3514 2751 3570 2760
rect 3516 2644 3568 2650
rect 3516 2586 3568 2592
rect 3422 2408 3478 2417
rect 3332 2372 3384 2378
rect 3422 2343 3478 2352
rect 3332 2314 3384 2320
rect 2778 1391 2834 1400
rect 3068 1414 3188 1442
rect 3068 800 3096 1414
rect 3528 800 3556 2586
rect 3620 2530 3648 3334
rect 3698 3295 3754 3304
rect 3804 2990 3832 3454
rect 3884 3392 3936 3398
rect 3884 3334 3936 3340
rect 3792 2984 3844 2990
rect 3896 2961 3924 3334
rect 3792 2926 3844 2932
rect 3882 2952 3938 2961
rect 3882 2887 3938 2896
rect 3988 2774 4016 4422
rect 4080 3058 4108 6616
rect 4160 5908 4212 5914
rect 4160 5850 4212 5856
rect 4172 5234 4200 5850
rect 4160 5228 4212 5234
rect 4160 5170 4212 5176
rect 4264 5098 4292 6718
rect 4356 5234 4384 7414
rect 4448 6882 4476 8327
rect 4540 8090 4568 8774
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4632 7342 4660 8792
rect 4698 8732 5006 8752
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8656 5006 8676
rect 4698 7644 5006 7664
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7568 5006 7588
rect 5092 7478 5120 12038
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5184 11665 5212 11834
rect 5170 11656 5226 11665
rect 5170 11591 5226 11600
rect 5276 11558 5304 12378
rect 5264 11552 5316 11558
rect 5264 11494 5316 11500
rect 5368 11506 5396 12406
rect 5540 12232 5592 12238
rect 5538 12200 5540 12209
rect 5592 12200 5594 12209
rect 5538 12135 5594 12144
rect 5448 12096 5500 12102
rect 5448 12038 5500 12044
rect 5460 11626 5488 12038
rect 5644 11762 5672 13654
rect 5736 13530 5764 14350
rect 5814 14311 5870 14320
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5828 13462 5856 14311
rect 5908 13932 5960 13938
rect 5908 13874 5960 13880
rect 5816 13456 5868 13462
rect 5816 13398 5868 13404
rect 5828 12434 5856 13398
rect 5736 12406 5856 12434
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5368 11478 5488 11506
rect 5460 10470 5488 11478
rect 5736 11336 5764 12406
rect 5816 12232 5868 12238
rect 5816 12174 5868 12180
rect 5644 11308 5764 11336
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5448 10464 5500 10470
rect 5448 10406 5500 10412
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 8294 5212 9862
rect 5276 9722 5304 10066
rect 5460 9994 5488 10406
rect 5552 10266 5580 10610
rect 5540 10260 5592 10266
rect 5540 10202 5592 10208
rect 5448 9988 5500 9994
rect 5448 9930 5500 9936
rect 5540 9920 5592 9926
rect 5540 9862 5592 9868
rect 5264 9716 5316 9722
rect 5264 9658 5316 9664
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5356 9512 5408 9518
rect 5276 9472 5356 9500
rect 5172 8288 5224 8294
rect 5172 8230 5224 8236
rect 5276 7954 5304 9472
rect 5356 9454 5408 9460
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5368 8634 5396 8842
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5264 7948 5316 7954
rect 5264 7890 5316 7896
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 5080 7472 5132 7478
rect 5080 7414 5132 7420
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4620 7336 4672 7342
rect 4620 7278 4672 7284
rect 4620 7200 4672 7206
rect 4620 7142 4672 7148
rect 4448 6854 4568 6882
rect 4632 6866 4660 7142
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4448 5234 4476 6666
rect 4540 6254 4568 6854
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4816 6644 4844 7346
rect 5080 7336 5132 7342
rect 5080 7278 5132 7284
rect 5092 6712 5120 7278
rect 5184 7274 5212 7754
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5172 7268 5224 7274
rect 5172 7210 5224 7216
rect 5184 7002 5212 7210
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5092 6684 5212 6712
rect 4816 6616 5120 6644
rect 4698 6556 5006 6576
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6480 5006 6500
rect 5092 6458 5120 6616
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4528 6248 4580 6254
rect 4528 6190 4580 6196
rect 4986 6216 5042 6225
rect 4986 6151 4988 6160
rect 5040 6151 5042 6160
rect 4988 6122 5040 6128
rect 5080 5636 5132 5642
rect 5080 5578 5132 5584
rect 4698 5468 5006 5488
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5392 5006 5412
rect 4344 5228 4396 5234
rect 4344 5170 4396 5176
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4528 5160 4580 5166
rect 4528 5102 4580 5108
rect 4252 5092 4304 5098
rect 4252 5034 4304 5040
rect 4160 5024 4212 5030
rect 4160 4966 4212 4972
rect 4172 3126 4200 4966
rect 4344 4548 4396 4554
rect 4344 4490 4396 4496
rect 4356 4146 4384 4490
rect 4436 4276 4488 4282
rect 4436 4218 4488 4224
rect 4344 4140 4396 4146
rect 4344 4082 4396 4088
rect 4448 3602 4476 4218
rect 4540 4214 4568 5102
rect 5092 4758 5120 5578
rect 5080 4752 5132 4758
rect 5080 4694 5132 4700
rect 5078 4584 5134 4593
rect 5184 4554 5212 6684
rect 5276 4622 5304 7686
rect 5460 7546 5488 9590
rect 5552 9586 5580 9862
rect 5644 9674 5672 11308
rect 5724 11212 5776 11218
rect 5828 11200 5856 12174
rect 5920 11830 5948 13874
rect 6012 13025 6040 15846
rect 6104 15162 6132 16390
rect 6196 16114 6224 16594
rect 6184 16108 6236 16114
rect 6184 16050 6236 16056
rect 6196 15706 6224 16050
rect 6288 15978 6316 19200
rect 6460 17672 6512 17678
rect 6460 17614 6512 17620
rect 6472 16998 6500 17614
rect 6748 17610 6776 19200
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 7116 17270 7144 19200
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7104 17264 7156 17270
rect 7104 17206 7156 17212
rect 7196 17196 7248 17202
rect 7196 17138 7248 17144
rect 6828 17060 6880 17066
rect 6880 17020 7052 17048
rect 6828 17002 6880 17008
rect 6460 16992 6512 16998
rect 6460 16934 6512 16940
rect 6572 16892 6880 16912
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16816 6880 16836
rect 6920 16720 6972 16726
rect 6920 16662 6972 16668
rect 6368 16584 6420 16590
rect 6368 16526 6420 16532
rect 6380 16250 6408 16526
rect 6460 16448 6512 16454
rect 6460 16390 6512 16396
rect 6368 16244 6420 16250
rect 6368 16186 6420 16192
rect 6276 15972 6328 15978
rect 6276 15914 6328 15920
rect 6184 15700 6236 15706
rect 6184 15642 6236 15648
rect 6092 15156 6144 15162
rect 6092 15098 6144 15104
rect 6380 14958 6408 16186
rect 6472 15162 6500 16390
rect 6572 15804 6880 15824
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15728 6880 15748
rect 6734 15464 6790 15473
rect 6734 15399 6790 15408
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6748 15026 6776 15399
rect 6932 15162 6960 16662
rect 7024 16250 7052 17020
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16794 7144 16934
rect 7104 16788 7156 16794
rect 7104 16730 7156 16736
rect 7012 16244 7064 16250
rect 7012 16186 7064 16192
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 6920 15156 6972 15162
rect 6920 15098 6972 15104
rect 6736 15020 6788 15026
rect 6736 14962 6788 14968
rect 7024 14958 7052 15574
rect 7104 15496 7156 15502
rect 7104 15438 7156 15444
rect 7116 15026 7144 15438
rect 7208 15144 7236 17138
rect 7300 15502 7328 17546
rect 7576 17270 7604 19200
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7380 17196 7432 17202
rect 7380 17138 7432 17144
rect 7392 15706 7420 17138
rect 7472 17128 7524 17134
rect 7472 17070 7524 17076
rect 7484 16114 7512 17070
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 7760 16114 7788 16526
rect 7840 16516 7892 16522
rect 7840 16458 7892 16464
rect 7852 16250 7880 16458
rect 7944 16250 7972 19200
rect 8404 17678 8432 19200
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8772 17524 8800 19200
rect 9036 17536 9088 17542
rect 8772 17496 8892 17524
rect 8446 17436 8754 17456
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17360 8754 17380
rect 8864 17338 8892 17496
rect 9036 17478 9088 17484
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 8024 16992 8076 16998
rect 8024 16934 8076 16940
rect 8036 16454 8064 16934
rect 8128 16658 8156 17070
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7932 16244 7984 16250
rect 7932 16186 7984 16192
rect 7472 16108 7524 16114
rect 7472 16050 7524 16056
rect 7748 16108 7800 16114
rect 7748 16050 7800 16056
rect 7380 15700 7432 15706
rect 7380 15642 7432 15648
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 7564 15496 7616 15502
rect 7564 15438 7616 15444
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7288 15156 7340 15162
rect 7208 15116 7288 15144
rect 7288 15098 7340 15104
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 7012 14952 7064 14958
rect 7012 14894 7064 14900
rect 6572 14716 6880 14736
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14640 6880 14660
rect 6092 14544 6144 14550
rect 6092 14486 6144 14492
rect 5998 13016 6054 13025
rect 5998 12951 6054 12960
rect 6104 12900 6132 14486
rect 6460 14340 6512 14346
rect 6460 14282 6512 14288
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6184 13796 6236 13802
rect 6184 13738 6236 13744
rect 6196 12918 6224 13738
rect 6368 13728 6420 13734
rect 6368 13670 6420 13676
rect 6380 13394 6408 13670
rect 6368 13388 6420 13394
rect 6368 13330 6420 13336
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6012 12872 6132 12900
rect 6184 12912 6236 12918
rect 6012 11898 6040 12872
rect 6184 12854 6236 12860
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6104 12170 6132 12582
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6000 11892 6052 11898
rect 6000 11834 6052 11840
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 5998 11792 6054 11801
rect 5998 11727 6000 11736
rect 6052 11727 6054 11736
rect 6000 11698 6052 11704
rect 5776 11172 5856 11200
rect 5724 11154 5776 11160
rect 5724 11008 5776 11014
rect 5724 10950 5776 10956
rect 5736 10033 5764 10950
rect 5828 10674 5856 11172
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 6012 10606 6040 11698
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 5722 10024 5778 10033
rect 5722 9959 5778 9968
rect 5644 9646 5764 9674
rect 5540 9580 5592 9586
rect 5540 9522 5592 9528
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5552 8566 5580 8910
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 5644 7886 5672 9454
rect 5736 9081 5764 9646
rect 6196 9625 6224 12854
rect 6288 12084 6316 13262
rect 6472 12850 6500 14282
rect 6840 13870 6868 14282
rect 6932 14006 6960 14894
rect 7012 14272 7064 14278
rect 7012 14214 7064 14220
rect 6920 14000 6972 14006
rect 6920 13942 6972 13948
rect 6828 13864 6880 13870
rect 6828 13806 6880 13812
rect 6572 13628 6880 13648
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13552 6880 13572
rect 6932 13308 6960 13942
rect 7024 13870 7052 14214
rect 7012 13864 7064 13870
rect 7064 13824 7144 13852
rect 7012 13806 7064 13812
rect 6734 13288 6790 13297
rect 6734 13223 6790 13232
rect 6840 13280 6960 13308
rect 6748 12986 6776 13223
rect 6840 13190 6868 13280
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 6828 13184 6880 13190
rect 6828 13126 6880 13132
rect 6920 13184 6972 13190
rect 6920 13126 6972 13132
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6460 12844 6512 12850
rect 6460 12786 6512 12792
rect 6828 12776 6880 12782
rect 6932 12764 6960 13126
rect 6880 12736 6960 12764
rect 6828 12718 6880 12724
rect 6460 12640 6512 12646
rect 6460 12582 6512 12588
rect 6368 12096 6420 12102
rect 6288 12056 6368 12084
rect 6368 12038 6420 12044
rect 6472 11898 6500 12582
rect 6572 12540 6880 12560
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12464 6880 12484
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6460 11892 6512 11898
rect 6460 11834 6512 11840
rect 6460 11756 6512 11762
rect 6460 11698 6512 11704
rect 6472 11354 6500 11698
rect 6840 11694 6868 12038
rect 6828 11688 6880 11694
rect 6828 11630 6880 11636
rect 6572 11452 6880 11472
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11376 6880 11396
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 11082 6500 11290
rect 6920 11144 6972 11150
rect 6920 11086 6972 11092
rect 6460 11076 6512 11082
rect 6460 11018 6512 11024
rect 6736 11008 6788 11014
rect 6736 10950 6788 10956
rect 6748 10810 6776 10950
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6932 10674 6960 11086
rect 7024 10674 7052 13194
rect 7116 12782 7144 13824
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 7104 11076 7156 11082
rect 7104 11018 7156 11024
rect 6920 10668 6972 10674
rect 6920 10610 6972 10616
rect 7012 10668 7064 10674
rect 7012 10610 7064 10616
rect 6572 10364 6880 10384
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10288 6880 10308
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6182 9616 6238 9625
rect 6182 9551 6238 9560
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5722 9072 5778 9081
rect 5722 9007 5778 9016
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5736 8090 5764 8570
rect 5724 8084 5776 8090
rect 5724 8026 5776 8032
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5356 7540 5408 7546
rect 5356 7482 5408 7488
rect 5448 7540 5500 7546
rect 5448 7482 5500 7488
rect 5368 6322 5396 7482
rect 5540 7472 5592 7478
rect 5540 7414 5592 7420
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5460 6866 5488 7142
rect 5448 6860 5500 6866
rect 5448 6802 5500 6808
rect 5552 6662 5580 7414
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5644 6662 5672 7346
rect 5816 6996 5868 7002
rect 5816 6938 5868 6944
rect 5828 6866 5856 6938
rect 5816 6860 5868 6866
rect 5816 6802 5868 6808
rect 5920 6798 5948 9114
rect 6274 9072 6330 9081
rect 6472 9042 6500 9998
rect 6932 9738 6960 10610
rect 6840 9710 6960 9738
rect 6840 9586 6868 9710
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 7116 9450 7144 11018
rect 7208 9926 7236 14962
rect 7288 14884 7340 14890
rect 7288 14826 7340 14832
rect 7300 13530 7328 14826
rect 7392 14074 7420 15302
rect 7470 15192 7526 15201
rect 7470 15127 7526 15136
rect 7380 14068 7432 14074
rect 7380 14010 7432 14016
rect 7484 13530 7512 15127
rect 7576 13938 7604 15438
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7668 14618 7696 14894
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7760 14414 7788 16050
rect 8036 14929 8064 16390
rect 8128 15910 8156 16594
rect 8116 15904 8168 15910
rect 8116 15846 8168 15852
rect 8116 15428 8168 15434
rect 8116 15370 8168 15376
rect 8022 14920 8078 14929
rect 8022 14855 8078 14864
rect 8128 14414 8156 15370
rect 8220 14958 8248 17002
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8852 16788 8904 16794
rect 8852 16730 8904 16736
rect 8300 16584 8352 16590
rect 8300 16526 8352 16532
rect 8312 16114 8340 16526
rect 8446 16348 8754 16368
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16272 8754 16292
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8208 14952 8260 14958
rect 8208 14894 8260 14900
rect 7748 14408 7800 14414
rect 7748 14350 7800 14356
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7472 13524 7524 13530
rect 7472 13466 7524 13472
rect 7484 12986 7512 13466
rect 7472 12980 7524 12986
rect 7472 12922 7524 12928
rect 7380 11620 7432 11626
rect 7380 11562 7432 11568
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 6920 9444 6972 9450
rect 6920 9386 6972 9392
rect 7104 9444 7156 9450
rect 7104 9386 7156 9392
rect 6932 9330 6960 9386
rect 6932 9302 7144 9330
rect 6572 9276 6880 9296
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9200 6880 9220
rect 6274 9007 6330 9016
rect 6460 9036 6512 9042
rect 6092 8832 6144 8838
rect 6092 8774 6144 8780
rect 6104 8566 6132 8774
rect 6092 8560 6144 8566
rect 6092 8502 6144 8508
rect 6288 8498 6316 9007
rect 6460 8978 6512 8984
rect 6276 8492 6328 8498
rect 6196 8452 6276 8480
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 7410 6040 8230
rect 6196 7886 6224 8452
rect 6276 8434 6328 8440
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6380 7954 6408 8298
rect 6472 8022 6500 8978
rect 6918 8936 6974 8945
rect 6918 8871 6974 8880
rect 6572 8188 6880 8208
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8112 6880 8132
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6184 7880 6236 7886
rect 6184 7822 6236 7828
rect 6000 7404 6052 7410
rect 6052 7364 6132 7392
rect 6000 7346 6052 7352
rect 6104 7313 6132 7364
rect 6090 7304 6146 7313
rect 6000 7268 6052 7274
rect 6090 7239 6146 7248
rect 6000 7210 6052 7216
rect 6012 6866 6040 7210
rect 6000 6860 6052 6866
rect 6000 6802 6052 6808
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5540 6656 5592 6662
rect 5632 6656 5684 6662
rect 5540 6598 5592 6604
rect 5630 6624 5632 6633
rect 5684 6624 5686 6633
rect 5630 6559 5686 6568
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5920 5914 5948 6734
rect 6196 6338 6224 7822
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6196 6310 6316 6338
rect 6000 6248 6052 6254
rect 6184 6248 6236 6254
rect 6000 6190 6052 6196
rect 6182 6216 6184 6225
rect 6236 6216 6238 6225
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 5354 5808 5410 5817
rect 5354 5743 5410 5752
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5078 4519 5134 4528
rect 5172 4548 5224 4554
rect 4698 4380 5006 4400
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4304 5006 4324
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4528 4208 4580 4214
rect 4528 4150 4580 4156
rect 4436 3596 4488 3602
rect 4488 3556 4568 3584
rect 4436 3538 4488 3544
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4250 3224 4306 3233
rect 4250 3159 4306 3168
rect 4160 3120 4212 3126
rect 4160 3062 4212 3068
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4264 2922 4292 3159
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 3988 2746 4108 2774
rect 4080 2666 4108 2746
rect 4080 2638 4200 2666
rect 4356 2650 4384 3334
rect 4448 3194 4476 3334
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4540 2689 4568 3556
rect 4526 2680 4582 2689
rect 3976 2576 4028 2582
rect 3620 2502 3740 2530
rect 3976 2518 4028 2524
rect 4066 2544 4122 2553
rect 3608 2440 3660 2446
rect 3608 2382 3660 2388
rect 3620 1970 3648 2382
rect 3608 1964 3660 1970
rect 3608 1906 3660 1912
rect 3712 1834 3740 2502
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3700 1828 3752 1834
rect 3700 1770 3752 1776
rect 3896 1630 3924 2246
rect 3884 1624 3936 1630
rect 3884 1566 3936 1572
rect 3988 800 4016 2518
rect 4066 2479 4122 2488
rect 4080 2446 4108 2479
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4172 2310 4200 2638
rect 4344 2644 4396 2650
rect 4526 2615 4582 2624
rect 4344 2586 4396 2592
rect 4632 2530 4660 4218
rect 4698 3292 5006 3312
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3216 5006 3236
rect 5092 3126 5120 4519
rect 5172 4490 5224 4496
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5276 3602 5304 4082
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5172 3392 5224 3398
rect 5172 3334 5224 3340
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5184 3194 5212 3334
rect 5172 3188 5224 3194
rect 5172 3130 5224 3136
rect 5080 3120 5132 3126
rect 5276 3097 5304 3334
rect 5080 3062 5132 3068
rect 5262 3088 5318 3097
rect 5262 3023 5318 3032
rect 4988 2916 5040 2922
rect 5172 2916 5224 2922
rect 5040 2876 5172 2904
rect 4988 2858 5040 2864
rect 5172 2858 5224 2864
rect 4344 2508 4396 2514
rect 4344 2450 4396 2456
rect 4540 2502 4660 2530
rect 5184 2514 5212 2858
rect 5264 2848 5316 2854
rect 5264 2790 5316 2796
rect 5172 2508 5224 2514
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4356 800 4384 2450
rect 4540 1902 4568 2502
rect 5172 2450 5224 2456
rect 5276 2446 5304 2790
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5368 2378 5396 5743
rect 5632 5704 5684 5710
rect 5632 5646 5684 5652
rect 5644 5302 5672 5646
rect 5920 5522 5948 5850
rect 6012 5846 6040 6190
rect 6182 6151 6238 6160
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 6196 5778 6224 6054
rect 6288 5817 6316 6310
rect 6274 5808 6330 5817
rect 6184 5772 6236 5778
rect 6274 5743 6330 5752
rect 6184 5714 6236 5720
rect 5736 5494 5948 5522
rect 6000 5568 6052 5574
rect 6000 5510 6052 5516
rect 5632 5296 5684 5302
rect 5632 5238 5684 5244
rect 5644 4758 5672 5238
rect 5632 4752 5684 4758
rect 5632 4694 5684 4700
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 5460 3670 5488 4422
rect 5644 4282 5672 4422
rect 5632 4276 5684 4282
rect 5632 4218 5684 4224
rect 5632 3936 5684 3942
rect 5632 3878 5684 3884
rect 5448 3664 5500 3670
rect 5448 3606 5500 3612
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 2990 5488 3402
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5552 3194 5580 3334
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5448 2984 5500 2990
rect 5448 2926 5500 2932
rect 5540 2576 5592 2582
rect 5540 2518 5592 2524
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 5356 2372 5408 2378
rect 5356 2314 5408 2320
rect 4528 1896 4580 1902
rect 4528 1838 4580 1844
rect 4632 1170 4660 2314
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 4698 2204 5006 2224
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2128 5006 2148
rect 5460 2106 5488 2246
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 5448 2100 5500 2106
rect 5448 2042 5500 2048
rect 4632 1142 4844 1170
rect 4816 800 4844 1142
rect 5184 800 5212 2042
rect 5552 1766 5580 2518
rect 5540 1760 5592 1766
rect 5540 1702 5592 1708
rect 5644 800 5672 3878
rect 5736 3534 5764 5494
rect 5816 5364 5868 5370
rect 5816 5306 5868 5312
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5724 3392 5776 3398
rect 5724 3334 5776 3340
rect 5736 3194 5764 3334
rect 5724 3188 5776 3194
rect 5724 3130 5776 3136
rect 5724 2984 5776 2990
rect 5724 2926 5776 2932
rect 5736 2689 5764 2926
rect 5722 2680 5778 2689
rect 5722 2615 5778 2624
rect 5828 2446 5856 5306
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5920 4146 5948 4626
rect 6012 4622 6040 5510
rect 6196 5234 6224 5714
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6288 5030 6316 5578
rect 6380 5234 6408 7686
rect 6460 7404 6512 7410
rect 6460 7346 6512 7352
rect 6472 7002 6500 7346
rect 6932 7342 6960 8871
rect 7116 8430 7144 9302
rect 7196 8900 7248 8906
rect 7196 8842 7248 8848
rect 7104 8424 7156 8430
rect 7104 8366 7156 8372
rect 6920 7336 6972 7342
rect 6920 7278 6972 7284
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6572 7100 6880 7120
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7024 6880 7044
rect 6460 6996 6512 7002
rect 6460 6938 6512 6944
rect 6572 6012 6880 6032
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5936 6880 5956
rect 6460 5840 6512 5846
rect 6460 5782 6512 5788
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6368 5092 6420 5098
rect 6368 5034 6420 5040
rect 6092 5024 6144 5030
rect 6092 4966 6144 4972
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6000 4616 6052 4622
rect 6000 4558 6052 4564
rect 5908 4140 5960 4146
rect 5908 4082 5960 4088
rect 6104 3942 6132 4966
rect 6288 4078 6316 4966
rect 6380 4282 6408 5034
rect 6368 4276 6420 4282
rect 6368 4218 6420 4224
rect 6472 4214 6500 5782
rect 6572 4924 6880 4944
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4848 6880 4868
rect 6460 4208 6512 4214
rect 6460 4150 6512 4156
rect 6276 4072 6328 4078
rect 6276 4014 6328 4020
rect 6092 3936 6144 3942
rect 6092 3878 6144 3884
rect 6572 3836 6880 3856
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3760 6880 3780
rect 6182 3632 6238 3641
rect 6182 3567 6238 3576
rect 6368 3596 6420 3602
rect 6196 3058 6224 3567
rect 6368 3538 6420 3544
rect 6184 3052 6236 3058
rect 6184 2994 6236 3000
rect 6196 2825 6224 2994
rect 6380 2922 6408 3538
rect 6460 3188 6512 3194
rect 6460 3130 6512 3136
rect 6368 2916 6420 2922
rect 6368 2858 6420 2864
rect 6182 2816 6238 2825
rect 6182 2751 6238 2760
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6368 2304 6420 2310
rect 6368 2246 6420 2252
rect 6000 2032 6052 2038
rect 6000 1974 6052 1980
rect 6012 800 6040 1974
rect 6380 1834 6408 2246
rect 6368 1828 6420 1834
rect 6368 1770 6420 1776
rect 6472 800 6500 3130
rect 6572 2748 6880 2768
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2672 6880 2692
rect 6932 2553 6960 7142
rect 7012 6656 7064 6662
rect 7012 6598 7064 6604
rect 7024 5710 7052 6598
rect 7012 5704 7064 5710
rect 7012 5646 7064 5652
rect 7116 5098 7144 8366
rect 7208 7886 7236 8842
rect 7288 8832 7340 8838
rect 7288 8774 7340 8780
rect 7300 8430 7328 8774
rect 7288 8424 7340 8430
rect 7288 8366 7340 8372
rect 7392 8294 7420 11562
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7484 10198 7512 11086
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7668 9738 7696 14010
rect 7760 13938 7788 14350
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 7748 13932 7800 13938
rect 7748 13874 7800 13880
rect 8024 13932 8076 13938
rect 8024 13874 8076 13880
rect 8036 13734 8064 13874
rect 8024 13728 8076 13734
rect 8024 13670 8076 13676
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7840 12776 7892 12782
rect 7840 12718 7892 12724
rect 7746 12200 7802 12209
rect 7746 12135 7802 12144
rect 7760 11898 7788 12135
rect 7748 11892 7800 11898
rect 7748 11834 7800 11840
rect 7852 11694 7880 12718
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7748 11212 7800 11218
rect 7748 11154 7800 11160
rect 7760 10810 7788 11154
rect 7932 11008 7984 11014
rect 7932 10950 7984 10956
rect 7748 10804 7800 10810
rect 7748 10746 7800 10752
rect 7484 9710 7696 9738
rect 7484 8430 7512 9710
rect 7944 9654 7972 10950
rect 8036 9674 8064 13126
rect 8128 12986 8156 14214
rect 8312 13938 8340 16050
rect 8446 15260 8754 15280
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15184 8754 15204
rect 8760 15020 8812 15026
rect 8760 14962 8812 14968
rect 8772 14346 8800 14962
rect 8864 14958 8892 16730
rect 8956 16182 8984 16934
rect 8944 16176 8996 16182
rect 8944 16118 8996 16124
rect 9048 15434 9076 17478
rect 9140 16250 9168 19200
rect 9600 17954 9628 19200
rect 9600 17926 9720 17954
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9588 17196 9640 17202
rect 9588 17138 9640 17144
rect 9220 17060 9272 17066
rect 9220 17002 9272 17008
rect 9232 16522 9260 17002
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9128 16244 9180 16250
rect 9128 16186 9180 16192
rect 9140 15502 9168 16186
rect 9232 16182 9260 16458
rect 9220 16176 9272 16182
rect 9220 16118 9272 16124
rect 9128 15496 9180 15502
rect 9128 15438 9180 15444
rect 9036 15428 9088 15434
rect 9036 15370 9088 15376
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 15026 8984 15302
rect 9048 15094 9076 15370
rect 9036 15088 9088 15094
rect 9036 15030 9088 15036
rect 8944 15020 8996 15026
rect 8944 14962 8996 14968
rect 8852 14952 8904 14958
rect 8852 14894 8904 14900
rect 8852 14816 8904 14822
rect 8852 14758 8904 14764
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8864 14278 8892 14758
rect 8852 14272 8904 14278
rect 8852 14214 8904 14220
rect 8446 14172 8754 14192
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14096 8754 14116
rect 8864 14056 8892 14214
rect 8680 14028 8892 14056
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8680 13258 8708 14028
rect 8760 13932 8812 13938
rect 8760 13874 8812 13880
rect 8772 13705 8800 13874
rect 8758 13696 8814 13705
rect 8758 13631 8814 13640
rect 8772 13394 8800 13631
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8760 13388 8812 13394
rect 8760 13330 8812 13336
rect 8668 13252 8720 13258
rect 8668 13194 8720 13200
rect 8446 13084 8754 13104
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13008 8754 13028
rect 8116 12980 8168 12986
rect 8116 12922 8168 12928
rect 8116 12844 8168 12850
rect 8116 12786 8168 12792
rect 8128 11218 8156 12786
rect 8300 12436 8352 12442
rect 8300 12378 8352 12384
rect 8312 11762 8340 12378
rect 8864 12102 8892 13466
rect 8956 12753 8984 14962
rect 9048 13002 9076 15030
rect 9324 14822 9352 17138
rect 9600 16794 9628 17138
rect 9692 17105 9720 17926
rect 9678 17096 9734 17105
rect 9678 17031 9734 17040
rect 9588 16788 9640 16794
rect 9588 16730 9640 16736
rect 9588 16516 9640 16522
rect 9588 16458 9640 16464
rect 9600 15910 9628 16458
rect 9968 16454 9996 19200
rect 10428 19122 10456 19200
rect 10520 19122 10548 19230
rect 10428 19094 10548 19122
rect 10048 17196 10100 17202
rect 10704 17184 10732 19230
rect 10782 19200 10838 20000
rect 11242 19200 11298 20000
rect 11610 19200 11666 20000
rect 12070 19200 12126 20000
rect 12438 19200 12494 20000
rect 12898 19200 12954 20000
rect 13266 19200 13322 20000
rect 13634 19200 13690 20000
rect 14094 19200 14150 20000
rect 14200 19230 14412 19258
rect 10796 17320 10824 19200
rect 10796 17292 11008 17320
rect 10704 17156 10824 17184
rect 10048 17138 10100 17144
rect 9956 16448 10008 16454
rect 9956 16390 10008 16396
rect 9956 15972 10008 15978
rect 9956 15914 10008 15920
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9772 15904 9824 15910
rect 9772 15846 9824 15852
rect 9784 15570 9812 15846
rect 9968 15706 9996 15914
rect 10060 15706 10088 17138
rect 10692 17060 10744 17066
rect 10692 17002 10744 17008
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 10152 16522 10180 16934
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 9956 15700 10008 15706
rect 9956 15642 10008 15648
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10046 15600 10102 15609
rect 9772 15564 9824 15570
rect 9772 15506 9824 15512
rect 9956 15564 10008 15570
rect 10046 15535 10102 15544
rect 9956 15506 10008 15512
rect 9496 15360 9548 15366
rect 9496 15302 9548 15308
rect 9508 15162 9536 15302
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9772 14952 9824 14958
rect 9772 14894 9824 14900
rect 9312 14816 9364 14822
rect 9312 14758 9364 14764
rect 9220 14476 9272 14482
rect 9220 14418 9272 14424
rect 9128 14340 9180 14346
rect 9128 14282 9180 14288
rect 9140 14249 9168 14282
rect 9126 14240 9182 14249
rect 9126 14175 9182 14184
rect 9126 14104 9182 14113
rect 9126 14039 9182 14048
rect 9140 13326 9168 14039
rect 9232 13802 9260 14418
rect 9496 14272 9548 14278
rect 9494 14240 9496 14249
rect 9680 14272 9732 14278
rect 9548 14240 9550 14249
rect 9680 14214 9732 14220
rect 9494 14175 9550 14184
rect 9586 14104 9642 14113
rect 9692 14090 9720 14214
rect 9642 14062 9720 14090
rect 9586 14039 9642 14048
rect 9579 14000 9631 14006
rect 9579 13942 9631 13948
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 9048 12974 9168 13002
rect 8942 12744 8998 12753
rect 9140 12730 9168 12974
rect 9232 12850 9260 13738
rect 9324 12986 9352 13874
rect 9591 13852 9619 13942
rect 9591 13824 9628 13852
rect 9600 13705 9628 13824
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9586 13560 9642 13569
rect 9586 13495 9588 13504
rect 9640 13495 9642 13504
rect 9588 13466 9640 13472
rect 9588 13252 9640 13258
rect 9588 13194 9640 13200
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 9312 12980 9364 12986
rect 9312 12922 9364 12928
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8942 12679 8998 12688
rect 9036 12708 9088 12714
rect 9140 12702 9260 12730
rect 9036 12650 9088 12656
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 8852 12096 8904 12102
rect 8852 12038 8904 12044
rect 8446 11996 8754 12016
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11920 8754 11940
rect 8850 11928 8906 11937
rect 8850 11863 8906 11872
rect 8300 11756 8352 11762
rect 8300 11698 8352 11704
rect 8300 11620 8352 11626
rect 8300 11562 8352 11568
rect 8116 11212 8168 11218
rect 8116 11154 8168 11160
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 7932 9648 7984 9654
rect 8036 9646 8156 9674
rect 7932 9590 7984 9596
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 9178 7604 9522
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7564 9172 7616 9178
rect 7564 9114 7616 9120
rect 7564 9036 7616 9042
rect 7564 8978 7616 8984
rect 7472 8424 7524 8430
rect 7472 8366 7524 8372
rect 7380 8288 7432 8294
rect 7380 8230 7432 8236
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 7392 7562 7420 8230
rect 7484 7750 7512 8366
rect 7576 8242 7604 8978
rect 7668 8362 7696 9454
rect 7748 8900 7800 8906
rect 7748 8842 7800 8848
rect 7760 8401 7788 8842
rect 7746 8392 7802 8401
rect 7656 8356 7708 8362
rect 7746 8327 7748 8336
rect 7656 8298 7708 8304
rect 7800 8327 7802 8336
rect 7748 8298 7800 8304
rect 7576 8214 7696 8242
rect 7562 8120 7618 8129
rect 7562 8055 7618 8064
rect 7472 7744 7524 7750
rect 7472 7686 7524 7692
rect 7300 7546 7420 7562
rect 7300 7540 7432 7546
rect 7300 7534 7380 7540
rect 7300 6798 7328 7534
rect 7380 7482 7432 7488
rect 7378 7440 7434 7449
rect 7378 7375 7380 7384
rect 7432 7375 7434 7384
rect 7380 7346 7432 7352
rect 7470 6896 7526 6905
rect 7470 6831 7472 6840
rect 7524 6831 7526 6840
rect 7472 6802 7524 6808
rect 7288 6792 7340 6798
rect 7288 6734 7340 6740
rect 7196 5160 7248 5166
rect 7196 5102 7248 5108
rect 7104 5092 7156 5098
rect 7104 5034 7156 5040
rect 7116 4826 7144 5034
rect 7208 4826 7236 5102
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7196 4820 7248 4826
rect 7196 4762 7248 4768
rect 7300 4570 7328 6734
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7392 5710 7420 6190
rect 7484 5846 7512 6802
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7576 5710 7604 8055
rect 7668 7206 7696 8214
rect 7852 7546 7880 9454
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 8022 7972 8910
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7944 7818 7972 7958
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7380 5704 7432 5710
rect 7380 5646 7432 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 7380 5160 7432 5166
rect 7380 5102 7432 5108
rect 7116 4542 7328 4570
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 3602 7052 4422
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6918 2544 6974 2553
rect 6918 2479 6974 2488
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 6564 1902 6592 2314
rect 7024 2310 7052 3538
rect 7116 3534 7144 4542
rect 7288 4480 7340 4486
rect 7288 4422 7340 4428
rect 7300 4146 7328 4422
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7300 3602 7328 4082
rect 7392 3738 7420 5102
rect 7564 4752 7616 4758
rect 7562 4720 7564 4729
rect 7616 4720 7618 4729
rect 7562 4655 7618 4664
rect 7564 4548 7616 4554
rect 7668 4536 7696 7142
rect 7932 6656 7984 6662
rect 7932 6598 7984 6604
rect 7944 6458 7972 6598
rect 7932 6452 7984 6458
rect 7932 6394 7984 6400
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7616 4508 7696 4536
rect 7564 4490 7616 4496
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 7380 3732 7432 3738
rect 7380 3674 7432 3680
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 7104 3528 7156 3534
rect 7104 3470 7156 3476
rect 7392 2774 7420 3674
rect 7484 3194 7512 4422
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7564 3528 7616 3534
rect 7564 3470 7616 3476
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7576 2774 7604 3470
rect 7668 3126 7696 3878
rect 7760 3398 7788 6326
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 5370 7880 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7944 3777 7972 6394
rect 8036 5370 8064 8502
rect 8128 5574 8156 9646
rect 8220 9042 8248 9862
rect 8208 9036 8260 9042
rect 8208 8978 8260 8984
rect 8312 8922 8340 11562
rect 8392 11552 8444 11558
rect 8392 11494 8444 11500
rect 8404 11218 8432 11494
rect 8864 11354 8892 11863
rect 8852 11348 8904 11354
rect 8852 11290 8904 11296
rect 8392 11212 8444 11218
rect 8392 11154 8444 11160
rect 8446 10908 8754 10928
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10832 8754 10852
rect 8446 9820 8754 9840
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9744 8754 9764
rect 8864 9674 8892 11290
rect 8956 10130 8984 12174
rect 9048 11812 9076 12650
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 9140 11937 9168 12582
rect 9126 11928 9182 11937
rect 9126 11863 9182 11872
rect 9048 11784 9168 11812
rect 9036 11212 9088 11218
rect 9036 11154 9088 11160
rect 9048 10130 9076 11154
rect 8944 10124 8996 10130
rect 8944 10066 8996 10072
rect 9036 10124 9088 10130
rect 9036 10066 9088 10072
rect 8772 9646 8892 9674
rect 8772 9110 8800 9646
rect 9048 9518 9076 10066
rect 9140 9994 9168 11784
rect 9128 9988 9180 9994
rect 9128 9930 9180 9936
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9036 9512 9088 9518
rect 9036 9454 9088 9460
rect 8944 9444 8996 9450
rect 8944 9386 8996 9392
rect 8760 9104 8812 9110
rect 8760 9046 8812 9052
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8220 8894 8340 8922
rect 8220 8616 8248 8894
rect 8446 8732 8754 8752
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8656 8754 8676
rect 8220 8588 8524 8616
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 6905 8248 8366
rect 8404 8090 8432 8434
rect 8496 8129 8524 8588
rect 8668 8424 8720 8430
rect 8668 8366 8720 8372
rect 8482 8120 8538 8129
rect 8392 8084 8444 8090
rect 8482 8055 8538 8064
rect 8392 8026 8444 8032
rect 8496 7954 8524 8055
rect 8484 7948 8536 7954
rect 8484 7890 8536 7896
rect 8680 7886 8708 8366
rect 8864 8090 8892 8978
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8446 7644 8754 7664
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7568 8754 7588
rect 8864 7478 8892 8026
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8206 6896 8262 6905
rect 8206 6831 8262 6840
rect 8852 6860 8904 6866
rect 8220 5710 8248 6831
rect 8852 6802 8904 6808
rect 8300 6724 8352 6730
rect 8300 6666 8352 6672
rect 8312 6390 8340 6666
rect 8446 6556 8754 6576
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6480 8754 6500
rect 8864 6458 8892 6802
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8312 5778 8340 6326
rect 8956 6066 8984 9386
rect 9140 9382 9168 9590
rect 9036 9376 9088 9382
rect 9036 9318 9088 9324
rect 9128 9376 9180 9382
rect 9128 9318 9180 9324
rect 9048 8945 9076 9318
rect 9034 8936 9090 8945
rect 9034 8871 9090 8880
rect 9036 8832 9088 8838
rect 9036 8774 9088 8780
rect 9048 8634 9076 8774
rect 9036 8628 9088 8634
rect 9036 8570 9088 8576
rect 9232 8566 9260 12702
rect 9312 12164 9364 12170
rect 9312 12106 9364 12112
rect 9324 11898 9352 12106
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9600 11014 9628 13194
rect 9692 11898 9720 13194
rect 9784 12850 9812 14894
rect 9864 14816 9916 14822
rect 9864 14758 9916 14764
rect 9876 12986 9904 14758
rect 9968 13462 9996 15506
rect 10060 15366 10088 15535
rect 10048 15360 10100 15366
rect 10048 15302 10100 15308
rect 10048 15156 10100 15162
rect 10048 15098 10100 15104
rect 9956 13456 10008 13462
rect 9956 13398 10008 13404
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9772 12708 9824 12714
rect 9772 12650 9824 12656
rect 9680 11892 9732 11898
rect 9680 11834 9732 11840
rect 9784 11218 9812 12650
rect 9772 11212 9824 11218
rect 9772 11154 9824 11160
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9416 10266 9444 10950
rect 9404 10260 9456 10266
rect 9404 10202 9456 10208
rect 9404 9988 9456 9994
rect 9404 9930 9456 9936
rect 9416 9722 9444 9930
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9404 9580 9456 9586
rect 9404 9522 9456 9528
rect 9416 9330 9444 9522
rect 9324 9302 9444 9330
rect 9324 9081 9352 9302
rect 9310 9072 9366 9081
rect 9310 9007 9366 9016
rect 9220 8560 9272 8566
rect 9220 8502 9272 8508
rect 9128 8492 9180 8498
rect 9128 8434 9180 8440
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 8864 6038 8984 6066
rect 8666 5808 8722 5817
rect 8300 5772 8352 5778
rect 8666 5743 8668 5752
rect 8300 5714 8352 5720
rect 8720 5743 8722 5752
rect 8668 5714 8720 5720
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8116 5568 8168 5574
rect 8116 5510 8168 5516
rect 8312 5370 8340 5714
rect 8446 5468 8754 5488
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5392 8754 5412
rect 8024 5364 8076 5370
rect 8024 5306 8076 5312
rect 8300 5364 8352 5370
rect 8352 5324 8524 5352
rect 8300 5306 8352 5312
rect 8024 5092 8076 5098
rect 8024 5034 8076 5040
rect 7930 3768 7986 3777
rect 7930 3703 7986 3712
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7852 3058 7880 3334
rect 8036 3058 8064 5034
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4690 8340 4966
rect 8496 4690 8524 5324
rect 8300 4684 8352 4690
rect 8300 4626 8352 4632
rect 8484 4684 8536 4690
rect 8484 4626 8536 4632
rect 8206 4584 8262 4593
rect 8206 4519 8262 4528
rect 8116 4004 8168 4010
rect 8116 3946 8168 3952
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7392 2746 7512 2774
rect 7576 2746 7696 2774
rect 7194 2544 7250 2553
rect 7194 2479 7250 2488
rect 7208 2378 7236 2479
rect 7484 2446 7512 2746
rect 7380 2440 7432 2446
rect 7380 2382 7432 2388
rect 7472 2440 7524 2446
rect 7472 2382 7524 2388
rect 7196 2372 7248 2378
rect 7196 2314 7248 2320
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6552 1896 6604 1902
rect 6552 1838 6604 1844
rect 7392 1766 7420 2382
rect 7668 2310 7696 2746
rect 7748 2644 7800 2650
rect 8128 2632 8156 3946
rect 8220 3058 8248 4519
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8208 3052 8260 3058
rect 8208 2994 8260 3000
rect 7748 2586 7800 2592
rect 8036 2604 8156 2632
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7288 1760 7340 1766
rect 7288 1702 7340 1708
rect 7380 1760 7432 1766
rect 7380 1702 7432 1708
rect 6828 1624 6880 1630
rect 6828 1566 6880 1572
rect 6840 800 6868 1566
rect 7300 800 7328 1702
rect 7760 800 7788 2586
rect 8036 2378 8064 2604
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 8024 2372 8076 2378
rect 8024 2314 8076 2320
rect 8128 800 8156 2450
rect 8220 1834 8248 2994
rect 8312 2582 8340 4422
rect 8446 4380 8754 4400
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4304 8754 4324
rect 8668 4208 8720 4214
rect 8668 4150 8720 4156
rect 8484 3936 8536 3942
rect 8484 3878 8536 3884
rect 8496 3534 8524 3878
rect 8680 3534 8708 4150
rect 8484 3528 8536 3534
rect 8484 3470 8536 3476
rect 8668 3528 8720 3534
rect 8668 3470 8720 3476
rect 8446 3292 8754 3312
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3216 8754 3236
rect 8390 2952 8446 2961
rect 8390 2887 8446 2896
rect 8300 2576 8352 2582
rect 8300 2518 8352 2524
rect 8208 1828 8260 1834
rect 8208 1770 8260 1776
rect 8312 1698 8340 2518
rect 8404 2446 8432 2887
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8446 2204 8754 2224
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2128 8754 2148
rect 8864 1902 8892 6038
rect 8944 5908 8996 5914
rect 8944 5850 8996 5856
rect 8956 4622 8984 5850
rect 8944 4616 8996 4622
rect 8944 4558 8996 4564
rect 9048 4486 9076 7958
rect 9140 7750 9168 8434
rect 9220 8356 9272 8362
rect 9220 8298 9272 8304
rect 9232 7886 9260 8298
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9140 5794 9168 7686
rect 9218 6352 9274 6361
rect 9218 6287 9274 6296
rect 9232 5914 9260 6287
rect 9324 5914 9352 9007
rect 9404 8832 9456 8838
rect 9404 8774 9456 8780
rect 9416 8090 9444 8774
rect 9600 8090 9628 10950
rect 9876 9722 9904 12922
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 9968 10826 9996 12786
rect 10060 12714 10088 15098
rect 10152 15076 10180 15982
rect 10244 15366 10272 16934
rect 10320 16892 10628 16912
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16816 10628 16836
rect 10704 16794 10732 17002
rect 10796 16998 10824 17156
rect 10784 16992 10836 16998
rect 10836 16952 10916 16980
rect 10784 16934 10836 16940
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10704 16114 10732 16730
rect 10784 16448 10836 16454
rect 10784 16390 10836 16396
rect 10796 16250 10824 16390
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10692 16108 10744 16114
rect 10692 16050 10744 16056
rect 10888 15994 10916 16952
rect 10980 16776 11008 17292
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 11072 16969 11100 17070
rect 11152 17060 11204 17066
rect 11152 17002 11204 17008
rect 11058 16960 11114 16969
rect 11058 16895 11114 16904
rect 11060 16788 11112 16794
rect 10980 16748 11060 16776
rect 11060 16730 11112 16736
rect 11060 16584 11112 16590
rect 11058 16552 11060 16561
rect 11112 16552 11114 16561
rect 11058 16487 11114 16496
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16153 11100 16390
rect 11058 16144 11114 16153
rect 11058 16079 11114 16088
rect 10704 15966 10916 15994
rect 11060 15972 11112 15978
rect 10320 15804 10628 15824
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15728 10628 15748
rect 10704 15586 10732 15966
rect 11060 15914 11112 15920
rect 10784 15904 10836 15910
rect 10784 15846 10836 15852
rect 10796 15638 10824 15846
rect 10336 15558 10732 15586
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10968 15564 11020 15570
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10232 15088 10284 15094
rect 10152 15048 10232 15076
rect 10232 15030 10284 15036
rect 10138 14920 10194 14929
rect 10336 14872 10364 15558
rect 10968 15506 11020 15512
rect 10692 15428 10744 15434
rect 10692 15370 10744 15376
rect 10138 14855 10194 14864
rect 10152 14074 10180 14855
rect 10244 14844 10364 14872
rect 10140 14068 10192 14074
rect 10140 14010 10192 14016
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 10152 13394 10180 13670
rect 10244 13410 10272 14844
rect 10320 14716 10628 14736
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14640 10628 14660
rect 10508 14544 10560 14550
rect 10322 14512 10378 14521
rect 10508 14486 10560 14492
rect 10322 14447 10324 14456
rect 10376 14447 10378 14456
rect 10324 14418 10376 14424
rect 10324 14272 10376 14278
rect 10324 14214 10376 14220
rect 10336 14074 10364 14214
rect 10324 14068 10376 14074
rect 10324 14010 10376 14016
rect 10520 13938 10548 14486
rect 10704 14278 10732 15370
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10520 13802 10548 13874
rect 10508 13796 10560 13802
rect 10508 13738 10560 13744
rect 10320 13628 10628 13648
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13552 10628 13572
rect 10140 13388 10192 13394
rect 10244 13382 10640 13410
rect 10140 13330 10192 13336
rect 10232 13252 10284 13258
rect 10232 13194 10284 13200
rect 10048 12708 10100 12714
rect 10048 12650 10100 12656
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10152 11898 10180 12582
rect 10140 11892 10192 11898
rect 10140 11834 10192 11840
rect 10140 11756 10192 11762
rect 10140 11698 10192 11704
rect 10152 11354 10180 11698
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9968 10798 10088 10826
rect 9956 10464 10008 10470
rect 9956 10406 10008 10412
rect 9968 10130 9996 10406
rect 9956 10124 10008 10130
rect 9956 10066 10008 10072
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9968 9722 9996 9862
rect 9864 9716 9916 9722
rect 9864 9658 9916 9664
rect 9956 9716 10008 9722
rect 9956 9658 10008 9664
rect 9680 9376 9732 9382
rect 9680 9318 9732 9324
rect 9692 9178 9720 9318
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9876 9058 9904 9658
rect 10060 9654 10088 10798
rect 10152 9654 10180 11086
rect 10244 10538 10272 13194
rect 10506 13152 10562 13161
rect 10506 13087 10562 13096
rect 10520 12850 10548 13087
rect 10612 12866 10640 13382
rect 10796 13274 10824 15302
rect 10980 15162 11008 15506
rect 11072 15337 11100 15914
rect 11058 15328 11114 15337
rect 11058 15263 11114 15272
rect 10876 15156 10928 15162
rect 10876 15098 10928 15104
rect 10968 15156 11020 15162
rect 10968 15098 11020 15104
rect 10888 15042 10916 15098
rect 10888 15014 11008 15042
rect 10980 14958 11008 15014
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14414 11008 14758
rect 11058 14648 11114 14657
rect 11058 14583 11114 14592
rect 10968 14408 11020 14414
rect 10968 14350 11020 14356
rect 10876 14272 10928 14278
rect 10876 14214 10928 14220
rect 10888 13462 10916 14214
rect 10980 14006 11008 14350
rect 11072 14249 11100 14583
rect 11058 14240 11114 14249
rect 11058 14175 11114 14184
rect 11058 14104 11114 14113
rect 11058 14039 11114 14048
rect 10968 14000 11020 14006
rect 10968 13942 11020 13948
rect 10980 13530 11008 13942
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10796 13246 10916 13274
rect 10508 12844 10560 12850
rect 10612 12838 10732 12866
rect 10508 12786 10560 12792
rect 10320 12540 10628 12560
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12464 10628 12484
rect 10704 12442 10732 12838
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10796 12374 10824 12718
rect 10784 12368 10836 12374
rect 10784 12310 10836 12316
rect 10796 12170 10824 12310
rect 10784 12164 10836 12170
rect 10784 12106 10836 12112
rect 10320 11452 10628 11472
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11376 10628 11396
rect 10796 11218 10824 12106
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10888 11150 10916 13246
rect 10966 13152 11022 13161
rect 10966 13087 11022 13096
rect 10980 12986 11008 13087
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10968 12640 11020 12646
rect 10968 12582 11020 12588
rect 10980 12442 11008 12582
rect 10968 12436 11020 12442
rect 10968 12378 11020 12384
rect 11072 12374 11100 14039
rect 11164 12646 11192 17002
rect 11256 16182 11284 19200
rect 11428 17536 11480 17542
rect 11428 17478 11480 17484
rect 11440 17134 11468 17478
rect 11520 17264 11572 17270
rect 11520 17206 11572 17212
rect 11428 17128 11480 17134
rect 11428 17070 11480 17076
rect 11336 16720 11388 16726
rect 11336 16662 11388 16668
rect 11244 16176 11296 16182
rect 11244 16118 11296 16124
rect 11256 14006 11284 16118
rect 11348 15978 11376 16662
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11348 15570 11376 15914
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11336 15360 11388 15366
rect 11336 15302 11388 15308
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11244 13728 11296 13734
rect 11244 13670 11296 13676
rect 11256 12986 11284 13670
rect 11348 13258 11376 15302
rect 11440 14521 11468 16390
rect 11532 16250 11560 17206
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11520 16040 11572 16046
rect 11520 15982 11572 15988
rect 11532 15910 11560 15982
rect 11520 15904 11572 15910
rect 11520 15846 11572 15852
rect 11532 15366 11560 15846
rect 11520 15360 11572 15366
rect 11518 15328 11520 15337
rect 11572 15328 11574 15337
rect 11518 15263 11574 15272
rect 11520 14884 11572 14890
rect 11520 14826 11572 14832
rect 11426 14512 11482 14521
rect 11426 14447 11482 14456
rect 11532 14396 11560 14826
rect 11440 14368 11560 14396
rect 11336 13252 11388 13258
rect 11336 13194 11388 13200
rect 11244 12980 11296 12986
rect 11244 12922 11296 12928
rect 11256 12889 11284 12922
rect 11242 12880 11298 12889
rect 11440 12832 11468 14368
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11532 12986 11560 13126
rect 11520 12980 11572 12986
rect 11520 12922 11572 12928
rect 11242 12815 11298 12824
rect 11348 12804 11468 12832
rect 11520 12844 11572 12850
rect 11152 12640 11204 12646
rect 11152 12582 11204 12588
rect 11060 12368 11112 12374
rect 11060 12310 11112 12316
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 10968 11552 11020 11558
rect 10966 11520 10968 11529
rect 11020 11520 11022 11529
rect 10966 11455 11022 11464
rect 11152 11280 11204 11286
rect 11152 11222 11204 11228
rect 10876 11144 10928 11150
rect 10876 11086 10928 11092
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10232 10532 10284 10538
rect 10232 10474 10284 10480
rect 10244 9994 10272 10474
rect 10320 10364 10628 10384
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10288 10628 10308
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 9692 9030 9904 9058
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9402 7984 9458 7993
rect 9402 7919 9404 7928
rect 9456 7919 9458 7928
rect 9404 7890 9456 7896
rect 9600 7818 9628 8026
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9416 7206 9444 7686
rect 9404 7200 9456 7206
rect 9404 7142 9456 7148
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9140 5766 9260 5794
rect 9128 5228 9180 5234
rect 9128 5170 9180 5176
rect 9036 4480 9088 4486
rect 9036 4422 9088 4428
rect 8942 4176 8998 4185
rect 8942 4111 8998 4120
rect 9036 4140 9088 4146
rect 8852 1896 8904 1902
rect 8852 1838 8904 1844
rect 8300 1692 8352 1698
rect 8300 1634 8352 1640
rect 8588 870 8708 898
rect 8588 800 8616 870
rect 1490 504 1546 513
rect 1490 439 1546 448
rect 1858 0 1914 800
rect 2226 0 2282 800
rect 2686 0 2742 800
rect 3054 0 3110 800
rect 3514 0 3570 800
rect 3974 0 4030 800
rect 4342 0 4398 800
rect 4802 0 4858 800
rect 5170 0 5226 800
rect 5630 0 5686 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6826 0 6882 800
rect 7286 0 7342 800
rect 7746 0 7802 800
rect 8114 0 8170 800
rect 8574 0 8630 800
rect 8680 762 8708 870
rect 8864 762 8892 1838
rect 8956 800 8984 4111
rect 9036 4082 9088 4088
rect 9048 2854 9076 4082
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9034 2680 9090 2689
rect 9034 2615 9036 2624
rect 9088 2615 9090 2624
rect 9036 2586 9088 2592
rect 9140 2582 9168 5170
rect 9232 4826 9260 5766
rect 9312 5568 9364 5574
rect 9312 5510 9364 5516
rect 9220 4820 9272 4826
rect 9220 4762 9272 4768
rect 9218 4720 9274 4729
rect 9218 4655 9220 4664
rect 9272 4655 9274 4664
rect 9220 4626 9272 4632
rect 9220 4480 9272 4486
rect 9220 4422 9272 4428
rect 9232 3505 9260 4422
rect 9324 4078 9352 5510
rect 9416 4486 9444 7142
rect 9692 6798 9720 9030
rect 9862 8936 9918 8945
rect 9862 8871 9918 8880
rect 9772 8832 9824 8838
rect 9772 8774 9824 8780
rect 9784 8566 9812 8774
rect 9876 8634 9904 8871
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9876 7562 9904 8026
rect 9784 7534 9904 7562
rect 9784 7206 9812 7534
rect 9864 7404 9916 7410
rect 9864 7346 9916 7352
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9876 6798 9904 7346
rect 9956 7336 10008 7342
rect 9956 7278 10008 7284
rect 9968 7002 9996 7278
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9864 6792 9916 6798
rect 9864 6734 9916 6740
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9600 6458 9628 6598
rect 9588 6452 9640 6458
rect 9588 6394 9640 6400
rect 9600 6100 9628 6394
rect 9692 6202 9720 6734
rect 9876 6304 9904 6734
rect 10060 6458 10088 9590
rect 10140 8968 10192 8974
rect 10140 8910 10192 8916
rect 10152 8566 10180 8910
rect 10140 8560 10192 8566
rect 10140 8502 10192 8508
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9956 6316 10008 6322
rect 9876 6276 9956 6304
rect 9956 6258 10008 6264
rect 10048 6248 10100 6254
rect 9692 6196 10048 6202
rect 9692 6190 10100 6196
rect 9692 6174 10088 6190
rect 9772 6112 9824 6118
rect 9600 6072 9720 6100
rect 9588 5908 9640 5914
rect 9588 5850 9640 5856
rect 9404 4480 9456 4486
rect 9404 4422 9456 4428
rect 9600 4282 9628 5850
rect 9692 4758 9720 6072
rect 9772 6054 9824 6060
rect 10048 6112 10100 6118
rect 10048 6054 10100 6060
rect 9784 5234 9812 6054
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9772 5228 9824 5234
rect 9772 5170 9824 5176
rect 9680 4752 9732 4758
rect 9680 4694 9732 4700
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9588 4276 9640 4282
rect 9588 4218 9640 4224
rect 9586 4176 9642 4185
rect 9404 4140 9456 4146
rect 9586 4111 9588 4120
rect 9404 4082 9456 4088
rect 9640 4111 9642 4120
rect 9588 4082 9640 4088
rect 9312 4072 9364 4078
rect 9312 4014 9364 4020
rect 9416 3738 9444 4082
rect 9692 4026 9720 4422
rect 9508 4010 9720 4026
rect 9496 4004 9720 4010
rect 9548 3998 9720 4004
rect 9496 3946 9548 3952
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9496 3528 9548 3534
rect 9218 3496 9274 3505
rect 9586 3496 9642 3505
rect 9548 3476 9586 3482
rect 9496 3470 9586 3476
rect 9508 3454 9586 3470
rect 9218 3431 9274 3440
rect 9586 3431 9642 3440
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 9232 1902 9260 2382
rect 9324 1970 9352 3334
rect 9588 2848 9640 2854
rect 9588 2790 9640 2796
rect 9402 2544 9458 2553
rect 9600 2514 9628 2790
rect 9402 2479 9458 2488
rect 9588 2508 9640 2514
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 9220 1896 9272 1902
rect 9220 1838 9272 1844
rect 9416 800 9444 2479
rect 9588 2450 9640 2456
rect 9692 2446 9720 3878
rect 9784 3670 9812 5170
rect 9876 4282 9904 5782
rect 10060 5710 10088 6054
rect 10152 5914 10180 7142
rect 10140 5908 10192 5914
rect 10140 5850 10192 5856
rect 10140 5772 10192 5778
rect 10140 5714 10192 5720
rect 10048 5704 10100 5710
rect 10048 5646 10100 5652
rect 9956 5568 10008 5574
rect 9956 5510 10008 5516
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9968 4010 9996 5510
rect 10152 5370 10180 5714
rect 10244 5642 10272 9930
rect 10796 9450 10824 10610
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10888 9518 10916 10066
rect 11060 9920 11112 9926
rect 11060 9862 11112 9868
rect 11072 9654 11100 9862
rect 11164 9654 11192 11222
rect 11256 11218 11284 12174
rect 11348 11830 11376 12804
rect 11520 12786 11572 12792
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 11336 11824 11388 11830
rect 11336 11766 11388 11772
rect 11440 11694 11468 12106
rect 11428 11688 11480 11694
rect 11428 11630 11480 11636
rect 11532 11234 11560 12786
rect 11624 11558 11652 19200
rect 11704 17264 11756 17270
rect 11702 17232 11704 17241
rect 11756 17232 11758 17241
rect 11702 17167 11758 17176
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 11704 17128 11756 17134
rect 11900 17105 11928 17138
rect 12084 17134 12112 19200
rect 12452 17762 12480 19200
rect 12452 17734 12664 17762
rect 12532 17604 12584 17610
rect 12532 17546 12584 17552
rect 12194 17436 12502 17456
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17360 12502 17380
rect 12072 17128 12124 17134
rect 11704 17070 11756 17076
rect 11886 17096 11942 17105
rect 11716 15570 11744 17070
rect 12072 17070 12124 17076
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 11886 17031 11942 17040
rect 11888 16992 11940 16998
rect 11888 16934 11940 16940
rect 11796 16652 11848 16658
rect 11796 16594 11848 16600
rect 11704 15564 11756 15570
rect 11704 15506 11756 15512
rect 11702 15464 11758 15473
rect 11702 15399 11758 15408
rect 11716 14414 11744 15399
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11704 13796 11756 13802
rect 11704 13738 11756 13744
rect 11716 12782 11744 13738
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11612 11552 11664 11558
rect 11612 11494 11664 11500
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11348 11206 11560 11234
rect 11256 10674 11284 11154
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11256 10266 11284 10610
rect 11244 10260 11296 10266
rect 11244 10202 11296 10208
rect 11348 9674 11376 11206
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11060 9648 11112 9654
rect 11060 9590 11112 9596
rect 11152 9648 11204 9654
rect 11152 9590 11204 9596
rect 11256 9646 11376 9674
rect 11440 9654 11468 11086
rect 11624 10810 11652 11086
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11532 9722 11560 9998
rect 11520 9716 11572 9722
rect 11520 9658 11572 9664
rect 11428 9648 11480 9654
rect 11256 9586 11284 9646
rect 11428 9590 11480 9596
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 11256 9382 11284 9522
rect 11244 9376 11296 9382
rect 11244 9318 11296 9324
rect 10320 9276 10628 9296
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9200 10628 9220
rect 10782 9208 10838 9217
rect 10782 9143 10838 9152
rect 10796 9042 10824 9143
rect 10784 9036 10836 9042
rect 10784 8978 10836 8984
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 10600 8900 10652 8906
rect 10600 8842 10652 8848
rect 10612 8634 10640 8842
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10980 8566 11008 8910
rect 10876 8560 10928 8566
rect 10876 8502 10928 8508
rect 10968 8560 11020 8566
rect 10968 8502 11020 8508
rect 10320 8188 10628 8208
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8112 10628 8132
rect 10888 7954 10916 8502
rect 10876 7948 10928 7954
rect 10876 7890 10928 7896
rect 10784 7880 10836 7886
rect 10322 7848 10378 7857
rect 10784 7822 10836 7828
rect 10322 7783 10378 7792
rect 10336 7750 10364 7783
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10416 7744 10468 7750
rect 10416 7686 10468 7692
rect 10428 7546 10456 7686
rect 10416 7540 10468 7546
rect 10416 7482 10468 7488
rect 10320 7100 10628 7120
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7024 10628 7044
rect 10796 6338 10824 7822
rect 10876 7200 10928 7206
rect 10876 7142 10928 7148
rect 10888 6458 10916 7142
rect 10876 6452 10928 6458
rect 10876 6394 10928 6400
rect 10796 6310 10916 6338
rect 10980 6322 11008 8502
rect 11060 7880 11112 7886
rect 11060 7822 11112 7828
rect 11072 7478 11100 7822
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11152 7472 11204 7478
rect 11152 7414 11204 7420
rect 11164 7342 11192 7414
rect 11152 7336 11204 7342
rect 11058 7304 11114 7313
rect 11152 7278 11204 7284
rect 11058 7239 11114 7248
rect 11072 6458 11100 7239
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 10320 6012 10628 6032
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5936 10628 5956
rect 10232 5636 10284 5642
rect 10232 5578 10284 5584
rect 10140 5364 10192 5370
rect 10140 5306 10192 5312
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 10060 4622 10088 4966
rect 10048 4616 10100 4622
rect 10048 4558 10100 4564
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10152 4282 10180 4558
rect 10140 4276 10192 4282
rect 10140 4218 10192 4224
rect 10046 4176 10102 4185
rect 10046 4111 10102 4120
rect 9864 4004 9916 4010
rect 9864 3946 9916 3952
rect 9956 4004 10008 4010
rect 9956 3946 10008 3952
rect 9772 3664 9824 3670
rect 9772 3606 9824 3612
rect 9784 3058 9812 3606
rect 9772 3052 9824 3058
rect 9772 2994 9824 3000
rect 9876 2922 9904 3946
rect 10060 3534 10088 4111
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10048 3392 10100 3398
rect 10152 3380 10180 4218
rect 10244 3534 10272 5578
rect 10692 5296 10744 5302
rect 10692 5238 10744 5244
rect 10320 4924 10628 4944
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4848 10628 4868
rect 10600 4684 10652 4690
rect 10704 4672 10732 5238
rect 10652 4644 10732 4672
rect 10600 4626 10652 4632
rect 10324 4480 10376 4486
rect 10324 4422 10376 4428
rect 10336 4185 10364 4422
rect 10322 4176 10378 4185
rect 10322 4111 10378 4120
rect 10704 4078 10732 4644
rect 10796 4146 10824 6190
rect 10888 4622 10916 6310
rect 10968 6316 11020 6322
rect 10968 6258 11020 6264
rect 10980 5914 11008 6258
rect 10968 5908 11020 5914
rect 10968 5850 11020 5856
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 10784 4140 10836 4146
rect 10784 4082 10836 4088
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10320 3836 10628 3856
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3760 10628 3780
rect 10324 3664 10376 3670
rect 10322 3632 10324 3641
rect 10376 3632 10378 3641
rect 10322 3567 10378 3576
rect 10232 3528 10284 3534
rect 10232 3470 10284 3476
rect 10152 3352 10272 3380
rect 10048 3334 10100 3340
rect 9864 2916 9916 2922
rect 9864 2858 9916 2864
rect 9876 2514 9904 2858
rect 10060 2774 10088 3334
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 9968 2746 10088 2774
rect 9864 2508 9916 2514
rect 9864 2450 9916 2456
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 9968 2258 9996 2746
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 10060 2446 10088 2586
rect 10048 2440 10100 2446
rect 10048 2382 10100 2388
rect 10048 2304 10100 2310
rect 9968 2252 10048 2258
rect 9968 2246 10100 2252
rect 9968 2230 10088 2246
rect 9772 2100 9824 2106
rect 9772 2042 9824 2048
rect 9784 800 9812 2042
rect 10152 1986 10180 3130
rect 10244 2530 10272 3352
rect 10320 2748 10628 2768
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2672 10628 2692
rect 10796 2650 10824 4082
rect 10980 3602 11008 5306
rect 11072 5030 11100 6394
rect 11060 5024 11112 5030
rect 11112 4984 11192 5012
rect 11060 4966 11112 4972
rect 11060 4140 11112 4146
rect 11060 4082 11112 4088
rect 10968 3596 11020 3602
rect 10968 3538 11020 3544
rect 10980 3058 11008 3538
rect 11072 3194 11100 4082
rect 11060 3188 11112 3194
rect 11060 3130 11112 3136
rect 10968 3052 11020 3058
rect 11164 3040 11192 4984
rect 11256 4865 11284 9318
rect 11336 8356 11388 8362
rect 11336 8298 11388 8304
rect 11348 7041 11376 8298
rect 11440 7154 11468 9590
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11520 8424 11572 8430
rect 11520 8366 11572 8372
rect 11532 7954 11560 8366
rect 11520 7948 11572 7954
rect 11520 7890 11572 7896
rect 11532 7274 11560 7890
rect 11624 7478 11652 9522
rect 11716 8294 11744 12718
rect 11808 10554 11836 16594
rect 11900 16522 11928 16934
rect 12452 16697 12480 17070
rect 12544 16998 12572 17546
rect 12636 17202 12664 17734
rect 12624 17196 12676 17202
rect 12676 17156 12756 17184
rect 12624 17138 12676 17144
rect 12532 16992 12584 16998
rect 12532 16934 12584 16940
rect 12438 16688 12494 16697
rect 12438 16623 12494 16632
rect 12070 16552 12126 16561
rect 11888 16516 11940 16522
rect 12070 16487 12126 16496
rect 12530 16552 12586 16561
rect 12530 16487 12586 16496
rect 11888 16458 11940 16464
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11900 14906 11928 16050
rect 11980 16040 12032 16046
rect 11980 15982 12032 15988
rect 11992 15881 12020 15982
rect 11978 15872 12034 15881
rect 11978 15807 12034 15816
rect 11978 15600 12034 15609
rect 11978 15535 12034 15544
rect 11992 15162 12020 15535
rect 11980 15156 12032 15162
rect 11980 15098 12032 15104
rect 11900 14878 12020 14906
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11900 14618 11928 14758
rect 11888 14612 11940 14618
rect 11888 14554 11940 14560
rect 11992 14362 12020 14878
rect 11900 14334 12020 14362
rect 11900 13734 11928 14334
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11992 14074 12020 14214
rect 11980 14068 12032 14074
rect 12084 14056 12112 16487
rect 12544 16454 12572 16487
rect 12532 16448 12584 16454
rect 12532 16390 12584 16396
rect 12194 16348 12502 16368
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16272 12502 16292
rect 12532 16244 12584 16250
rect 12532 16186 12584 16192
rect 12194 15260 12502 15280
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15184 12502 15204
rect 12164 15088 12216 15094
rect 12544 15042 12572 16186
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 12164 15030 12216 15036
rect 12176 14793 12204 15030
rect 12268 15026 12572 15042
rect 12636 15026 12664 16079
rect 12256 15020 12572 15026
rect 12308 15014 12572 15020
rect 12624 15020 12676 15026
rect 12256 14962 12308 14968
rect 12624 14962 12676 14968
rect 12440 14952 12492 14958
rect 12438 14920 12440 14929
rect 12492 14920 12494 14929
rect 12438 14855 12494 14864
rect 12162 14784 12218 14793
rect 12162 14719 12218 14728
rect 12728 14482 12756 17156
rect 12912 16182 12940 19200
rect 13084 16992 13136 16998
rect 13084 16934 13136 16940
rect 12990 16416 13046 16425
rect 12990 16351 13046 16360
rect 12900 16176 12952 16182
rect 12900 16118 12952 16124
rect 13004 15502 13032 16351
rect 12992 15496 13044 15502
rect 12992 15438 13044 15444
rect 13096 15366 13124 16934
rect 13176 16516 13228 16522
rect 13176 16458 13228 16464
rect 13188 16425 13216 16458
rect 13174 16416 13230 16425
rect 13174 16351 13230 16360
rect 13280 16114 13308 19200
rect 13452 17128 13504 17134
rect 13452 17070 13504 17076
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13176 16108 13228 16114
rect 13176 16050 13228 16056
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 12900 15360 12952 15366
rect 12900 15302 12952 15308
rect 13084 15360 13136 15366
rect 13084 15302 13136 15308
rect 12912 15162 12940 15302
rect 12808 15156 12860 15162
rect 12808 15098 12860 15104
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12716 14476 12768 14482
rect 12716 14418 12768 14424
rect 12194 14172 12502 14192
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14096 12502 14116
rect 12084 14028 12204 14056
rect 11980 14010 12032 14016
rect 12176 13802 12204 14028
rect 12544 13954 12572 14418
rect 12714 14376 12770 14385
rect 12714 14311 12716 14320
rect 12768 14311 12770 14320
rect 12716 14282 12768 14288
rect 12820 14074 12848 15098
rect 13096 15042 13124 15302
rect 13004 15014 13124 15042
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12912 14346 12940 14826
rect 13004 14482 13032 15014
rect 13084 14952 13136 14958
rect 13084 14894 13136 14900
rect 12992 14476 13044 14482
rect 12992 14418 13044 14424
rect 12990 14376 13046 14385
rect 12900 14340 12952 14346
rect 12990 14311 13046 14320
rect 12900 14282 12952 14288
rect 12808 14068 12860 14074
rect 12808 14010 12860 14016
rect 12900 14068 12952 14074
rect 12900 14010 12952 14016
rect 12452 13926 12572 13954
rect 12624 14000 12676 14006
rect 12624 13942 12676 13948
rect 12164 13796 12216 13802
rect 12164 13738 12216 13744
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 12254 13696 12310 13705
rect 12254 13631 12310 13640
rect 12268 13462 12296 13631
rect 12072 13456 12124 13462
rect 12072 13398 12124 13404
rect 12256 13456 12308 13462
rect 12256 13398 12308 13404
rect 12084 12986 12112 13398
rect 12452 13258 12480 13926
rect 12532 13864 12584 13870
rect 12532 13806 12584 13812
rect 12544 13705 12572 13806
rect 12530 13696 12586 13705
rect 12530 13631 12586 13640
rect 12636 13376 12664 13942
rect 12544 13348 12664 13376
rect 12440 13252 12492 13258
rect 12440 13194 12492 13200
rect 12194 13084 12502 13104
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13008 12502 13028
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12544 12832 12572 13348
rect 12808 13320 12860 13326
rect 12728 13280 12808 13308
rect 12624 13252 12676 13258
rect 12624 13194 12676 13200
rect 12452 12804 12572 12832
rect 11980 12776 12032 12782
rect 11980 12718 12032 12724
rect 11992 12322 12020 12718
rect 12452 12442 12480 12804
rect 12532 12708 12584 12714
rect 12636 12696 12664 13194
rect 12584 12668 12664 12696
rect 12532 12650 12584 12656
rect 12440 12436 12492 12442
rect 12440 12378 12492 12384
rect 11900 12294 12020 12322
rect 12544 12306 12572 12650
rect 12532 12300 12584 12306
rect 11900 11898 11928 12294
rect 12532 12242 12584 12248
rect 12544 12102 12572 12242
rect 12532 12096 12584 12102
rect 12532 12038 12584 12044
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12728 12050 12756 13280
rect 12808 13262 12860 13268
rect 12808 12776 12860 12782
rect 12808 12718 12860 12724
rect 12820 12238 12848 12718
rect 12808 12232 12860 12238
rect 12912 12220 12940 14010
rect 13004 13870 13032 14311
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13004 12918 13032 13806
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 13004 12345 13032 12854
rect 12990 12336 13046 12345
rect 12990 12271 13046 12280
rect 12912 12192 13032 12220
rect 12808 12174 12860 12180
rect 12194 11996 12502 12016
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11920 12502 11940
rect 11888 11892 11940 11898
rect 11888 11834 11940 11840
rect 11978 11792 12034 11801
rect 11888 11756 11940 11762
rect 11978 11727 11980 11736
rect 11888 11698 11940 11704
rect 12032 11727 12034 11736
rect 11980 11698 12032 11704
rect 11900 10713 11928 11698
rect 12348 11688 12400 11694
rect 12348 11630 12400 11636
rect 12360 11558 12388 11630
rect 12544 11626 12572 12038
rect 12532 11620 12584 11626
rect 12532 11562 12584 11568
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12440 11552 12492 11558
rect 12636 11506 12664 12038
rect 12728 12022 12940 12050
rect 12714 11928 12770 11937
rect 12714 11863 12770 11872
rect 12492 11500 12664 11506
rect 12440 11494 12664 11500
rect 12452 11478 12664 11494
rect 12452 11098 12480 11478
rect 12452 11070 12572 11098
rect 12194 10908 12502 10928
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10832 12502 10852
rect 11886 10704 11942 10713
rect 11886 10639 11942 10648
rect 11808 10526 11928 10554
rect 11796 8424 11848 8430
rect 11796 8366 11848 8372
rect 11704 8288 11756 8294
rect 11704 8230 11756 8236
rect 11704 8084 11756 8090
rect 11704 8026 11756 8032
rect 11612 7472 11664 7478
rect 11612 7414 11664 7420
rect 11520 7268 11572 7274
rect 11520 7210 11572 7216
rect 11440 7126 11652 7154
rect 11334 7032 11390 7041
rect 11334 6967 11390 6976
rect 11520 6996 11572 7002
rect 11520 6938 11572 6944
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11348 5234 11376 5850
rect 11336 5228 11388 5234
rect 11336 5170 11388 5176
rect 11334 5128 11390 5137
rect 11334 5063 11390 5072
rect 11242 4856 11298 4865
rect 11242 4791 11298 4800
rect 11348 4758 11376 5063
rect 11428 4820 11480 4826
rect 11428 4762 11480 4768
rect 11336 4752 11388 4758
rect 11242 4720 11298 4729
rect 11336 4694 11388 4700
rect 11242 4655 11298 4664
rect 11256 3194 11284 4655
rect 11440 4282 11468 4762
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11336 4072 11388 4078
rect 11334 4040 11336 4049
rect 11388 4040 11390 4049
rect 11334 3975 11390 3984
rect 11244 3188 11296 3194
rect 11244 3130 11296 3136
rect 10968 2994 11020 3000
rect 11072 3012 11192 3040
rect 11072 2938 11100 3012
rect 10980 2910 11100 2938
rect 11150 2952 11206 2961
rect 10980 2650 11008 2910
rect 11150 2887 11206 2896
rect 11164 2836 11192 2887
rect 11072 2808 11192 2836
rect 11244 2848 11296 2854
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10692 2576 10744 2582
rect 10244 2502 10364 2530
rect 10692 2518 10744 2524
rect 10232 2440 10284 2446
rect 10232 2382 10284 2388
rect 10244 2106 10272 2382
rect 10232 2100 10284 2106
rect 10232 2042 10284 2048
rect 10152 1958 10272 1986
rect 10244 800 10272 1958
rect 10336 1766 10364 2502
rect 10324 1760 10376 1766
rect 10324 1702 10376 1708
rect 10704 800 10732 2518
rect 11072 800 11100 2808
rect 11244 2790 11296 2796
rect 11256 2446 11284 2790
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11440 2038 11468 4218
rect 11532 2938 11560 6938
rect 11624 6662 11652 7126
rect 11612 6656 11664 6662
rect 11612 6598 11664 6604
rect 11624 6458 11652 6598
rect 11612 6452 11664 6458
rect 11612 6394 11664 6400
rect 11716 5794 11744 8026
rect 11624 5766 11744 5794
rect 11624 4690 11652 5766
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 11612 3936 11664 3942
rect 11612 3878 11664 3884
rect 11624 3398 11652 3878
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11624 3126 11652 3334
rect 11612 3120 11664 3126
rect 11612 3062 11664 3068
rect 11716 3058 11744 5646
rect 11808 5137 11836 8366
rect 11900 8090 11928 10526
rect 12544 10266 12572 11070
rect 12624 10804 12676 10810
rect 12624 10746 12676 10752
rect 12532 10260 12584 10266
rect 12532 10202 12584 10208
rect 12544 10169 12572 10202
rect 12530 10160 12586 10169
rect 12072 10124 12124 10130
rect 12530 10095 12586 10104
rect 12072 10066 12124 10072
rect 12084 9518 12112 10066
rect 12194 9820 12502 9840
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9744 12502 9764
rect 12636 9518 12664 10746
rect 12072 9512 12124 9518
rect 12624 9512 12676 9518
rect 12072 9454 12124 9460
rect 12346 9480 12402 9489
rect 12624 9454 12676 9460
rect 12346 9415 12348 9424
rect 12400 9415 12402 9424
rect 12532 9444 12584 9450
rect 12348 9386 12400 9392
rect 12532 9386 12584 9392
rect 12072 9036 12124 9042
rect 12072 8978 12124 8984
rect 11980 8832 12032 8838
rect 11980 8774 12032 8780
rect 11992 8430 12020 8774
rect 11980 8424 12032 8430
rect 11980 8366 12032 8372
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 11978 7984 12034 7993
rect 11978 7919 12034 7928
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11900 6458 11928 7686
rect 11888 6452 11940 6458
rect 11888 6394 11940 6400
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11794 5128 11850 5137
rect 11794 5063 11850 5072
rect 11796 4616 11848 4622
rect 11796 4558 11848 4564
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 11532 2910 11744 2938
rect 11612 2848 11664 2854
rect 11532 2808 11612 2836
rect 11428 2032 11480 2038
rect 11428 1974 11480 1980
rect 11532 800 11560 2808
rect 11612 2790 11664 2796
rect 11716 2514 11744 2910
rect 11704 2508 11756 2514
rect 11704 2450 11756 2456
rect 11808 2258 11836 4558
rect 11900 3534 11928 6287
rect 11992 5522 12020 7919
rect 12084 7528 12112 8978
rect 12194 8732 12502 8752
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8656 12502 8676
rect 12544 8634 12572 9386
rect 12728 8786 12756 11863
rect 12808 11824 12860 11830
rect 12808 11766 12860 11772
rect 12820 11558 12848 11766
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 9602 12848 11494
rect 12912 11150 12940 12022
rect 13004 11937 13032 12192
rect 12990 11928 13046 11937
rect 12990 11863 13046 11872
rect 12990 11792 13046 11801
rect 12990 11727 13046 11736
rect 13004 11626 13032 11727
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13096 11558 13124 14894
rect 13188 14521 13216 16050
rect 13268 15700 13320 15706
rect 13268 15642 13320 15648
rect 13280 15366 13308 15642
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13174 14512 13230 14521
rect 13174 14447 13230 14456
rect 13176 14408 13228 14414
rect 13176 14350 13228 14356
rect 13188 12209 13216 14350
rect 13280 14074 13308 15302
rect 13372 14385 13400 16390
rect 13358 14376 13414 14385
rect 13358 14311 13414 14320
rect 13268 14068 13320 14074
rect 13268 14010 13320 14016
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13266 13968 13322 13977
rect 13266 13903 13268 13912
rect 13320 13903 13322 13912
rect 13268 13874 13320 13880
rect 13372 13870 13400 14010
rect 13360 13864 13412 13870
rect 13360 13806 13412 13812
rect 13358 13696 13414 13705
rect 13358 13631 13414 13640
rect 13266 13424 13322 13433
rect 13266 13359 13322 13368
rect 13280 13258 13308 13359
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13268 12776 13320 12782
rect 13268 12718 13320 12724
rect 13174 12200 13230 12209
rect 13174 12135 13230 12144
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13188 11898 13216 12038
rect 13176 11892 13228 11898
rect 13176 11834 13228 11840
rect 13084 11552 13136 11558
rect 13084 11494 13136 11500
rect 12900 11144 12952 11150
rect 12952 11092 13124 11098
rect 12900 11086 13124 11092
rect 12912 11070 13124 11086
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12912 10130 12940 10950
rect 13096 10674 13124 11070
rect 13176 11008 13228 11014
rect 13176 10950 13228 10956
rect 12992 10668 13044 10674
rect 12992 10610 13044 10616
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 13004 10130 13032 10610
rect 13188 10452 13216 10950
rect 13280 10742 13308 12718
rect 13372 11898 13400 13631
rect 13464 12306 13492 17070
rect 13542 16552 13598 16561
rect 13542 16487 13544 16496
rect 13596 16487 13598 16496
rect 13544 16458 13596 16464
rect 13544 16108 13596 16114
rect 13544 16050 13596 16056
rect 13452 12300 13504 12306
rect 13452 12242 13504 12248
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13464 11830 13492 12106
rect 13452 11824 13504 11830
rect 13452 11766 13504 11772
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13268 10736 13320 10742
rect 13268 10678 13320 10684
rect 13188 10424 13308 10452
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12992 10124 13044 10130
rect 12992 10066 13044 10072
rect 13280 9994 13308 10424
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9722 13124 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 12820 9574 13124 9602
rect 12992 9376 13044 9382
rect 12992 9318 13044 9324
rect 12900 8900 12952 8906
rect 12900 8842 12952 8848
rect 12636 8758 12756 8786
rect 12532 8628 12584 8634
rect 12532 8570 12584 8576
rect 12636 8022 12664 8758
rect 12714 8664 12770 8673
rect 12714 8599 12770 8608
rect 12728 8566 12756 8599
rect 12716 8560 12768 8566
rect 12716 8502 12768 8508
rect 12716 8288 12768 8294
rect 12716 8230 12768 8236
rect 12624 8016 12676 8022
rect 12624 7958 12676 7964
rect 12728 7886 12756 8230
rect 12716 7880 12768 7886
rect 12716 7822 12768 7828
rect 12624 7744 12676 7750
rect 12624 7686 12676 7692
rect 12194 7644 12502 7664
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7568 12502 7588
rect 12084 7500 12204 7528
rect 12176 7002 12204 7500
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12532 7472 12584 7478
rect 12532 7414 12584 7420
rect 12256 7404 12308 7410
rect 12256 7346 12308 7352
rect 12164 6996 12216 7002
rect 12164 6938 12216 6944
rect 12268 6730 12296 7346
rect 12360 6866 12388 7414
rect 12544 7002 12572 7414
rect 12636 7206 12664 7686
rect 12624 7200 12676 7206
rect 12624 7142 12676 7148
rect 12532 6996 12584 7002
rect 12532 6938 12584 6944
rect 12624 6996 12676 7002
rect 12624 6938 12676 6944
rect 12348 6860 12400 6866
rect 12348 6802 12400 6808
rect 12256 6724 12308 6730
rect 12256 6666 12308 6672
rect 12194 6556 12502 6576
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6480 12502 6500
rect 12440 6384 12492 6390
rect 12346 6352 12402 6361
rect 12440 6326 12492 6332
rect 12346 6287 12348 6296
rect 12400 6287 12402 6296
rect 12348 6258 12400 6264
rect 12452 6100 12480 6326
rect 12544 6254 12572 6938
rect 12636 6390 12664 6938
rect 12728 6662 12756 7822
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12820 7002 12848 7754
rect 12912 7410 12940 8842
rect 13004 8634 13032 9318
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 13004 7018 13032 7686
rect 12808 6996 12860 7002
rect 12808 6938 12860 6944
rect 12912 6990 13032 7018
rect 12716 6656 12768 6662
rect 12716 6598 12768 6604
rect 12728 6458 12756 6598
rect 12716 6452 12768 6458
rect 12716 6394 12768 6400
rect 12912 6390 12940 6990
rect 12990 6896 13046 6905
rect 12990 6831 13046 6840
rect 13004 6390 13032 6831
rect 12624 6384 12676 6390
rect 12624 6326 12676 6332
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12992 6384 13044 6390
rect 12992 6326 13044 6332
rect 12532 6248 12584 6254
rect 12532 6190 12584 6196
rect 12900 6248 12952 6254
rect 12900 6190 12952 6196
rect 12624 6180 12676 6186
rect 12624 6122 12676 6128
rect 12452 6072 12572 6100
rect 11992 5494 12112 5522
rect 11980 5364 12032 5370
rect 11980 5306 12032 5312
rect 11992 4146 12020 5306
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11888 3528 11940 3534
rect 11886 3496 11888 3505
rect 11940 3496 11942 3505
rect 11886 3431 11942 3440
rect 11888 3392 11940 3398
rect 11888 3334 11940 3340
rect 11978 3360 12034 3369
rect 11900 2378 11928 3334
rect 12084 3346 12112 5494
rect 12194 5468 12502 5488
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5392 12502 5412
rect 12544 5137 12572 6072
rect 12636 5710 12664 6122
rect 12912 5817 12940 6190
rect 12898 5808 12954 5817
rect 12808 5772 12860 5778
rect 12898 5743 12954 5752
rect 12808 5714 12860 5720
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12530 5128 12586 5137
rect 12530 5063 12586 5072
rect 12532 5024 12584 5030
rect 12532 4966 12584 4972
rect 12544 4622 12572 4966
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12194 4380 12502 4400
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4304 12502 4324
rect 12544 4078 12572 4558
rect 12624 4548 12676 4554
rect 12624 4490 12676 4496
rect 12636 4282 12664 4490
rect 12728 4282 12756 5510
rect 12820 5302 12848 5714
rect 13096 5658 13124 9574
rect 13174 8120 13230 8129
rect 13174 8055 13230 8064
rect 13188 7818 13216 8055
rect 13176 7812 13228 7818
rect 13176 7754 13228 7760
rect 13174 7032 13230 7041
rect 13174 6967 13230 6976
rect 13188 6662 13216 6967
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13176 6452 13228 6458
rect 13176 6394 13228 6400
rect 12912 5630 13124 5658
rect 12808 5296 12860 5302
rect 12808 5238 12860 5244
rect 12806 5128 12862 5137
rect 12806 5063 12862 5072
rect 12624 4276 12676 4282
rect 12624 4218 12676 4224
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12532 4072 12584 4078
rect 12532 4014 12584 4020
rect 12820 3942 12848 5063
rect 12808 3936 12860 3942
rect 12808 3878 12860 3884
rect 12622 3632 12678 3641
rect 12622 3567 12678 3576
rect 12162 3496 12218 3505
rect 12162 3431 12164 3440
rect 12216 3431 12218 3440
rect 12164 3402 12216 3408
rect 12636 3398 12664 3567
rect 12034 3318 12112 3346
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 11978 3295 12034 3304
rect 12084 3194 12112 3318
rect 12194 3292 12502 3312
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3216 12502 3236
rect 12072 3188 12124 3194
rect 12072 3130 12124 3136
rect 12716 3120 12768 3126
rect 12714 3088 12716 3097
rect 12912 3108 12940 5630
rect 12992 5568 13044 5574
rect 13188 5522 13216 6394
rect 12992 5510 13044 5516
rect 13004 4593 13032 5510
rect 13096 5494 13216 5522
rect 12990 4584 13046 4593
rect 12990 4519 13046 4528
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 13004 3126 13032 3674
rect 13096 3602 13124 5494
rect 13174 5400 13230 5409
rect 13174 5335 13176 5344
rect 13228 5335 13230 5344
rect 13176 5306 13228 5312
rect 13188 4185 13216 5306
rect 13174 4176 13230 4185
rect 13174 4111 13230 4120
rect 13084 3596 13136 3602
rect 13084 3538 13136 3544
rect 13176 3596 13228 3602
rect 13176 3538 13228 3544
rect 13084 3188 13136 3194
rect 13084 3130 13136 3136
rect 12768 3088 12940 3108
rect 12770 3080 12940 3088
rect 12992 3120 13044 3126
rect 12992 3062 13044 3068
rect 13096 3058 13124 3130
rect 12714 3023 12770 3032
rect 13084 3052 13136 3058
rect 13084 2994 13136 3000
rect 12716 2984 12768 2990
rect 12714 2952 12716 2961
rect 12768 2952 12770 2961
rect 12714 2887 12770 2896
rect 12532 2508 12584 2514
rect 12532 2450 12584 2456
rect 11888 2372 11940 2378
rect 11888 2314 11940 2320
rect 11808 2230 11928 2258
rect 11900 800 11928 2230
rect 12194 2204 12502 2224
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2128 12502 2148
rect 12544 2088 12572 2450
rect 12992 2440 13044 2446
rect 12990 2408 12992 2417
rect 13044 2408 13046 2417
rect 12716 2372 12768 2378
rect 12990 2343 13046 2352
rect 12716 2314 12768 2320
rect 12360 2060 12572 2088
rect 12360 800 12388 2060
rect 12728 800 12756 2314
rect 13188 800 13216 3538
rect 13280 2417 13308 9930
rect 13372 9489 13400 11494
rect 13556 11354 13584 16050
rect 13648 15570 13676 19200
rect 14108 19122 14136 19200
rect 14200 19122 14228 19230
rect 14108 19094 14228 19122
rect 13820 17128 13872 17134
rect 13820 17070 13872 17076
rect 13832 16658 13860 17070
rect 14384 16980 14412 19230
rect 14462 19200 14518 20000
rect 14922 19200 14978 20000
rect 15290 19200 15346 20000
rect 15750 19200 15806 20000
rect 16118 19200 16174 20000
rect 16578 19200 16634 20000
rect 16946 19200 17002 20000
rect 14476 17184 14504 19200
rect 14936 17354 14964 19200
rect 14752 17326 14964 17354
rect 14476 17156 14596 17184
rect 14384 16952 14504 16980
rect 14068 16892 14376 16912
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16816 14376 16836
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13728 15632 13780 15638
rect 13728 15574 13780 15580
rect 13636 15564 13688 15570
rect 13636 15506 13688 15512
rect 13636 15360 13688 15366
rect 13636 15302 13688 15308
rect 13648 12646 13676 15302
rect 13740 14958 13768 15574
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13740 14550 13768 14894
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13740 14346 13768 14486
rect 13832 14414 13860 16594
rect 13910 16008 13966 16017
rect 13910 15943 13912 15952
rect 13964 15943 13966 15952
rect 13912 15914 13964 15920
rect 14068 15804 14376 15824
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15728 14376 15748
rect 14476 15586 14504 16952
rect 14568 16250 14596 17156
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14384 15558 14504 15586
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13924 14521 13952 14962
rect 14200 14929 14228 15438
rect 14384 15026 14412 15558
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14186 14920 14242 14929
rect 14186 14855 14242 14864
rect 14068 14716 14376 14736
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14640 14376 14660
rect 13910 14512 13966 14521
rect 13910 14447 13966 14456
rect 13820 14408 13872 14414
rect 13820 14350 13872 14356
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13740 14074 13768 14282
rect 13728 14068 13780 14074
rect 13728 14010 13780 14016
rect 13832 13530 13860 14350
rect 14004 14000 14056 14006
rect 14004 13942 14056 13948
rect 13912 13864 13964 13870
rect 13910 13832 13912 13841
rect 13964 13832 13966 13841
rect 13910 13767 13966 13776
rect 14016 13716 14044 13942
rect 13924 13688 14044 13716
rect 13924 13530 13952 13688
rect 14068 13628 14376 13648
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13552 14376 13572
rect 13820 13524 13872 13530
rect 13820 13466 13872 13472
rect 13912 13524 13964 13530
rect 13912 13466 13964 13472
rect 14280 13456 14332 13462
rect 14280 13398 14332 13404
rect 14370 13424 14426 13433
rect 14096 13320 14148 13326
rect 13910 13288 13966 13297
rect 14096 13262 14148 13268
rect 13910 13223 13912 13232
rect 13964 13223 13966 13232
rect 13912 13194 13964 13200
rect 14108 12986 14136 13262
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14096 12980 14148 12986
rect 14096 12922 14148 12928
rect 14200 12889 14228 13126
rect 13726 12880 13782 12889
rect 14186 12880 14242 12889
rect 13726 12815 13782 12824
rect 13912 12844 13964 12850
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13636 12300 13688 12306
rect 13636 12242 13688 12248
rect 13544 11348 13596 11354
rect 13544 11290 13596 11296
rect 13648 11218 13676 12242
rect 13740 11694 13768 12815
rect 14186 12815 14242 12824
rect 13912 12786 13964 12792
rect 13820 12776 13872 12782
rect 13820 12718 13872 12724
rect 13832 12481 13860 12718
rect 13818 12472 13874 12481
rect 13818 12407 13874 12416
rect 13728 11688 13780 11694
rect 13728 11630 13780 11636
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13464 10062 13492 11154
rect 13832 10674 13860 11154
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13452 9920 13504 9926
rect 13452 9862 13504 9868
rect 13544 9920 13596 9926
rect 13544 9862 13596 9868
rect 13464 9722 13492 9862
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13450 9616 13506 9625
rect 13450 9551 13452 9560
rect 13504 9551 13506 9560
rect 13452 9522 13504 9528
rect 13358 9480 13414 9489
rect 13358 9415 13414 9424
rect 13372 8974 13400 9415
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13450 8664 13506 8673
rect 13556 8634 13584 9862
rect 13832 9518 13860 10610
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13728 9444 13780 9450
rect 13648 9404 13728 9432
rect 13450 8599 13506 8608
rect 13544 8628 13596 8634
rect 13464 8498 13492 8599
rect 13544 8570 13596 8576
rect 13452 8492 13504 8498
rect 13452 8434 13504 8440
rect 13648 8106 13676 9404
rect 13728 9386 13780 9392
rect 13728 8968 13780 8974
rect 13728 8910 13780 8916
rect 13464 8078 13676 8106
rect 13360 7744 13412 7750
rect 13360 7686 13412 7692
rect 13372 6798 13400 7686
rect 13360 6792 13412 6798
rect 13360 6734 13412 6740
rect 13360 6656 13412 6662
rect 13360 6598 13412 6604
rect 13266 2408 13322 2417
rect 13266 2343 13322 2352
rect 13372 1902 13400 6598
rect 13464 2774 13492 8078
rect 13740 8004 13768 8910
rect 13832 8838 13860 9454
rect 13820 8832 13872 8838
rect 13820 8774 13872 8780
rect 13832 8566 13860 8774
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 13648 7976 13768 8004
rect 13818 7984 13874 7993
rect 13648 7750 13676 7976
rect 13818 7919 13874 7928
rect 13728 7812 13780 7818
rect 13728 7754 13780 7760
rect 13636 7744 13688 7750
rect 13556 7704 13636 7732
rect 13556 5914 13584 7704
rect 13636 7686 13688 7692
rect 13740 6934 13768 7754
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13832 6780 13860 7919
rect 13924 7546 13952 12786
rect 14292 12782 14320 13398
rect 14370 13359 14372 13368
rect 14424 13359 14426 13368
rect 14372 13330 14424 13336
rect 14280 12776 14332 12782
rect 14280 12718 14332 12724
rect 14068 12540 14376 12560
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12464 14376 12484
rect 14476 12434 14504 15438
rect 14648 15020 14700 15026
rect 14648 14962 14700 14968
rect 14556 14952 14608 14958
rect 14556 14894 14608 14900
rect 14568 13190 14596 14894
rect 14556 13184 14608 13190
rect 14554 13152 14556 13161
rect 14608 13152 14610 13161
rect 14554 13087 14610 13096
rect 14660 12696 14688 14962
rect 14752 14958 14780 17326
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14740 14952 14792 14958
rect 14740 14894 14792 14900
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 14752 12986 14780 14758
rect 14844 12986 14872 17138
rect 15014 15600 15070 15609
rect 14924 15564 14976 15570
rect 15014 15535 15070 15544
rect 14924 15506 14976 15512
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14832 12980 14884 12986
rect 14832 12922 14884 12928
rect 14936 12866 14964 15506
rect 15028 15502 15056 15535
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15106 15056 15162 15065
rect 15028 13818 15056 15030
rect 15106 14991 15108 15000
rect 15160 14991 15162 15000
rect 15108 14962 15160 14968
rect 15108 14884 15160 14890
rect 15108 14826 15160 14832
rect 15120 14550 15148 14826
rect 15108 14544 15160 14550
rect 15108 14486 15160 14492
rect 15028 13790 15148 13818
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14384 12406 14504 12434
rect 14568 12668 14688 12696
rect 14752 12838 14964 12866
rect 15028 12850 15056 13670
rect 15120 13025 15148 13790
rect 15106 13016 15162 13025
rect 15106 12951 15162 12960
rect 15016 12844 15068 12850
rect 14094 12336 14150 12345
rect 14094 12271 14096 12280
rect 14148 12271 14150 12280
rect 14096 12242 14148 12248
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14108 11898 14136 12038
rect 14096 11892 14148 11898
rect 14096 11834 14148 11840
rect 14108 11665 14136 11834
rect 14384 11778 14412 12406
rect 14568 12288 14596 12668
rect 14752 12594 14780 12838
rect 15016 12786 15068 12792
rect 15108 12844 15160 12850
rect 15108 12786 15160 12792
rect 14830 12744 14886 12753
rect 14830 12679 14886 12688
rect 14476 12260 14596 12288
rect 14660 12566 14780 12594
rect 14476 11898 14504 12260
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14384 11750 14596 11778
rect 14660 11762 14688 12566
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14752 11898 14780 12174
rect 14844 11898 14872 12679
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14832 11892 14884 11898
rect 14832 11834 14884 11840
rect 14464 11688 14516 11694
rect 14094 11656 14150 11665
rect 14464 11630 14516 11636
rect 14094 11591 14150 11600
rect 14068 11452 14376 11472
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11376 14376 11396
rect 14476 10849 14504 11630
rect 14568 11218 14596 11750
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14556 11212 14608 11218
rect 14556 11154 14608 11160
rect 14556 11008 14608 11014
rect 14556 10950 14608 10956
rect 14462 10840 14518 10849
rect 14462 10775 14518 10784
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14068 10364 14376 10384
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10288 14376 10308
rect 14476 10062 14504 10474
rect 14568 10130 14596 10950
rect 14752 10554 14780 11834
rect 15028 10810 15056 12582
rect 15120 12170 15148 12786
rect 15108 12164 15160 12170
rect 15108 12106 15160 12112
rect 15120 12073 15148 12106
rect 15106 12064 15162 12073
rect 15106 11999 15162 12008
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 14844 10606 14872 10746
rect 15016 10668 15068 10674
rect 15016 10610 15068 10616
rect 14660 10526 14780 10554
rect 14832 10600 14884 10606
rect 14832 10542 14884 10548
rect 14556 10124 14608 10130
rect 14556 10066 14608 10072
rect 14464 10056 14516 10062
rect 14464 9998 14516 10004
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9654 14136 9862
rect 14096 9648 14148 9654
rect 14096 9590 14148 9596
rect 14464 9648 14516 9654
rect 14464 9590 14516 9596
rect 14280 9512 14332 9518
rect 14278 9480 14280 9489
rect 14332 9480 14334 9489
rect 14278 9415 14334 9424
rect 14476 9382 14504 9590
rect 14556 9512 14608 9518
rect 14556 9454 14608 9460
rect 14464 9376 14516 9382
rect 14464 9318 14516 9324
rect 14068 9276 14376 9296
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9200 14376 9220
rect 14568 8906 14596 9454
rect 14660 9110 14688 10526
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10198 14780 10406
rect 14740 10192 14792 10198
rect 14740 10134 14792 10140
rect 14844 10010 14872 10542
rect 15028 10130 15056 10610
rect 15016 10124 15068 10130
rect 15016 10066 15068 10072
rect 14752 9982 14872 10010
rect 14648 9104 14700 9110
rect 14648 9046 14700 9052
rect 14648 8968 14700 8974
rect 14752 8945 14780 9982
rect 14830 9888 14886 9897
rect 14830 9823 14886 9832
rect 14844 9586 14872 9823
rect 14832 9580 14884 9586
rect 14832 9522 14884 9528
rect 14648 8910 14700 8916
rect 14738 8936 14794 8945
rect 14556 8900 14608 8906
rect 14556 8842 14608 8848
rect 14372 8832 14424 8838
rect 14372 8774 14424 8780
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14384 8634 14412 8774
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14068 8188 14376 8208
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8112 14376 8132
rect 14280 8016 14332 8022
rect 14280 7958 14332 7964
rect 14370 7984 14426 7993
rect 13912 7540 13964 7546
rect 13912 7482 13964 7488
rect 13912 7336 13964 7342
rect 13912 7278 13964 7284
rect 13740 6752 13860 6780
rect 13636 6724 13688 6730
rect 13636 6666 13688 6672
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13542 5808 13598 5817
rect 13542 5743 13544 5752
rect 13596 5743 13598 5752
rect 13544 5714 13596 5720
rect 13556 5166 13584 5714
rect 13544 5160 13596 5166
rect 13544 5102 13596 5108
rect 13556 3738 13584 5102
rect 13544 3732 13596 3738
rect 13544 3674 13596 3680
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 13556 2961 13584 3470
rect 13542 2952 13598 2961
rect 13542 2887 13598 2896
rect 13464 2746 13584 2774
rect 13556 2378 13584 2746
rect 13544 2372 13596 2378
rect 13544 2314 13596 2320
rect 13544 2100 13596 2106
rect 13544 2042 13596 2048
rect 13360 1896 13412 1902
rect 13360 1838 13412 1844
rect 13556 800 13584 2042
rect 13648 2009 13676 6666
rect 13740 6390 13768 6752
rect 13728 6384 13780 6390
rect 13728 6326 13780 6332
rect 13820 6248 13872 6254
rect 13740 6196 13820 6202
rect 13740 6190 13872 6196
rect 13740 6174 13860 6190
rect 13740 4826 13768 6174
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 4826 13860 6054
rect 13924 5642 13952 7278
rect 14292 7274 14320 7958
rect 14370 7919 14426 7928
rect 14384 7886 14412 7919
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14372 7472 14424 7478
rect 14370 7440 14372 7449
rect 14424 7440 14426 7449
rect 14370 7375 14426 7384
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 14068 7100 14376 7120
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7024 14376 7044
rect 14280 6792 14332 6798
rect 14476 6746 14504 8774
rect 14568 7954 14596 8842
rect 14556 7948 14608 7954
rect 14556 7890 14608 7896
rect 14554 7848 14610 7857
rect 14554 7783 14610 7792
rect 14568 7546 14596 7783
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 14556 7268 14608 7274
rect 14556 7210 14608 7216
rect 14280 6734 14332 6740
rect 14292 6458 14320 6734
rect 14384 6718 14504 6746
rect 14568 6730 14596 7210
rect 14556 6724 14608 6730
rect 14280 6452 14332 6458
rect 14280 6394 14332 6400
rect 14384 6202 14412 6718
rect 14556 6666 14608 6672
rect 14568 6458 14596 6666
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 14384 6174 14596 6202
rect 14464 6112 14516 6118
rect 14464 6054 14516 6060
rect 14068 6012 14376 6032
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5936 14376 5956
rect 14278 5672 14334 5681
rect 13912 5636 13964 5642
rect 14278 5607 14334 5616
rect 13912 5578 13964 5584
rect 14292 5574 14320 5607
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13912 5364 13964 5370
rect 13912 5306 13964 5312
rect 13728 4820 13780 4826
rect 13728 4762 13780 4768
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 4282 13860 4558
rect 13820 4276 13872 4282
rect 13820 4218 13872 4224
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13740 3126 13768 4082
rect 13832 3602 13860 4082
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 13728 3120 13780 3126
rect 13728 3062 13780 3068
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 13726 2952 13782 2961
rect 13726 2887 13782 2896
rect 13740 2650 13768 2887
rect 13728 2644 13780 2650
rect 13728 2586 13780 2592
rect 13740 2310 13768 2586
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13832 2258 13860 2994
rect 13924 2446 13952 5306
rect 14068 4924 14376 4944
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4848 14376 4868
rect 14476 4554 14504 6054
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14476 4010 14504 4490
rect 14568 4214 14596 6174
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14464 4004 14516 4010
rect 14464 3946 14516 3952
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14068 3836 14376 3856
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3760 14376 3780
rect 14464 3596 14516 3602
rect 14464 3538 14516 3544
rect 14096 3528 14148 3534
rect 14094 3496 14096 3505
rect 14148 3496 14150 3505
rect 14094 3431 14150 3440
rect 14068 2748 14376 2768
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2672 14376 2692
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14188 2304 14240 2310
rect 13832 2230 14044 2258
rect 14188 2246 14240 2252
rect 13634 2000 13690 2009
rect 13634 1935 13690 1944
rect 14016 800 14044 2230
rect 14200 2038 14228 2246
rect 14188 2032 14240 2038
rect 14188 1974 14240 1980
rect 14476 800 14504 3538
rect 14568 2446 14596 3878
rect 14660 3602 14688 8910
rect 14738 8871 14794 8880
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14752 5250 14780 8774
rect 14844 7342 14872 9522
rect 14924 9376 14976 9382
rect 14922 9344 14924 9353
rect 14976 9344 14978 9353
rect 14922 9279 14978 9288
rect 14924 9104 14976 9110
rect 14924 9046 14976 9052
rect 14936 8090 14964 9046
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14924 8084 14976 8090
rect 14924 8026 14976 8032
rect 14924 7744 14976 7750
rect 14924 7686 14976 7692
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14936 6361 14964 7686
rect 14922 6352 14978 6361
rect 14832 6316 14884 6322
rect 14922 6287 14978 6296
rect 14832 6258 14884 6264
rect 14844 5574 14872 6258
rect 14924 6248 14976 6254
rect 14924 6190 14976 6196
rect 14936 5914 14964 6190
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14752 5222 14872 5250
rect 14740 5092 14792 5098
rect 14740 5034 14792 5040
rect 14752 4826 14780 5034
rect 14740 4820 14792 4826
rect 14740 4762 14792 4768
rect 14738 4720 14794 4729
rect 14738 4655 14794 4664
rect 14648 3596 14700 3602
rect 14648 3538 14700 3544
rect 14752 3058 14780 4655
rect 14844 4146 14872 5222
rect 14832 4140 14884 4146
rect 14832 4082 14884 4088
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14830 2680 14886 2689
rect 14830 2615 14886 2624
rect 14844 2446 14872 2615
rect 14556 2440 14608 2446
rect 14556 2382 14608 2388
rect 14832 2440 14884 2446
rect 14832 2382 14884 2388
rect 14568 2106 14596 2382
rect 14936 2258 14964 3470
rect 15028 2582 15056 8978
rect 15120 5370 15148 11698
rect 15212 11150 15240 15098
rect 15304 15094 15332 19200
rect 15658 17912 15714 17921
rect 15658 17847 15714 17856
rect 15384 16992 15436 16998
rect 15384 16934 15436 16940
rect 15396 15706 15424 16934
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15384 15700 15436 15706
rect 15384 15642 15436 15648
rect 15292 15088 15344 15094
rect 15292 15030 15344 15036
rect 15290 14920 15346 14929
rect 15290 14855 15346 14864
rect 15304 14346 15332 14855
rect 15292 14340 15344 14346
rect 15292 14282 15344 14288
rect 15304 13462 15332 14282
rect 15384 14272 15436 14278
rect 15384 14214 15436 14220
rect 15488 14226 15516 16390
rect 15672 16182 15700 17847
rect 15764 17270 15792 19200
rect 15752 17264 15804 17270
rect 15752 17206 15804 17212
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15660 16176 15712 16182
rect 15660 16118 15712 16124
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15580 15162 15608 15982
rect 15658 15464 15714 15473
rect 15658 15399 15660 15408
rect 15712 15399 15714 15408
rect 15660 15370 15712 15376
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15856 14890 15884 17002
rect 16028 16516 16080 16522
rect 16028 16458 16080 16464
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15292 13456 15344 13462
rect 15292 13398 15344 13404
rect 15292 12708 15344 12714
rect 15292 12650 15344 12656
rect 15304 12238 15332 12650
rect 15292 12232 15344 12238
rect 15292 12174 15344 12180
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15200 11144 15252 11150
rect 15200 11086 15252 11092
rect 15212 10062 15240 11086
rect 15304 11014 15332 12038
rect 15396 11830 15424 14214
rect 15488 14198 15608 14226
rect 15476 13864 15528 13870
rect 15476 13806 15528 13812
rect 15384 11824 15436 11830
rect 15384 11766 15436 11772
rect 15384 11688 15436 11694
rect 15384 11630 15436 11636
rect 15396 11354 15424 11630
rect 15488 11354 15516 13806
rect 15580 13394 15608 14198
rect 15752 13864 15804 13870
rect 15752 13806 15804 13812
rect 15568 13388 15620 13394
rect 15568 13330 15620 13336
rect 15580 12850 15608 13330
rect 15660 13252 15712 13258
rect 15660 13194 15712 13200
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 15672 12442 15700 13194
rect 15660 12436 15712 12442
rect 15660 12378 15712 12384
rect 15764 11898 15792 13806
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15384 11348 15436 11354
rect 15384 11290 15436 11296
rect 15476 11348 15528 11354
rect 15476 11290 15528 11296
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15292 11008 15344 11014
rect 15292 10950 15344 10956
rect 15290 10840 15346 10849
rect 15290 10775 15346 10784
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15304 8634 15332 10775
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15292 7812 15344 7818
rect 15292 7754 15344 7760
rect 15200 7336 15252 7342
rect 15200 7278 15252 7284
rect 15212 6730 15240 7278
rect 15304 7002 15332 7754
rect 15292 6996 15344 7002
rect 15292 6938 15344 6944
rect 15396 6934 15424 11018
rect 15568 9920 15620 9926
rect 15566 9888 15568 9897
rect 15620 9888 15622 9897
rect 15566 9823 15622 9832
rect 15856 9602 15884 14826
rect 15948 11286 15976 15438
rect 16040 12306 16068 16458
rect 16132 15502 16160 19200
rect 16592 16250 16620 19200
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 16960 14618 16988 19200
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16118 13968 16174 13977
rect 16118 13903 16174 13912
rect 16028 12300 16080 12306
rect 16028 12242 16080 12248
rect 16132 11694 16160 13903
rect 16304 12776 16356 12782
rect 16304 12718 16356 12724
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 16120 11552 16172 11558
rect 16120 11494 16172 11500
rect 15936 11280 15988 11286
rect 15936 11222 15988 11228
rect 15488 9574 15884 9602
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15488 6798 15516 9574
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15752 8832 15804 8838
rect 15752 8774 15804 8780
rect 15660 8288 15712 8294
rect 15660 8230 15712 8236
rect 15568 7744 15620 7750
rect 15568 7686 15620 7692
rect 15476 6792 15528 6798
rect 15476 6734 15528 6740
rect 15580 6730 15608 7686
rect 15672 7410 15700 8230
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 15568 6724 15620 6730
rect 15568 6666 15620 6672
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15212 2774 15240 6666
rect 15384 6656 15436 6662
rect 15384 6598 15436 6604
rect 15292 6452 15344 6458
rect 15292 6394 15344 6400
rect 15304 5710 15332 6394
rect 15396 6322 15424 6598
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15384 6316 15436 6322
rect 15384 6258 15436 6264
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15292 5704 15344 5710
rect 15292 5646 15344 5652
rect 15292 5568 15344 5574
rect 15292 5510 15344 5516
rect 15304 3602 15332 5510
rect 15396 4146 15424 5782
rect 15488 4282 15516 6326
rect 15568 6112 15620 6118
rect 15568 6054 15620 6060
rect 15580 5953 15608 6054
rect 15566 5944 15622 5953
rect 15566 5879 15622 5888
rect 15568 5772 15620 5778
rect 15568 5714 15620 5720
rect 15476 4276 15528 4282
rect 15476 4218 15528 4224
rect 15384 4140 15436 4146
rect 15384 4082 15436 4088
rect 15580 4078 15608 5714
rect 15672 5302 15700 7346
rect 15660 5296 15712 5302
rect 15660 5238 15712 5244
rect 15764 4690 15792 8774
rect 15752 4684 15804 4690
rect 15752 4626 15804 4632
rect 15660 4548 15712 4554
rect 15660 4490 15712 4496
rect 15568 4072 15620 4078
rect 15568 4014 15620 4020
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15580 3194 15608 4014
rect 15672 3641 15700 4490
rect 15658 3632 15714 3641
rect 15658 3567 15714 3576
rect 15568 3188 15620 3194
rect 15568 3130 15620 3136
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15212 2746 15332 2774
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 14844 2230 14964 2258
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14844 800 14872 2230
rect 15304 800 15332 2746
rect 15488 2514 15516 2994
rect 15764 2774 15792 4626
rect 15856 3942 15884 9318
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 15936 8900 15988 8906
rect 15936 8842 15988 8848
rect 15844 3936 15896 3942
rect 15844 3878 15896 3884
rect 15948 3534 15976 8842
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16040 2990 16068 8910
rect 16132 7206 16160 11494
rect 16212 7812 16264 7818
rect 16212 7754 16264 7760
rect 16120 7200 16172 7206
rect 16120 7142 16172 7148
rect 16120 6724 16172 6730
rect 16120 6666 16172 6672
rect 16028 2984 16080 2990
rect 16028 2926 16080 2932
rect 15672 2746 15792 2774
rect 15476 2508 15528 2514
rect 15476 2450 15528 2456
rect 15672 800 15700 2746
rect 16132 800 16160 6666
rect 16224 2922 16252 7754
rect 16316 7546 16344 12718
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16396 8628 16448 8634
rect 16396 8570 16448 8576
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16316 5234 16344 7482
rect 16304 5228 16356 5234
rect 16304 5170 16356 5176
rect 16408 4554 16436 8570
rect 16500 5710 16528 10950
rect 16580 7200 16632 7206
rect 16580 7142 16632 7148
rect 16488 5704 16540 5710
rect 16488 5646 16540 5652
rect 16396 4548 16448 4554
rect 16396 4490 16448 4496
rect 16592 4434 16620 7142
rect 16408 4406 16620 4434
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 16408 2310 16436 4406
rect 16488 4004 16540 4010
rect 16488 3946 16540 3952
rect 16396 2304 16448 2310
rect 16396 2246 16448 2252
rect 16500 800 16528 3946
rect 16948 2848 17000 2854
rect 16948 2790 17000 2796
rect 16960 800 16988 2790
rect 8680 734 8892 762
rect 8942 0 8998 800
rect 9402 0 9458 800
rect 9770 0 9826 800
rect 10230 0 10286 800
rect 10690 0 10746 800
rect 11058 0 11114 800
rect 11518 0 11574 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12714 0 12770 800
rect 13174 0 13230 800
rect 13542 0 13598 800
rect 14002 0 14058 800
rect 14462 0 14518 800
rect 14830 0 14886 800
rect 15290 0 15346 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< via2 >>
rect 1858 17584 1914 17640
rect 2778 19080 2834 19136
rect 1490 16668 1492 16688
rect 1492 16668 1544 16688
rect 1544 16668 1546 16688
rect 1490 16632 1546 16668
rect 1490 15680 1546 15736
rect 3330 18536 3386 18592
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 1490 14728 1546 14784
rect 1950 14048 2006 14104
rect 1490 13796 1546 13832
rect 1490 13776 1492 13796
rect 1492 13776 1544 13796
rect 1544 13776 1546 13796
rect 2318 15544 2374 15600
rect 2226 13640 2282 13696
rect 1490 12824 1546 12880
rect 1582 12416 1638 12472
rect 1490 10956 1492 10976
rect 1492 10956 1544 10976
rect 1544 10956 1546 10976
rect 1490 10920 1546 10956
rect 1858 10648 1914 10704
rect 1490 9968 1546 10024
rect 1858 9868 1860 9888
rect 1860 9868 1912 9888
rect 1912 9868 1914 9888
rect 1858 9832 1914 9868
rect 1490 9016 1546 9072
rect 1490 8064 1546 8120
rect 1490 7148 1492 7168
rect 1492 7148 1544 7168
rect 1544 7148 1546 7168
rect 1490 7112 1546 7148
rect 1490 6180 1546 6216
rect 1490 6160 1492 6180
rect 1492 6160 1544 6180
rect 1544 6160 1546 6180
rect 1490 5208 1546 5264
rect 1490 4256 1546 4312
rect 1398 3984 1454 4040
rect 1950 9424 2006 9480
rect 1858 7792 1914 7848
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 3238 13948 3240 13968
rect 3240 13948 3292 13968
rect 3292 13948 3294 13968
rect 3238 13912 3294 13948
rect 3422 13368 3478 13424
rect 3606 15952 3662 16008
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 3974 16632 4030 16688
rect 3790 16516 3846 16552
rect 3790 16496 3792 16516
rect 3792 16496 3844 16516
rect 3844 16496 3846 16516
rect 4066 16088 4122 16144
rect 3606 15700 3662 15736
rect 3606 15680 3608 15700
rect 3608 15680 3660 15700
rect 3660 15680 3662 15700
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2410 12144 2466 12200
rect 2318 11872 2374 11928
rect 2410 10004 2412 10024
rect 2412 10004 2464 10024
rect 2464 10004 2466 10024
rect 2410 9968 2466 10004
rect 3330 12436 3386 12472
rect 3330 12416 3332 12436
rect 3332 12416 3384 12436
rect 3384 12416 3386 12436
rect 3606 12688 3662 12744
rect 3606 12552 3662 12608
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 3882 13912 3938 13968
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4250 15272 4306 15328
rect 4342 14864 4398 14920
rect 4158 14320 4214 14376
rect 3790 12416 3846 12472
rect 4710 15408 4766 15464
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4526 14048 4582 14104
rect 3974 11736 4030 11792
rect 3330 9868 3332 9888
rect 3332 9868 3384 9888
rect 3384 9868 3386 9888
rect 3330 9832 3386 9868
rect 2502 9596 2504 9616
rect 2504 9596 2556 9616
rect 2556 9596 2558 9616
rect 2502 9560 2558 9596
rect 2226 8608 2282 8664
rect 2502 9016 2558 9072
rect 2502 8336 2558 8392
rect 2134 5228 2190 5264
rect 2134 5208 2136 5228
rect 2136 5208 2188 5228
rect 2188 5208 2190 5228
rect 1950 3052 2006 3088
rect 2410 6432 2466 6488
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2594 7384 2650 7440
rect 1950 3032 1952 3052
rect 1952 3032 2004 3052
rect 2004 3032 2006 3052
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 3054 6160 3110 6216
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 3330 6160 3386 6216
rect 4066 10512 4122 10568
rect 3606 6160 3662 6216
rect 3514 5480 3570 5536
rect 3422 5208 3478 5264
rect 3238 4564 3240 4584
rect 3240 4564 3292 4584
rect 3292 4564 3294 4584
rect 3238 4528 3294 4564
rect 3238 3984 3294 4040
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 2778 1400 2834 1456
rect 3882 8880 3938 8936
rect 4158 9016 4214 9072
rect 4158 8628 4214 8664
rect 4158 8608 4160 8628
rect 4160 8608 4212 8628
rect 4212 8608 4214 8628
rect 4066 7520 4122 7576
rect 4066 7384 4122 7440
rect 4710 14340 4766 14376
rect 4710 14320 4712 14340
rect 4712 14320 4764 14340
rect 4764 14320 4766 14340
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 5538 16088 5594 16144
rect 4986 12688 5042 12744
rect 5078 12280 5134 12336
rect 5538 15680 5594 15736
rect 5354 15136 5410 15192
rect 5538 14456 5594 14512
rect 5538 13912 5594 13968
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4710 8880 4766 8936
rect 4434 8744 4490 8800
rect 4986 9288 5042 9344
rect 4434 8336 4490 8392
rect 3514 2760 3570 2816
rect 3422 2352 3478 2408
rect 3698 3304 3754 3360
rect 3882 2896 3938 2952
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 5170 11600 5226 11656
rect 5538 12180 5540 12200
rect 5540 12180 5592 12200
rect 5592 12180 5594 12200
rect 5538 12144 5594 12180
rect 5814 14320 5870 14376
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4986 6180 5042 6216
rect 4986 6160 4988 6180
rect 4988 6160 5040 6180
rect 5040 6160 5042 6180
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 5078 4528 5134 4584
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6734 15408 6790 15464
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 5998 12960 6054 13016
rect 5998 11756 6054 11792
rect 5998 11736 6000 11756
rect 6000 11736 6052 11756
rect 6052 11736 6054 11756
rect 5722 9968 5778 10024
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6734 13232 6790 13288
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6182 9560 6238 9616
rect 5722 9016 5778 9072
rect 6274 9016 6330 9072
rect 7470 15136 7526 15192
rect 8022 14864 8078 14920
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6918 8880 6974 8936
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6090 7248 6146 7304
rect 5630 6604 5632 6624
rect 5632 6604 5684 6624
rect 5684 6604 5686 6624
rect 5630 6568 5686 6604
rect 6182 6196 6184 6216
rect 6184 6196 6236 6216
rect 6236 6196 6238 6216
rect 5354 5752 5410 5808
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 4250 3168 4306 3224
rect 4066 2488 4122 2544
rect 4526 2624 4582 2680
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 5262 3032 5318 3088
rect 6182 6160 6238 6196
rect 6274 5752 6330 5808
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 5722 2624 5778 2680
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 6182 3576 6238 3632
rect 6182 2760 6238 2816
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 7746 12144 7802 12200
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8758 13640 8814 13696
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 9678 17040 9734 17096
rect 10046 15544 10102 15600
rect 9126 14184 9182 14240
rect 9126 14048 9182 14104
rect 9494 14220 9496 14240
rect 9496 14220 9548 14240
rect 9548 14220 9550 14240
rect 9494 14184 9550 14220
rect 9586 14048 9642 14104
rect 8942 12688 8998 12744
rect 9586 13640 9642 13696
rect 9586 13524 9642 13560
rect 9586 13504 9588 13524
rect 9588 13504 9640 13524
rect 9640 13504 9642 13524
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8850 11872 8906 11928
rect 7746 8356 7802 8392
rect 7746 8336 7748 8356
rect 7748 8336 7800 8356
rect 7800 8336 7802 8356
rect 7562 8064 7618 8120
rect 7378 7404 7434 7440
rect 7378 7384 7380 7404
rect 7380 7384 7432 7404
rect 7432 7384 7434 7404
rect 7470 6860 7526 6896
rect 7470 6840 7472 6860
rect 7472 6840 7524 6860
rect 7524 6840 7526 6860
rect 6918 2488 6974 2544
rect 7562 4700 7564 4720
rect 7564 4700 7616 4720
rect 7616 4700 7618 4720
rect 7562 4664 7618 4700
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 9126 11872 9182 11928
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8482 8064 8538 8120
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8206 6840 8262 6896
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 9034 8880 9090 8936
rect 9310 9016 9366 9072
rect 8666 5772 8722 5808
rect 8666 5752 8668 5772
rect 8668 5752 8720 5772
rect 8720 5752 8722 5772
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 7930 3712 7986 3768
rect 8206 4528 8262 4584
rect 7194 2488 7250 2544
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8390 2896 8446 2952
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 9218 6296 9274 6352
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 11058 16904 11114 16960
rect 11058 16532 11060 16552
rect 11060 16532 11112 16552
rect 11112 16532 11114 16552
rect 11058 16496 11114 16532
rect 11058 16088 11114 16144
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 10138 14864 10194 14920
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10322 14476 10378 14512
rect 10322 14456 10324 14476
rect 10324 14456 10376 14476
rect 10376 14456 10378 14476
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10506 13096 10562 13152
rect 11058 15272 11114 15328
rect 11058 14592 11114 14648
rect 11058 14184 11114 14240
rect 11058 14048 11114 14104
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 10966 13096 11022 13152
rect 11518 15308 11520 15328
rect 11520 15308 11572 15328
rect 11572 15308 11574 15328
rect 11518 15272 11574 15308
rect 11426 14456 11482 14512
rect 11242 12824 11298 12880
rect 10966 11500 10968 11520
rect 10968 11500 11020 11520
rect 11020 11500 11022 11520
rect 10966 11464 11022 11500
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 9402 7948 9458 7984
rect 9402 7928 9404 7948
rect 9404 7928 9456 7948
rect 9456 7928 9458 7948
rect 8942 4120 8998 4176
rect 1490 448 1546 504
rect 9034 2644 9090 2680
rect 9034 2624 9036 2644
rect 9036 2624 9088 2644
rect 9088 2624 9090 2644
rect 9218 4684 9274 4720
rect 9218 4664 9220 4684
rect 9220 4664 9272 4684
rect 9272 4664 9274 4684
rect 9862 8880 9918 8936
rect 9586 4140 9642 4176
rect 9586 4120 9588 4140
rect 9588 4120 9640 4140
rect 9640 4120 9642 4140
rect 9218 3440 9274 3496
rect 9586 3440 9642 3496
rect 9402 2488 9458 2544
rect 11702 17212 11704 17232
rect 11704 17212 11756 17232
rect 11756 17212 11758 17232
rect 11702 17176 11758 17212
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 11886 17040 11942 17096
rect 11702 15408 11758 15464
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 10782 9152 10838 9208
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10322 7792 10378 7848
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 11058 7248 11114 7304
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 10046 4120 10102 4176
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 10322 4120 10378 4176
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10322 3612 10324 3632
rect 10324 3612 10376 3632
rect 10376 3612 10378 3632
rect 10322 3576 10378 3612
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 12438 16632 12494 16688
rect 12070 16496 12126 16552
rect 12530 16496 12586 16552
rect 11978 15816 12034 15872
rect 11978 15544 12034 15600
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12622 16088 12678 16144
rect 12438 14900 12440 14920
rect 12440 14900 12492 14920
rect 12492 14900 12494 14920
rect 12438 14864 12494 14900
rect 12162 14728 12218 14784
rect 12990 16360 13046 16416
rect 13174 16360 13230 16416
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12714 14340 12770 14376
rect 12714 14320 12716 14340
rect 12716 14320 12768 14340
rect 12768 14320 12770 14340
rect 12990 14320 13046 14376
rect 12254 13640 12310 13696
rect 12530 13640 12586 13696
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12990 12280 13046 12336
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 11978 11756 12034 11792
rect 11978 11736 11980 11756
rect 11980 11736 12032 11756
rect 12032 11736 12034 11756
rect 12714 11872 12770 11928
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 11886 10648 11942 10704
rect 11334 6976 11390 7032
rect 11334 5072 11390 5128
rect 11242 4800 11298 4856
rect 11242 4664 11298 4720
rect 11334 4020 11336 4040
rect 11336 4020 11388 4040
rect 11388 4020 11390 4040
rect 11334 3984 11390 4020
rect 11150 2896 11206 2952
rect 12530 10104 12586 10160
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12346 9444 12402 9480
rect 12346 9424 12348 9444
rect 12348 9424 12400 9444
rect 12400 9424 12402 9444
rect 11978 7928 12034 7984
rect 11886 6296 11942 6352
rect 11794 5072 11850 5128
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12990 11872 13046 11928
rect 12990 11736 13046 11792
rect 13174 14456 13230 14512
rect 13358 14320 13414 14376
rect 13266 13932 13322 13968
rect 13266 13912 13268 13932
rect 13268 13912 13320 13932
rect 13320 13912 13322 13932
rect 13358 13640 13414 13696
rect 13266 13368 13322 13424
rect 13174 12144 13230 12200
rect 13542 16516 13598 16552
rect 13542 16496 13544 16516
rect 13544 16496 13596 16516
rect 13596 16496 13598 16516
rect 12714 8608 12770 8664
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12346 6316 12402 6352
rect 12346 6296 12348 6316
rect 12348 6296 12400 6316
rect 12400 6296 12402 6316
rect 12990 6840 13046 6896
rect 11886 3476 11888 3496
rect 11888 3476 11940 3496
rect 11940 3476 11942 3496
rect 11886 3440 11942 3476
rect 11978 3304 12034 3360
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 12898 5752 12954 5808
rect 12530 5072 12586 5128
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 13174 8064 13230 8120
rect 13174 6976 13230 7032
rect 12806 5072 12862 5128
rect 12622 3576 12678 3632
rect 12162 3460 12218 3496
rect 12162 3440 12164 3460
rect 12164 3440 12216 3460
rect 12216 3440 12218 3460
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12990 4528 13046 4584
rect 13174 5364 13230 5400
rect 13174 5344 13176 5364
rect 13176 5344 13228 5364
rect 13228 5344 13230 5364
rect 13174 4120 13230 4176
rect 12714 3068 12716 3088
rect 12716 3068 12768 3088
rect 12768 3068 12770 3088
rect 12714 3032 12770 3068
rect 12714 2932 12716 2952
rect 12716 2932 12768 2952
rect 12768 2932 12770 2952
rect 12714 2896 12770 2932
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 12990 2388 12992 2408
rect 12992 2388 13044 2408
rect 13044 2388 13046 2408
rect 12990 2352 13046 2388
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 13910 15972 13966 16008
rect 13910 15952 13912 15972
rect 13912 15952 13964 15972
rect 13964 15952 13966 15972
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14186 14864 14242 14920
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 13910 14456 13966 14512
rect 13910 13812 13912 13832
rect 13912 13812 13964 13832
rect 13964 13812 13966 13832
rect 13910 13776 13966 13812
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 13910 13252 13966 13288
rect 13910 13232 13912 13252
rect 13912 13232 13964 13252
rect 13964 13232 13966 13252
rect 13726 12824 13782 12880
rect 14186 12824 14242 12880
rect 13818 12416 13874 12472
rect 13450 9580 13506 9616
rect 13450 9560 13452 9580
rect 13452 9560 13504 9580
rect 13504 9560 13506 9580
rect 13358 9424 13414 9480
rect 13450 8608 13506 8664
rect 13266 2352 13322 2408
rect 13818 7928 13874 7984
rect 14370 13388 14426 13424
rect 14370 13368 14372 13388
rect 14372 13368 14424 13388
rect 14424 13368 14426 13388
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14554 13132 14556 13152
rect 14556 13132 14608 13152
rect 14608 13132 14610 13152
rect 14554 13096 14610 13132
rect 15014 15544 15070 15600
rect 15106 15020 15162 15056
rect 15106 15000 15108 15020
rect 15108 15000 15160 15020
rect 15160 15000 15162 15020
rect 15106 12960 15162 13016
rect 14094 12300 14150 12336
rect 14094 12280 14096 12300
rect 14096 12280 14148 12300
rect 14148 12280 14150 12300
rect 14830 12688 14886 12744
rect 14094 11600 14150 11656
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14462 10784 14518 10840
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 15106 12008 15162 12064
rect 14278 9460 14280 9480
rect 14280 9460 14332 9480
rect 14332 9460 14334 9480
rect 14278 9424 14334 9460
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 14830 9832 14886 9888
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 13542 5772 13598 5808
rect 13542 5752 13544 5772
rect 13544 5752 13596 5772
rect 13596 5752 13598 5772
rect 13542 2896 13598 2952
rect 14370 7928 14426 7984
rect 14370 7420 14372 7440
rect 14372 7420 14424 7440
rect 14424 7420 14426 7440
rect 14370 7384 14426 7420
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 14554 7792 14610 7848
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 14278 5616 14334 5672
rect 13726 2896 13782 2952
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14094 3476 14096 3496
rect 14096 3476 14148 3496
rect 14148 3476 14150 3496
rect 14094 3440 14150 3476
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 13634 1944 13690 2000
rect 14738 8880 14794 8936
rect 14922 9324 14924 9344
rect 14924 9324 14976 9344
rect 14976 9324 14978 9344
rect 14922 9288 14978 9324
rect 14922 6296 14978 6352
rect 14738 4664 14794 4720
rect 14830 2624 14886 2680
rect 15658 17856 15714 17912
rect 15290 14864 15346 14920
rect 15658 15428 15714 15464
rect 15658 15408 15660 15428
rect 15660 15408 15712 15428
rect 15712 15408 15714 15428
rect 15290 10784 15346 10840
rect 15566 9868 15568 9888
rect 15568 9868 15620 9888
rect 15620 9868 15622 9888
rect 15566 9832 15622 9868
rect 16118 13912 16174 13968
rect 15566 5888 15622 5944
rect 15658 3576 15714 3632
<< metal3 >>
rect 0 19546 800 19576
rect 0 19486 2698 19546
rect 0 19456 800 19486
rect 2638 19138 2698 19486
rect 2773 19138 2839 19141
rect 2638 19136 2839 19138
rect 2638 19080 2778 19136
rect 2834 19080 2839 19136
rect 2638 19078 2839 19080
rect 2773 19075 2839 19078
rect 0 18594 800 18624
rect 3325 18594 3391 18597
rect 0 18592 3391 18594
rect 0 18536 3330 18592
rect 3386 18536 3391 18592
rect 0 18534 3391 18536
rect 0 18504 800 18534
rect 3325 18531 3391 18534
rect 15653 17914 15719 17917
rect 16400 17914 17200 17944
rect 15653 17912 17200 17914
rect 15653 17856 15658 17912
rect 15714 17856 17200 17912
rect 15653 17854 17200 17856
rect 15653 17851 15719 17854
rect 16400 17824 17200 17854
rect 0 17642 800 17672
rect 1853 17642 1919 17645
rect 0 17640 1919 17642
rect 0 17584 1858 17640
rect 1914 17584 1919 17640
rect 0 17582 1919 17584
rect 0 17552 800 17582
rect 1853 17579 1919 17582
rect 4692 17440 5012 17441
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 17375 5012 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 12188 17440 12508 17441
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 17375 12508 17376
rect 11697 17236 11763 17237
rect 11646 17172 11652 17236
rect 11716 17234 11763 17236
rect 11716 17232 11808 17234
rect 11758 17176 11808 17232
rect 11716 17174 11808 17176
rect 11716 17172 11763 17174
rect 11697 17171 11763 17172
rect 9673 17098 9739 17101
rect 11462 17098 11468 17100
rect 9673 17096 11468 17098
rect 9673 17040 9678 17096
rect 9734 17040 11468 17096
rect 9673 17038 11468 17040
rect 9673 17035 9739 17038
rect 11462 17036 11468 17038
rect 11532 17098 11538 17100
rect 11881 17098 11947 17101
rect 11532 17096 11947 17098
rect 11532 17040 11886 17096
rect 11942 17040 11947 17096
rect 11532 17038 11947 17040
rect 11532 17036 11538 17038
rect 11881 17035 11947 17038
rect 11053 16962 11119 16965
rect 12566 16962 12572 16964
rect 11053 16960 12572 16962
rect 11053 16904 11058 16960
rect 11114 16904 12572 16960
rect 11053 16902 12572 16904
rect 11053 16899 11119 16902
rect 12566 16900 12572 16902
rect 12636 16900 12642 16964
rect 2818 16896 3138 16897
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 16831 3138 16832
rect 6566 16896 6886 16897
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 16831 6886 16832
rect 10314 16896 10634 16897
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 16831 10634 16832
rect 14062 16896 14382 16897
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 16831 14382 16832
rect 0 16690 800 16720
rect 1485 16690 1551 16693
rect 0 16688 1551 16690
rect 0 16632 1490 16688
rect 1546 16632 1551 16688
rect 0 16630 1551 16632
rect 0 16600 800 16630
rect 1485 16627 1551 16630
rect 3969 16690 4035 16693
rect 4102 16690 4108 16692
rect 3969 16688 4108 16690
rect 3969 16632 3974 16688
rect 4030 16632 4108 16688
rect 3969 16630 4108 16632
rect 3969 16627 4035 16630
rect 4102 16628 4108 16630
rect 4172 16628 4178 16692
rect 12433 16690 12499 16693
rect 13486 16690 13492 16692
rect 12433 16688 13492 16690
rect 12433 16632 12438 16688
rect 12494 16632 13492 16688
rect 12433 16630 13492 16632
rect 12433 16627 12499 16630
rect 13486 16628 13492 16630
rect 13556 16628 13562 16692
rect 3785 16556 3851 16557
rect 3734 16554 3740 16556
rect 3658 16494 3740 16554
rect 3804 16554 3851 16556
rect 11053 16554 11119 16557
rect 12065 16554 12131 16557
rect 3804 16552 12131 16554
rect 3846 16496 11058 16552
rect 11114 16496 12070 16552
rect 12126 16496 12131 16552
rect 3734 16492 3740 16494
rect 3804 16494 12131 16496
rect 3804 16492 3851 16494
rect 3785 16491 3851 16492
rect 11053 16491 11119 16494
rect 12065 16491 12131 16494
rect 12525 16554 12591 16557
rect 13537 16554 13603 16557
rect 12525 16552 13603 16554
rect 12525 16496 12530 16552
rect 12586 16496 13542 16552
rect 13598 16496 13603 16552
rect 12525 16494 13603 16496
rect 12525 16491 12591 16494
rect 13537 16491 13603 16494
rect 12985 16418 13051 16421
rect 13169 16418 13235 16421
rect 12985 16416 13235 16418
rect 12985 16360 12990 16416
rect 13046 16360 13174 16416
rect 13230 16360 13235 16416
rect 12985 16358 13235 16360
rect 12985 16355 13051 16358
rect 13169 16355 13235 16358
rect 4692 16352 5012 16353
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 16287 5012 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 12188 16352 12508 16353
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 16287 12508 16288
rect 4061 16146 4127 16149
rect 5533 16146 5599 16149
rect 9070 16146 9076 16148
rect 4061 16144 9076 16146
rect 4061 16088 4066 16144
rect 4122 16088 5538 16144
rect 5594 16088 9076 16144
rect 4061 16086 9076 16088
rect 4061 16083 4127 16086
rect 5533 16083 5599 16086
rect 9070 16084 9076 16086
rect 9140 16084 9146 16148
rect 11053 16146 11119 16149
rect 12617 16146 12683 16149
rect 11053 16144 12683 16146
rect 11053 16088 11058 16144
rect 11114 16088 12622 16144
rect 12678 16088 12683 16144
rect 11053 16086 12683 16088
rect 11053 16083 11119 16086
rect 12617 16083 12683 16086
rect 3601 16010 3667 16013
rect 13905 16010 13971 16013
rect 3601 16008 13971 16010
rect 3601 15952 3606 16008
rect 3662 15952 13910 16008
rect 13966 15952 13971 16008
rect 3601 15950 13971 15952
rect 3601 15947 3667 15950
rect 13905 15947 13971 15950
rect 11830 15812 11836 15876
rect 11900 15874 11906 15876
rect 11973 15874 12039 15877
rect 11900 15872 12039 15874
rect 11900 15816 11978 15872
rect 12034 15816 12039 15872
rect 11900 15814 12039 15816
rect 11900 15812 11906 15814
rect 11973 15811 12039 15814
rect 2818 15808 3138 15809
rect 0 15738 800 15768
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 15743 3138 15744
rect 6566 15808 6886 15809
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 15743 6886 15744
rect 10314 15808 10634 15809
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 15743 10634 15744
rect 14062 15808 14382 15809
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 15743 14382 15744
rect 1485 15738 1551 15741
rect 0 15736 1551 15738
rect 0 15680 1490 15736
rect 1546 15680 1551 15736
rect 0 15678 1551 15680
rect 0 15648 800 15678
rect 1485 15675 1551 15678
rect 3601 15738 3667 15741
rect 5533 15738 5599 15741
rect 3601 15736 5599 15738
rect 3601 15680 3606 15736
rect 3662 15680 5538 15736
rect 5594 15680 5599 15736
rect 3601 15678 5599 15680
rect 3601 15675 3667 15678
rect 5533 15675 5599 15678
rect 2313 15602 2379 15605
rect 10041 15602 10107 15605
rect 2313 15600 10107 15602
rect 2313 15544 2318 15600
rect 2374 15544 10046 15600
rect 10102 15544 10107 15600
rect 2313 15542 10107 15544
rect 2313 15539 2379 15542
rect 10041 15539 10107 15542
rect 11973 15602 12039 15605
rect 15009 15602 15075 15605
rect 11973 15600 15075 15602
rect 11973 15544 11978 15600
rect 12034 15544 15014 15600
rect 15070 15544 15075 15600
rect 11973 15542 15075 15544
rect 11973 15539 12039 15542
rect 15009 15539 15075 15542
rect 4705 15466 4771 15469
rect 6729 15466 6795 15469
rect 4705 15464 6795 15466
rect 4705 15408 4710 15464
rect 4766 15408 6734 15464
rect 6790 15408 6795 15464
rect 4705 15406 6795 15408
rect 4705 15403 4771 15406
rect 6729 15403 6795 15406
rect 11697 15466 11763 15469
rect 15653 15466 15719 15469
rect 11697 15464 15719 15466
rect 11697 15408 11702 15464
rect 11758 15408 15658 15464
rect 15714 15408 15719 15464
rect 11697 15406 15719 15408
rect 11697 15403 11763 15406
rect 15653 15403 15719 15406
rect 4245 15330 4311 15333
rect 11053 15332 11119 15333
rect 4470 15330 4476 15332
rect 4245 15328 4476 15330
rect 4245 15272 4250 15328
rect 4306 15272 4476 15328
rect 4245 15270 4476 15272
rect 4245 15267 4311 15270
rect 4470 15268 4476 15270
rect 4540 15268 4546 15332
rect 11053 15328 11100 15332
rect 11164 15330 11170 15332
rect 11053 15272 11058 15328
rect 11053 15268 11100 15272
rect 11164 15270 11210 15330
rect 11164 15268 11170 15270
rect 11278 15268 11284 15332
rect 11348 15330 11354 15332
rect 11513 15330 11579 15333
rect 11348 15328 11579 15330
rect 11348 15272 11518 15328
rect 11574 15272 11579 15328
rect 11348 15270 11579 15272
rect 11348 15268 11354 15270
rect 11053 15267 11119 15268
rect 11513 15267 11579 15270
rect 4692 15264 5012 15265
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 15199 5012 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 12188 15264 12508 15265
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 15199 12508 15200
rect 5349 15194 5415 15197
rect 7465 15194 7531 15197
rect 5349 15192 7531 15194
rect 5349 15136 5354 15192
rect 5410 15136 7470 15192
rect 7526 15136 7531 15192
rect 5349 15134 7531 15136
rect 5349 15131 5415 15134
rect 7465 15131 7531 15134
rect 4102 14996 4108 15060
rect 4172 15058 4178 15060
rect 15101 15058 15167 15061
rect 4172 15056 15167 15058
rect 4172 15000 15106 15056
rect 15162 15000 15167 15056
rect 4172 14998 15167 15000
rect 4172 14996 4178 14998
rect 15101 14995 15167 14998
rect 4337 14922 4403 14925
rect 8017 14922 8083 14925
rect 4337 14920 8083 14922
rect 4337 14864 4342 14920
rect 4398 14864 8022 14920
rect 8078 14864 8083 14920
rect 4337 14862 8083 14864
rect 4337 14859 4403 14862
rect 8017 14859 8083 14862
rect 10133 14922 10199 14925
rect 12433 14922 12499 14925
rect 14181 14922 14247 14925
rect 15285 14922 15351 14925
rect 10133 14920 12220 14922
rect 10133 14864 10138 14920
rect 10194 14864 12220 14920
rect 10133 14862 12220 14864
rect 10133 14859 10199 14862
rect 0 14786 800 14816
rect 12160 14789 12220 14862
rect 12433 14920 15351 14922
rect 12433 14864 12438 14920
rect 12494 14864 14186 14920
rect 14242 14864 15290 14920
rect 15346 14864 15351 14920
rect 12433 14862 15351 14864
rect 12433 14859 12499 14862
rect 14181 14859 14247 14862
rect 15285 14859 15351 14862
rect 1485 14786 1551 14789
rect 0 14784 1551 14786
rect 0 14728 1490 14784
rect 1546 14728 1551 14784
rect 0 14726 1551 14728
rect 0 14696 800 14726
rect 1485 14723 1551 14726
rect 12157 14786 12223 14789
rect 12750 14786 12756 14788
rect 12157 14784 12756 14786
rect 12157 14728 12162 14784
rect 12218 14728 12756 14784
rect 12157 14726 12756 14728
rect 12157 14723 12223 14726
rect 12750 14724 12756 14726
rect 12820 14724 12826 14788
rect 2818 14720 3138 14721
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 14655 3138 14656
rect 6566 14720 6886 14721
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 14655 6886 14656
rect 10314 14720 10634 14721
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 14655 10634 14656
rect 14062 14720 14382 14721
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 14655 14382 14656
rect 11053 14650 11119 14653
rect 11053 14648 13968 14650
rect 11053 14592 11058 14648
rect 11114 14592 13968 14648
rect 11053 14590 13968 14592
rect 11053 14587 11119 14590
rect 13908 14517 13968 14590
rect 5533 14514 5599 14517
rect 8886 14514 8892 14516
rect 5533 14512 8892 14514
rect 5533 14456 5538 14512
rect 5594 14456 8892 14512
rect 5533 14454 8892 14456
rect 5533 14451 5599 14454
rect 8886 14452 8892 14454
rect 8956 14452 8962 14516
rect 10317 14514 10383 14517
rect 11421 14514 11487 14517
rect 13169 14516 13235 14517
rect 13118 14514 13124 14516
rect 10317 14512 11487 14514
rect 10317 14456 10322 14512
rect 10378 14456 11426 14512
rect 11482 14456 11487 14512
rect 10317 14454 11487 14456
rect 13078 14454 13124 14514
rect 13188 14512 13235 14516
rect 13230 14456 13235 14512
rect 10317 14451 10383 14454
rect 11421 14451 11487 14454
rect 13118 14452 13124 14454
rect 13188 14452 13235 14456
rect 13169 14451 13235 14452
rect 13905 14514 13971 14517
rect 14958 14514 14964 14516
rect 13905 14512 14964 14514
rect 13905 14456 13910 14512
rect 13966 14456 14964 14512
rect 13905 14454 14964 14456
rect 13905 14451 13971 14454
rect 14958 14452 14964 14454
rect 15028 14452 15034 14516
rect 4153 14378 4219 14381
rect 4705 14378 4771 14381
rect 4153 14376 4771 14378
rect 4153 14320 4158 14376
rect 4214 14320 4710 14376
rect 4766 14320 4771 14376
rect 4153 14318 4771 14320
rect 4153 14315 4219 14318
rect 4705 14315 4771 14318
rect 5809 14378 5875 14381
rect 12709 14378 12775 14381
rect 5809 14376 12775 14378
rect 5809 14320 5814 14376
rect 5870 14320 12714 14376
rect 12770 14320 12775 14376
rect 5809 14318 12775 14320
rect 5809 14315 5875 14318
rect 12709 14315 12775 14318
rect 12985 14378 13051 14381
rect 13353 14378 13419 14381
rect 12985 14376 13419 14378
rect 12985 14320 12990 14376
rect 13046 14320 13358 14376
rect 13414 14320 13419 14376
rect 12985 14318 13419 14320
rect 12985 14315 13051 14318
rect 13353 14315 13419 14318
rect 9121 14242 9187 14245
rect 9254 14242 9260 14244
rect 9121 14240 9260 14242
rect 9121 14184 9126 14240
rect 9182 14184 9260 14240
rect 9121 14182 9260 14184
rect 9121 14179 9187 14182
rect 9254 14180 9260 14182
rect 9324 14180 9330 14244
rect 9489 14242 9555 14245
rect 11053 14242 11119 14245
rect 9489 14240 11119 14242
rect 9489 14184 9494 14240
rect 9550 14184 11058 14240
rect 11114 14184 11119 14240
rect 9489 14182 11119 14184
rect 9489 14179 9555 14182
rect 11053 14179 11119 14182
rect 4692 14176 5012 14177
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 14111 5012 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 12188 14176 12508 14177
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 14111 12508 14112
rect 1945 14106 2011 14109
rect 4521 14106 4587 14109
rect 1945 14104 4587 14106
rect 1945 14048 1950 14104
rect 2006 14048 4526 14104
rect 4582 14048 4587 14104
rect 1945 14046 4587 14048
rect 1945 14043 2011 14046
rect 4521 14043 4587 14046
rect 9121 14106 9187 14109
rect 9581 14106 9647 14109
rect 9121 14104 9647 14106
rect 9121 14048 9126 14104
rect 9182 14048 9586 14104
rect 9642 14048 9647 14104
rect 9121 14046 9647 14048
rect 9121 14043 9187 14046
rect 9581 14043 9647 14046
rect 11053 14106 11119 14109
rect 11462 14106 11468 14108
rect 11053 14104 11468 14106
rect 11053 14048 11058 14104
rect 11114 14048 11468 14104
rect 11053 14046 11468 14048
rect 11053 14043 11119 14046
rect 11462 14044 11468 14046
rect 11532 14044 11538 14108
rect 3233 13970 3299 13973
rect 3877 13970 3943 13973
rect 5533 13970 5599 13973
rect 13261 13972 13327 13973
rect 13261 13970 13308 13972
rect 3233 13968 5599 13970
rect 3233 13912 3238 13968
rect 3294 13912 3882 13968
rect 3938 13912 5538 13968
rect 5594 13912 5599 13968
rect 3233 13910 5599 13912
rect 13216 13968 13308 13970
rect 13216 13912 13266 13968
rect 13216 13910 13308 13912
rect 3233 13907 3299 13910
rect 3877 13907 3943 13910
rect 5533 13907 5599 13910
rect 13261 13908 13308 13910
rect 13372 13908 13378 13972
rect 16113 13970 16179 13973
rect 16400 13970 17200 14000
rect 16113 13968 17200 13970
rect 16113 13912 16118 13968
rect 16174 13912 17200 13968
rect 16113 13910 17200 13912
rect 13261 13907 13327 13908
rect 16113 13907 16179 13910
rect 16400 13880 17200 13910
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 13905 13834 13971 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 2638 13832 13971 13834
rect 2638 13776 13910 13832
rect 13966 13776 13971 13832
rect 2638 13774 13971 13776
rect 2221 13698 2287 13701
rect 2638 13698 2698 13774
rect 13905 13771 13971 13774
rect 2221 13696 2698 13698
rect 2221 13640 2226 13696
rect 2282 13640 2698 13696
rect 2221 13638 2698 13640
rect 8753 13698 8819 13701
rect 9581 13698 9647 13701
rect 8753 13696 9647 13698
rect 8753 13640 8758 13696
rect 8814 13640 9586 13696
rect 9642 13640 9647 13696
rect 8753 13638 9647 13640
rect 2221 13635 2287 13638
rect 8753 13635 8819 13638
rect 9581 13635 9647 13638
rect 12249 13698 12315 13701
rect 12525 13698 12591 13701
rect 12249 13696 12591 13698
rect 12249 13640 12254 13696
rect 12310 13640 12530 13696
rect 12586 13640 12591 13696
rect 12249 13638 12591 13640
rect 12249 13635 12315 13638
rect 12525 13635 12591 13638
rect 13118 13636 13124 13700
rect 13188 13698 13194 13700
rect 13353 13698 13419 13701
rect 13188 13696 13419 13698
rect 13188 13640 13358 13696
rect 13414 13640 13419 13696
rect 13188 13638 13419 13640
rect 13188 13636 13194 13638
rect 13353 13635 13419 13638
rect 2818 13632 3138 13633
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 13567 3138 13568
rect 6566 13632 6886 13633
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 13567 6886 13568
rect 10314 13632 10634 13633
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 13567 10634 13568
rect 14062 13632 14382 13633
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 13567 14382 13568
rect 9254 13500 9260 13564
rect 9324 13562 9330 13564
rect 9581 13562 9647 13565
rect 9324 13560 9647 13562
rect 9324 13504 9586 13560
rect 9642 13504 9647 13560
rect 9324 13502 9647 13504
rect 9324 13500 9330 13502
rect 9581 13499 9647 13502
rect 3417 13426 3483 13429
rect 13261 13426 13327 13429
rect 14365 13426 14431 13429
rect 3417 13424 11346 13426
rect 3417 13368 3422 13424
rect 3478 13368 11346 13424
rect 3417 13366 11346 13368
rect 3417 13363 3483 13366
rect 6310 13228 6316 13292
rect 6380 13290 6386 13292
rect 6729 13290 6795 13293
rect 11094 13290 11100 13292
rect 6380 13288 11100 13290
rect 6380 13232 6734 13288
rect 6790 13232 11100 13288
rect 6380 13230 11100 13232
rect 6380 13228 6386 13230
rect 6729 13227 6795 13230
rect 11094 13228 11100 13230
rect 11164 13228 11170 13292
rect 11286 13290 11346 13366
rect 13261 13424 14431 13426
rect 13261 13368 13266 13424
rect 13322 13368 14370 13424
rect 14426 13368 14431 13424
rect 13261 13366 14431 13368
rect 13261 13363 13327 13366
rect 14365 13363 14431 13366
rect 13905 13290 13971 13293
rect 11286 13288 13971 13290
rect 11286 13232 13910 13288
rect 13966 13232 13971 13288
rect 11286 13230 13971 13232
rect 13905 13227 13971 13230
rect 8886 13092 8892 13156
rect 8956 13154 8962 13156
rect 10501 13154 10567 13157
rect 8956 13152 10567 13154
rect 8956 13096 10506 13152
rect 10562 13096 10567 13152
rect 8956 13094 10567 13096
rect 8956 13092 8962 13094
rect 10501 13091 10567 13094
rect 10961 13154 11027 13157
rect 14549 13156 14615 13157
rect 11646 13154 11652 13156
rect 10961 13152 11652 13154
rect 10961 13096 10966 13152
rect 11022 13096 11652 13152
rect 10961 13094 11652 13096
rect 10961 13091 11027 13094
rect 11646 13092 11652 13094
rect 11716 13092 11722 13156
rect 14549 13154 14596 13156
rect 14504 13152 14596 13154
rect 14504 13096 14554 13152
rect 14504 13094 14596 13096
rect 14549 13092 14596 13094
rect 14660 13092 14666 13156
rect 14549 13091 14615 13092
rect 4692 13088 5012 13089
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 13023 5012 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 12188 13088 12508 13089
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 13023 12508 13024
rect 5574 12956 5580 13020
rect 5644 13018 5650 13020
rect 5993 13018 6059 13021
rect 5644 13016 6059 13018
rect 5644 12960 5998 13016
rect 6054 12960 6059 13016
rect 5644 12958 6059 12960
rect 5644 12956 5650 12958
rect 5993 12955 6059 12958
rect 9070 12956 9076 13020
rect 9140 13018 9146 13020
rect 9140 12958 12128 13018
rect 9140 12956 9146 12958
rect 0 12882 800 12912
rect 1485 12882 1551 12885
rect 0 12880 1551 12882
rect 0 12824 1490 12880
rect 1546 12824 1551 12880
rect 0 12822 1551 12824
rect 0 12792 800 12822
rect 1485 12819 1551 12822
rect 11094 12820 11100 12884
rect 11164 12882 11170 12884
rect 11237 12882 11303 12885
rect 11164 12880 11303 12882
rect 11164 12824 11242 12880
rect 11298 12824 11303 12880
rect 11164 12822 11303 12824
rect 12068 12882 12128 12958
rect 15101 13016 15167 13021
rect 15101 12960 15106 13016
rect 15162 12960 15167 13016
rect 15101 12955 15167 12960
rect 13721 12882 13787 12885
rect 14181 12882 14247 12885
rect 12068 12880 14247 12882
rect 12068 12824 13726 12880
rect 13782 12824 14186 12880
rect 14242 12824 14247 12880
rect 12068 12822 14247 12824
rect 11164 12820 11170 12822
rect 11237 12819 11303 12822
rect 13721 12819 13787 12822
rect 14181 12819 14247 12822
rect 3601 12746 3667 12749
rect 2270 12744 3667 12746
rect 2270 12688 3606 12744
rect 3662 12688 3667 12744
rect 2270 12686 3667 12688
rect 1577 12474 1643 12477
rect 2270 12476 2330 12686
rect 3601 12683 3667 12686
rect 4981 12746 5047 12749
rect 8937 12746 9003 12749
rect 4981 12744 9003 12746
rect 4981 12688 4986 12744
rect 5042 12688 8942 12744
rect 8998 12688 9003 12744
rect 4981 12686 9003 12688
rect 4981 12683 5047 12686
rect 8937 12683 9003 12686
rect 14825 12746 14891 12749
rect 15104 12746 15164 12955
rect 14825 12744 15164 12746
rect 14825 12688 14830 12744
rect 14886 12688 15164 12744
rect 14825 12686 15164 12688
rect 14825 12683 14891 12686
rect 3601 12610 3667 12613
rect 3734 12610 3740 12612
rect 3601 12608 3740 12610
rect 3601 12552 3606 12608
rect 3662 12552 3740 12608
rect 3601 12550 3740 12552
rect 3601 12547 3667 12550
rect 3734 12548 3740 12550
rect 3804 12548 3810 12612
rect 2818 12544 3138 12545
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 12479 3138 12480
rect 6566 12544 6886 12545
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 12479 6886 12480
rect 10314 12544 10634 12545
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 12479 10634 12480
rect 14062 12544 14382 12545
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 12479 14382 12480
rect 2262 12474 2268 12476
rect 1577 12472 2268 12474
rect 1577 12416 1582 12472
rect 1638 12416 2268 12472
rect 1577 12414 2268 12416
rect 1577 12411 1643 12414
rect 2262 12412 2268 12414
rect 2332 12412 2338 12476
rect 3325 12474 3391 12477
rect 3785 12474 3851 12477
rect 3325 12472 3851 12474
rect 3325 12416 3330 12472
rect 3386 12416 3790 12472
rect 3846 12416 3851 12472
rect 3325 12414 3851 12416
rect 3325 12411 3391 12414
rect 3785 12411 3851 12414
rect 13813 12474 13879 12477
rect 13813 12472 13922 12474
rect 13813 12416 13818 12472
rect 13874 12416 13922 12472
rect 13813 12411 13922 12416
rect 4470 12276 4476 12340
rect 4540 12338 4546 12340
rect 5073 12338 5139 12341
rect 12985 12338 13051 12341
rect 4540 12336 5139 12338
rect 4540 12280 5078 12336
rect 5134 12280 5139 12336
rect 4540 12278 5139 12280
rect 4540 12276 4546 12278
rect 5073 12275 5139 12278
rect 5766 12336 13051 12338
rect 5766 12280 12990 12336
rect 13046 12280 13051 12336
rect 5766 12278 13051 12280
rect 13862 12338 13922 12411
rect 14089 12338 14155 12341
rect 13862 12336 14155 12338
rect 13862 12280 14094 12336
rect 14150 12280 14155 12336
rect 13862 12278 14155 12280
rect 2405 12202 2471 12205
rect 5533 12202 5599 12205
rect 2405 12200 5599 12202
rect 2405 12144 2410 12200
rect 2466 12144 5538 12200
rect 5594 12144 5599 12200
rect 2405 12142 5599 12144
rect 2405 12139 2471 12142
rect 5533 12139 5599 12142
rect 4692 12000 5012 12001
rect 0 11930 800 11960
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 11935 5012 11936
rect 2313 11930 2379 11933
rect 0 11928 2379 11930
rect 0 11872 2318 11928
rect 2374 11872 2379 11928
rect 0 11870 2379 11872
rect 0 11840 800 11870
rect 2313 11867 2379 11870
rect 3969 11794 4035 11797
rect 5766 11794 5826 12278
rect 12985 12275 13051 12278
rect 14089 12275 14155 12278
rect 7414 12140 7420 12204
rect 7484 12202 7490 12204
rect 7741 12202 7807 12205
rect 13169 12202 13235 12205
rect 13854 12202 13860 12204
rect 7484 12200 13048 12202
rect 7484 12144 7746 12200
rect 7802 12144 13048 12200
rect 7484 12142 13048 12144
rect 7484 12140 7490 12142
rect 7741 12139 7807 12142
rect 12988 12066 13048 12142
rect 13169 12200 13860 12202
rect 13169 12144 13174 12200
rect 13230 12144 13860 12200
rect 13169 12142 13860 12144
rect 13169 12139 13235 12142
rect 13854 12140 13860 12142
rect 13924 12140 13930 12204
rect 15101 12066 15167 12069
rect 12988 12064 15167 12066
rect 12988 12008 15106 12064
rect 15162 12008 15167 12064
rect 12988 12006 15167 12008
rect 15101 12003 15167 12006
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 12188 12000 12508 12001
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 11935 12508 11936
rect 8845 11930 8911 11933
rect 9121 11930 9187 11933
rect 8845 11928 9187 11930
rect 8845 11872 8850 11928
rect 8906 11872 9126 11928
rect 9182 11872 9187 11928
rect 8845 11870 9187 11872
rect 8845 11867 8911 11870
rect 9121 11867 9187 11870
rect 12709 11930 12775 11933
rect 12985 11930 13051 11933
rect 12709 11928 13051 11930
rect 12709 11872 12714 11928
rect 12770 11872 12990 11928
rect 13046 11872 13051 11928
rect 12709 11870 13051 11872
rect 12709 11867 12775 11870
rect 12985 11867 13051 11870
rect 3969 11792 5826 11794
rect 3969 11736 3974 11792
rect 4030 11736 5826 11792
rect 3969 11734 5826 11736
rect 5993 11794 6059 11797
rect 11973 11794 12039 11797
rect 5993 11792 12039 11794
rect 5993 11736 5998 11792
rect 6054 11736 11978 11792
rect 12034 11736 12039 11792
rect 5993 11734 12039 11736
rect 3969 11731 4035 11734
rect 5993 11731 6059 11734
rect 11973 11731 12039 11734
rect 12750 11732 12756 11796
rect 12820 11794 12826 11796
rect 12985 11794 13051 11797
rect 12820 11792 13051 11794
rect 12820 11736 12990 11792
rect 13046 11736 13051 11792
rect 12820 11734 13051 11736
rect 12820 11732 12826 11734
rect 12985 11731 13051 11734
rect 5165 11658 5231 11661
rect 5758 11658 5764 11660
rect 5165 11656 5764 11658
rect 5165 11600 5170 11656
rect 5226 11600 5764 11656
rect 5165 11598 5764 11600
rect 5165 11595 5231 11598
rect 5758 11596 5764 11598
rect 5828 11658 5834 11660
rect 6310 11658 6316 11660
rect 5828 11598 6316 11658
rect 5828 11596 5834 11598
rect 6310 11596 6316 11598
rect 6380 11596 6386 11660
rect 14089 11658 14155 11661
rect 14774 11658 14780 11660
rect 14089 11656 14780 11658
rect 14089 11600 14094 11656
rect 14150 11600 14780 11656
rect 14089 11598 14780 11600
rect 14089 11595 14155 11598
rect 14774 11596 14780 11598
rect 14844 11596 14850 11660
rect 10961 11522 11027 11525
rect 11278 11522 11284 11524
rect 10961 11520 11284 11522
rect 10961 11464 10966 11520
rect 11022 11464 11284 11520
rect 10961 11462 11284 11464
rect 10961 11459 11027 11462
rect 11278 11460 11284 11462
rect 11348 11460 11354 11524
rect 2818 11456 3138 11457
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 11391 3138 11392
rect 6566 11456 6886 11457
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 11391 6886 11392
rect 10314 11456 10634 11457
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 11391 10634 11392
rect 14062 11456 14382 11457
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 11391 14382 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 4692 10912 5012 10913
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 10847 5012 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 12188 10912 12508 10913
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 10847 12508 10848
rect 14457 10842 14523 10845
rect 15285 10842 15351 10845
rect 14457 10840 15351 10842
rect 14457 10784 14462 10840
rect 14518 10784 15290 10840
rect 15346 10784 15351 10840
rect 14457 10782 15351 10784
rect 14457 10779 14523 10782
rect 15285 10779 15351 10782
rect 1853 10706 1919 10709
rect 5574 10706 5580 10708
rect 1853 10704 5580 10706
rect 1853 10648 1858 10704
rect 1914 10648 5580 10704
rect 1853 10646 5580 10648
rect 1853 10643 1919 10646
rect 5574 10644 5580 10646
rect 5644 10644 5650 10708
rect 11881 10706 11947 10709
rect 11838 10704 11947 10706
rect 11838 10648 11886 10704
rect 11942 10648 11947 10704
rect 11838 10643 11947 10648
rect 4061 10570 4127 10573
rect 11838 10570 11898 10643
rect 4061 10568 11898 10570
rect 4061 10512 4066 10568
rect 4122 10512 11898 10568
rect 4061 10510 11898 10512
rect 4061 10507 4127 10510
rect 2818 10368 3138 10369
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 10303 3138 10304
rect 6566 10368 6886 10369
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 10303 6886 10304
rect 10314 10368 10634 10369
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 10303 10634 10304
rect 14062 10368 14382 10369
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 10303 14382 10304
rect 12525 10164 12591 10165
rect 12525 10162 12572 10164
rect 12480 10160 12572 10162
rect 12480 10104 12530 10160
rect 12480 10102 12572 10104
rect 12525 10100 12572 10102
rect 12636 10100 12642 10164
rect 12525 10099 12591 10100
rect 0 10026 800 10056
rect 1485 10026 1551 10029
rect 0 10024 1551 10026
rect 0 9968 1490 10024
rect 1546 9968 1551 10024
rect 0 9966 1551 9968
rect 0 9936 800 9966
rect 1485 9963 1551 9966
rect 2405 10026 2471 10029
rect 5717 10026 5783 10029
rect 2405 10024 5783 10026
rect 2405 9968 2410 10024
rect 2466 9968 5722 10024
rect 5778 9968 5783 10024
rect 2405 9966 5783 9968
rect 2405 9963 2471 9966
rect 5717 9963 5783 9966
rect 1526 9828 1532 9892
rect 1596 9890 1602 9892
rect 1853 9890 1919 9893
rect 1596 9888 1919 9890
rect 1596 9832 1858 9888
rect 1914 9832 1919 9888
rect 1596 9830 1919 9832
rect 1596 9828 1602 9830
rect 1853 9827 1919 9830
rect 2262 9828 2268 9892
rect 2332 9890 2338 9892
rect 3325 9890 3391 9893
rect 2332 9888 3391 9890
rect 2332 9832 3330 9888
rect 3386 9832 3391 9888
rect 2332 9830 3391 9832
rect 2332 9828 2338 9830
rect 3325 9827 3391 9830
rect 14825 9890 14891 9893
rect 14958 9890 14964 9892
rect 14825 9888 14964 9890
rect 14825 9832 14830 9888
rect 14886 9832 14964 9888
rect 14825 9830 14964 9832
rect 14825 9827 14891 9830
rect 14958 9828 14964 9830
rect 15028 9828 15034 9892
rect 15561 9890 15627 9893
rect 16400 9890 17200 9920
rect 15561 9888 17200 9890
rect 15561 9832 15566 9888
rect 15622 9832 17200 9888
rect 15561 9830 17200 9832
rect 15561 9827 15627 9830
rect 4692 9824 5012 9825
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 9759 5012 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 12188 9824 12508 9825
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 16400 9800 17200 9830
rect 12188 9759 12508 9760
rect 2497 9618 2563 9621
rect 3366 9618 3372 9620
rect 2497 9616 3372 9618
rect 2497 9560 2502 9616
rect 2558 9560 3372 9616
rect 2497 9558 3372 9560
rect 2497 9555 2563 9558
rect 3366 9556 3372 9558
rect 3436 9556 3442 9620
rect 6177 9618 6243 9621
rect 13445 9618 13511 9621
rect 6177 9616 13511 9618
rect 6177 9560 6182 9616
rect 6238 9560 13450 9616
rect 13506 9560 13511 9616
rect 6177 9558 13511 9560
rect 6177 9555 6243 9558
rect 13445 9555 13511 9558
rect 1945 9482 2011 9485
rect 12341 9482 12407 9485
rect 1945 9480 12407 9482
rect 1945 9424 1950 9480
rect 2006 9424 12346 9480
rect 12402 9424 12407 9480
rect 1945 9422 12407 9424
rect 1945 9419 2011 9422
rect 12341 9419 12407 9422
rect 13353 9482 13419 9485
rect 14273 9482 14339 9485
rect 13353 9480 14339 9482
rect 13353 9424 13358 9480
rect 13414 9424 14278 9480
rect 14334 9424 14339 9480
rect 13353 9422 14339 9424
rect 13353 9419 13419 9422
rect 14273 9419 14339 9422
rect 4981 9346 5047 9349
rect 14917 9348 14983 9349
rect 5206 9346 5212 9348
rect 4981 9344 5212 9346
rect 4981 9288 4986 9344
rect 5042 9288 5212 9344
rect 4981 9286 5212 9288
rect 4981 9283 5047 9286
rect 5206 9284 5212 9286
rect 5276 9284 5282 9348
rect 14917 9346 14964 9348
rect 14872 9344 14964 9346
rect 14872 9288 14922 9344
rect 14872 9286 14964 9288
rect 14917 9284 14964 9286
rect 15028 9284 15034 9348
rect 14917 9283 14983 9284
rect 2818 9280 3138 9281
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 9215 3138 9216
rect 6566 9280 6886 9281
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 9215 6886 9216
rect 10314 9280 10634 9281
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 9215 10634 9216
rect 14062 9280 14382 9281
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 9215 14382 9216
rect 10777 9210 10843 9213
rect 11094 9210 11100 9212
rect 10777 9208 11100 9210
rect 10777 9152 10782 9208
rect 10838 9152 11100 9208
rect 10777 9150 11100 9152
rect 10777 9147 10843 9150
rect 11094 9148 11100 9150
rect 11164 9148 11170 9212
rect 0 9074 800 9104
rect 1485 9074 1551 9077
rect 0 9072 1551 9074
rect 0 9016 1490 9072
rect 1546 9016 1551 9072
rect 0 9014 1551 9016
rect 0 8984 800 9014
rect 1485 9011 1551 9014
rect 2497 9074 2563 9077
rect 4153 9074 4219 9077
rect 5717 9074 5783 9077
rect 6269 9074 6335 9077
rect 2497 9072 2790 9074
rect 2497 9016 2502 9072
rect 2558 9016 2790 9072
rect 2497 9014 2790 9016
rect 2497 9011 2563 9014
rect 2730 8802 2790 9014
rect 4153 9072 6335 9074
rect 4153 9016 4158 9072
rect 4214 9016 5722 9072
rect 5778 9016 6274 9072
rect 6330 9016 6335 9072
rect 4153 9014 6335 9016
rect 4153 9011 4219 9014
rect 5717 9011 5783 9014
rect 6269 9011 6335 9014
rect 9305 9074 9371 9077
rect 14590 9074 14596 9076
rect 9305 9072 14596 9074
rect 9305 9016 9310 9072
rect 9366 9016 14596 9072
rect 9305 9014 14596 9016
rect 9305 9011 9371 9014
rect 14590 9012 14596 9014
rect 14660 9012 14666 9076
rect 3877 8938 3943 8941
rect 4705 8938 4771 8941
rect 6913 8938 6979 8941
rect 3877 8936 6979 8938
rect 3877 8880 3882 8936
rect 3938 8880 4710 8936
rect 4766 8880 6918 8936
rect 6974 8880 6979 8936
rect 3877 8878 6979 8880
rect 3877 8875 3943 8878
rect 4705 8875 4771 8878
rect 6913 8875 6979 8878
rect 8886 8876 8892 8940
rect 8956 8938 8962 8940
rect 9029 8938 9095 8941
rect 8956 8936 9095 8938
rect 8956 8880 9034 8936
rect 9090 8880 9095 8936
rect 8956 8878 9095 8880
rect 8956 8876 8962 8878
rect 9029 8875 9095 8878
rect 9857 8938 9923 8941
rect 14733 8938 14799 8941
rect 9857 8936 14799 8938
rect 9857 8880 9862 8936
rect 9918 8880 14738 8936
rect 14794 8880 14799 8936
rect 9857 8878 14799 8880
rect 9857 8875 9923 8878
rect 14733 8875 14799 8878
rect 4429 8802 4495 8805
rect 2730 8800 4495 8802
rect 2730 8744 4434 8800
rect 4490 8744 4495 8800
rect 2730 8742 4495 8744
rect 4429 8739 4495 8742
rect 4692 8736 5012 8737
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 8671 5012 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 12188 8736 12508 8737
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 8671 12508 8672
rect 2221 8666 2287 8669
rect 4153 8666 4219 8669
rect 2221 8664 4219 8666
rect 2221 8608 2226 8664
rect 2282 8608 4158 8664
rect 4214 8608 4219 8664
rect 2221 8606 4219 8608
rect 2221 8603 2287 8606
rect 4153 8603 4219 8606
rect 12709 8666 12775 8669
rect 13445 8668 13511 8669
rect 13445 8666 13492 8668
rect 12709 8664 13492 8666
rect 12709 8608 12714 8664
rect 12770 8608 13450 8664
rect 12709 8606 13492 8608
rect 12709 8603 12775 8606
rect 13445 8604 13492 8606
rect 13556 8604 13562 8668
rect 13445 8603 13511 8604
rect 8150 8530 8156 8532
rect 4294 8470 8156 8530
rect 2497 8394 2563 8397
rect 4294 8394 4354 8470
rect 8150 8468 8156 8470
rect 8220 8468 8226 8532
rect 2497 8392 4354 8394
rect 2497 8336 2502 8392
rect 2558 8336 4354 8392
rect 2497 8334 4354 8336
rect 4429 8394 4495 8397
rect 7741 8394 7807 8397
rect 4429 8392 7807 8394
rect 4429 8336 4434 8392
rect 4490 8336 7746 8392
rect 7802 8336 7807 8392
rect 4429 8334 7807 8336
rect 2497 8331 2563 8334
rect 4429 8331 4495 8334
rect 7741 8331 7807 8334
rect 2818 8192 3138 8193
rect 0 8122 800 8152
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 8127 3138 8128
rect 6566 8192 6886 8193
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 8127 6886 8128
rect 10314 8192 10634 8193
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 8127 10634 8128
rect 14062 8192 14382 8193
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 8127 14382 8128
rect 1485 8122 1551 8125
rect 0 8120 1551 8122
rect 0 8064 1490 8120
rect 1546 8064 1551 8120
rect 0 8062 1551 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 7557 8122 7623 8125
rect 8477 8122 8543 8125
rect 7557 8120 8543 8122
rect 7557 8064 7562 8120
rect 7618 8064 8482 8120
rect 8538 8064 8543 8120
rect 7557 8062 8543 8064
rect 7557 8059 7623 8062
rect 8477 8059 8543 8062
rect 11094 8060 11100 8124
rect 11164 8122 11170 8124
rect 13169 8122 13235 8125
rect 11164 8120 13235 8122
rect 11164 8064 13174 8120
rect 13230 8064 13235 8120
rect 11164 8062 13235 8064
rect 11164 8060 11170 8062
rect 13169 8059 13235 8062
rect 1526 7924 1532 7988
rect 1596 7986 1602 7988
rect 9397 7986 9463 7989
rect 11973 7986 12039 7989
rect 13813 7988 13879 7989
rect 12566 7986 12572 7988
rect 1596 7984 11898 7986
rect 1596 7928 9402 7984
rect 9458 7928 11898 7984
rect 1596 7926 11898 7928
rect 1596 7924 1602 7926
rect 9397 7923 9463 7926
rect 1853 7850 1919 7853
rect 10317 7850 10383 7853
rect 1853 7848 10383 7850
rect 1853 7792 1858 7848
rect 1914 7792 10322 7848
rect 10378 7792 10383 7848
rect 1853 7790 10383 7792
rect 11838 7850 11898 7926
rect 11973 7984 12572 7986
rect 11973 7928 11978 7984
rect 12034 7928 12572 7984
rect 11973 7926 12572 7928
rect 11973 7923 12039 7926
rect 12566 7924 12572 7926
rect 12636 7924 12642 7988
rect 13813 7986 13860 7988
rect 13732 7984 13860 7986
rect 13924 7986 13930 7988
rect 14365 7986 14431 7989
rect 13924 7984 14431 7986
rect 13732 7928 13818 7984
rect 13924 7928 14370 7984
rect 14426 7928 14431 7984
rect 13732 7926 13860 7928
rect 13813 7924 13860 7926
rect 13924 7926 14431 7928
rect 13924 7924 13930 7926
rect 13813 7923 13879 7924
rect 14365 7923 14431 7926
rect 14549 7852 14615 7853
rect 14549 7850 14596 7852
rect 11838 7848 14596 7850
rect 14660 7850 14666 7852
rect 11838 7792 14554 7848
rect 11838 7790 14596 7792
rect 1853 7787 1919 7790
rect 10317 7787 10383 7790
rect 14549 7788 14596 7790
rect 14660 7790 14742 7850
rect 14660 7788 14666 7790
rect 14549 7787 14615 7788
rect 4692 7648 5012 7649
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 7583 5012 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 12188 7648 12508 7649
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 7583 12508 7584
rect 4061 7580 4127 7581
rect 4061 7576 4108 7580
rect 4172 7578 4178 7580
rect 4061 7520 4066 7576
rect 4061 7516 4108 7520
rect 4172 7518 4218 7578
rect 4172 7516 4178 7518
rect 4061 7515 4127 7516
rect 2589 7442 2655 7445
rect 4061 7442 4127 7445
rect 7373 7444 7439 7445
rect 7373 7442 7420 7444
rect 2589 7440 4127 7442
rect 2589 7384 2594 7440
rect 2650 7384 4066 7440
rect 4122 7384 4127 7440
rect 2589 7382 4127 7384
rect 7328 7440 7420 7442
rect 7328 7384 7378 7440
rect 7328 7382 7420 7384
rect 2589 7379 2655 7382
rect 4061 7379 4127 7382
rect 7373 7380 7420 7382
rect 7484 7380 7490 7444
rect 13302 7380 13308 7444
rect 13372 7442 13378 7444
rect 14365 7442 14431 7445
rect 13372 7440 14431 7442
rect 13372 7384 14370 7440
rect 14426 7384 14431 7440
rect 13372 7382 14431 7384
rect 13372 7380 13378 7382
rect 7373 7379 7439 7380
rect 14365 7379 14431 7382
rect 6085 7306 6151 7309
rect 11053 7306 11119 7309
rect 6085 7304 11119 7306
rect 6085 7248 6090 7304
rect 6146 7248 11058 7304
rect 11114 7248 11119 7304
rect 6085 7246 11119 7248
rect 6085 7243 6151 7246
rect 11053 7243 11119 7246
rect 0 7170 800 7200
rect 1485 7170 1551 7173
rect 0 7168 1551 7170
rect 0 7112 1490 7168
rect 1546 7112 1551 7168
rect 0 7110 1551 7112
rect 0 7080 800 7110
rect 1485 7107 1551 7110
rect 11278 7108 11284 7172
rect 11348 7170 11354 7172
rect 11348 7110 12450 7170
rect 11348 7108 11354 7110
rect 2818 7104 3138 7105
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 7039 3138 7040
rect 6566 7104 6886 7105
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 7039 6886 7040
rect 10314 7104 10634 7105
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 7039 10634 7040
rect 11094 6972 11100 7036
rect 11164 7034 11170 7036
rect 11329 7034 11395 7037
rect 11164 7032 11395 7034
rect 11164 6976 11334 7032
rect 11390 6976 11395 7032
rect 11164 6974 11395 6976
rect 12390 7034 12450 7110
rect 14062 7104 14382 7105
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 7039 14382 7040
rect 13169 7034 13235 7037
rect 12390 7032 13235 7034
rect 12390 6976 13174 7032
rect 13230 6976 13235 7032
rect 12390 6974 13235 6976
rect 11164 6972 11170 6974
rect 11329 6971 11395 6974
rect 13169 6971 13235 6974
rect 5758 6836 5764 6900
rect 5828 6898 5834 6900
rect 7465 6898 7531 6901
rect 5828 6896 7531 6898
rect 5828 6840 7470 6896
rect 7526 6840 7531 6896
rect 5828 6838 7531 6840
rect 5828 6836 5834 6838
rect 7465 6835 7531 6838
rect 8201 6898 8267 6901
rect 12985 6898 13051 6901
rect 8201 6896 13051 6898
rect 8201 6840 8206 6896
rect 8262 6840 12990 6896
rect 13046 6840 13051 6896
rect 8201 6838 13051 6840
rect 8201 6835 8267 6838
rect 12985 6835 13051 6838
rect 5625 6626 5691 6629
rect 5758 6626 5764 6628
rect 5625 6624 5764 6626
rect 5625 6568 5630 6624
rect 5686 6568 5764 6624
rect 5625 6566 5764 6568
rect 5625 6563 5691 6566
rect 5758 6564 5764 6566
rect 5828 6564 5834 6628
rect 4692 6560 5012 6561
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 6495 5012 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 12188 6560 12508 6561
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 6495 12508 6496
rect 2405 6490 2471 6493
rect 2405 6488 2514 6490
rect 2405 6432 2410 6488
rect 2466 6432 2514 6488
rect 2405 6427 2514 6432
rect 2454 6354 2514 6427
rect 9213 6354 9279 6357
rect 11881 6356 11947 6357
rect 11830 6354 11836 6356
rect 2454 6352 9279 6354
rect 2454 6296 9218 6352
rect 9274 6296 9279 6352
rect 2454 6294 9279 6296
rect 11754 6294 11836 6354
rect 11900 6354 11947 6356
rect 12341 6354 12407 6357
rect 11900 6352 12407 6354
rect 11942 6296 12346 6352
rect 12402 6296 12407 6352
rect 9213 6291 9279 6294
rect 11830 6292 11836 6294
rect 11900 6294 12407 6296
rect 11900 6292 11947 6294
rect 11881 6291 11947 6292
rect 12341 6291 12407 6294
rect 12750 6292 12756 6356
rect 12820 6354 12826 6356
rect 14917 6354 14983 6357
rect 12820 6352 14983 6354
rect 12820 6296 14922 6352
rect 14978 6296 14983 6352
rect 12820 6294 14983 6296
rect 12820 6292 12826 6294
rect 14917 6291 14983 6294
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 3049 6218 3115 6221
rect 3325 6218 3391 6221
rect 3049 6216 3391 6218
rect 3049 6160 3054 6216
rect 3110 6160 3330 6216
rect 3386 6160 3391 6216
rect 3049 6158 3391 6160
rect 3049 6155 3115 6158
rect 3325 6155 3391 6158
rect 3601 6216 3667 6221
rect 3601 6160 3606 6216
rect 3662 6160 3667 6216
rect 3601 6155 3667 6160
rect 4981 6218 5047 6221
rect 6177 6218 6243 6221
rect 4981 6216 6243 6218
rect 4981 6160 4986 6216
rect 5042 6160 6182 6216
rect 6238 6160 6243 6216
rect 4981 6158 6243 6160
rect 4981 6155 5047 6158
rect 6177 6155 6243 6158
rect 2818 6016 3138 6017
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 5951 3138 5952
rect 3604 5674 3664 6155
rect 6566 6016 6886 6017
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 5951 6886 5952
rect 10314 6016 10634 6017
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 5951 10634 5952
rect 14062 6016 14382 6017
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 5951 14382 5952
rect 15561 5946 15627 5949
rect 16400 5946 17200 5976
rect 15561 5944 17200 5946
rect 15561 5888 15566 5944
rect 15622 5888 17200 5944
rect 15561 5886 17200 5888
rect 15561 5883 15627 5886
rect 16400 5856 17200 5886
rect 5349 5810 5415 5813
rect 6269 5810 6335 5813
rect 8661 5810 8727 5813
rect 5349 5808 8727 5810
rect 5349 5752 5354 5808
rect 5410 5752 6274 5808
rect 6330 5752 8666 5808
rect 8722 5752 8727 5808
rect 5349 5750 8727 5752
rect 5349 5747 5415 5750
rect 6269 5747 6335 5750
rect 8661 5747 8727 5750
rect 12893 5810 12959 5813
rect 13537 5810 13603 5813
rect 12893 5808 13603 5810
rect 12893 5752 12898 5808
rect 12954 5752 13542 5808
rect 13598 5752 13603 5808
rect 12893 5750 13603 5752
rect 12893 5747 12959 5750
rect 13537 5747 13603 5750
rect 3558 5614 3664 5674
rect 14273 5674 14339 5677
rect 14590 5674 14596 5676
rect 14273 5672 14596 5674
rect 14273 5616 14278 5672
rect 14334 5616 14596 5672
rect 14273 5614 14596 5616
rect 3558 5541 3618 5614
rect 14273 5611 14339 5614
rect 14590 5612 14596 5614
rect 14660 5612 14666 5676
rect 3509 5536 3618 5541
rect 3509 5480 3514 5536
rect 3570 5480 3618 5536
rect 3509 5478 3618 5480
rect 3509 5475 3575 5478
rect 4692 5472 5012 5473
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 5407 5012 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 12188 5472 12508 5473
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 5407 12508 5408
rect 13169 5402 13235 5405
rect 13302 5402 13308 5404
rect 13169 5400 13308 5402
rect 13169 5344 13174 5400
rect 13230 5344 13308 5400
rect 13169 5342 13308 5344
rect 13169 5339 13235 5342
rect 13302 5340 13308 5342
rect 13372 5340 13378 5404
rect 0 5266 800 5296
rect 1485 5266 1551 5269
rect 0 5264 1551 5266
rect 0 5208 1490 5264
rect 1546 5208 1551 5264
rect 0 5206 1551 5208
rect 0 5176 800 5206
rect 1485 5203 1551 5206
rect 2129 5266 2195 5269
rect 2262 5266 2268 5268
rect 2129 5264 2268 5266
rect 2129 5208 2134 5264
rect 2190 5208 2268 5264
rect 2129 5206 2268 5208
rect 2129 5203 2195 5206
rect 2262 5204 2268 5206
rect 2332 5266 2338 5268
rect 3417 5266 3483 5269
rect 11094 5266 11100 5268
rect 2332 5206 2790 5266
rect 2332 5204 2338 5206
rect 2730 5130 2790 5206
rect 3417 5264 11100 5266
rect 3417 5208 3422 5264
rect 3478 5208 11100 5264
rect 3417 5206 11100 5208
rect 3417 5203 3483 5206
rect 11094 5204 11100 5206
rect 11164 5204 11170 5268
rect 11329 5130 11395 5133
rect 11789 5130 11855 5133
rect 2730 5128 11855 5130
rect 2730 5072 11334 5128
rect 11390 5072 11794 5128
rect 11850 5072 11855 5128
rect 2730 5070 11855 5072
rect 11329 5067 11395 5070
rect 11789 5067 11855 5070
rect 12525 5130 12591 5133
rect 12801 5130 12867 5133
rect 12525 5128 12867 5130
rect 12525 5072 12530 5128
rect 12586 5072 12806 5128
rect 12862 5072 12867 5128
rect 12525 5070 12867 5072
rect 12525 5067 12591 5070
rect 12801 5067 12867 5070
rect 2818 4928 3138 4929
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 4863 3138 4864
rect 6566 4928 6886 4929
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 4863 6886 4864
rect 10314 4928 10634 4929
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 4863 10634 4864
rect 14062 4928 14382 4929
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 4863 14382 4864
rect 11237 4858 11303 4861
rect 11237 4856 11530 4858
rect 11237 4800 11242 4856
rect 11298 4800 11530 4856
rect 11237 4798 11530 4800
rect 11237 4795 11303 4798
rect 4102 4660 4108 4724
rect 4172 4722 4178 4724
rect 7557 4722 7623 4725
rect 4172 4720 7623 4722
rect 4172 4664 7562 4720
rect 7618 4664 7623 4720
rect 4172 4662 7623 4664
rect 4172 4660 4178 4662
rect 7557 4659 7623 4662
rect 9213 4722 9279 4725
rect 11237 4722 11303 4725
rect 9213 4720 11303 4722
rect 9213 4664 9218 4720
rect 9274 4664 11242 4720
rect 11298 4664 11303 4720
rect 9213 4662 11303 4664
rect 11470 4722 11530 4798
rect 14733 4722 14799 4725
rect 11470 4720 14799 4722
rect 11470 4664 14738 4720
rect 14794 4664 14799 4720
rect 11470 4662 14799 4664
rect 9213 4659 9279 4662
rect 11237 4659 11303 4662
rect 14733 4659 14799 4662
rect 3233 4586 3299 4589
rect 3366 4586 3372 4588
rect 3233 4584 3372 4586
rect 3233 4528 3238 4584
rect 3294 4528 3372 4584
rect 3233 4526 3372 4528
rect 3233 4523 3299 4526
rect 3366 4524 3372 4526
rect 3436 4524 3442 4588
rect 5073 4586 5139 4589
rect 5206 4586 5212 4588
rect 5073 4584 5212 4586
rect 5073 4528 5078 4584
rect 5134 4528 5212 4584
rect 5073 4526 5212 4528
rect 5073 4523 5139 4526
rect 5206 4524 5212 4526
rect 5276 4524 5282 4588
rect 8201 4586 8267 4589
rect 12985 4586 13051 4589
rect 8201 4584 13051 4586
rect 8201 4528 8206 4584
rect 8262 4528 12990 4584
rect 13046 4528 13051 4584
rect 8201 4526 13051 4528
rect 8201 4523 8267 4526
rect 12985 4523 13051 4526
rect 4692 4384 5012 4385
rect 0 4314 800 4344
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 4319 5012 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 12188 4384 12508 4385
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 4319 12508 4320
rect 1485 4314 1551 4317
rect 0 4312 1551 4314
rect 0 4256 1490 4312
rect 1546 4256 1551 4312
rect 0 4254 1551 4256
rect 0 4224 800 4254
rect 1485 4251 1551 4254
rect 8937 4178 9003 4181
rect 9581 4178 9647 4181
rect 8937 4176 9647 4178
rect 8937 4120 8942 4176
rect 8998 4120 9586 4176
rect 9642 4120 9647 4176
rect 8937 4118 9647 4120
rect 8937 4115 9003 4118
rect 9581 4115 9647 4118
rect 10041 4178 10107 4181
rect 10317 4178 10383 4181
rect 13169 4178 13235 4181
rect 10041 4176 10383 4178
rect 10041 4120 10046 4176
rect 10102 4120 10322 4176
rect 10378 4120 10383 4176
rect 10041 4118 10383 4120
rect 10041 4115 10107 4118
rect 10317 4115 10383 4118
rect 12390 4176 13235 4178
rect 12390 4120 13174 4176
rect 13230 4120 13235 4176
rect 12390 4118 13235 4120
rect 1393 4042 1459 4045
rect 1526 4042 1532 4044
rect 1393 4040 1532 4042
rect 1393 3984 1398 4040
rect 1454 3984 1532 4040
rect 1393 3982 1532 3984
rect 1393 3979 1459 3982
rect 1526 3980 1532 3982
rect 1596 3980 1602 4044
rect 3233 4042 3299 4045
rect 11329 4042 11395 4045
rect 12390 4042 12450 4118
rect 13169 4115 13235 4118
rect 3233 4040 12450 4042
rect 3233 3984 3238 4040
rect 3294 3984 11334 4040
rect 11390 3984 12450 4040
rect 3233 3982 12450 3984
rect 3233 3979 3299 3982
rect 11329 3979 11395 3982
rect 2818 3840 3138 3841
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 3775 3138 3776
rect 6566 3840 6886 3841
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 3775 6886 3776
rect 10314 3840 10634 3841
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10314 3775 10634 3776
rect 14062 3840 14382 3841
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 3775 14382 3776
rect 7925 3770 7991 3773
rect 7925 3768 9690 3770
rect 7925 3712 7930 3768
rect 7986 3712 9690 3768
rect 7925 3710 9690 3712
rect 7925 3707 7991 3710
rect 6177 3634 6243 3637
rect 9630 3634 9690 3710
rect 10317 3634 10383 3637
rect 6177 3632 9506 3634
rect 6177 3576 6182 3632
rect 6238 3576 9506 3632
rect 6177 3574 9506 3576
rect 9630 3632 10383 3634
rect 9630 3576 10322 3632
rect 10378 3576 10383 3632
rect 9630 3574 10383 3576
rect 6177 3571 6243 3574
rect 9213 3498 9279 3501
rect 4478 3496 9279 3498
rect 4478 3440 9218 3496
rect 9274 3440 9279 3496
rect 4478 3438 9279 3440
rect 0 3362 800 3392
rect 3693 3362 3759 3365
rect 0 3360 3759 3362
rect 0 3304 3698 3360
rect 3754 3304 3759 3360
rect 0 3302 3759 3304
rect 0 3272 800 3302
rect 3693 3299 3759 3302
rect 4102 3164 4108 3228
rect 4172 3226 4178 3228
rect 4245 3226 4311 3229
rect 4172 3224 4311 3226
rect 4172 3168 4250 3224
rect 4306 3168 4311 3224
rect 4172 3166 4311 3168
rect 4172 3164 4178 3166
rect 4245 3163 4311 3166
rect 1945 3090 2011 3093
rect 4478 3090 4538 3438
rect 9213 3435 9279 3438
rect 9446 3362 9506 3574
rect 10317 3571 10383 3574
rect 12617 3634 12683 3637
rect 15653 3634 15719 3637
rect 12617 3632 15719 3634
rect 12617 3576 12622 3632
rect 12678 3576 15658 3632
rect 15714 3576 15719 3632
rect 12617 3574 15719 3576
rect 12617 3571 12683 3574
rect 15653 3571 15719 3574
rect 9581 3498 9647 3501
rect 11881 3498 11947 3501
rect 9581 3496 11947 3498
rect 9581 3440 9586 3496
rect 9642 3440 11886 3496
rect 11942 3440 11947 3496
rect 9581 3438 11947 3440
rect 9581 3435 9647 3438
rect 11881 3435 11947 3438
rect 12157 3498 12223 3501
rect 14089 3498 14155 3501
rect 12157 3496 14155 3498
rect 12157 3440 12162 3496
rect 12218 3440 14094 3496
rect 14150 3440 14155 3496
rect 12157 3438 14155 3440
rect 12157 3435 12223 3438
rect 14089 3435 14155 3438
rect 11973 3362 12039 3365
rect 9446 3360 12039 3362
rect 9446 3304 11978 3360
rect 12034 3304 12039 3360
rect 9446 3302 12039 3304
rect 11973 3299 12039 3302
rect 4692 3296 5012 3297
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 3231 5012 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 12188 3296 12508 3297
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 3231 12508 3232
rect 1945 3088 4538 3090
rect 1945 3032 1950 3088
rect 2006 3032 4538 3088
rect 1945 3030 4538 3032
rect 5257 3090 5323 3093
rect 12709 3090 12775 3093
rect 5257 3088 12775 3090
rect 5257 3032 5262 3088
rect 5318 3032 12714 3088
rect 12770 3032 12775 3088
rect 5257 3030 12775 3032
rect 1945 3027 2011 3030
rect 5257 3027 5323 3030
rect 12709 3027 12775 3030
rect 3877 2954 3943 2957
rect 8385 2954 8451 2957
rect 3877 2952 8451 2954
rect 3877 2896 3882 2952
rect 3938 2896 8390 2952
rect 8446 2896 8451 2952
rect 3877 2894 8451 2896
rect 3877 2891 3943 2894
rect 8385 2891 8451 2894
rect 11145 2954 11211 2957
rect 12709 2956 12775 2957
rect 12709 2954 12756 2956
rect 11145 2952 12756 2954
rect 11145 2896 11150 2952
rect 11206 2896 12714 2952
rect 11145 2894 12756 2896
rect 11145 2891 11211 2894
rect 12709 2892 12756 2894
rect 12820 2892 12826 2956
rect 13537 2954 13603 2957
rect 13721 2954 13787 2957
rect 13537 2952 13787 2954
rect 13537 2896 13542 2952
rect 13598 2896 13726 2952
rect 13782 2896 13787 2952
rect 13537 2894 13787 2896
rect 12709 2891 12775 2892
rect 13537 2891 13603 2894
rect 13721 2891 13787 2894
rect 3509 2818 3575 2821
rect 6177 2818 6243 2821
rect 3509 2816 6243 2818
rect 3509 2760 3514 2816
rect 3570 2760 6182 2816
rect 6238 2760 6243 2816
rect 3509 2758 6243 2760
rect 3509 2755 3575 2758
rect 6177 2755 6243 2758
rect 2818 2752 3138 2753
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2687 3138 2688
rect 6566 2752 6886 2753
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2687 6886 2688
rect 10314 2752 10634 2753
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2687 10634 2688
rect 14062 2752 14382 2753
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2687 14382 2688
rect 4521 2682 4587 2685
rect 5717 2682 5783 2685
rect 4521 2680 5783 2682
rect 4521 2624 4526 2680
rect 4582 2624 5722 2680
rect 5778 2624 5783 2680
rect 4521 2622 5783 2624
rect 4521 2619 4587 2622
rect 5717 2619 5783 2622
rect 8150 2620 8156 2684
rect 8220 2682 8226 2684
rect 9029 2682 9095 2685
rect 8220 2680 9095 2682
rect 8220 2624 9034 2680
rect 9090 2624 9095 2680
rect 8220 2622 9095 2624
rect 8220 2620 8226 2622
rect 9029 2619 9095 2622
rect 14825 2682 14891 2685
rect 14958 2682 14964 2684
rect 14825 2680 14964 2682
rect 14825 2624 14830 2680
rect 14886 2624 14964 2680
rect 14825 2622 14964 2624
rect 14825 2619 14891 2622
rect 14958 2620 14964 2622
rect 15028 2620 15034 2684
rect 4061 2546 4127 2549
rect 6913 2546 6979 2549
rect 4061 2544 6979 2546
rect 4061 2488 4066 2544
rect 4122 2488 6918 2544
rect 6974 2488 6979 2544
rect 4061 2486 6979 2488
rect 4061 2483 4127 2486
rect 6913 2483 6979 2486
rect 7189 2546 7255 2549
rect 8886 2546 8892 2548
rect 7189 2544 8892 2546
rect 7189 2488 7194 2544
rect 7250 2488 8892 2544
rect 7189 2486 8892 2488
rect 7189 2483 7255 2486
rect 8886 2484 8892 2486
rect 8956 2546 8962 2548
rect 9397 2546 9463 2549
rect 8956 2544 9463 2546
rect 8956 2488 9402 2544
rect 9458 2488 9463 2544
rect 8956 2486 9463 2488
rect 8956 2484 8962 2486
rect 9397 2483 9463 2486
rect 0 2410 800 2440
rect 3417 2410 3483 2413
rect 0 2408 3483 2410
rect 0 2352 3422 2408
rect 3478 2352 3483 2408
rect 0 2350 3483 2352
rect 0 2320 800 2350
rect 3417 2347 3483 2350
rect 5758 2348 5764 2412
rect 5828 2410 5834 2412
rect 12985 2410 13051 2413
rect 13261 2410 13327 2413
rect 5828 2408 13327 2410
rect 5828 2352 12990 2408
rect 13046 2352 13266 2408
rect 13322 2352 13327 2408
rect 5828 2350 13327 2352
rect 5828 2348 5834 2350
rect 12985 2347 13051 2350
rect 13261 2347 13327 2350
rect 4692 2208 5012 2209
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2143 5012 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 12188 2208 12508 2209
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2143 12508 2144
rect 13629 2002 13695 2005
rect 16400 2002 17200 2032
rect 13629 2000 17200 2002
rect 13629 1944 13634 2000
rect 13690 1944 17200 2000
rect 13629 1942 17200 1944
rect 13629 1939 13695 1942
rect 16400 1912 17200 1942
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 0 506 800 536
rect 1485 506 1551 509
rect 0 504 1551 506
rect 0 448 1490 504
rect 1546 448 1551 504
rect 0 446 1551 448
rect 0 416 800 446
rect 1485 443 1551 446
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 11652 17232 11716 17236
rect 11652 17176 11702 17232
rect 11702 17176 11716 17232
rect 11652 17172 11716 17176
rect 11468 17036 11532 17100
rect 12572 16900 12636 16964
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 4108 16628 4172 16692
rect 13492 16628 13556 16692
rect 3740 16552 3804 16556
rect 3740 16496 3790 16552
rect 3790 16496 3804 16552
rect 3740 16492 3804 16496
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 9076 16084 9140 16148
rect 11836 15812 11900 15876
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 4476 15268 4540 15332
rect 11100 15328 11164 15332
rect 11100 15272 11114 15328
rect 11114 15272 11164 15328
rect 11100 15268 11164 15272
rect 11284 15268 11348 15332
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 4108 14996 4172 15060
rect 12756 14724 12820 14788
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 8892 14452 8956 14516
rect 13124 14512 13188 14516
rect 13124 14456 13174 14512
rect 13174 14456 13188 14512
rect 13124 14452 13188 14456
rect 14964 14452 15028 14516
rect 9260 14180 9324 14244
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 11468 14044 11532 14108
rect 13308 13968 13372 13972
rect 13308 13912 13322 13968
rect 13322 13912 13372 13968
rect 13308 13908 13372 13912
rect 13124 13636 13188 13700
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 9260 13500 9324 13564
rect 6316 13228 6380 13292
rect 11100 13228 11164 13292
rect 8892 13092 8956 13156
rect 11652 13092 11716 13156
rect 14596 13152 14660 13156
rect 14596 13096 14610 13152
rect 14610 13096 14660 13152
rect 14596 13092 14660 13096
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 5580 12956 5644 13020
rect 9076 12956 9140 13020
rect 11100 12820 11164 12884
rect 3740 12548 3804 12612
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 2268 12412 2332 12476
rect 4476 12276 4540 12340
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 7420 12140 7484 12204
rect 13860 12140 13924 12204
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 12756 11732 12820 11796
rect 5764 11596 5828 11660
rect 6316 11596 6380 11660
rect 14780 11596 14844 11660
rect 11284 11460 11348 11524
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 5580 10644 5644 10708
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 12572 10160 12636 10164
rect 12572 10104 12586 10160
rect 12586 10104 12636 10160
rect 12572 10100 12636 10104
rect 1532 9828 1596 9892
rect 2268 9828 2332 9892
rect 14964 9828 15028 9892
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 3372 9556 3436 9620
rect 5212 9284 5276 9348
rect 14964 9344 15028 9348
rect 14964 9288 14978 9344
rect 14978 9288 15028 9344
rect 14964 9284 15028 9288
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 11100 9148 11164 9212
rect 14596 9012 14660 9076
rect 8892 8876 8956 8940
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 13492 8664 13556 8668
rect 13492 8608 13506 8664
rect 13506 8608 13556 8664
rect 13492 8604 13556 8608
rect 8156 8468 8220 8532
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 11100 8060 11164 8124
rect 1532 7924 1596 7988
rect 12572 7924 12636 7988
rect 13860 7984 13924 7988
rect 13860 7928 13874 7984
rect 13874 7928 13924 7984
rect 13860 7924 13924 7928
rect 14596 7848 14660 7852
rect 14596 7792 14610 7848
rect 14610 7792 14660 7848
rect 14596 7788 14660 7792
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 4108 7576 4172 7580
rect 4108 7520 4122 7576
rect 4122 7520 4172 7576
rect 4108 7516 4172 7520
rect 7420 7440 7484 7444
rect 7420 7384 7434 7440
rect 7434 7384 7484 7440
rect 7420 7380 7484 7384
rect 13308 7380 13372 7444
rect 11284 7108 11348 7172
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 11100 6972 11164 7036
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 5764 6836 5828 6900
rect 5764 6564 5828 6628
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 11836 6352 11900 6356
rect 11836 6296 11886 6352
rect 11886 6296 11900 6352
rect 11836 6292 11900 6296
rect 12756 6292 12820 6356
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 14596 5612 14660 5676
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 13308 5340 13372 5404
rect 2268 5204 2332 5268
rect 11100 5204 11164 5268
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 4108 4660 4172 4724
rect 3372 4524 3436 4588
rect 5212 4524 5276 4588
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 1532 3980 1596 4044
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 4108 3164 4172 3228
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 12756 2952 12820 2956
rect 12756 2896 12770 2952
rect 12770 2896 12820 2952
rect 12756 2892 12820 2896
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 8156 2620 8220 2684
rect 14964 2620 15028 2684
rect 8892 2484 8956 2548
rect 5764 2348 5828 2412
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4107 16692 4173 16693
rect 4107 16628 4108 16692
rect 4172 16628 4173 16692
rect 4107 16627 4173 16628
rect 3739 16556 3805 16557
rect 3739 16492 3740 16556
rect 3804 16492 3805 16556
rect 3739 16491 3805 16492
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 3742 12613 3802 16491
rect 4110 15061 4170 16627
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4475 15332 4541 15333
rect 4475 15268 4476 15332
rect 4540 15268 4541 15332
rect 4475 15267 4541 15268
rect 4107 15060 4173 15061
rect 4107 14996 4108 15060
rect 4172 14996 4173 15060
rect 4107 14995 4173 14996
rect 3739 12612 3805 12613
rect 3739 12548 3740 12612
rect 3804 12548 3805 12612
rect 3739 12547 3805 12548
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2267 12476 2333 12477
rect 2267 12412 2268 12476
rect 2332 12412 2333 12476
rect 2267 12411 2333 12412
rect 2270 9893 2330 12411
rect 2818 11456 3138 12480
rect 4478 12341 4538 15267
rect 4692 15264 5012 16288
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6315 13292 6381 13293
rect 6315 13228 6316 13292
rect 6380 13228 6381 13292
rect 6315 13227 6381 13228
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4475 12340 4541 12341
rect 4475 12276 4476 12340
rect 4540 12276 4541 12340
rect 4475 12275 4541 12276
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 1531 9892 1597 9893
rect 1531 9828 1532 9892
rect 1596 9828 1597 9892
rect 1531 9827 1597 9828
rect 2267 9892 2333 9893
rect 2267 9828 2268 9892
rect 2332 9828 2333 9892
rect 2267 9827 2333 9828
rect 1534 7989 1594 9827
rect 1531 7988 1597 7989
rect 1531 7924 1532 7988
rect 1596 7924 1597 7988
rect 1531 7923 1597 7924
rect 1534 4045 1594 7923
rect 2270 5269 2330 9827
rect 2818 9280 3138 10304
rect 4692 12000 5012 13024
rect 5579 13020 5645 13021
rect 5579 12956 5580 13020
rect 5644 12956 5645 13020
rect 5579 12955 5645 12956
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 5582 10709 5642 12955
rect 6318 11661 6378 13227
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 5763 11660 5829 11661
rect 5763 11596 5764 11660
rect 5828 11596 5829 11660
rect 5763 11595 5829 11596
rect 6315 11660 6381 11661
rect 6315 11596 6316 11660
rect 6380 11596 6381 11660
rect 6315 11595 6381 11596
rect 5579 10708 5645 10709
rect 5579 10644 5580 10708
rect 5644 10644 5645 10708
rect 5579 10643 5645 10644
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 3371 9620 3437 9621
rect 3371 9556 3372 9620
rect 3436 9556 3437 9620
rect 3371 9555 3437 9556
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2267 5268 2333 5269
rect 2267 5204 2268 5268
rect 2332 5204 2333 5268
rect 2267 5203 2333 5204
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 1531 4044 1597 4045
rect 1531 3980 1532 4044
rect 1596 3980 1597 4044
rect 1531 3979 1597 3980
rect 2818 3840 3138 4864
rect 3374 4589 3434 9555
rect 4692 8736 5012 9760
rect 5211 9348 5277 9349
rect 5211 9284 5212 9348
rect 5276 9284 5277 9348
rect 5211 9283 5277 9284
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4107 7580 4173 7581
rect 4107 7516 4108 7580
rect 4172 7516 4173 7580
rect 4107 7515 4173 7516
rect 4110 4725 4170 7515
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4107 4724 4173 4725
rect 4107 4660 4108 4724
rect 4172 4660 4173 4724
rect 4107 4659 4173 4660
rect 3371 4588 3437 4589
rect 3371 4524 3372 4588
rect 3436 4524 3437 4588
rect 3371 4523 3437 4524
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 4110 3229 4170 4659
rect 4692 4384 5012 5408
rect 5214 4589 5274 9283
rect 5766 6901 5826 11595
rect 6566 11456 6886 12480
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 10314 16896 10634 17456
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 11651 17236 11717 17237
rect 11651 17172 11652 17236
rect 11716 17172 11717 17236
rect 11651 17171 11717 17172
rect 11467 17100 11533 17101
rect 11467 17036 11468 17100
rect 11532 17036 11533 17100
rect 11467 17035 11533 17036
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 9075 16148 9141 16149
rect 9075 16084 9076 16148
rect 9140 16084 9141 16148
rect 9075 16083 9141 16084
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8891 14516 8957 14517
rect 8891 14452 8892 14516
rect 8956 14452 8957 14516
rect 8891 14451 8957 14452
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8894 13157 8954 14451
rect 8891 13156 8957 13157
rect 8891 13092 8892 13156
rect 8956 13092 8957 13156
rect 8891 13091 8957 13092
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 7419 12204 7485 12205
rect 7419 12140 7420 12204
rect 7484 12140 7485 12204
rect 7419 12139 7485 12140
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 7422 7445 7482 12139
rect 8440 12000 8760 13024
rect 9078 13021 9138 16083
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 14720 10634 15744
rect 11099 15332 11165 15333
rect 11099 15268 11100 15332
rect 11164 15268 11165 15332
rect 11099 15267 11165 15268
rect 11283 15332 11349 15333
rect 11283 15268 11284 15332
rect 11348 15268 11349 15332
rect 11283 15267 11349 15268
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 9259 14244 9325 14245
rect 9259 14180 9260 14244
rect 9324 14180 9325 14244
rect 9259 14179 9325 14180
rect 9262 13565 9322 14179
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 9259 13564 9325 13565
rect 9259 13500 9260 13564
rect 9324 13500 9325 13564
rect 9259 13499 9325 13500
rect 9075 13020 9141 13021
rect 9075 12956 9076 13020
rect 9140 12956 9141 13020
rect 9075 12955 9141 12956
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 10314 12544 10634 13568
rect 11102 13293 11162 15267
rect 11099 13292 11165 13293
rect 11099 13228 11100 13292
rect 11164 13228 11165 13292
rect 11099 13227 11165 13228
rect 11099 12884 11165 12885
rect 11099 12820 11100 12884
rect 11164 12820 11165 12884
rect 11099 12819 11165 12820
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 8891 8940 8957 8941
rect 8891 8876 8892 8940
rect 8956 8876 8957 8940
rect 8891 8875 8957 8876
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8155 8532 8221 8533
rect 8155 8468 8156 8532
rect 8220 8468 8221 8532
rect 8155 8467 8221 8468
rect 7419 7444 7485 7445
rect 7419 7380 7420 7444
rect 7484 7380 7485 7444
rect 7419 7379 7485 7380
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 5763 6900 5829 6901
rect 5763 6836 5764 6900
rect 5828 6836 5829 6900
rect 5763 6835 5829 6836
rect 5763 6628 5829 6629
rect 5763 6564 5764 6628
rect 5828 6564 5829 6628
rect 5763 6563 5829 6564
rect 5211 4588 5277 4589
rect 5211 4524 5212 4588
rect 5276 4524 5277 4588
rect 5211 4523 5277 4524
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4107 3228 4173 3229
rect 4107 3164 4108 3228
rect 4172 3164 4173 3228
rect 4107 3163 4173 3164
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 4692 2208 5012 3232
rect 5766 2413 5826 6563
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 5763 2412 5829 2413
rect 5763 2348 5764 2412
rect 5828 2348 5829 2412
rect 5763 2347 5829 2348
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 2128 6886 2688
rect 8158 2685 8218 8467
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 8440 2208 8760 3232
rect 8894 2549 8954 8875
rect 10314 8192 10634 9216
rect 11102 9213 11162 12819
rect 11286 11525 11346 15267
rect 11470 14109 11530 17035
rect 11467 14108 11533 14109
rect 11467 14044 11468 14108
rect 11532 14044 11533 14108
rect 11467 14043 11533 14044
rect 11654 13157 11714 17171
rect 12188 16352 12508 17376
rect 12571 16964 12637 16965
rect 12571 16900 12572 16964
rect 12636 16900 12637 16964
rect 12571 16899 12637 16900
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 11835 15876 11901 15877
rect 11835 15812 11836 15876
rect 11900 15812 11901 15876
rect 11835 15811 11901 15812
rect 11651 13156 11717 13157
rect 11651 13092 11652 13156
rect 11716 13092 11717 13156
rect 11651 13091 11717 13092
rect 11283 11524 11349 11525
rect 11283 11460 11284 11524
rect 11348 11460 11349 11524
rect 11283 11459 11349 11460
rect 11099 9212 11165 9213
rect 11099 9148 11100 9212
rect 11164 9148 11165 9212
rect 11099 9147 11165 9148
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 11102 8125 11162 9147
rect 11099 8124 11165 8125
rect 11099 8060 11100 8124
rect 11164 8060 11165 8124
rect 11099 8059 11165 8060
rect 11286 7173 11346 11459
rect 11283 7172 11349 7173
rect 11283 7108 11284 7172
rect 11348 7108 11349 7172
rect 11283 7107 11349 7108
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 11099 7036 11165 7037
rect 11099 6972 11100 7036
rect 11164 6972 11165 7036
rect 11099 6971 11165 6972
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 4928 10634 5952
rect 11102 5269 11162 6971
rect 11838 6357 11898 15811
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12574 10165 12634 16899
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 13491 16692 13557 16693
rect 13491 16628 13492 16692
rect 13556 16628 13557 16692
rect 13491 16627 13557 16628
rect 12755 14788 12821 14789
rect 12755 14724 12756 14788
rect 12820 14724 12821 14788
rect 12755 14723 12821 14724
rect 12758 11797 12818 14723
rect 13123 14516 13189 14517
rect 13123 14452 13124 14516
rect 13188 14452 13189 14516
rect 13123 14451 13189 14452
rect 13126 13701 13186 14451
rect 13307 13972 13373 13973
rect 13307 13908 13308 13972
rect 13372 13908 13373 13972
rect 13307 13907 13373 13908
rect 13123 13700 13189 13701
rect 13123 13636 13124 13700
rect 13188 13636 13189 13700
rect 13123 13635 13189 13636
rect 12755 11796 12821 11797
rect 12755 11732 12756 11796
rect 12820 11732 12821 11796
rect 12755 11731 12821 11732
rect 12571 10164 12637 10165
rect 12571 10100 12572 10164
rect 12636 10100 12637 10164
rect 12571 10099 12637 10100
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12574 7989 12634 10099
rect 12571 7988 12637 7989
rect 12571 7924 12572 7988
rect 12636 7924 12637 7988
rect 12571 7923 12637 7924
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 13310 7445 13370 13907
rect 13494 8669 13554 16627
rect 14062 15808 14382 16832
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14963 14516 15029 14517
rect 14963 14452 14964 14516
rect 15028 14452 15029 14516
rect 14963 14451 15029 14452
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14595 13156 14661 13157
rect 14595 13092 14596 13156
rect 14660 13092 14661 13156
rect 14595 13091 14661 13092
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 13859 12204 13925 12205
rect 13859 12140 13860 12204
rect 13924 12140 13925 12204
rect 13859 12139 13925 12140
rect 13491 8668 13557 8669
rect 13491 8604 13492 8668
rect 13556 8604 13557 8668
rect 13491 8603 13557 8604
rect 13862 7989 13922 12139
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 8192 14382 9216
rect 14598 9077 14658 13091
rect 14779 11660 14845 11661
rect 14779 11596 14780 11660
rect 14844 11596 14845 11660
rect 14779 11595 14845 11596
rect 14595 9076 14661 9077
rect 14595 9012 14596 9076
rect 14660 9012 14661 9076
rect 14595 9011 14661 9012
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 13859 7988 13925 7989
rect 13859 7924 13860 7988
rect 13924 7924 13925 7988
rect 13859 7923 13925 7924
rect 13307 7444 13373 7445
rect 13307 7380 13308 7444
rect 13372 7380 13373 7444
rect 13307 7379 13373 7380
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 11835 6356 11901 6357
rect 11835 6292 11836 6356
rect 11900 6292 11901 6356
rect 11835 6291 11901 6292
rect 12188 5472 12508 6496
rect 12755 6356 12821 6357
rect 12755 6292 12756 6356
rect 12820 6292 12821 6356
rect 12755 6291 12821 6292
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 11099 5268 11165 5269
rect 11099 5204 11100 5268
rect 11164 5204 11165 5268
rect 11099 5203 11165 5204
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10314 2752 10634 3776
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 8891 2548 8957 2549
rect 8891 2484 8892 2548
rect 8956 2484 8957 2548
rect 8891 2483 8957 2484
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 10314 2128 10634 2688
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 3296 12508 4320
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 2208 12508 3232
rect 12758 2957 12818 6291
rect 13310 5405 13370 7379
rect 14062 7104 14382 8128
rect 14595 7852 14661 7853
rect 14595 7788 14596 7852
rect 14660 7850 14661 7852
rect 14782 7850 14842 11595
rect 14966 9893 15026 14451
rect 14963 9892 15029 9893
rect 14963 9828 14964 9892
rect 15028 9828 15029 9892
rect 14963 9827 15029 9828
rect 14963 9348 15029 9349
rect 14963 9284 14964 9348
rect 15028 9284 15029 9348
rect 14963 9283 15029 9284
rect 14660 7790 14842 7850
rect 14660 7788 14661 7790
rect 14595 7787 14661 7788
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 13307 5404 13373 5405
rect 13307 5340 13308 5404
rect 13372 5340 13373 5404
rect 13307 5339 13373 5340
rect 14062 4928 14382 5952
rect 14598 5677 14658 7787
rect 14595 5676 14661 5677
rect 14595 5612 14596 5676
rect 14660 5612 14661 5676
rect 14595 5611 14661 5612
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 12755 2956 12821 2957
rect 12755 2892 12756 2956
rect 12820 2892 12821 2956
rect 12755 2891 12821 2892
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2128 14382 2688
rect 14966 2685 15026 9283
rect 14963 2684 15029 2685
rect 14963 2620 14964 2684
rect 15028 2620 15029 2684
rect 14963 2619 15029 2620
use sky130_fd_sc_hd__diode_2  ANTENNA__38__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__39__A
timestamp 1649977179
transform 1 0 2576 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__41__A
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__42__A
timestamp 1649977179
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__43__A
timestamp 1649977179
transform -1 0 2760 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__44__A
timestamp 1649977179
transform 1 0 2024 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__46__A
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__48__A
timestamp 1649977179
transform -1 0 2484 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__49__A
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__51__A
timestamp 1649977179
transform 1 0 7176 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__52__A
timestamp 1649977179
transform 1 0 7544 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__53__A
timestamp 1649977179
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__57__A
timestamp 1649977179
transform 1 0 3220 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__58__A
timestamp 1649977179
transform 1 0 5612 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__59__A
timestamp 1649977179
transform -1 0 1840 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__60__A
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__61__A
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__62__A
timestamp 1649977179
transform -1 0 1656 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__63__A
timestamp 1649977179
transform 1 0 4600 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__64__A
timestamp 1649977179
transform -1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__65__A
timestamp 1649977179
transform -1 0 3036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__66__A
timestamp 1649977179
transform 1 0 7544 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__67__A
timestamp 1649977179
transform -1 0 3680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__68__A
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__69__A
timestamp 1649977179
transform -1 0 1564 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__70__A
timestamp 1649977179
transform -1 0 3956 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__71__A
timestamp 1649977179
transform -1 0 4140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__72__A
timestamp 1649977179
transform -1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__73__A
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_prog_clk_0_W_in_A
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 3956 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 14812 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 14996 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 15364 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15732 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 15180 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 11684 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 9200 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 5520 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 6532 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 12512 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 14628 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 8832 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 14260 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform 1 0 12696 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 15732 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 13984 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 10948 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 8004 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 10764 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 15732 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 11684 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 9384 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 15272 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 3220 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 15732 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 15364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 15088 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_ipin_0.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15180 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11132 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14260 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_0.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 3680 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_1.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 8372 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 7912 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 3680 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_2.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 2208 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 3128 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2760 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 3680 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 7728 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6532 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_4.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_5.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9752 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12972 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_6.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 13892 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13616 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11592 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_2__A1
timestamp 1649977179
transform -1 0 15456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_7.mux_l2_in_3__A1
timestamp 1649977179
transform -1 0 15640 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 13524 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8832 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 9384 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5520 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_9.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 3956 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_10.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 4232 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 7176 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 5152 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_11.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 8832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12328 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_12.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 12420 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 7176 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_13.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 7360 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_14.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 15732 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 12880 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_ipin_15.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater114_A
timestamp 1649977179
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_repeater120_A
timestamp 1649977179
transform 1 0 9292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_133
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_158
timestamp 1649977179
transform 1 0 15640 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_18
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_145
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_66
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1649977179
transform 1 0 9476 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_95
timestamp 1649977179
transform 1 0 9844 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_138
timestamp 1649977179
transform 1 0 13800 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1649977179
transform 1 0 9476 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_116
timestamp 1649977179
transform 1 0 11776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_144
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_154
timestamp 1649977179
transform 1 0 15272 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_63
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_75
timestamp 1649977179
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_11
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_81
timestamp 1649977179
transform 1 0 8556 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_111
timestamp 1649977179
transform 1 0 11316 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_156
timestamp 1649977179
transform 1 0 15456 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_22
timestamp 1649977179
transform 1 0 3128 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_136
timestamp 1649977179
transform 1 0 13616 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_90
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_155 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_12
timestamp 1649977179
transform 1 0 2208 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_100
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_153 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_7 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_94
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_18
timestamp 1649977179
transform 1 0 2760 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_59
timestamp 1649977179
transform 1 0 6532 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_70
timestamp 1649977179
transform 1 0 7544 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_135
timestamp 1649977179
transform 1 0 13524 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_79 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_92
timestamp 1649977179
transform 1 0 9568 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_104
timestamp 1649977179
transform 1 0 10672 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_122
timestamp 1649977179
transform 1 0 12328 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_158
timestamp 1649977179
transform 1 0 15640 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_25
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_101
timestamp 1649977179
transform 1 0 10396 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_40
timestamp 1649977179
transform 1 0 4784 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_86
timestamp 1649977179
transform 1 0 9016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_95
timestamp 1649977179
transform 1 0 9844 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_124
timestamp 1649977179
transform 1 0 12512 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_87
timestamp 1649977179
transform 1 0 9108 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_10
timestamp 1649977179
transform 1 0 2024 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_54
timestamp 1649977179
transform 1 0 6072 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_71
timestamp 1649977179
transform 1 0 7636 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_81
timestamp 1649977179
transform 1 0 8556 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_87
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_46
timestamp 1649977179
transform 1 0 5336 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_75
timestamp 1649977179
transform 1 0 8004 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_95
timestamp 1649977179
transform 1 0 9844 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_10
timestamp 1649977179
transform 1 0 2024 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_57
timestamp 1649977179
transform 1 0 6348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_106
timestamp 1649977179
transform 1 0 10856 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_116
timestamp 1649977179
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_18
timestamp 1649977179
transform 1 0 2760 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_31
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_35
timestamp 1649977179
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_79
timestamp 1649977179
transform 1 0 8372 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_118
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _34_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 2576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform -1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform -1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform -1 0 2576 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform 1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _43_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _44_
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _45_
timestamp 1649977179
transform 1 0 9292 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _46_
timestamp 1649977179
transform 1 0 5612 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _47_
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _48_
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _49_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform 1 0 3220 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform 1 0 2944 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform 1 0 3680 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform 1 0 2852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform 1 0 4324 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 3680 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform 1 0 4416 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 4876 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 4968 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform -1 0 5428 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 5704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform -1 0 6624 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform 1 0 8464 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform 1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9752 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_prog_clk_0_W_in
timestamp 1649977179
transform 1 0 13892 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_prog_clk_0_W_in
timestamp 1649977179
transform -1 0 15732 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_prog_clk_0_W_in
timestamp 1649977179
transform -1 0 14812 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform -1 0 9660 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 7268 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform 1 0 8096 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform -1 0 3496 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 8648 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform -1 0 5428 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform -1 0 2668 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 8096 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 10120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform -1 0 6164 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 3680 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform -1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 3128 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform 1 0 14996 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 5336 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 1472 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 10672 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform -1 0 11684 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform -1 0 15732 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 4048 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13984 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1649977179
transform 1 0 14536 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform 1 0 14536 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1649977179
transform -1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1649977179
transform -1 0 15364 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input11
timestamp 1649977179
transform -1 0 15732 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform -1 0 15732 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1649977179
transform -1 0 14904 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 10120 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1649977179
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform -1 0 12696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform -1 0 13064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1649977179
transform -1 0 11684 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1649977179
transform -1 0 13340 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform -1 0 11868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1649977179
transform -1 0 9292 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform -1 0 13800 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform 1 0 14168 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input28
timestamp 1649977179
transform -1 0 11868 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1649977179
transform -1 0 13064 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform -1 0 14168 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform -1 0 11408 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 13892 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1649977179
transform -1 0 12696 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 12144 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 8832 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1649977179
transform 1 0 13524 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 11960 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 11408 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 13892 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input41
timestamp 1649977179
transform 1 0 12144 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1649977179
transform 1 0 13064 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 15088 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 3680 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2024 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 13064 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12512 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11316 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9844 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8832 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9844 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8464 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5888 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8004 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5888 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2208 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5428 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3496 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2208 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5244 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2208 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 4692 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4968 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6440 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6900 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 9292 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10028 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12972 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_6.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 11408 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_7.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 13156 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11684 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11408 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7176 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5888 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5244 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 2852 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 1840 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3312 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_10.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3036 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4416 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6164 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 5796 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_11.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7268 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13708 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_12.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9200 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8832 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_13.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 7820 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 6900 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8372 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 9292 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_14.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 9936 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 13524 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_15.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13892 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13524 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12972 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12512 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_ipin_0.mux_l2_in_3__129 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12512 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 14352 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14444 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10120 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 10396 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9568 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_0.mux_l2_in_3__130
timestamp 1649977179
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9844 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 10488 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9016 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8372 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7912 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6992 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_1.mux_l2_in_3__131
timestamp 1649977179
transform -1 0 6992 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l3_in_1_
timestamp 1649977179
transform -1 0 6992 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_1.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5704 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 5704 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_2.mux_l2_in_3__138
timestamp 1649977179
transform -1 0 2024 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 4508 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_2.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2024 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 2208 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 1932 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_3.mux_l2_in_3__139
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5428 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2208 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4600 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 5428 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6072 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4784 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_4.mux_l2_in_3__123
timestamp 1649977179
transform 1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l3_in_1_
timestamp 1649977179
transform 1 0 4140 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_4.mux_l4_in_0_
timestamp 1649977179
transform 1 0 3864 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6716 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_5.mux_l2_in_3__124
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 6256 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l3_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11224 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11868 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_6.mux_l2_in_3__125
timestamp 1649977179
transform -1 0 13432 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10488 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11408 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_6.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10304 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13984 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12604 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13432 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_1_
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14628 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_7.mux_l2_in_3__126
timestamp 1649977179
transform -1 0 15180 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l3_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_7.mux_l4_in_0_
timestamp 1649977179
transform 1 0 12328 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9476 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 8004 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_8.mux_l2_in_3__127
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7912 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 7176 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_8.mux_l4_in_0_
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3312 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3680 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_9.mux_l2_in_3__128
timestamp 1649977179
transform 1 0 6072 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l2_in_3_
timestamp 1649977179
transform 1 0 5244 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2852 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l3_in_1_
timestamp 1649977179
transform 1 0 3864 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_9.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2760 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2576 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_1_
timestamp 1649977179
transform 1 0 2944 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_2_
timestamp 1649977179
transform 1 0 4508 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_10.mux_l2_in_3__132
timestamp 1649977179
transform 1 0 4140 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2852 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2852 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_10.mux_l4_in_0_
timestamp 1649977179
transform -1 0 2944 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_0_
timestamp 1649977179
transform -1 0 5428 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6256 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l1_in_2_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_1_
timestamp 1649977179
transform 1 0 5336 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7268 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_11.mux_l2_in_3__133
timestamp 1649977179
transform 1 0 8096 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l2_in_3_
timestamp 1649977179
transform 1 0 7268 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 5244 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6440 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_11.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4784 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9936 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_2_
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_12.mux_l2_in_3__134
timestamp 1649977179
transform -1 0 12880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l2_in_3_
timestamp 1649977179
transform 1 0 12604 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_0_
timestamp 1649977179
transform 1 0 9568 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l3_in_1_
timestamp 1649977179
transform 1 0 11960 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_12.mux_l4_in_0_
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_2_
timestamp 1649977179
transform 1 0 7820 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_13.mux_l2_in_3__135
timestamp 1649977179
transform 1 0 8556 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l2_in_3_
timestamp 1649977179
transform -1 0 7268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6072 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l3_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_13.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5428 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1472 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10028 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_1_
timestamp 1649977179
transform 1 0 10764 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l2_in_3_
timestamp 1649977179
transform 1 0 10948 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_14.mux_l2_in_3__136
timestamp 1649977179
transform 1 0 13708 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10856 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l3_in_1_
timestamp 1649977179
transform -1 0 10488 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_14.mux_l4_in_0_
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 12696 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l1_in_2_
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11868 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11868 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_15.mux_l2_in_3__137
timestamp 1649977179
transform -1 0 11960 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l2_in_3_
timestamp 1649977179
transform -1 0 14996 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_0_
timestamp 1649977179
transform -1 0 10948 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l3_in_1_
timestamp 1649977179
transform -1 0 15732 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_15.mux_l4_in_0_
timestamp 1649977179
transform 1 0 14904 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output45 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform 1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 3680 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 6256 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 7728 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 6256 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 2116 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 1932 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 2576 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 2024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 1840 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 2944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 4968 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 5704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 6992 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 3680 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 1748 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1748 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 2576 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 2484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output104
timestamp 1649977179
transform -1 0 12696 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  output105
timestamp 1649977179
transform -1 0 15732 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 15364 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14168 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_N_FTB01 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  prog_clk_0_S_FTB01
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater107
timestamp 1649977179
transform 1 0 10488 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater108
timestamp 1649977179
transform 1 0 12696 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater109
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater110
timestamp 1649977179
transform 1 0 13064 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater111
timestamp 1649977179
transform 1 0 10212 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  repeater112
timestamp 1649977179
transform -1 0 9844 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater113
timestamp 1649977179
transform -1 0 6256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater114
timestamp 1649977179
transform -1 0 8372 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater115
timestamp 1649977179
transform -1 0 8464 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  repeater116
timestamp 1649977179
transform -1 0 8556 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  repeater117
timestamp 1649977179
transform -1 0 11776 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  repeater118
timestamp 1649977179
transform -1 0 10212 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater119
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater120
timestamp 1649977179
transform -1 0 8832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater121
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater122
timestamp 1649977179
transform -1 0 7084 0 1 2176
box -38 -48 406 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal4 s 4692 2128 5012 17456 6 VGND
port 1 nsew ground input
rlabel metal4 s 8440 2128 8760 17456 6 VGND
port 1 nsew ground input
rlabel metal4 s 12188 2128 12508 17456 6 VGND
port 1 nsew ground input
rlabel metal4 s 2818 2128 3138 17456 6 VPWR
port 2 nsew power input
rlabel metal4 s 6566 2128 6886 17456 6 VPWR
port 2 nsew power input
rlabel metal4 s 10314 2128 10634 17456 6 VPWR
port 2 nsew power input
rlabel metal4 s 14062 2128 14382 17456 6 VPWR
port 2 nsew power input
rlabel metal3 s 0 1368 800 1488 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 16400 1912 17200 2032 6 ccff_tail
port 4 nsew signal tristate
rlabel metal2 s 8574 0 8630 800 6 chany_bottom_in[0]
port 5 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_in[10]
port 6 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 chany_bottom_in[11]
port 7 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 chany_bottom_in[12]
port 8 nsew signal input
rlabel metal2 s 14002 0 14058 800 6 chany_bottom_in[13]
port 9 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 chany_bottom_in[14]
port 10 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 chany_bottom_in[15]
port 11 nsew signal input
rlabel metal2 s 15290 0 15346 800 6 chany_bottom_in[16]
port 12 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[17]
port 13 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 chany_bottom_in[18]
port 14 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[19]
port 15 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[1]
port 16 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 chany_bottom_in[2]
port 17 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 chany_bottom_in[3]
port 18 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 chany_bottom_in[4]
port 19 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 chany_bottom_in[5]
port 20 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 chany_bottom_in[6]
port 21 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 chany_bottom_in[7]
port 22 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[8]
port 23 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[9]
port 24 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 25 nsew signal tristate
rlabel metal2 s 4342 0 4398 800 6 chany_bottom_out[10]
port 26 nsew signal tristate
rlabel metal2 s 4802 0 4858 800 6 chany_bottom_out[11]
port 27 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 chany_bottom_out[12]
port 28 nsew signal tristate
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_out[13]
port 29 nsew signal tristate
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_out[14]
port 30 nsew signal tristate
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_out[15]
port 31 nsew signal tristate
rlabel metal2 s 6826 0 6882 800 6 chany_bottom_out[16]
port 32 nsew signal tristate
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_out[17]
port 33 nsew signal tristate
rlabel metal2 s 7746 0 7802 800 6 chany_bottom_out[18]
port 34 nsew signal tristate
rlabel metal2 s 8114 0 8170 800 6 chany_bottom_out[19]
port 35 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 36 nsew signal tristate
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 37 nsew signal tristate
rlabel metal2 s 1398 0 1454 800 6 chany_bottom_out[3]
port 38 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 39 nsew signal tristate
rlabel metal2 s 2226 0 2282 800 6 chany_bottom_out[5]
port 40 nsew signal tristate
rlabel metal2 s 2686 0 2742 800 6 chany_bottom_out[6]
port 41 nsew signal tristate
rlabel metal2 s 3054 0 3110 800 6 chany_bottom_out[7]
port 42 nsew signal tristate
rlabel metal2 s 3514 0 3570 800 6 chany_bottom_out[8]
port 43 nsew signal tristate
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_out[9]
port 44 nsew signal tristate
rlabel metal2 s 8758 19200 8814 20000 6 chany_top_in[0]
port 45 nsew signal input
rlabel metal2 s 12898 19200 12954 20000 6 chany_top_in[10]
port 46 nsew signal input
rlabel metal2 s 13266 19200 13322 20000 6 chany_top_in[11]
port 47 nsew signal input
rlabel metal2 s 13634 19200 13690 20000 6 chany_top_in[12]
port 48 nsew signal input
rlabel metal2 s 14094 19200 14150 20000 6 chany_top_in[13]
port 49 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[14]
port 50 nsew signal input
rlabel metal2 s 14922 19200 14978 20000 6 chany_top_in[15]
port 51 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[16]
port 52 nsew signal input
rlabel metal2 s 15750 19200 15806 20000 6 chany_top_in[17]
port 53 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[18]
port 54 nsew signal input
rlabel metal2 s 16578 19200 16634 20000 6 chany_top_in[19]
port 55 nsew signal input
rlabel metal2 s 9126 19200 9182 20000 6 chany_top_in[1]
port 56 nsew signal input
rlabel metal2 s 9586 19200 9642 20000 6 chany_top_in[2]
port 57 nsew signal input
rlabel metal2 s 9954 19200 10010 20000 6 chany_top_in[3]
port 58 nsew signal input
rlabel metal2 s 10414 19200 10470 20000 6 chany_top_in[4]
port 59 nsew signal input
rlabel metal2 s 10782 19200 10838 20000 6 chany_top_in[5]
port 60 nsew signal input
rlabel metal2 s 11242 19200 11298 20000 6 chany_top_in[6]
port 61 nsew signal input
rlabel metal2 s 11610 19200 11666 20000 6 chany_top_in[7]
port 62 nsew signal input
rlabel metal2 s 12070 19200 12126 20000 6 chany_top_in[8]
port 63 nsew signal input
rlabel metal2 s 12438 19200 12494 20000 6 chany_top_in[9]
port 64 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 65 nsew signal tristate
rlabel metal2 s 4618 19200 4674 20000 6 chany_top_out[10]
port 66 nsew signal tristate
rlabel metal2 s 5078 19200 5134 20000 6 chany_top_out[11]
port 67 nsew signal tristate
rlabel metal2 s 5446 19200 5502 20000 6 chany_top_out[12]
port 68 nsew signal tristate
rlabel metal2 s 5906 19200 5962 20000 6 chany_top_out[13]
port 69 nsew signal tristate
rlabel metal2 s 6274 19200 6330 20000 6 chany_top_out[14]
port 70 nsew signal tristate
rlabel metal2 s 6734 19200 6790 20000 6 chany_top_out[15]
port 71 nsew signal tristate
rlabel metal2 s 7102 19200 7158 20000 6 chany_top_out[16]
port 72 nsew signal tristate
rlabel metal2 s 7562 19200 7618 20000 6 chany_top_out[17]
port 73 nsew signal tristate
rlabel metal2 s 7930 19200 7986 20000 6 chany_top_out[18]
port 74 nsew signal tristate
rlabel metal2 s 8390 19200 8446 20000 6 chany_top_out[19]
port 75 nsew signal tristate
rlabel metal2 s 938 19200 994 20000 6 chany_top_out[1]
port 76 nsew signal tristate
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 77 nsew signal tristate
rlabel metal2 s 1766 19200 1822 20000 6 chany_top_out[3]
port 78 nsew signal tristate
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 79 nsew signal tristate
rlabel metal2 s 2594 19200 2650 20000 6 chany_top_out[5]
port 80 nsew signal tristate
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 81 nsew signal tristate
rlabel metal2 s 3422 19200 3478 20000 6 chany_top_out[7]
port 82 nsew signal tristate
rlabel metal2 s 3882 19200 3938 20000 6 chany_top_out[8]
port 83 nsew signal tristate
rlabel metal2 s 4250 19200 4306 20000 6 chany_top_out[9]
port 84 nsew signal tristate
rlabel metal3 s 16400 9800 17200 9920 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 85 nsew signal tristate
rlabel metal3 s 16400 13880 17200 14000 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 86 nsew signal input
rlabel metal3 s 16400 17824 17200 17944 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 87 nsew signal tristate
rlabel metal3 s 0 3272 800 3392 6 left_grid_pin_16_
port 88 nsew signal tristate
rlabel metal3 s 0 4224 800 4344 6 left_grid_pin_17_
port 89 nsew signal tristate
rlabel metal3 s 0 5176 800 5296 6 left_grid_pin_18_
port 90 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 left_grid_pin_19_
port 91 nsew signal tristate
rlabel metal3 s 0 7080 800 7200 6 left_grid_pin_20_
port 92 nsew signal tristate
rlabel metal3 s 0 8032 800 8152 6 left_grid_pin_21_
port 93 nsew signal tristate
rlabel metal3 s 0 8984 800 9104 6 left_grid_pin_22_
port 94 nsew signal tristate
rlabel metal3 s 0 9936 800 10056 6 left_grid_pin_23_
port 95 nsew signal tristate
rlabel metal3 s 0 10888 800 11008 6 left_grid_pin_24_
port 96 nsew signal tristate
rlabel metal3 s 0 11840 800 11960 6 left_grid_pin_25_
port 97 nsew signal tristate
rlabel metal3 s 0 12792 800 12912 6 left_grid_pin_26_
port 98 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 left_grid_pin_27_
port 99 nsew signal tristate
rlabel metal3 s 0 14696 800 14816 6 left_grid_pin_28_
port 100 nsew signal tristate
rlabel metal3 s 0 15648 800 15768 6 left_grid_pin_29_
port 101 nsew signal tristate
rlabel metal3 s 0 16600 800 16720 6 left_grid_pin_30_
port 102 nsew signal tristate
rlabel metal3 s 0 17552 800 17672 6 left_grid_pin_31_
port 103 nsew signal tristate
rlabel metal3 s 0 18504 800 18624 6 left_width_0_height_0__pin_0_
port 104 nsew signal input
rlabel metal3 s 0 416 800 536 6 left_width_0_height_0__pin_1_lower
port 105 nsew signal tristate
rlabel metal3 s 0 19456 800 19576 6 left_width_0_height_0__pin_1_upper
port 106 nsew signal tristate
rlabel metal2 s 16946 19200 17002 20000 6 prog_clk_0_N_out
port 107 nsew signal tristate
rlabel metal2 s 16946 0 17002 800 6 prog_clk_0_S_out
port 108 nsew signal tristate
rlabel metal3 s 0 2320 800 2440 6 prog_clk_0_W_in
port 109 nsew signal input
rlabel metal3 s 16400 5856 17200 5976 6 right_grid_pin_0_
port 110 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
