magic
tech sky130A
magscale 1 2
timestamp 1650893698
<< viali >>
rect 1501 20553 1535 20587
rect 2053 20553 2087 20587
rect 4261 20553 4295 20587
rect 5181 20553 5215 20587
rect 17509 20553 17543 20587
rect 19625 20553 19659 20587
rect 20177 20553 20211 20587
rect 1685 20417 1719 20451
rect 2237 20417 2271 20451
rect 2789 20417 2823 20451
rect 3249 20417 3283 20451
rect 3985 20417 4019 20451
rect 4445 20417 4479 20451
rect 4721 20417 4755 20451
rect 5825 20417 5859 20451
rect 6377 20417 6411 20451
rect 17325 20417 17359 20451
rect 18429 20417 18463 20451
rect 18705 20417 18739 20451
rect 19441 20417 19475 20451
rect 19993 20417 20027 20451
rect 20545 20417 20579 20451
rect 21097 20417 21131 20451
rect 6745 20349 6779 20383
rect 2605 20281 2639 20315
rect 3065 20281 3099 20315
rect 6009 20281 6043 20315
rect 20729 20281 20763 20315
rect 3801 20213 3835 20247
rect 4905 20213 4939 20247
rect 18889 20213 18923 20247
rect 21281 20213 21315 20247
rect 2605 20009 2639 20043
rect 7573 20009 7607 20043
rect 10333 20009 10367 20043
rect 18429 20009 18463 20043
rect 18889 20009 18923 20043
rect 19717 20009 19751 20043
rect 20177 19941 20211 19975
rect 8217 19873 8251 19907
rect 1685 19805 1719 19839
rect 2237 19805 2271 19839
rect 2789 19805 2823 19839
rect 3249 19805 3283 19839
rect 5181 19805 5215 19839
rect 5457 19805 5491 19839
rect 8953 19805 8987 19839
rect 11161 19805 11195 19839
rect 11417 19805 11451 19839
rect 18245 19805 18279 19839
rect 18705 19805 18739 19839
rect 19533 19805 19567 19839
rect 19993 19805 20027 19839
rect 20545 19805 20579 19839
rect 21097 19805 21131 19839
rect 4914 19737 4948 19771
rect 6377 19737 6411 19771
rect 9220 19737 9254 19771
rect 17601 19737 17635 19771
rect 1501 19669 1535 19703
rect 2053 19669 2087 19703
rect 3065 19669 3099 19703
rect 3801 19669 3835 19703
rect 6101 19669 6135 19703
rect 7941 19669 7975 19703
rect 8033 19669 8067 19703
rect 12541 19669 12575 19703
rect 17969 19669 18003 19703
rect 20729 19669 20763 19703
rect 21281 19669 21315 19703
rect 2053 19465 2087 19499
rect 2513 19465 2547 19499
rect 2973 19465 3007 19499
rect 5365 19465 5399 19499
rect 7757 19465 7791 19499
rect 9413 19465 9447 19499
rect 19349 19465 19383 19499
rect 20085 19465 20119 19499
rect 21281 19465 21315 19499
rect 8125 19397 8159 19431
rect 9689 19397 9723 19431
rect 1685 19329 1719 19363
rect 2237 19329 2271 19363
rect 2697 19329 2731 19363
rect 3157 19329 3191 19363
rect 3709 19329 3743 19363
rect 3965 19329 3999 19363
rect 8217 19329 8251 19363
rect 8769 19329 8803 19363
rect 12541 19329 12575 19363
rect 12797 19329 12831 19363
rect 14197 19329 14231 19363
rect 14464 19329 14498 19363
rect 18889 19329 18923 19363
rect 19165 19329 19199 19363
rect 19625 19329 19659 19363
rect 20269 19329 20303 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 8401 19261 8435 19295
rect 18429 19193 18463 19227
rect 19809 19193 19843 19227
rect 20729 19193 20763 19227
rect 1501 19125 1535 19159
rect 5089 19125 5123 19159
rect 5825 19125 5859 19159
rect 13921 19125 13955 19159
rect 15577 19125 15611 19159
rect 1961 18921 1995 18955
rect 2421 18921 2455 18955
rect 2881 18921 2915 18955
rect 8953 18921 8987 18955
rect 17969 18921 18003 18955
rect 19441 18921 19475 18955
rect 19901 18921 19935 18955
rect 8585 18853 8619 18887
rect 20361 18853 20395 18887
rect 20821 18853 20855 18887
rect 3893 18785 3927 18819
rect 9505 18785 9539 18819
rect 17601 18785 17635 18819
rect 1685 18717 1719 18751
rect 2145 18717 2179 18751
rect 2605 18717 2639 18751
rect 3065 18717 3099 18751
rect 5181 18717 5215 18751
rect 5448 18717 5482 18751
rect 7205 18717 7239 18751
rect 14565 18717 14599 18751
rect 14832 18717 14866 18751
rect 16221 18717 16255 18751
rect 19257 18717 19291 18751
rect 19717 18717 19751 18751
rect 20177 18717 20211 18751
rect 20637 18717 20671 18751
rect 21097 18717 21131 18751
rect 3433 18649 3467 18683
rect 7472 18649 7506 18683
rect 1501 18581 1535 18615
rect 4169 18581 4203 18615
rect 4629 18581 4663 18615
rect 6561 18581 6595 18615
rect 9321 18581 9355 18615
rect 9413 18581 9447 18615
rect 15945 18581 15979 18615
rect 16865 18581 16899 18615
rect 18337 18581 18371 18615
rect 18889 18581 18923 18615
rect 21281 18581 21315 18615
rect 2421 18377 2455 18411
rect 3985 18377 4019 18411
rect 4629 18377 4663 18411
rect 9413 18377 9447 18411
rect 9781 18377 9815 18411
rect 19441 18377 19475 18411
rect 20361 18377 20395 18411
rect 6377 18309 6411 18343
rect 8953 18309 8987 18343
rect 14105 18309 14139 18343
rect 15761 18309 15795 18343
rect 1685 18241 1719 18275
rect 2145 18241 2179 18275
rect 2605 18241 2639 18275
rect 3617 18241 3651 18275
rect 9045 18241 9079 18275
rect 11989 18241 12023 18275
rect 14013 18241 14047 18275
rect 15117 18241 15151 18275
rect 17877 18241 17911 18275
rect 19165 18241 19199 18275
rect 20177 18241 20211 18275
rect 20637 18241 20671 18275
rect 21097 18241 21131 18275
rect 3341 18173 3375 18207
rect 3525 18173 3559 18207
rect 4721 18173 4755 18207
rect 4905 18173 4939 18207
rect 8769 18173 8803 18207
rect 12909 18173 12943 18207
rect 13921 18173 13955 18207
rect 14841 18173 14875 18207
rect 15025 18173 15059 18207
rect 17969 18173 18003 18207
rect 18153 18173 18187 18207
rect 1961 18105 1995 18139
rect 5641 18105 5675 18139
rect 8401 18105 8435 18139
rect 1501 18037 1535 18071
rect 2881 18037 2915 18071
rect 4261 18037 4295 18071
rect 5273 18037 5307 18071
rect 12633 18037 12667 18071
rect 13461 18037 13495 18071
rect 14473 18037 14507 18071
rect 15485 18037 15519 18071
rect 17509 18037 17543 18071
rect 18521 18037 18555 18071
rect 19809 18037 19843 18071
rect 20821 18037 20855 18071
rect 21281 18037 21315 18071
rect 4445 17833 4479 17867
rect 7849 17833 7883 17867
rect 13645 17833 13679 17867
rect 15117 17833 15151 17867
rect 19349 17833 19383 17867
rect 19717 17833 19751 17867
rect 20361 17833 20395 17867
rect 1961 17765 1995 17799
rect 3433 17765 3467 17799
rect 10333 17765 10367 17799
rect 4997 17697 5031 17731
rect 12817 17697 12851 17731
rect 14289 17697 14323 17731
rect 15669 17697 15703 17731
rect 16681 17697 16715 17731
rect 1685 17629 1719 17663
rect 2145 17629 2179 17663
rect 2605 17629 2639 17663
rect 3065 17629 3099 17663
rect 7205 17629 7239 17663
rect 8033 17629 8067 17663
rect 8953 17629 8987 17663
rect 10609 17629 10643 17663
rect 10876 17629 10910 17663
rect 15485 17629 15519 17663
rect 18889 17629 18923 17663
rect 19901 17629 19935 17663
rect 20177 17629 20211 17663
rect 20637 17629 20671 17663
rect 21097 17629 21131 17663
rect 3801 17561 3835 17595
rect 4813 17561 4847 17595
rect 6938 17561 6972 17595
rect 9220 17561 9254 17595
rect 12725 17561 12759 17595
rect 16589 17561 16623 17595
rect 18622 17561 18656 17595
rect 1501 17493 1535 17527
rect 2421 17493 2455 17527
rect 2881 17493 2915 17527
rect 4905 17493 4939 17527
rect 5549 17493 5583 17527
rect 5825 17493 5859 17527
rect 7481 17493 7515 17527
rect 11989 17493 12023 17527
rect 12265 17493 12299 17527
rect 12633 17493 12667 17527
rect 14381 17493 14415 17527
rect 14473 17493 14507 17527
rect 14841 17493 14875 17527
rect 15577 17493 15611 17527
rect 16129 17493 16163 17527
rect 16497 17493 16531 17527
rect 17509 17493 17543 17527
rect 20821 17493 20855 17527
rect 21281 17493 21315 17527
rect 2421 17289 2455 17323
rect 3893 17289 3927 17323
rect 4997 17289 5031 17323
rect 5733 17289 5767 17323
rect 6377 17289 6411 17323
rect 6929 17289 6963 17323
rect 8217 17289 8251 17323
rect 8677 17289 8711 17323
rect 9137 17289 9171 17323
rect 10793 17289 10827 17323
rect 11989 17289 12023 17323
rect 12357 17289 12391 17323
rect 14381 17289 14415 17323
rect 14749 17289 14783 17323
rect 15117 17289 15151 17323
rect 15209 17289 15243 17323
rect 16681 17289 16715 17323
rect 18153 17289 18187 17323
rect 20085 17289 20119 17323
rect 3433 17221 3467 17255
rect 5641 17221 5675 17255
rect 19288 17221 19322 17255
rect 1685 17153 1719 17187
rect 2145 17153 2179 17187
rect 2605 17153 2639 17187
rect 3525 17153 3559 17187
rect 4629 17153 4663 17187
rect 7297 17153 7331 17187
rect 8309 17153 8343 17187
rect 9505 17153 9539 17187
rect 11713 17153 11747 17187
rect 12449 17153 12483 17187
rect 13369 17153 13403 17187
rect 14013 17153 14047 17187
rect 17049 17153 17083 17187
rect 19533 17153 19567 17187
rect 19901 17153 19935 17187
rect 20637 17153 20671 17187
rect 21097 17153 21131 17187
rect 3341 17085 3375 17119
rect 4445 17085 4479 17119
rect 4537 17085 4571 17119
rect 5825 17085 5859 17119
rect 7389 17085 7423 17119
rect 7481 17085 7515 17119
rect 8125 17085 8159 17119
rect 9597 17085 9631 17119
rect 9689 17085 9723 17119
rect 10609 17085 10643 17119
rect 10701 17085 10735 17119
rect 12633 17085 12667 17119
rect 13829 17085 13863 17119
rect 13921 17085 13955 17119
rect 15393 17085 15427 17119
rect 17141 17085 17175 17119
rect 17233 17085 17267 17119
rect 1501 17017 1535 17051
rect 5273 17017 5307 17051
rect 1961 16949 1995 16983
rect 11161 16949 11195 16983
rect 17693 16949 17727 16983
rect 20821 16949 20855 16983
rect 21281 16949 21315 16983
rect 5825 16745 5859 16779
rect 8585 16745 8619 16779
rect 8953 16745 8987 16779
rect 10609 16745 10643 16779
rect 13737 16745 13771 16779
rect 14841 16745 14875 16779
rect 16405 16745 16439 16779
rect 18429 16745 18463 16779
rect 20361 16745 20395 16779
rect 20821 16745 20855 16779
rect 8217 16677 8251 16711
rect 16037 16677 16071 16711
rect 17417 16677 17451 16711
rect 2881 16609 2915 16643
rect 2973 16609 3007 16643
rect 3801 16609 3835 16643
rect 4445 16609 4479 16643
rect 7297 16609 7331 16643
rect 10333 16609 10367 16643
rect 11529 16609 11563 16643
rect 13277 16609 13311 16643
rect 14289 16609 14323 16643
rect 15117 16609 15151 16643
rect 16957 16609 16991 16643
rect 17877 16609 17911 16643
rect 17969 16609 18003 16643
rect 1685 16541 1719 16575
rect 1961 16541 1995 16575
rect 3065 16541 3099 16575
rect 6101 16541 6135 16575
rect 6745 16541 6779 16575
rect 7389 16541 7423 16575
rect 11713 16541 11747 16575
rect 14381 16541 14415 16575
rect 16773 16541 16807 16575
rect 19257 16541 19291 16575
rect 19901 16541 19935 16575
rect 20177 16541 20211 16575
rect 20637 16541 20671 16575
rect 21097 16541 21131 16575
rect 4712 16473 4746 16507
rect 10088 16473 10122 16507
rect 11621 16473 11655 16507
rect 1501 16405 1535 16439
rect 2145 16405 2179 16439
rect 3433 16405 3467 16439
rect 7481 16405 7515 16439
rect 7849 16405 7883 16439
rect 12081 16405 12115 16439
rect 14473 16405 14507 16439
rect 16865 16405 16899 16439
rect 17785 16405 17819 16439
rect 18797 16405 18831 16439
rect 21281 16405 21315 16439
rect 1961 16201 1995 16235
rect 2605 16201 2639 16235
rect 8033 16201 8067 16235
rect 11529 16201 11563 16235
rect 19441 16201 19475 16235
rect 20177 16201 20211 16235
rect 3985 16133 4019 16167
rect 17233 16133 17267 16167
rect 1685 16065 1719 16099
rect 2145 16065 2179 16099
rect 2421 16065 2455 16099
rect 8401 16065 8435 16099
rect 9137 16065 9171 16099
rect 11897 16065 11931 16099
rect 14565 16065 14599 16099
rect 15209 16065 15243 16099
rect 17509 16065 17543 16099
rect 17776 16065 17810 16099
rect 19993 16065 20027 16099
rect 20637 16065 20671 16099
rect 21097 16065 21131 16099
rect 3249 15997 3283 16031
rect 3709 15997 3743 16031
rect 4997 15997 5031 16031
rect 7297 15997 7331 16031
rect 7757 15997 7791 16031
rect 10241 15997 10275 16031
rect 11989 15997 12023 16031
rect 12173 15997 12207 16031
rect 14657 15997 14691 16031
rect 14749 15997 14783 16031
rect 2973 15929 3007 15963
rect 5549 15929 5583 15963
rect 6469 15929 6503 15963
rect 20821 15929 20855 15963
rect 1501 15861 1535 15895
rect 4353 15861 4387 15895
rect 5825 15861 5859 15895
rect 7021 15861 7055 15895
rect 8769 15861 8803 15895
rect 9505 15861 9539 15895
rect 9873 15861 9907 15895
rect 10701 15861 10735 15895
rect 11069 15861 11103 15895
rect 13829 15861 13863 15895
rect 14197 15861 14231 15895
rect 15853 15861 15887 15895
rect 16221 15861 16255 15895
rect 16865 15861 16899 15895
rect 18889 15861 18923 15895
rect 21281 15861 21315 15895
rect 2421 15657 2455 15691
rect 3341 15657 3375 15691
rect 7573 15657 7607 15691
rect 10333 15657 10367 15691
rect 12817 15657 12851 15691
rect 18797 15657 18831 15691
rect 19901 15657 19935 15691
rect 16957 15589 16991 15623
rect 18429 15589 18463 15623
rect 14197 15521 14231 15555
rect 15117 15521 15151 15555
rect 1685 15453 1719 15487
rect 1961 15453 1995 15487
rect 2605 15453 2639 15487
rect 3801 15453 3835 15487
rect 7297 15453 7331 15487
rect 7941 15453 7975 15487
rect 9689 15453 9723 15487
rect 11437 15453 11471 15487
rect 11704 15453 11738 15487
rect 14473 15453 14507 15487
rect 15577 15453 15611 15487
rect 18061 15453 18095 15487
rect 19717 15453 19751 15487
rect 20177 15453 20211 15487
rect 20637 15453 20671 15487
rect 21097 15453 21131 15487
rect 4046 15385 4080 15419
rect 5549 15385 5583 15419
rect 7030 15385 7064 15419
rect 9321 15385 9355 15419
rect 15844 15385 15878 15419
rect 17417 15385 17451 15419
rect 1501 15317 1535 15351
rect 2145 15317 2179 15351
rect 2973 15317 3007 15351
rect 5181 15317 5215 15351
rect 5917 15317 5951 15351
rect 8585 15317 8619 15351
rect 8953 15317 8987 15351
rect 10609 15317 10643 15351
rect 14381 15317 14415 15351
rect 14841 15317 14875 15351
rect 17693 15317 17727 15351
rect 19441 15317 19475 15351
rect 20361 15317 20395 15351
rect 20821 15317 20855 15351
rect 21281 15317 21315 15351
rect 5825 15113 5859 15147
rect 9321 15113 9355 15147
rect 13369 15113 13403 15147
rect 15025 15113 15059 15147
rect 15669 15113 15703 15147
rect 16037 15113 16071 15147
rect 18061 15113 18095 15147
rect 19717 15113 19751 15147
rect 20545 15113 20579 15147
rect 8208 15045 8242 15079
rect 13912 15045 13946 15079
rect 1685 14977 1719 15011
rect 2145 14977 2179 15011
rect 3729 14977 3763 15011
rect 5181 14977 5215 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 10710 14977 10744 15011
rect 11989 14977 12023 15011
rect 12256 14977 12290 15011
rect 13645 14977 13679 15011
rect 16681 14977 16715 15011
rect 16948 14977 16982 15011
rect 18705 14977 18739 15011
rect 20361 14977 20395 15011
rect 21097 14977 21131 15011
rect 3985 14909 4019 14943
rect 7021 14909 7055 14943
rect 7941 14909 7975 14943
rect 10977 14909 11011 14943
rect 15393 14909 15427 14943
rect 15577 14909 15611 14943
rect 18521 14909 18555 14943
rect 18613 14909 18647 14943
rect 19809 14909 19843 14943
rect 19901 14909 19935 14943
rect 4261 14841 4295 14875
rect 6377 14841 6411 14875
rect 19073 14841 19107 14875
rect 1501 14773 1535 14807
rect 1961 14773 1995 14807
rect 2605 14773 2639 14807
rect 4629 14773 4663 14807
rect 7481 14773 7515 14807
rect 9597 14773 9631 14807
rect 19349 14773 19383 14807
rect 21281 14773 21315 14807
rect 1961 14569 1995 14603
rect 2697 14569 2731 14603
rect 7941 14569 7975 14603
rect 12173 14569 12207 14603
rect 14841 14569 14875 14603
rect 17141 14569 17175 14603
rect 18889 14569 18923 14603
rect 19533 14569 19567 14603
rect 6193 14501 6227 14535
rect 17417 14501 17451 14535
rect 17785 14501 17819 14535
rect 3341 14433 3375 14467
rect 4353 14433 4387 14467
rect 6561 14433 6595 14467
rect 11621 14433 11655 14467
rect 14289 14433 14323 14467
rect 18245 14433 18279 14467
rect 18429 14433 18463 14467
rect 19993 14433 20027 14467
rect 20177 14433 20211 14467
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 9137 14365 9171 14399
rect 11161 14365 11195 14399
rect 11805 14365 11839 14399
rect 13737 14365 13771 14399
rect 15761 14365 15795 14399
rect 20637 14365 20671 14399
rect 21097 14365 21131 14399
rect 4261 14297 4295 14331
rect 5181 14297 5215 14331
rect 6828 14297 6862 14331
rect 9404 14297 9438 14331
rect 14473 14297 14507 14331
rect 16028 14297 16062 14331
rect 18521 14297 18555 14331
rect 19901 14297 19935 14331
rect 1501 14229 1535 14263
rect 3065 14229 3099 14263
rect 3157 14229 3191 14263
rect 3801 14229 3835 14263
rect 4169 14229 4203 14263
rect 4813 14229 4847 14263
rect 5733 14229 5767 14263
rect 8217 14229 8251 14263
rect 10517 14229 10551 14263
rect 11713 14229 11747 14263
rect 13369 14229 13403 14263
rect 14381 14229 14415 14263
rect 15485 14229 15519 14263
rect 20821 14229 20855 14263
rect 21281 14229 21315 14263
rect 3157 14025 3191 14059
rect 4721 14025 4755 14059
rect 6009 14025 6043 14059
rect 7481 14025 7515 14059
rect 8217 14025 8251 14059
rect 8585 14025 8619 14059
rect 11805 14025 11839 14059
rect 11897 14025 11931 14059
rect 12265 14025 12299 14059
rect 14473 14025 14507 14059
rect 16865 14025 16899 14059
rect 17601 14025 17635 14059
rect 18429 14025 18463 14059
rect 18797 14025 18831 14059
rect 19073 14025 19107 14059
rect 19533 14025 19567 14059
rect 20085 14025 20119 14059
rect 20545 14025 20579 14059
rect 21281 14025 21315 14059
rect 11069 13957 11103 13991
rect 14933 13957 14967 13991
rect 17233 13957 17267 13991
rect 20453 13957 20487 13991
rect 1685 13889 1719 13923
rect 2789 13889 2823 13923
rect 3617 13889 3651 13923
rect 4629 13889 4663 13923
rect 5549 13889 5583 13923
rect 5641 13889 5675 13923
rect 8953 13889 8987 13923
rect 9965 13889 9999 13923
rect 10057 13889 10091 13923
rect 10609 13889 10643 13923
rect 14197 13889 14231 13923
rect 14841 13889 14875 13923
rect 16313 13889 16347 13923
rect 19441 13889 19475 13923
rect 21097 13889 21131 13923
rect 2145 13821 2179 13855
rect 2605 13821 2639 13855
rect 2697 13821 2731 13855
rect 3433 13821 3467 13855
rect 4813 13821 4847 13855
rect 5457 13821 5491 13855
rect 6469 13821 6503 13855
rect 6745 13821 6779 13855
rect 7205 13821 7239 13855
rect 7389 13821 7423 13855
rect 9045 13821 9079 13855
rect 9137 13821 9171 13855
rect 10149 13821 10183 13855
rect 11713 13821 11747 13855
rect 12541 13821 12575 13855
rect 13093 13821 13127 13855
rect 13461 13821 13495 13855
rect 13829 13821 13863 13855
rect 15025 13821 15059 13855
rect 16037 13821 16071 13855
rect 18153 13821 18187 13855
rect 18337 13821 18371 13855
rect 19625 13821 19659 13855
rect 20637 13821 20671 13855
rect 1501 13753 1535 13787
rect 4261 13685 4295 13719
rect 7849 13685 7883 13719
rect 9597 13685 9631 13719
rect 3065 13481 3099 13515
rect 3801 13481 3835 13515
rect 4997 13481 5031 13515
rect 7297 13481 7331 13515
rect 9229 13481 9263 13515
rect 10425 13481 10459 13515
rect 16957 13481 16991 13515
rect 18429 13481 18463 13515
rect 18889 13413 18923 13447
rect 20545 13413 20579 13447
rect 2513 13345 2547 13379
rect 4353 13345 4387 13379
rect 7757 13345 7791 13379
rect 7849 13345 7883 13379
rect 9689 13345 9723 13379
rect 9781 13345 9815 13379
rect 12265 13345 12299 13379
rect 17877 13345 17911 13379
rect 19809 13345 19843 13379
rect 1685 13277 1719 13311
rect 2697 13277 2731 13311
rect 4169 13277 4203 13311
rect 7021 13277 7055 13311
rect 11253 13277 11287 13311
rect 14105 13277 14139 13311
rect 18705 13277 18739 13311
rect 21097 13277 21131 13311
rect 5273 13209 5307 13243
rect 15025 13209 15059 13243
rect 15669 13209 15703 13243
rect 18061 13209 18095 13243
rect 19625 13209 19659 13243
rect 20361 13209 20395 13243
rect 1501 13141 1535 13175
rect 1961 13141 1995 13175
rect 2605 13141 2639 13175
rect 3341 13141 3375 13175
rect 4261 13141 4295 13175
rect 7665 13141 7699 13175
rect 8309 13141 8343 13175
rect 9597 13141 9631 13175
rect 10793 13141 10827 13175
rect 11529 13141 11563 13175
rect 11897 13141 11931 13175
rect 12725 13141 12759 13175
rect 13277 13141 13311 13175
rect 13645 13141 13679 13175
rect 14749 13141 14783 13175
rect 17969 13141 18003 13175
rect 19257 13141 19291 13175
rect 19717 13141 19751 13175
rect 21281 13141 21315 13175
rect 2513 12937 2547 12971
rect 2881 12937 2915 12971
rect 3893 12937 3927 12971
rect 4169 12937 4203 12971
rect 4629 12937 4663 12971
rect 6377 12937 6411 12971
rect 6745 12937 6779 12971
rect 10057 12937 10091 12971
rect 10425 12937 10459 12971
rect 10517 12937 10551 12971
rect 11069 12937 11103 12971
rect 11989 12937 12023 12971
rect 15945 12937 15979 12971
rect 16957 12937 16991 12971
rect 17417 12937 17451 12971
rect 18153 12937 18187 12971
rect 19441 12937 19475 12971
rect 20453 12937 20487 12971
rect 4537 12869 4571 12903
rect 7389 12869 7423 12903
rect 7849 12869 7883 12903
rect 13001 12869 13035 12903
rect 15485 12869 15519 12903
rect 18061 12869 18095 12903
rect 20821 12869 20855 12903
rect 20913 12869 20947 12903
rect 1685 12801 1719 12835
rect 2421 12801 2455 12835
rect 3525 12801 3559 12835
rect 15577 12801 15611 12835
rect 17049 12801 17083 12835
rect 18981 12801 19015 12835
rect 19809 12801 19843 12835
rect 2329 12733 2363 12767
rect 3249 12733 3283 12767
rect 3433 12733 3467 12767
rect 4813 12733 4847 12767
rect 5733 12733 5767 12767
rect 6009 12733 6043 12767
rect 6837 12733 6871 12767
rect 7021 12733 7055 12767
rect 10609 12733 10643 12767
rect 11805 12733 11839 12767
rect 11897 12733 11931 12767
rect 15393 12733 15427 12767
rect 16865 12733 16899 12767
rect 18245 12733 18279 12767
rect 19901 12733 19935 12767
rect 20085 12733 20119 12767
rect 21005 12733 21039 12767
rect 1869 12665 1903 12699
rect 19165 12665 19199 12699
rect 9137 12597 9171 12631
rect 12357 12597 12391 12631
rect 12725 12597 12759 12631
rect 14289 12597 14323 12631
rect 16221 12597 16255 12631
rect 17693 12597 17727 12631
rect 4721 12393 4755 12427
rect 7021 12393 7055 12427
rect 7389 12393 7423 12427
rect 8585 12393 8619 12427
rect 13737 12393 13771 12427
rect 16221 12393 16255 12427
rect 5733 12325 5767 12359
rect 19441 12325 19475 12359
rect 5273 12257 5307 12291
rect 6285 12257 6319 12291
rect 7941 12257 7975 12291
rect 9137 12257 9171 12291
rect 10149 12257 10183 12291
rect 10241 12257 10275 12291
rect 18705 12257 18739 12291
rect 20085 12257 20119 12291
rect 3433 12189 3467 12223
rect 6101 12189 6135 12223
rect 7757 12189 7791 12223
rect 10701 12189 10735 12223
rect 12357 12189 12391 12223
rect 14841 12189 14875 12223
rect 15097 12189 15131 12223
rect 17877 12189 17911 12223
rect 20637 12189 20671 12223
rect 1593 12121 1627 12155
rect 1777 12121 1811 12155
rect 3166 12121 3200 12155
rect 3801 12121 3835 12155
rect 4445 12121 4479 12155
rect 10968 12121 11002 12155
rect 12624 12121 12658 12155
rect 17632 12121 17666 12155
rect 18613 12121 18647 12155
rect 19809 12121 19843 12155
rect 2053 12053 2087 12087
rect 5089 12053 5123 12087
rect 5181 12053 5215 12087
rect 6193 12053 6227 12087
rect 7849 12053 7883 12087
rect 9689 12053 9723 12087
rect 10057 12053 10091 12087
rect 12081 12053 12115 12087
rect 14289 12053 14323 12087
rect 16497 12053 16531 12087
rect 18153 12053 18187 12087
rect 18521 12053 18555 12087
rect 19901 12053 19935 12087
rect 21281 12053 21315 12087
rect 3065 11849 3099 11883
rect 5641 11849 5675 11883
rect 6469 11849 6503 11883
rect 7205 11849 7239 11883
rect 9045 11849 9079 11883
rect 9505 11849 9539 11883
rect 12725 11849 12759 11883
rect 13369 11849 13403 11883
rect 14105 11849 14139 11883
rect 14473 11849 14507 11883
rect 15577 11849 15611 11883
rect 16957 11849 16991 11883
rect 17325 11849 17359 11883
rect 17417 11849 17451 11883
rect 21005 11849 21039 11883
rect 21097 11849 21131 11883
rect 1869 11781 1903 11815
rect 12357 11781 12391 11815
rect 16313 11781 16347 11815
rect 20269 11781 20303 11815
rect 1685 11713 1719 11747
rect 2697 11713 2731 11747
rect 3341 11713 3375 11747
rect 3801 11713 3835 11747
rect 4261 11713 4295 11747
rect 4528 11713 4562 11747
rect 7573 11713 7607 11747
rect 7665 11713 7699 11747
rect 9413 11713 9447 11747
rect 10425 11713 10459 11747
rect 15485 11713 15519 11747
rect 18337 11713 18371 11747
rect 18613 11713 18647 11747
rect 19073 11713 19107 11747
rect 20085 11713 20119 11747
rect 2421 11645 2455 11679
rect 2605 11645 2639 11679
rect 5917 11645 5951 11679
rect 6929 11645 6963 11679
rect 7757 11645 7791 11679
rect 9597 11645 9631 11679
rect 10241 11645 10275 11679
rect 10333 11645 10367 11679
rect 12173 11645 12207 11679
rect 12265 11645 12299 11679
rect 13093 11645 13127 11679
rect 13277 11645 13311 11679
rect 14565 11645 14599 11679
rect 14749 11645 14783 11679
rect 15669 11645 15703 11679
rect 17509 11645 17543 11679
rect 21189 11645 21223 11679
rect 8309 11577 8343 11611
rect 10793 11577 10827 11611
rect 15117 11577 15151 11611
rect 18797 11577 18831 11611
rect 3525 11509 3559 11543
rect 8585 11509 8619 11543
rect 11161 11509 11195 11543
rect 11713 11509 11747 11543
rect 13737 11509 13771 11543
rect 19717 11509 19751 11543
rect 20637 11509 20671 11543
rect 1685 11305 1719 11339
rect 2513 11305 2547 11339
rect 9781 11305 9815 11339
rect 10241 11305 10275 11339
rect 11069 11305 11103 11339
rect 12265 11305 12299 11339
rect 20637 11305 20671 11339
rect 21189 11305 21223 11339
rect 2145 11237 2179 11271
rect 4813 11237 4847 11271
rect 5917 11237 5951 11271
rect 7113 11237 7147 11271
rect 16681 11237 16715 11271
rect 3157 11169 3191 11203
rect 5365 11169 5399 11203
rect 6469 11169 6503 11203
rect 8493 11169 8527 11203
rect 9229 11169 9263 11203
rect 15853 11169 15887 11203
rect 18245 11169 18279 11203
rect 1501 11101 1535 11135
rect 1961 11101 1995 11135
rect 2881 11101 2915 11135
rect 3893 11101 3927 11135
rect 4537 11101 4571 11135
rect 5181 11101 5215 11135
rect 9413 11101 9447 11135
rect 15597 11101 15631 11135
rect 17325 11101 17359 11135
rect 19257 11101 19291 11135
rect 19524 11101 19558 11135
rect 21281 11101 21315 11135
rect 2973 11033 3007 11067
rect 6285 11033 6319 11067
rect 8226 11033 8260 11067
rect 9321 11033 9355 11067
rect 10609 11033 10643 11067
rect 13553 11033 13587 11067
rect 14197 11033 14231 11067
rect 16129 11033 16163 11067
rect 18061 11033 18095 11067
rect 18705 11033 18739 11067
rect 5273 10965 5307 10999
rect 6377 10965 6411 10999
rect 11345 10965 11379 10999
rect 14473 10965 14507 10999
rect 16957 10965 16991 10999
rect 17693 10965 17727 10999
rect 18153 10965 18187 10999
rect 2145 10761 2179 10795
rect 2513 10761 2547 10795
rect 2881 10761 2915 10795
rect 3801 10761 3835 10795
rect 6745 10761 6779 10795
rect 7113 10761 7147 10795
rect 7205 10761 7239 10795
rect 11897 10761 11931 10795
rect 12265 10761 12299 10795
rect 14841 10761 14875 10795
rect 17049 10761 17083 10795
rect 4936 10693 4970 10727
rect 8401 10693 8435 10727
rect 9505 10693 9539 10727
rect 17960 10693 17994 10727
rect 21128 10693 21162 10727
rect 1685 10625 1719 10659
rect 2973 10625 3007 10659
rect 5641 10625 5675 10659
rect 7757 10625 7791 10659
rect 10793 10625 10827 10659
rect 11805 10625 11839 10659
rect 13093 10625 13127 10659
rect 14749 10625 14783 10659
rect 3157 10557 3191 10591
rect 5181 10557 5215 10591
rect 7297 10557 7331 10591
rect 9137 10557 9171 10591
rect 9965 10557 9999 10591
rect 10517 10557 10551 10591
rect 10701 10557 10735 10591
rect 11621 10557 11655 10591
rect 15025 10557 15059 10591
rect 15669 10557 15703 10591
rect 17141 10557 17175 10591
rect 17325 10557 17359 10591
rect 17693 10557 17727 10591
rect 19717 10557 19751 10591
rect 21373 10557 21407 10591
rect 1869 10489 1903 10523
rect 6469 10489 6503 10523
rect 12817 10489 12851 10523
rect 14105 10489 14139 10523
rect 5457 10421 5491 10455
rect 5917 10421 5951 10455
rect 8861 10421 8895 10455
rect 11161 10421 11195 10455
rect 13737 10421 13771 10455
rect 14381 10421 14415 10455
rect 15945 10421 15979 10455
rect 16681 10421 16715 10455
rect 19073 10421 19107 10455
rect 19993 10421 20027 10455
rect 2145 10217 2179 10251
rect 4905 10217 4939 10251
rect 5457 10217 5491 10251
rect 6469 10217 6503 10251
rect 9781 10217 9815 10251
rect 11437 10217 11471 10251
rect 17785 10217 17819 10251
rect 19533 10217 19567 10251
rect 3065 10149 3099 10183
rect 13737 10149 13771 10183
rect 1869 10081 1903 10115
rect 6009 10081 6043 10115
rect 7021 10081 7055 10115
rect 8033 10081 8067 10115
rect 9229 10081 9263 10115
rect 9321 10081 9355 10115
rect 16313 10081 16347 10115
rect 17325 10081 17359 10115
rect 18337 10081 18371 10115
rect 20545 10081 20579 10115
rect 21097 10081 21131 10115
rect 2329 10013 2363 10047
rect 2881 10013 2915 10047
rect 3801 10013 3835 10047
rect 4721 10013 4755 10047
rect 6929 10013 6963 10047
rect 9413 10013 9447 10047
rect 10057 10013 10091 10047
rect 12357 10013 12391 10047
rect 12624 10013 12658 10047
rect 15485 10013 15519 10047
rect 18889 10013 18923 10047
rect 19625 10013 19659 10047
rect 20361 10013 20395 10047
rect 21281 10013 21315 10047
rect 1685 9945 1719 9979
rect 5917 9945 5951 9979
rect 8493 9945 8527 9979
rect 10302 9945 10336 9979
rect 15218 9945 15252 9979
rect 17141 9945 17175 9979
rect 17233 9945 17267 9979
rect 18153 9945 18187 9979
rect 20453 9945 20487 9979
rect 3433 9877 3467 9911
rect 4445 9877 4479 9911
rect 5825 9877 5859 9911
rect 6837 9877 6871 9911
rect 7481 9877 7515 9911
rect 7849 9877 7883 9911
rect 7941 9877 7975 9911
rect 11989 9877 12023 9911
rect 14105 9877 14139 9911
rect 15761 9877 15795 9911
rect 16129 9877 16163 9911
rect 16221 9877 16255 9911
rect 16773 9877 16807 9911
rect 18245 9877 18279 9911
rect 19993 9877 20027 9911
rect 8677 9673 8711 9707
rect 8953 9673 8987 9707
rect 14105 9673 14139 9707
rect 14749 9673 14783 9707
rect 15761 9673 15795 9707
rect 15853 9673 15887 9707
rect 18153 9673 18187 9707
rect 4252 9605 4286 9639
rect 8217 9605 8251 9639
rect 14657 9605 14691 9639
rect 19257 9605 19291 9639
rect 1593 9537 1627 9571
rect 2053 9537 2087 9571
rect 2320 9537 2354 9571
rect 3985 9537 4019 9571
rect 6377 9537 6411 9571
rect 7297 9537 7331 9571
rect 8309 9537 8343 9571
rect 10077 9537 10111 9571
rect 10701 9537 10735 9571
rect 11713 9537 11747 9571
rect 11980 9537 12014 9571
rect 13461 9537 13495 9571
rect 16773 9537 16807 9571
rect 17040 9537 17074 9571
rect 18613 9537 18647 9571
rect 19349 9537 19383 9571
rect 21106 9537 21140 9571
rect 5641 9469 5675 9503
rect 7389 9469 7423 9503
rect 7481 9469 7515 9503
rect 8125 9469 8159 9503
rect 10333 9469 10367 9503
rect 14473 9469 14507 9503
rect 16037 9469 16071 9503
rect 19165 9469 19199 9503
rect 21373 9469 21407 9503
rect 6561 9401 6595 9435
rect 6929 9401 6963 9435
rect 15117 9401 15151 9435
rect 15393 9401 15427 9435
rect 18429 9401 18463 9435
rect 1685 9333 1719 9367
rect 3433 9333 3467 9367
rect 5365 9333 5399 9367
rect 11161 9333 11195 9367
rect 13093 9333 13127 9367
rect 19717 9333 19751 9367
rect 19993 9333 20027 9367
rect 3065 9129 3099 9163
rect 6653 9129 6687 9163
rect 7665 9129 7699 9163
rect 10517 9129 10551 9163
rect 11161 9129 11195 9163
rect 12081 9129 12115 9163
rect 21005 9129 21039 9163
rect 8309 9061 8343 9095
rect 17141 9061 17175 9095
rect 19349 9061 19383 9095
rect 2513 8993 2547 9027
rect 4537 8993 4571 9027
rect 4721 8993 4755 9027
rect 7021 8993 7055 9027
rect 9873 8993 9907 9027
rect 19809 8993 19843 9027
rect 19993 8993 20027 9027
rect 5273 8925 5307 8959
rect 5529 8925 5563 8959
rect 7297 8925 7331 8959
rect 10057 8925 10091 8959
rect 11437 8925 11471 8959
rect 14197 8925 14231 8959
rect 15485 8925 15519 8959
rect 15761 8925 15795 8959
rect 17417 8925 17451 8959
rect 18613 8925 18647 8959
rect 19717 8925 19751 8959
rect 20361 8925 20395 8959
rect 1685 8857 1719 8891
rect 1869 8857 1903 8891
rect 2605 8857 2639 8891
rect 10149 8857 10183 8891
rect 16028 8857 16062 8891
rect 18797 8857 18831 8891
rect 2697 8789 2731 8823
rect 3341 8789 3375 8823
rect 4077 8789 4111 8823
rect 4445 8789 4479 8823
rect 7205 8789 7239 8823
rect 8033 8789 8067 8823
rect 8953 8789 8987 8823
rect 9413 8789 9447 8823
rect 12725 8789 12759 8823
rect 13093 8789 13127 8823
rect 13645 8789 13679 8823
rect 14841 8789 14875 8823
rect 15301 8789 15335 8823
rect 18061 8789 18095 8823
rect 21373 8789 21407 8823
rect 1961 8585 1995 8619
rect 3617 8585 3651 8619
rect 3985 8585 4019 8619
rect 5273 8585 5307 8619
rect 6561 8585 6595 8619
rect 7573 8585 7607 8619
rect 9045 8585 9079 8619
rect 9781 8585 9815 8619
rect 10149 8585 10183 8619
rect 7205 8517 7239 8551
rect 8677 8517 8711 8551
rect 14648 8517 14682 8551
rect 16957 8517 16991 8551
rect 1501 8449 1535 8483
rect 1685 8449 1719 8483
rect 3085 8449 3119 8483
rect 5089 8449 5123 8483
rect 5549 8449 5583 8483
rect 6377 8449 6411 8483
rect 7113 8449 7147 8483
rect 7849 8449 7883 8483
rect 12541 8449 12575 8483
rect 13553 8449 13587 8483
rect 13645 8449 13679 8483
rect 14381 8449 14415 8483
rect 16129 8449 16163 8483
rect 17049 8449 17083 8483
rect 18061 8449 18095 8483
rect 18889 8449 18923 8483
rect 19156 8449 19190 8483
rect 20545 8449 20579 8483
rect 3341 8381 3375 8415
rect 4077 8381 4111 8415
rect 4169 8381 4203 8415
rect 4629 8381 4663 8415
rect 7021 8381 7055 8415
rect 8309 8381 8343 8415
rect 9597 8381 9631 8415
rect 9689 8381 9723 8415
rect 11897 8381 11931 8415
rect 12265 8381 12299 8415
rect 12449 8381 12483 8415
rect 13737 8381 13771 8415
rect 16773 8381 16807 8415
rect 18153 8381 18187 8415
rect 18245 8381 18279 8415
rect 21189 8381 21223 8415
rect 5733 8313 5767 8347
rect 12909 8313 12943 8347
rect 15761 8313 15795 8347
rect 16313 8313 16347 8347
rect 17417 8313 17451 8347
rect 8033 8245 8067 8279
rect 10517 8245 10551 8279
rect 11161 8245 11195 8279
rect 13185 8245 13219 8279
rect 17693 8245 17727 8279
rect 20269 8245 20303 8279
rect 2513 8041 2547 8075
rect 11253 8041 11287 8075
rect 12909 8041 12943 8075
rect 7297 7973 7331 8007
rect 14749 7973 14783 8007
rect 3065 7905 3099 7939
rect 4353 7905 4387 7939
rect 8953 7905 8987 7939
rect 13369 7905 13403 7939
rect 13461 7905 13495 7939
rect 17417 7905 17451 7939
rect 18153 7905 18187 7939
rect 18337 7905 18371 7939
rect 18705 7905 18739 7939
rect 20269 7905 20303 7939
rect 1961 7837 1995 7871
rect 2237 7837 2271 7871
rect 4169 7837 4203 7871
rect 7481 7837 7515 7871
rect 7757 7837 7791 7871
rect 9597 7837 9631 7871
rect 12633 7837 12667 7871
rect 14933 7837 14967 7871
rect 15393 7837 15427 7871
rect 15669 7837 15703 7871
rect 18061 7837 18095 7871
rect 19441 7837 19475 7871
rect 20177 7837 20211 7871
rect 20729 7837 20763 7871
rect 2973 7769 3007 7803
rect 5273 7769 5307 7803
rect 7021 7769 7055 7803
rect 9864 7769 9898 7803
rect 12388 7769 12422 7803
rect 2881 7701 2915 7735
rect 3801 7701 3835 7735
rect 4261 7701 4295 7735
rect 4813 7701 4847 7735
rect 8401 7701 8435 7735
rect 10977 7701 11011 7735
rect 13277 7701 13311 7735
rect 14473 7701 14507 7735
rect 15209 7701 15243 7735
rect 17693 7701 17727 7735
rect 19257 7701 19291 7735
rect 19717 7701 19751 7735
rect 20085 7701 20119 7735
rect 21373 7701 21407 7735
rect 2513 7497 2547 7531
rect 2881 7497 2915 7531
rect 4537 7497 4571 7531
rect 4629 7497 4663 7531
rect 4997 7497 5031 7531
rect 5641 7497 5675 7531
rect 6009 7497 6043 7531
rect 9413 7497 9447 7531
rect 10333 7497 10367 7531
rect 11897 7497 11931 7531
rect 12265 7497 12299 7531
rect 12817 7497 12851 7531
rect 18061 7497 18095 7531
rect 21189 7497 21223 7531
rect 1869 7429 1903 7463
rect 8300 7429 8334 7463
rect 11805 7429 11839 7463
rect 14206 7429 14240 7463
rect 20576 7429 20610 7463
rect 1685 7361 1719 7395
rect 2973 7361 3007 7395
rect 3709 7361 3743 7395
rect 6633 7361 6667 7395
rect 9689 7361 9723 7395
rect 14473 7361 14507 7395
rect 15393 7361 15427 7395
rect 15669 7361 15703 7395
rect 16681 7361 16715 7395
rect 16948 7361 16982 7395
rect 19165 7361 19199 7395
rect 21281 7361 21315 7395
rect 3157 7293 3191 7327
rect 4445 7293 4479 7327
rect 5365 7293 5399 7327
rect 5549 7293 5583 7327
rect 6377 7293 6411 7327
rect 8033 7293 8067 7327
rect 11069 7293 11103 7327
rect 11713 7293 11747 7327
rect 14933 7293 14967 7327
rect 16313 7293 16347 7327
rect 20821 7293 20855 7327
rect 13093 7225 13127 7259
rect 18521 7225 18555 7259
rect 2237 7157 2271 7191
rect 3525 7157 3559 7191
rect 7757 7157 7791 7191
rect 10609 7157 10643 7191
rect 15209 7157 15243 7191
rect 15853 7157 15887 7191
rect 19441 7157 19475 7191
rect 11069 6953 11103 6987
rect 16957 6953 16991 6987
rect 17417 6953 17451 6987
rect 8953 6885 8987 6919
rect 18061 6885 18095 6919
rect 2329 6817 2363 6851
rect 7021 6817 7055 6851
rect 8493 6817 8527 6851
rect 11345 6817 11379 6851
rect 12449 6817 12483 6851
rect 15117 6817 15151 6851
rect 1685 6749 1719 6783
rect 3249 6749 3283 6783
rect 4169 6749 4203 6783
rect 4629 6749 4663 6783
rect 6285 6749 6319 6783
rect 7205 6749 7239 6783
rect 10066 6749 10100 6783
rect 10333 6749 10367 6783
rect 11989 6749 12023 6783
rect 13093 6749 13127 6783
rect 13553 6749 13587 6783
rect 14105 6749 14139 6783
rect 15393 6749 15427 6783
rect 15853 6749 15887 6783
rect 16313 6749 16347 6783
rect 17233 6749 17267 6783
rect 18245 6749 18279 6783
rect 18797 6749 18831 6783
rect 19625 6749 19659 6783
rect 21106 6749 21140 6783
rect 21373 6749 21407 6783
rect 1869 6681 1903 6715
rect 2513 6681 2547 6715
rect 3893 6681 3927 6715
rect 4896 6681 4930 6715
rect 18613 6681 18647 6715
rect 19441 6681 19475 6715
rect 2421 6613 2455 6647
rect 2881 6613 2915 6647
rect 3433 6613 3467 6647
rect 4353 6613 4387 6647
rect 6009 6613 6043 6647
rect 6469 6613 6503 6647
rect 7113 6613 7147 6647
rect 7573 6613 7607 6647
rect 7849 6613 7883 6647
rect 8217 6613 8251 6647
rect 8309 6613 8343 6647
rect 10609 6613 10643 6647
rect 12817 6613 12851 6647
rect 13277 6613 13311 6647
rect 13737 6613 13771 6647
rect 14749 6613 14783 6647
rect 15577 6613 15611 6647
rect 16037 6613 16071 6647
rect 17693 6613 17727 6647
rect 19993 6613 20027 6647
rect 1869 6409 1903 6443
rect 2237 6409 2271 6443
rect 2513 6409 2547 6443
rect 2881 6409 2915 6443
rect 6009 6409 6043 6443
rect 6837 6409 6871 6443
rect 7665 6409 7699 6443
rect 7941 6409 7975 6443
rect 8861 6409 8895 6443
rect 9229 6409 9263 6443
rect 9321 6409 9355 6443
rect 10057 6409 10091 6443
rect 10701 6409 10735 6443
rect 13369 6409 13403 6443
rect 14657 6409 14691 6443
rect 17049 6409 17083 6443
rect 17693 6409 17727 6443
rect 19441 6409 19475 6443
rect 19901 6409 19935 6443
rect 20821 6409 20855 6443
rect 1777 6341 1811 6375
rect 2973 6341 3007 6375
rect 18061 6341 18095 6375
rect 3525 6273 3559 6307
rect 4813 6273 4847 6307
rect 5549 6273 5583 6307
rect 5641 6273 5675 6307
rect 7481 6273 7515 6307
rect 8125 6273 8159 6307
rect 8401 6273 8435 6307
rect 9873 6273 9907 6307
rect 10793 6273 10827 6307
rect 11897 6273 11931 6307
rect 12633 6273 12667 6307
rect 13461 6273 13495 6307
rect 15200 6273 15234 6307
rect 18889 6273 18923 6307
rect 19073 6273 19107 6307
rect 19809 6273 19843 6307
rect 1685 6205 1719 6239
rect 3065 6205 3099 6239
rect 5457 6205 5491 6239
rect 6929 6205 6963 6239
rect 7021 6205 7055 6239
rect 9505 6205 9539 6239
rect 10609 6205 10643 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 13277 6205 13311 6239
rect 14289 6205 14323 6239
rect 14933 6205 14967 6239
rect 17141 6205 17175 6239
rect 17233 6205 17267 6239
rect 18153 6205 18187 6239
rect 18337 6205 18371 6239
rect 19993 6205 20027 6239
rect 20913 6205 20947 6239
rect 21005 6205 21039 6239
rect 4537 6137 4571 6171
rect 8585 6137 8619 6171
rect 16313 6137 16347 6171
rect 4169 6069 4203 6103
rect 4997 6069 5031 6103
rect 6469 6069 6503 6103
rect 11161 6069 11195 6103
rect 11529 6069 11563 6103
rect 12817 6069 12851 6103
rect 13829 6069 13863 6103
rect 16681 6069 16715 6103
rect 20453 6069 20487 6103
rect 1685 5865 1719 5899
rect 5181 5865 5215 5899
rect 7113 5865 7147 5899
rect 9045 5865 9079 5899
rect 18889 5865 18923 5899
rect 20269 5865 20303 5899
rect 21281 5865 21315 5899
rect 5641 5797 5675 5831
rect 6101 5797 6135 5831
rect 7389 5797 7423 5831
rect 8309 5797 8343 5831
rect 11989 5797 12023 5831
rect 13737 5797 13771 5831
rect 15117 5797 15151 5831
rect 6469 5729 6503 5763
rect 6653 5729 6687 5763
rect 9505 5729 9539 5763
rect 9597 5729 9631 5763
rect 12357 5729 12391 5763
rect 14565 5729 14599 5763
rect 14657 5729 14691 5763
rect 15669 5729 15703 5763
rect 16221 5729 16255 5763
rect 16405 5729 16439 5763
rect 19809 5729 19843 5763
rect 20821 5729 20855 5763
rect 1593 5661 1627 5695
rect 2053 5661 2087 5695
rect 3801 5661 3835 5695
rect 5457 5661 5491 5695
rect 5917 5661 5951 5695
rect 7573 5661 7607 5695
rect 8033 5661 8067 5695
rect 8493 5661 8527 5695
rect 10333 5661 10367 5695
rect 10600 5661 10634 5695
rect 15485 5661 15519 5695
rect 17509 5661 17543 5695
rect 17776 5661 17810 5695
rect 19625 5661 19659 5695
rect 20637 5661 20671 5695
rect 2298 5593 2332 5627
rect 4068 5593 4102 5627
rect 12624 5593 12658 5627
rect 14473 5593 14507 5627
rect 16497 5593 16531 5627
rect 20729 5593 20763 5627
rect 3433 5525 3467 5559
rect 6745 5525 6779 5559
rect 7849 5525 7883 5559
rect 9413 5525 9447 5559
rect 11713 5525 11747 5559
rect 14105 5525 14139 5559
rect 15577 5525 15611 5559
rect 16865 5525 16899 5559
rect 17233 5525 17267 5559
rect 19257 5525 19291 5559
rect 19717 5525 19751 5559
rect 2421 5321 2455 5355
rect 2973 5321 3007 5355
rect 3065 5321 3099 5355
rect 3709 5321 3743 5355
rect 4077 5321 4111 5355
rect 6469 5321 6503 5355
rect 6929 5321 6963 5355
rect 10701 5321 10735 5355
rect 17417 5321 17451 5355
rect 18337 5321 18371 5355
rect 18705 5321 18739 5355
rect 20361 5321 20395 5355
rect 2053 5253 2087 5287
rect 5733 5253 5767 5287
rect 9597 5253 9631 5287
rect 10793 5253 10827 5287
rect 13001 5253 13035 5287
rect 14749 5253 14783 5287
rect 17049 5253 17083 5287
rect 4721 5185 4755 5219
rect 6837 5185 6871 5219
rect 7573 5185 7607 5219
rect 9873 5185 9907 5219
rect 11713 5185 11747 5219
rect 15209 5185 15243 5219
rect 15669 5185 15703 5219
rect 15945 5185 15979 5219
rect 18245 5185 18279 5219
rect 18981 5185 19015 5219
rect 19248 5185 19282 5219
rect 20637 5185 20671 5219
rect 1777 5117 1811 5151
rect 1961 5117 1995 5151
rect 2881 5117 2915 5151
rect 4169 5117 4203 5151
rect 4261 5117 4295 5151
rect 7021 5117 7055 5151
rect 10609 5117 10643 5151
rect 16865 5117 16899 5151
rect 16957 5117 16991 5151
rect 18153 5117 18187 5151
rect 10057 5049 10091 5083
rect 15485 5049 15519 5083
rect 3433 4981 3467 5015
rect 5365 4981 5399 5015
rect 5825 4981 5859 5015
rect 8309 4981 8343 5015
rect 11161 4981 11195 5015
rect 12357 4981 12391 5015
rect 12633 4981 12667 5015
rect 15025 4981 15059 5015
rect 16129 4981 16163 5015
rect 21281 4981 21315 5015
rect 2513 4777 2547 4811
rect 6285 4777 6319 4811
rect 10333 4777 10367 4811
rect 12909 4777 12943 4811
rect 13369 4777 13403 4811
rect 17233 4777 17267 4811
rect 17693 4777 17727 4811
rect 7205 4709 7239 4743
rect 18061 4709 18095 4743
rect 19441 4709 19475 4743
rect 2237 4641 2271 4675
rect 3065 4641 3099 4675
rect 4353 4641 4387 4675
rect 4445 4641 4479 4675
rect 5641 4641 5675 4675
rect 5825 4641 5859 4675
rect 7941 4641 7975 4675
rect 9413 4641 9447 4675
rect 9597 4641 9631 4675
rect 14105 4641 14139 4675
rect 21189 4641 21223 4675
rect 1961 4573 1995 4607
rect 2973 4573 3007 4607
rect 7021 4573 7055 4607
rect 7481 4573 7515 4607
rect 8585 4573 8619 4607
rect 10149 4573 10183 4607
rect 10609 4573 10643 4607
rect 11529 4573 11563 4607
rect 13185 4573 13219 4607
rect 14372 4573 14406 4607
rect 15761 4573 15795 4607
rect 16313 4573 16347 4607
rect 17417 4573 17451 4607
rect 18889 4573 18923 4607
rect 19257 4573 19291 4607
rect 20933 4573 20967 4607
rect 5549 4505 5583 4539
rect 6745 4505 6779 4539
rect 9321 4505 9355 4539
rect 11796 4505 11830 4539
rect 18245 4505 18279 4539
rect 2881 4437 2915 4471
rect 3893 4437 3927 4471
rect 4537 4437 4571 4471
rect 4905 4437 4939 4471
rect 5181 4437 5215 4471
rect 7665 4437 7699 4471
rect 8953 4437 8987 4471
rect 10793 4437 10827 4471
rect 11253 4437 11287 4471
rect 13737 4437 13771 4471
rect 15485 4437 15519 4471
rect 15945 4437 15979 4471
rect 16957 4437 16991 4471
rect 18705 4437 18739 4471
rect 19809 4437 19843 4471
rect 1501 4233 1535 4267
rect 3341 4233 3375 4267
rect 6745 4233 6779 4267
rect 8401 4233 8435 4267
rect 10701 4233 10735 4267
rect 11989 4233 12023 4267
rect 18061 4233 18095 4267
rect 4997 4165 5031 4199
rect 6653 4165 6687 4199
rect 20177 4165 20211 4199
rect 2614 4097 2648 4131
rect 3985 4097 4019 4131
rect 5825 4097 5859 4131
rect 7389 4097 7423 4131
rect 9413 4097 9447 4131
rect 10609 4097 10643 4131
rect 11529 4097 11563 4131
rect 12173 4097 12207 4131
rect 12449 4097 12483 4131
rect 13093 4097 13127 4131
rect 13553 4097 13587 4131
rect 14013 4097 14047 4131
rect 14473 4097 14507 4131
rect 14933 4097 14967 4131
rect 15200 4097 15234 4131
rect 16681 4097 16715 4131
rect 16948 4097 16982 4131
rect 18613 4097 18647 4131
rect 19165 4097 19199 4131
rect 20821 4097 20855 4131
rect 2881 4029 2915 4063
rect 3709 4029 3743 4063
rect 3893 4029 3927 4063
rect 5089 4029 5123 4063
rect 5181 4029 5215 4063
rect 6561 4029 6595 4063
rect 8493 4029 8527 4063
rect 8677 4029 8711 4063
rect 9137 4029 9171 4063
rect 9321 4029 9355 4063
rect 10885 4029 10919 4063
rect 20545 4029 20579 4063
rect 4629 3961 4663 3995
rect 6009 3961 6043 3995
rect 9781 3961 9815 3995
rect 12633 3961 12667 3995
rect 13277 3961 13311 3995
rect 18797 3961 18831 3995
rect 4353 3893 4387 3927
rect 7113 3893 7147 3927
rect 7573 3893 7607 3927
rect 8033 3893 8067 3927
rect 10241 3893 10275 3927
rect 11713 3893 11747 3927
rect 13737 3893 13771 3927
rect 14197 3893 14231 3927
rect 14657 3893 14691 3927
rect 16313 3893 16347 3927
rect 19349 3893 19383 3927
rect 20085 3893 20119 3927
rect 6561 3689 6595 3723
rect 8585 3689 8619 3723
rect 6285 3621 6319 3655
rect 13645 3621 13679 3655
rect 18245 3621 18279 3655
rect 1961 3553 1995 3587
rect 2237 3553 2271 3587
rect 3065 3553 3099 3587
rect 4353 3553 4387 3587
rect 4629 3553 4663 3587
rect 5733 3553 5767 3587
rect 7021 3553 7055 3587
rect 7113 3553 7147 3587
rect 7941 3553 7975 3587
rect 8125 3553 8159 3587
rect 11161 3553 11195 3587
rect 14841 3553 14875 3587
rect 16221 3553 16255 3587
rect 19441 3553 19475 3587
rect 20821 3553 20855 3587
rect 3341 3485 3375 3519
rect 5825 3485 5859 3519
rect 5917 3485 5951 3519
rect 10333 3485 10367 3519
rect 10977 3485 11011 3519
rect 11621 3485 11655 3519
rect 12173 3485 12207 3519
rect 12817 3485 12851 3519
rect 13185 3485 13219 3519
rect 14197 3485 14231 3519
rect 15025 3485 15059 3519
rect 16957 3485 16991 3519
rect 17509 3485 17543 3519
rect 18061 3485 18095 3519
rect 18613 3485 18647 3519
rect 19717 3485 19751 3519
rect 20545 3485 20579 3519
rect 4997 3417 5031 3451
rect 6929 3417 6963 3451
rect 8217 3417 8251 3451
rect 10088 3417 10122 3451
rect 5089 3349 5123 3383
rect 8953 3349 8987 3383
rect 10609 3349 10643 3383
rect 11069 3349 11103 3383
rect 11805 3349 11839 3383
rect 12357 3349 12391 3383
rect 12633 3349 12667 3383
rect 13369 3349 13403 3383
rect 14381 3349 14415 3383
rect 14933 3349 14967 3383
rect 15393 3349 15427 3383
rect 15669 3349 15703 3383
rect 16037 3349 16071 3383
rect 16129 3349 16163 3383
rect 17141 3349 17175 3383
rect 17693 3349 17727 3383
rect 18797 3349 18831 3383
rect 3985 3145 4019 3179
rect 5733 3145 5767 3179
rect 7481 3145 7515 3179
rect 9321 3145 9355 3179
rect 9689 3145 9723 3179
rect 10057 3145 10091 3179
rect 14105 3145 14139 3179
rect 15485 3145 15519 3179
rect 16129 3145 16163 3179
rect 2872 3077 2906 3111
rect 10149 3077 10183 3111
rect 15577 3077 15611 3111
rect 1961 3009 1995 3043
rect 2237 3009 2271 3043
rect 4620 3009 4654 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7665 3009 7699 3043
rect 8208 3009 8242 3043
rect 10977 3009 11011 3043
rect 11529 3009 11563 3043
rect 11989 3009 12023 3043
rect 12449 3009 12483 3043
rect 12909 3009 12943 3043
rect 13369 3009 13403 3043
rect 14289 3009 14323 3043
rect 14565 3009 14599 3043
rect 16681 3009 16715 3043
rect 17417 3009 17451 3043
rect 18061 3009 18095 3043
rect 18337 3009 18371 3043
rect 19717 3009 19751 3043
rect 19993 3009 20027 3043
rect 21097 3009 21131 3043
rect 2605 2941 2639 2975
rect 4353 2941 4387 2975
rect 7941 2941 7975 2975
rect 10241 2941 10275 2975
rect 15761 2941 15795 2975
rect 20729 2941 20763 2975
rect 11713 2873 11747 2907
rect 13093 2873 13127 2907
rect 11161 2805 11195 2839
rect 12173 2805 12207 2839
rect 12633 2805 12667 2839
rect 13553 2805 13587 2839
rect 14749 2805 14783 2839
rect 15117 2805 15151 2839
rect 16865 2805 16899 2839
rect 17601 2805 17635 2839
rect 18521 2805 18555 2839
rect 1593 2601 1627 2635
rect 6377 2601 6411 2635
rect 8401 2601 8435 2635
rect 9413 2601 9447 2635
rect 10057 2601 10091 2635
rect 11759 2601 11793 2635
rect 14841 2533 14875 2567
rect 15945 2533 15979 2567
rect 17417 2533 17451 2567
rect 18521 2533 18555 2567
rect 2973 2465 3007 2499
rect 5457 2465 5491 2499
rect 5733 2465 5767 2499
rect 7757 2465 7791 2499
rect 8033 2465 8067 2499
rect 10333 2465 10367 2499
rect 21097 2465 21131 2499
rect 2717 2397 2751 2431
rect 3249 2397 3283 2431
rect 4353 2397 4387 2431
rect 4629 2397 4663 2431
rect 7490 2397 7524 2431
rect 8585 2397 8619 2431
rect 8953 2397 8987 2431
rect 9597 2397 9631 2431
rect 9873 2397 9907 2431
rect 11529 2397 11563 2431
rect 12909 2397 12943 2431
rect 13461 2397 13495 2431
rect 14105 2397 14139 2431
rect 14657 2397 14691 2431
rect 15209 2397 15243 2431
rect 15761 2397 15795 2431
rect 16681 2397 16715 2431
rect 17233 2397 17267 2431
rect 17785 2397 17819 2431
rect 18337 2397 18371 2431
rect 19993 2397 20027 2431
rect 20269 2397 20303 2431
rect 21373 2397 21407 2431
rect 3433 2261 3467 2295
rect 9137 2261 9171 2295
rect 10563 2261 10597 2295
rect 13093 2261 13127 2295
rect 13645 2261 13679 2295
rect 14289 2261 14323 2295
rect 15393 2261 15427 2295
rect 16865 2261 16899 2295
rect 17969 2261 18003 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 1486 20584 1492 20596
rect 1447 20556 1492 20584
rect 1486 20544 1492 20556
rect 1544 20544 1550 20596
rect 2038 20584 2044 20596
rect 1999 20556 2044 20584
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 2958 20544 2964 20596
rect 3016 20584 3022 20596
rect 4249 20587 4307 20593
rect 4249 20584 4261 20587
rect 3016 20556 4261 20584
rect 3016 20544 3022 20556
rect 4249 20553 4261 20556
rect 4295 20553 4307 20587
rect 5169 20587 5227 20593
rect 5169 20584 5181 20587
rect 4249 20547 4307 20553
rect 4448 20556 5181 20584
rect 1673 20451 1731 20457
rect 1673 20417 1685 20451
rect 1719 20448 1731 20451
rect 2225 20451 2283 20457
rect 1719 20420 2176 20448
rect 1719 20417 1731 20420
rect 1673 20411 1731 20417
rect 2148 20244 2176 20420
rect 2225 20417 2237 20451
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 3237 20451 3295 20457
rect 2823 20420 3096 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 2240 20380 2268 20411
rect 2958 20380 2964 20392
rect 2240 20352 2964 20380
rect 2958 20340 2964 20352
rect 3016 20340 3022 20392
rect 2593 20315 2651 20321
rect 2593 20281 2605 20315
rect 2639 20312 2651 20315
rect 2774 20312 2780 20324
rect 2639 20284 2780 20312
rect 2639 20281 2651 20284
rect 2593 20275 2651 20281
rect 2774 20272 2780 20284
rect 2832 20272 2838 20324
rect 3068 20321 3096 20420
rect 3237 20417 3249 20451
rect 3283 20448 3295 20451
rect 3878 20448 3884 20460
rect 3283 20420 3884 20448
rect 3283 20417 3295 20420
rect 3237 20411 3295 20417
rect 3878 20408 3884 20420
rect 3936 20408 3942 20460
rect 4448 20457 4476 20556
rect 5169 20553 5181 20556
rect 5215 20584 5227 20587
rect 9950 20584 9956 20596
rect 5215 20556 9956 20584
rect 5215 20553 5227 20556
rect 5169 20547 5227 20553
rect 9950 20544 9956 20556
rect 10008 20544 10014 20596
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17497 20587 17555 20593
rect 17497 20584 17509 20587
rect 17276 20556 17509 20584
rect 17276 20544 17282 20556
rect 17497 20553 17509 20556
rect 17543 20553 17555 20587
rect 19610 20584 19616 20596
rect 19571 20556 19616 20584
rect 17497 20547 17555 20553
rect 19610 20544 19616 20556
rect 19668 20544 19674 20596
rect 20162 20584 20168 20596
rect 20123 20556 20168 20584
rect 20162 20544 20168 20556
rect 20220 20544 20226 20596
rect 3973 20451 4031 20457
rect 3973 20417 3985 20451
rect 4019 20417 4031 20451
rect 3973 20411 4031 20417
rect 4433 20451 4491 20457
rect 4433 20417 4445 20451
rect 4479 20417 4491 20451
rect 4433 20411 4491 20417
rect 3988 20380 4016 20411
rect 4522 20408 4528 20460
rect 4580 20448 4586 20460
rect 4709 20451 4767 20457
rect 4709 20448 4721 20451
rect 4580 20420 4721 20448
rect 4580 20408 4586 20420
rect 4709 20417 4721 20420
rect 4755 20417 4767 20451
rect 4709 20411 4767 20417
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5776 20420 5825 20448
rect 5776 20408 5782 20420
rect 5813 20417 5825 20420
rect 5859 20448 5871 20451
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 5859 20420 6377 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 17313 20451 17371 20457
rect 17313 20448 17325 20451
rect 10376 20420 17325 20448
rect 10376 20408 10382 20420
rect 17313 20417 17325 20420
rect 17359 20417 17371 20451
rect 17313 20411 17371 20417
rect 18417 20451 18475 20457
rect 18417 20417 18429 20451
rect 18463 20448 18475 20451
rect 18690 20448 18696 20460
rect 18463 20420 18696 20448
rect 18463 20417 18475 20420
rect 18417 20411 18475 20417
rect 18690 20408 18696 20420
rect 18748 20408 18754 20460
rect 18782 20408 18788 20460
rect 18840 20448 18846 20460
rect 19429 20451 19487 20457
rect 19429 20448 19441 20451
rect 18840 20420 19441 20448
rect 18840 20408 18846 20420
rect 19429 20417 19441 20420
rect 19475 20417 19487 20451
rect 19429 20411 19487 20417
rect 19518 20408 19524 20460
rect 19576 20448 19582 20460
rect 19981 20451 20039 20457
rect 19981 20448 19993 20451
rect 19576 20420 19993 20448
rect 19576 20408 19582 20420
rect 19981 20417 19993 20420
rect 20027 20417 20039 20451
rect 20530 20448 20536 20460
rect 20491 20420 20536 20448
rect 19981 20411 20039 20417
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 21085 20451 21143 20457
rect 21085 20417 21097 20451
rect 21131 20417 21143 20451
rect 21085 20411 21143 20417
rect 6546 20380 6552 20392
rect 3988 20352 6552 20380
rect 6546 20340 6552 20352
rect 6604 20380 6610 20392
rect 6733 20383 6791 20389
rect 6733 20380 6745 20383
rect 6604 20352 6745 20380
rect 6604 20340 6610 20352
rect 6733 20349 6745 20352
rect 6779 20349 6791 20383
rect 6733 20343 6791 20349
rect 20438 20340 20444 20392
rect 20496 20380 20502 20392
rect 21100 20380 21128 20411
rect 20496 20352 21128 20380
rect 20496 20340 20502 20352
rect 3053 20315 3111 20321
rect 3053 20281 3065 20315
rect 3099 20281 3111 20315
rect 3053 20275 3111 20281
rect 5997 20315 6055 20321
rect 5997 20281 6009 20315
rect 6043 20312 6055 20315
rect 11238 20312 11244 20324
rect 6043 20284 11244 20312
rect 6043 20281 6055 20284
rect 5997 20275 6055 20281
rect 11238 20272 11244 20284
rect 11296 20272 11302 20324
rect 20714 20312 20720 20324
rect 20675 20284 20720 20312
rect 20714 20272 20720 20284
rect 20772 20272 20778 20324
rect 3789 20247 3847 20253
rect 3789 20244 3801 20247
rect 2148 20216 3801 20244
rect 3789 20213 3801 20216
rect 3835 20213 3847 20247
rect 3789 20207 3847 20213
rect 4893 20247 4951 20253
rect 4893 20213 4905 20247
rect 4939 20244 4951 20247
rect 4982 20244 4988 20256
rect 4939 20216 4988 20244
rect 4939 20213 4951 20216
rect 4893 20207 4951 20213
rect 4982 20204 4988 20216
rect 5040 20204 5046 20256
rect 18046 20204 18052 20256
rect 18104 20244 18110 20256
rect 18877 20247 18935 20253
rect 18877 20244 18889 20247
rect 18104 20216 18889 20244
rect 18104 20204 18110 20216
rect 18877 20213 18889 20216
rect 18923 20213 18935 20247
rect 18877 20207 18935 20213
rect 21269 20247 21327 20253
rect 21269 20213 21281 20247
rect 21315 20244 21327 20247
rect 21358 20244 21364 20256
rect 21315 20216 21364 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 2593 20043 2651 20049
rect 2593 20009 2605 20043
rect 2639 20040 2651 20043
rect 2866 20040 2872 20052
rect 2639 20012 2872 20040
rect 2639 20009 2651 20012
rect 2593 20003 2651 20009
rect 2866 20000 2872 20012
rect 2924 20000 2930 20052
rect 7561 20043 7619 20049
rect 7561 20040 7573 20043
rect 3252 20012 7573 20040
rect 1673 19839 1731 19845
rect 1673 19805 1685 19839
rect 1719 19836 1731 19839
rect 2130 19836 2136 19848
rect 1719 19808 2136 19836
rect 1719 19805 1731 19808
rect 1673 19799 1731 19805
rect 2130 19796 2136 19808
rect 2188 19796 2194 19848
rect 2225 19839 2283 19845
rect 2225 19805 2237 19839
rect 2271 19836 2283 19839
rect 2498 19836 2504 19848
rect 2271 19808 2504 19836
rect 2271 19805 2283 19808
rect 2225 19799 2283 19805
rect 2498 19796 2504 19808
rect 2556 19796 2562 19848
rect 2774 19796 2780 19848
rect 2832 19836 2838 19848
rect 3252 19845 3280 20012
rect 7561 20009 7573 20012
rect 7607 20009 7619 20043
rect 10318 20040 10324 20052
rect 7561 20003 7619 20009
rect 8220 20012 10324 20040
rect 8220 19913 8248 20012
rect 10318 20000 10324 20012
rect 10376 20000 10382 20052
rect 18417 20043 18475 20049
rect 18417 20009 18429 20043
rect 18463 20040 18475 20043
rect 18782 20040 18788 20052
rect 18463 20012 18788 20040
rect 18463 20009 18475 20012
rect 18417 20003 18475 20009
rect 18782 20000 18788 20012
rect 18840 20000 18846 20052
rect 18877 20043 18935 20049
rect 18877 20009 18889 20043
rect 18923 20040 18935 20043
rect 19518 20040 19524 20052
rect 18923 20012 19524 20040
rect 18923 20009 18935 20012
rect 18877 20003 18935 20009
rect 19518 20000 19524 20012
rect 19576 20000 19582 20052
rect 19705 20043 19763 20049
rect 19705 20009 19717 20043
rect 19751 20040 19763 20043
rect 20530 20040 20536 20052
rect 19751 20012 20536 20040
rect 19751 20009 19763 20012
rect 19705 20003 19763 20009
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 20165 19975 20223 19981
rect 20165 19941 20177 19975
rect 20211 19972 20223 19975
rect 20254 19972 20260 19984
rect 20211 19944 20260 19972
rect 20211 19941 20223 19944
rect 20165 19935 20223 19941
rect 20254 19932 20260 19944
rect 20312 19932 20318 19984
rect 8205 19907 8263 19913
rect 8205 19873 8217 19907
rect 8251 19873 8263 19907
rect 8205 19867 8263 19873
rect 3237 19839 3295 19845
rect 2832 19808 2877 19836
rect 2832 19796 2838 19808
rect 3237 19805 3249 19839
rect 3283 19805 3295 19839
rect 3237 19799 3295 19805
rect 4338 19796 4344 19848
rect 4396 19836 4402 19848
rect 5169 19839 5227 19845
rect 5169 19836 5181 19839
rect 4396 19808 5181 19836
rect 4396 19796 4402 19808
rect 5169 19805 5181 19808
rect 5215 19805 5227 19839
rect 5169 19799 5227 19805
rect 5258 19796 5264 19848
rect 5316 19836 5322 19848
rect 5445 19839 5503 19845
rect 5445 19836 5457 19839
rect 5316 19808 5457 19836
rect 5316 19796 5322 19808
rect 5445 19805 5457 19808
rect 5491 19805 5503 19839
rect 5445 19799 5503 19805
rect 8941 19839 8999 19845
rect 8941 19805 8953 19839
rect 8987 19836 8999 19839
rect 9490 19836 9496 19848
rect 8987 19808 9496 19836
rect 8987 19805 8999 19808
rect 8941 19799 8999 19805
rect 9490 19796 9496 19808
rect 9548 19836 9554 19848
rect 11149 19839 11207 19845
rect 11149 19836 11161 19839
rect 9548 19808 11161 19836
rect 9548 19796 9554 19808
rect 11149 19805 11161 19808
rect 11195 19805 11207 19839
rect 11149 19799 11207 19805
rect 11238 19796 11244 19848
rect 11296 19836 11302 19848
rect 11405 19839 11463 19845
rect 11405 19836 11417 19839
rect 11296 19808 11417 19836
rect 11296 19796 11302 19808
rect 11405 19805 11417 19808
rect 11451 19805 11463 19839
rect 11405 19799 11463 19805
rect 18233 19839 18291 19845
rect 18233 19805 18245 19839
rect 18279 19836 18291 19839
rect 18322 19836 18328 19848
rect 18279 19808 18328 19836
rect 18279 19805 18291 19808
rect 18233 19799 18291 19805
rect 18322 19796 18328 19808
rect 18380 19796 18386 19848
rect 18690 19836 18696 19848
rect 18651 19808 18696 19836
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 19518 19836 19524 19848
rect 19479 19808 19524 19836
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 19978 19836 19984 19848
rect 19939 19808 19984 19836
rect 19978 19796 19984 19808
rect 20036 19796 20042 19848
rect 20070 19796 20076 19848
rect 20128 19836 20134 19848
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20128 19808 20545 19836
rect 20128 19796 20134 19808
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 21085 19839 21143 19845
rect 21085 19805 21097 19839
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 4798 19728 4804 19780
rect 4856 19768 4862 19780
rect 4902 19771 4960 19777
rect 4902 19768 4914 19771
rect 4856 19740 4914 19768
rect 4856 19728 4862 19740
rect 4902 19737 4914 19740
rect 4948 19737 4960 19771
rect 6365 19771 6423 19777
rect 6365 19768 6377 19771
rect 4902 19731 4960 19737
rect 5000 19740 6377 19768
rect 1486 19700 1492 19712
rect 1447 19672 1492 19700
rect 1486 19660 1492 19672
rect 1544 19660 1550 19712
rect 2038 19700 2044 19712
rect 1999 19672 2044 19700
rect 2038 19660 2044 19672
rect 2096 19660 2102 19712
rect 3053 19703 3111 19709
rect 3053 19669 3065 19703
rect 3099 19700 3111 19703
rect 3142 19700 3148 19712
rect 3099 19672 3148 19700
rect 3099 19669 3111 19672
rect 3053 19663 3111 19669
rect 3142 19660 3148 19672
rect 3200 19660 3206 19712
rect 3326 19660 3332 19712
rect 3384 19700 3390 19712
rect 3789 19703 3847 19709
rect 3789 19700 3801 19703
rect 3384 19672 3801 19700
rect 3384 19660 3390 19672
rect 3789 19669 3801 19672
rect 3835 19669 3847 19703
rect 3789 19663 3847 19669
rect 3878 19660 3884 19712
rect 3936 19700 3942 19712
rect 4062 19700 4068 19712
rect 3936 19672 4068 19700
rect 3936 19660 3942 19672
rect 4062 19660 4068 19672
rect 4120 19700 4126 19712
rect 5000 19700 5028 19740
rect 6365 19737 6377 19740
rect 6411 19737 6423 19771
rect 6365 19731 6423 19737
rect 9208 19771 9266 19777
rect 9208 19737 9220 19771
rect 9254 19768 9266 19771
rect 9398 19768 9404 19780
rect 9254 19740 9404 19768
rect 9254 19737 9266 19740
rect 9208 19731 9266 19737
rect 9398 19728 9404 19740
rect 9456 19728 9462 19780
rect 17589 19771 17647 19777
rect 17589 19737 17601 19771
rect 17635 19768 17647 19771
rect 17635 19740 19334 19768
rect 17635 19737 17647 19740
rect 17589 19731 17647 19737
rect 4120 19672 5028 19700
rect 4120 19660 4126 19672
rect 5718 19660 5724 19712
rect 5776 19700 5782 19712
rect 6089 19703 6147 19709
rect 6089 19700 6101 19703
rect 5776 19672 6101 19700
rect 5776 19660 5782 19672
rect 6089 19669 6101 19672
rect 6135 19669 6147 19703
rect 6089 19663 6147 19669
rect 7742 19660 7748 19712
rect 7800 19700 7806 19712
rect 7929 19703 7987 19709
rect 7929 19700 7941 19703
rect 7800 19672 7941 19700
rect 7800 19660 7806 19672
rect 7929 19669 7941 19672
rect 7975 19669 7987 19703
rect 7929 19663 7987 19669
rect 8021 19703 8079 19709
rect 8021 19669 8033 19703
rect 8067 19700 8079 19703
rect 8386 19700 8392 19712
rect 8067 19672 8392 19700
rect 8067 19669 8079 19672
rect 8021 19663 8079 19669
rect 8386 19660 8392 19672
rect 8444 19660 8450 19712
rect 12529 19703 12587 19709
rect 12529 19669 12541 19703
rect 12575 19700 12587 19703
rect 12618 19700 12624 19712
rect 12575 19672 12624 19700
rect 12575 19669 12587 19672
rect 12529 19663 12587 19669
rect 12618 19660 12624 19672
rect 12676 19660 12682 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18322 19700 18328 19712
rect 18003 19672 18328 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18322 19660 18328 19672
rect 18380 19660 18386 19712
rect 19306 19700 19334 19740
rect 19610 19728 19616 19780
rect 19668 19768 19674 19780
rect 21100 19768 21128 19799
rect 19668 19740 21128 19768
rect 19668 19728 19674 19740
rect 19518 19700 19524 19712
rect 19306 19672 19524 19700
rect 19518 19660 19524 19672
rect 19576 19660 19582 19712
rect 20714 19700 20720 19712
rect 20675 19672 20720 19700
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 21266 19700 21272 19712
rect 21227 19672 21272 19700
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 1946 19456 1952 19508
rect 2004 19496 2010 19508
rect 2041 19499 2099 19505
rect 2041 19496 2053 19499
rect 2004 19468 2053 19496
rect 2004 19456 2010 19468
rect 2041 19465 2053 19468
rect 2087 19465 2099 19499
rect 2498 19496 2504 19508
rect 2459 19468 2504 19496
rect 2041 19459 2099 19465
rect 2498 19456 2504 19468
rect 2556 19456 2562 19508
rect 2961 19499 3019 19505
rect 2961 19496 2973 19499
rect 2746 19468 2973 19496
rect 2746 19428 2774 19468
rect 2961 19465 2973 19468
rect 3007 19465 3019 19499
rect 2961 19459 3019 19465
rect 4522 19456 4528 19508
rect 4580 19496 4586 19508
rect 5353 19499 5411 19505
rect 5353 19496 5365 19499
rect 4580 19468 5365 19496
rect 4580 19456 4586 19468
rect 5353 19465 5365 19468
rect 5399 19465 5411 19499
rect 7742 19496 7748 19508
rect 7703 19468 7748 19496
rect 5353 19459 5411 19465
rect 7742 19456 7748 19468
rect 7800 19456 7806 19508
rect 9398 19496 9404 19508
rect 9359 19468 9404 19496
rect 9398 19456 9404 19468
rect 9456 19456 9462 19508
rect 19337 19499 19395 19505
rect 19337 19465 19349 19499
rect 19383 19496 19395 19499
rect 19978 19496 19984 19508
rect 19383 19468 19984 19496
rect 19383 19465 19395 19468
rect 19337 19459 19395 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 20073 19499 20131 19505
rect 20073 19465 20085 19499
rect 20119 19465 20131 19499
rect 20073 19459 20131 19465
rect 4338 19428 4344 19440
rect 2240 19400 2774 19428
rect 3712 19400 4344 19428
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 2240 19369 2268 19400
rect 2225 19363 2283 19369
rect 2225 19329 2237 19363
rect 2271 19329 2283 19363
rect 2682 19360 2688 19372
rect 2643 19332 2688 19360
rect 2225 19323 2283 19329
rect 2682 19320 2688 19332
rect 2740 19320 2746 19372
rect 3142 19360 3148 19372
rect 3103 19332 3148 19360
rect 3142 19320 3148 19332
rect 3200 19320 3206 19372
rect 3712 19369 3740 19400
rect 4338 19388 4344 19400
rect 4396 19388 4402 19440
rect 8113 19431 8171 19437
rect 8113 19397 8125 19431
rect 8159 19428 8171 19431
rect 9677 19431 9735 19437
rect 9677 19428 9689 19431
rect 8159 19400 9689 19428
rect 8159 19397 8171 19400
rect 8113 19391 8171 19397
rect 9677 19397 9689 19400
rect 9723 19397 9735 19431
rect 9677 19391 9735 19397
rect 12544 19400 14228 19428
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 3953 19363 4011 19369
rect 3953 19360 3965 19363
rect 3697 19323 3755 19329
rect 3804 19332 3965 19360
rect 3326 19252 3332 19304
rect 3384 19292 3390 19304
rect 3804 19292 3832 19332
rect 3953 19329 3965 19332
rect 3999 19329 4011 19363
rect 3953 19323 4011 19329
rect 7834 19320 7840 19372
rect 7892 19360 7898 19372
rect 8205 19363 8263 19369
rect 8205 19360 8217 19363
rect 7892 19332 8217 19360
rect 7892 19320 7898 19332
rect 8205 19329 8217 19332
rect 8251 19329 8263 19363
rect 8205 19323 8263 19329
rect 8662 19320 8668 19372
rect 8720 19360 8726 19372
rect 12544 19369 12572 19400
rect 8757 19363 8815 19369
rect 8757 19360 8769 19363
rect 8720 19332 8769 19360
rect 8720 19320 8726 19332
rect 8757 19329 8769 19332
rect 8803 19329 8815 19363
rect 8757 19323 8815 19329
rect 12529 19363 12587 19369
rect 12529 19329 12541 19363
rect 12575 19329 12587 19363
rect 12529 19323 12587 19329
rect 12618 19320 12624 19372
rect 12676 19360 12682 19372
rect 12785 19363 12843 19369
rect 12785 19360 12797 19363
rect 12676 19332 12797 19360
rect 12676 19320 12682 19332
rect 12785 19329 12797 19332
rect 12831 19360 12843 19363
rect 13630 19360 13636 19372
rect 12831 19332 13636 19360
rect 12831 19329 12843 19332
rect 12785 19323 12843 19329
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 14200 19369 14228 19400
rect 18690 19388 18696 19440
rect 18748 19428 18754 19440
rect 20088 19428 20116 19459
rect 20530 19456 20536 19508
rect 20588 19456 20594 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 21269 19499 21327 19505
rect 21269 19496 21281 19499
rect 20680 19468 21281 19496
rect 20680 19456 20686 19468
rect 21269 19465 21281 19468
rect 21315 19465 21327 19499
rect 21269 19459 21327 19465
rect 18748 19400 20116 19428
rect 20548 19428 20576 19456
rect 20548 19400 20760 19428
rect 18748 19388 18754 19400
rect 14185 19363 14243 19369
rect 14185 19329 14197 19363
rect 14231 19360 14243 19363
rect 14274 19360 14280 19372
rect 14231 19332 14280 19360
rect 14231 19329 14243 19332
rect 14185 19323 14243 19329
rect 14274 19320 14280 19332
rect 14332 19320 14338 19372
rect 14458 19369 14464 19372
rect 14452 19360 14464 19369
rect 14419 19332 14464 19360
rect 14452 19323 14464 19332
rect 14458 19320 14464 19323
rect 14516 19320 14522 19372
rect 17954 19320 17960 19372
rect 18012 19360 18018 19372
rect 18877 19363 18935 19369
rect 18877 19360 18889 19363
rect 18012 19332 18889 19360
rect 18012 19320 18018 19332
rect 18877 19329 18889 19332
rect 18923 19360 18935 19363
rect 19153 19363 19211 19369
rect 19153 19360 19165 19363
rect 18923 19332 19165 19360
rect 18923 19329 18935 19332
rect 18877 19323 18935 19329
rect 19153 19329 19165 19332
rect 19199 19329 19211 19363
rect 19153 19323 19211 19329
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 20070 19360 20076 19372
rect 19613 19323 19671 19329
rect 19812 19332 20076 19360
rect 3384 19264 3832 19292
rect 8389 19295 8447 19301
rect 3384 19252 3390 19264
rect 8389 19261 8401 19295
rect 8435 19292 8447 19295
rect 8680 19292 8708 19320
rect 19628 19292 19656 19323
rect 8435 19264 8708 19292
rect 18432 19264 19656 19292
rect 8435 19261 8447 19264
rect 8389 19255 8447 19261
rect 18432 19233 18460 19264
rect 19812 19233 19840 19332
rect 20070 19320 20076 19332
rect 20128 19320 20134 19372
rect 20254 19360 20260 19372
rect 20215 19332 20260 19360
rect 20254 19320 20260 19332
rect 20312 19320 20318 19372
rect 20530 19360 20536 19372
rect 20491 19332 20536 19360
rect 20530 19320 20536 19332
rect 20588 19320 20594 19372
rect 20732 19233 20760 19400
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20824 19332 21097 19360
rect 18417 19227 18475 19233
rect 18417 19224 18429 19227
rect 15120 19196 18429 19224
rect 15120 19168 15148 19196
rect 18417 19193 18429 19196
rect 18463 19193 18475 19227
rect 18417 19187 18475 19193
rect 19797 19227 19855 19233
rect 19797 19193 19809 19227
rect 19843 19193 19855 19227
rect 19797 19187 19855 19193
rect 20717 19227 20775 19233
rect 20717 19193 20729 19227
rect 20763 19193 20775 19227
rect 20717 19187 20775 19193
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 4890 19116 4896 19168
rect 4948 19156 4954 19168
rect 5077 19159 5135 19165
rect 5077 19156 5089 19159
rect 4948 19128 5089 19156
rect 4948 19116 4954 19128
rect 5077 19125 5089 19128
rect 5123 19156 5135 19159
rect 5258 19156 5264 19168
rect 5123 19128 5264 19156
rect 5123 19125 5135 19128
rect 5077 19119 5135 19125
rect 5258 19116 5264 19128
rect 5316 19116 5322 19168
rect 5810 19156 5816 19168
rect 5723 19128 5816 19156
rect 5810 19116 5816 19128
rect 5868 19156 5874 19168
rect 12894 19156 12900 19168
rect 5868 19128 12900 19156
rect 5868 19116 5874 19128
rect 12894 19116 12900 19128
rect 12952 19116 12958 19168
rect 13909 19159 13967 19165
rect 13909 19125 13921 19159
rect 13955 19156 13967 19159
rect 14366 19156 14372 19168
rect 13955 19128 14372 19156
rect 13955 19125 13967 19128
rect 13909 19119 13967 19125
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 15102 19116 15108 19168
rect 15160 19116 15166 19168
rect 15562 19156 15568 19168
rect 15523 19128 15568 19156
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 20346 19116 20352 19168
rect 20404 19156 20410 19168
rect 20824 19156 20852 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 20404 19128 20852 19156
rect 20404 19116 20410 19128
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1670 18912 1676 18964
rect 1728 18952 1734 18964
rect 1949 18955 2007 18961
rect 1949 18952 1961 18955
rect 1728 18924 1961 18952
rect 1728 18912 1734 18924
rect 1949 18921 1961 18924
rect 1995 18921 2007 18955
rect 1949 18915 2007 18921
rect 2130 18912 2136 18964
rect 2188 18952 2194 18964
rect 2409 18955 2467 18961
rect 2409 18952 2421 18955
rect 2188 18924 2421 18952
rect 2188 18912 2194 18924
rect 2409 18921 2421 18924
rect 2455 18921 2467 18955
rect 2409 18915 2467 18921
rect 2774 18912 2780 18964
rect 2832 18952 2838 18964
rect 2869 18955 2927 18961
rect 2869 18952 2881 18955
rect 2832 18924 2881 18952
rect 2832 18912 2838 18924
rect 2869 18921 2881 18924
rect 2915 18921 2927 18955
rect 2869 18915 2927 18921
rect 8386 18912 8392 18964
rect 8444 18952 8450 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8444 18924 8953 18952
rect 8444 18912 8450 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 8941 18915 8999 18921
rect 13446 18912 13452 18964
rect 13504 18952 13510 18964
rect 17957 18955 18015 18961
rect 17957 18952 17969 18955
rect 13504 18924 17969 18952
rect 13504 18912 13510 18924
rect 17957 18921 17969 18924
rect 18003 18921 18015 18955
rect 17957 18915 18015 18921
rect 19429 18955 19487 18961
rect 19429 18921 19441 18955
rect 19475 18952 19487 18955
rect 19610 18952 19616 18964
rect 19475 18924 19616 18952
rect 19475 18921 19487 18924
rect 19429 18915 19487 18921
rect 4614 18884 4620 18896
rect 3712 18856 4620 18884
rect 3712 18816 3740 18856
rect 4614 18844 4620 18856
rect 4672 18844 4678 18896
rect 8573 18887 8631 18893
rect 8573 18853 8585 18887
rect 8619 18853 8631 18887
rect 17972 18884 18000 18915
rect 19610 18912 19616 18924
rect 19668 18912 19674 18964
rect 19889 18955 19947 18961
rect 19889 18921 19901 18955
rect 19935 18952 19947 18955
rect 20530 18952 20536 18964
rect 19935 18924 20536 18952
rect 19935 18921 19947 18924
rect 19889 18915 19947 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 20349 18887 20407 18893
rect 17972 18856 20208 18884
rect 8573 18847 8631 18853
rect 2608 18788 3740 18816
rect 3881 18819 3939 18825
rect 1670 18748 1676 18760
rect 1631 18720 1676 18748
rect 1670 18708 1676 18720
rect 1728 18708 1734 18760
rect 2130 18748 2136 18760
rect 2091 18720 2136 18748
rect 2130 18708 2136 18720
rect 2188 18708 2194 18760
rect 2608 18757 2636 18788
rect 3881 18785 3893 18819
rect 3927 18816 3939 18819
rect 8588 18816 8616 18847
rect 8662 18816 8668 18828
rect 3927 18788 5304 18816
rect 8575 18788 8668 18816
rect 3927 18785 3939 18788
rect 3881 18779 3939 18785
rect 2593 18751 2651 18757
rect 2593 18717 2605 18751
rect 2639 18717 2651 18751
rect 2593 18711 2651 18717
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3896 18748 3924 18779
rect 5276 18760 5304 18788
rect 8662 18776 8668 18788
rect 8720 18816 8726 18828
rect 9493 18819 9551 18825
rect 9493 18816 9505 18819
rect 8720 18788 9505 18816
rect 8720 18776 8726 18788
rect 9493 18785 9505 18788
rect 9539 18785 9551 18819
rect 17589 18819 17647 18825
rect 17589 18816 17601 18819
rect 9493 18779 9551 18785
rect 15856 18788 17601 18816
rect 3099 18720 3924 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 4338 18708 4344 18760
rect 4396 18748 4402 18760
rect 5169 18751 5227 18757
rect 5169 18748 5181 18751
rect 4396 18720 5181 18748
rect 4396 18708 4402 18720
rect 5169 18717 5181 18720
rect 5215 18717 5227 18751
rect 5169 18711 5227 18717
rect 5258 18708 5264 18760
rect 5316 18708 5322 18760
rect 5436 18751 5494 18757
rect 5436 18717 5448 18751
rect 5482 18748 5494 18751
rect 5718 18748 5724 18760
rect 5482 18720 5724 18748
rect 5482 18717 5494 18720
rect 5436 18711 5494 18717
rect 5718 18708 5724 18720
rect 5776 18708 5782 18760
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 14274 18708 14280 18760
rect 14332 18748 14338 18760
rect 14553 18751 14611 18757
rect 14553 18748 14565 18751
rect 14332 18720 14565 18748
rect 14332 18708 14338 18720
rect 14553 18717 14565 18720
rect 14599 18717 14611 18751
rect 14553 18711 14611 18717
rect 14820 18751 14878 18757
rect 14820 18717 14832 18751
rect 14866 18748 14878 18751
rect 15562 18748 15568 18760
rect 14866 18720 15568 18748
rect 14866 18717 14878 18720
rect 14820 18711 14878 18717
rect 15562 18708 15568 18720
rect 15620 18708 15626 18760
rect 1302 18640 1308 18692
rect 1360 18680 1366 18692
rect 1360 18652 1624 18680
rect 1360 18640 1366 18652
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 1596 18612 1624 18652
rect 2682 18640 2688 18692
rect 2740 18680 2746 18692
rect 3421 18683 3479 18689
rect 3421 18680 3433 18683
rect 2740 18652 3433 18680
rect 2740 18640 2746 18652
rect 3421 18649 3433 18652
rect 3467 18680 3479 18683
rect 6638 18680 6644 18692
rect 3467 18652 6644 18680
rect 3467 18649 3479 18652
rect 3421 18643 3479 18649
rect 6638 18640 6644 18652
rect 6696 18640 6702 18692
rect 7460 18683 7518 18689
rect 7460 18649 7472 18683
rect 7506 18680 7518 18683
rect 8662 18680 8668 18692
rect 7506 18652 8668 18680
rect 7506 18649 7518 18652
rect 7460 18643 7518 18649
rect 8662 18640 8668 18652
rect 8720 18640 8726 18692
rect 11238 18640 11244 18692
rect 11296 18680 11302 18692
rect 15856 18680 15884 18788
rect 17589 18785 17601 18788
rect 17635 18816 17647 18819
rect 17635 18788 20116 18816
rect 17635 18785 17647 18788
rect 17589 18779 17647 18785
rect 16209 18751 16267 18757
rect 16209 18748 16221 18751
rect 11296 18652 15884 18680
rect 15948 18720 16221 18748
rect 11296 18640 11302 18652
rect 3234 18612 3240 18624
rect 1596 18584 3240 18612
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 3878 18572 3884 18624
rect 3936 18612 3942 18624
rect 4157 18615 4215 18621
rect 4157 18612 4169 18615
rect 3936 18584 4169 18612
rect 3936 18572 3942 18584
rect 4157 18581 4169 18584
rect 4203 18581 4215 18615
rect 4614 18612 4620 18624
rect 4527 18584 4620 18612
rect 4157 18575 4215 18581
rect 4614 18572 4620 18584
rect 4672 18612 4678 18624
rect 5442 18612 5448 18624
rect 4672 18584 5448 18612
rect 4672 18572 4678 18584
rect 5442 18572 5448 18584
rect 5500 18572 5506 18624
rect 6549 18615 6607 18621
rect 6549 18581 6561 18615
rect 6595 18612 6607 18615
rect 7006 18612 7012 18624
rect 6595 18584 7012 18612
rect 6595 18581 6607 18584
rect 6549 18575 6607 18581
rect 7006 18572 7012 18584
rect 7064 18572 7070 18624
rect 9306 18612 9312 18624
rect 9267 18584 9312 18612
rect 9306 18572 9312 18584
rect 9364 18572 9370 18624
rect 9398 18572 9404 18624
rect 9456 18612 9462 18624
rect 9456 18584 9501 18612
rect 9456 18572 9462 18584
rect 14918 18572 14924 18624
rect 14976 18612 14982 18624
rect 15948 18621 15976 18720
rect 16209 18717 16221 18720
rect 16255 18717 16267 18751
rect 16209 18711 16267 18717
rect 19245 18751 19303 18757
rect 19245 18717 19257 18751
rect 19291 18748 19303 18751
rect 19518 18748 19524 18760
rect 19291 18720 19524 18748
rect 19291 18717 19303 18720
rect 19245 18711 19303 18717
rect 19518 18708 19524 18720
rect 19576 18708 19582 18760
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 19720 18680 19748 18711
rect 18984 18652 19748 18680
rect 20088 18680 20116 18788
rect 20180 18757 20208 18856
rect 20349 18853 20361 18887
rect 20395 18884 20407 18887
rect 20438 18884 20444 18896
rect 20395 18856 20444 18884
rect 20395 18853 20407 18856
rect 20349 18847 20407 18853
rect 20438 18844 20444 18856
rect 20496 18844 20502 18896
rect 20809 18887 20867 18893
rect 20809 18853 20821 18887
rect 20855 18853 20867 18887
rect 20809 18847 20867 18853
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 20625 18751 20683 18757
rect 20625 18717 20637 18751
rect 20671 18717 20683 18751
rect 20824 18748 20852 18847
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 20824 18720 21097 18748
rect 20625 18711 20683 18717
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 20640 18680 20668 18711
rect 20088 18652 20668 18680
rect 18984 18624 19012 18652
rect 15933 18615 15991 18621
rect 15933 18612 15945 18615
rect 14976 18584 15945 18612
rect 14976 18572 14982 18584
rect 15933 18581 15945 18584
rect 15979 18581 15991 18615
rect 15933 18575 15991 18581
rect 16853 18615 16911 18621
rect 16853 18581 16865 18615
rect 16899 18612 16911 18615
rect 17034 18612 17040 18624
rect 16899 18584 17040 18612
rect 16899 18581 16911 18584
rect 16853 18575 16911 18581
rect 17034 18572 17040 18584
rect 17092 18572 17098 18624
rect 17862 18572 17868 18624
rect 17920 18612 17926 18624
rect 18325 18615 18383 18621
rect 18325 18612 18337 18615
rect 17920 18584 18337 18612
rect 17920 18572 17926 18584
rect 18325 18581 18337 18584
rect 18371 18581 18383 18615
rect 18325 18575 18383 18581
rect 18877 18615 18935 18621
rect 18877 18581 18889 18615
rect 18923 18612 18935 18615
rect 18966 18612 18972 18624
rect 18923 18584 18972 18612
rect 18923 18581 18935 18584
rect 18877 18575 18935 18581
rect 18966 18572 18972 18584
rect 19024 18572 19030 18624
rect 21266 18612 21272 18624
rect 21227 18584 21272 18612
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 1670 18368 1676 18420
rect 1728 18408 1734 18420
rect 2409 18411 2467 18417
rect 2409 18408 2421 18411
rect 1728 18380 2421 18408
rect 1728 18368 1734 18380
rect 2409 18377 2421 18380
rect 2455 18377 2467 18411
rect 3878 18408 3884 18420
rect 2409 18371 2467 18377
rect 2746 18380 3884 18408
rect 2746 18340 2774 18380
rect 3878 18368 3884 18380
rect 3936 18368 3942 18420
rect 3973 18411 4031 18417
rect 3973 18377 3985 18411
rect 4019 18408 4031 18411
rect 4617 18411 4675 18417
rect 4617 18408 4629 18411
rect 4019 18380 4629 18408
rect 4019 18377 4031 18380
rect 3973 18371 4031 18377
rect 4617 18377 4629 18380
rect 4663 18377 4675 18411
rect 9398 18408 9404 18420
rect 9359 18380 9404 18408
rect 4617 18371 4675 18377
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 9769 18411 9827 18417
rect 9769 18377 9781 18411
rect 9815 18408 9827 18411
rect 13170 18408 13176 18420
rect 9815 18380 13176 18408
rect 9815 18377 9827 18380
rect 9769 18371 9827 18377
rect 2148 18312 2774 18340
rect 2148 18281 2176 18312
rect 3234 18300 3240 18352
rect 3292 18340 3298 18352
rect 6365 18343 6423 18349
rect 6365 18340 6377 18343
rect 3292 18312 6377 18340
rect 3292 18300 3298 18312
rect 6365 18309 6377 18312
rect 6411 18309 6423 18343
rect 6365 18303 6423 18309
rect 6638 18300 6644 18352
rect 6696 18340 6702 18352
rect 8941 18343 8999 18349
rect 8941 18340 8953 18343
rect 6696 18312 8953 18340
rect 6696 18300 6702 18312
rect 8941 18309 8953 18312
rect 8987 18340 8999 18343
rect 9784 18340 9812 18371
rect 13170 18368 13176 18380
rect 13228 18368 13234 18420
rect 13354 18368 13360 18420
rect 13412 18408 13418 18420
rect 19429 18411 19487 18417
rect 19429 18408 19441 18411
rect 13412 18380 19441 18408
rect 13412 18368 13418 18380
rect 19429 18377 19441 18380
rect 19475 18377 19487 18411
rect 20346 18408 20352 18420
rect 20307 18380 20352 18408
rect 19429 18371 19487 18377
rect 8987 18312 9812 18340
rect 14093 18343 14151 18349
rect 8987 18309 8999 18312
rect 8941 18303 8999 18309
rect 14093 18309 14105 18343
rect 14139 18340 14151 18343
rect 15749 18343 15807 18349
rect 15749 18340 15761 18343
rect 14139 18312 15761 18340
rect 14139 18309 14151 18312
rect 14093 18303 14151 18309
rect 15749 18309 15761 18312
rect 15795 18309 15807 18343
rect 15749 18303 15807 18309
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18272 1731 18275
rect 2133 18275 2191 18281
rect 1719 18244 1992 18272
rect 1719 18241 1731 18244
rect 1673 18235 1731 18241
rect 1964 18145 1992 18244
rect 2133 18241 2145 18275
rect 2179 18241 2191 18275
rect 2133 18235 2191 18241
rect 2593 18275 2651 18281
rect 2593 18241 2605 18275
rect 2639 18272 2651 18275
rect 2682 18272 2688 18284
rect 2639 18244 2688 18272
rect 2639 18241 2651 18244
rect 2593 18235 2651 18241
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 3418 18232 3424 18284
rect 3476 18272 3482 18284
rect 3605 18275 3663 18281
rect 3605 18272 3617 18275
rect 3476 18244 3617 18272
rect 3476 18232 3482 18244
rect 3605 18241 3617 18244
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 3970 18232 3976 18284
rect 4028 18272 4034 18284
rect 9033 18275 9091 18281
rect 4028 18244 8064 18272
rect 4028 18232 4034 18244
rect 3326 18204 3332 18216
rect 3287 18176 3332 18204
rect 3326 18164 3332 18176
rect 3384 18164 3390 18216
rect 3513 18207 3571 18213
rect 3513 18173 3525 18207
rect 3559 18204 3571 18207
rect 3878 18204 3884 18216
rect 3559 18176 3884 18204
rect 3559 18173 3571 18176
rect 3513 18167 3571 18173
rect 3878 18164 3884 18176
rect 3936 18164 3942 18216
rect 4706 18204 4712 18216
rect 4667 18176 4712 18204
rect 4706 18164 4712 18176
rect 4764 18164 4770 18216
rect 4890 18204 4896 18216
rect 4851 18176 4896 18204
rect 4890 18164 4896 18176
rect 4948 18164 4954 18216
rect 1949 18139 2007 18145
rect 1949 18105 1961 18139
rect 1995 18105 2007 18139
rect 1949 18099 2007 18105
rect 2314 18096 2320 18148
rect 2372 18136 2378 18148
rect 5629 18139 5687 18145
rect 5629 18136 5641 18139
rect 2372 18108 5641 18136
rect 2372 18096 2378 18108
rect 5629 18105 5641 18108
rect 5675 18105 5687 18139
rect 5629 18099 5687 18105
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 2774 18028 2780 18080
rect 2832 18068 2838 18080
rect 2869 18071 2927 18077
rect 2869 18068 2881 18071
rect 2832 18040 2881 18068
rect 2832 18028 2838 18040
rect 2869 18037 2881 18040
rect 2915 18037 2927 18071
rect 4246 18068 4252 18080
rect 4207 18040 4252 18068
rect 2869 18031 2927 18037
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 5258 18068 5264 18080
rect 5219 18040 5264 18068
rect 5258 18028 5264 18040
rect 5316 18028 5322 18080
rect 8036 18068 8064 18244
rect 9033 18241 9045 18275
rect 9079 18241 9091 18275
rect 11974 18272 11980 18284
rect 11935 18244 11980 18272
rect 9033 18235 9091 18241
rect 8662 18164 8668 18216
rect 8720 18204 8726 18216
rect 8757 18207 8815 18213
rect 8757 18204 8769 18207
rect 8720 18176 8769 18204
rect 8720 18164 8726 18176
rect 8757 18173 8769 18176
rect 8803 18173 8815 18207
rect 8757 18167 8815 18173
rect 8389 18139 8447 18145
rect 8389 18105 8401 18139
rect 8435 18136 8447 18139
rect 9048 18136 9076 18235
rect 11974 18232 11980 18244
rect 12032 18232 12038 18284
rect 13446 18232 13452 18284
rect 13504 18272 13510 18284
rect 14001 18275 14059 18281
rect 14001 18272 14013 18275
rect 13504 18244 14013 18272
rect 13504 18232 13510 18244
rect 14001 18241 14013 18244
rect 14047 18241 14059 18275
rect 15102 18272 15108 18284
rect 15063 18244 15108 18272
rect 14001 18235 14059 18241
rect 15102 18232 15108 18244
rect 15160 18232 15166 18284
rect 17126 18232 17132 18284
rect 17184 18272 17190 18284
rect 17862 18272 17868 18284
rect 17184 18244 17868 18272
rect 17184 18232 17190 18244
rect 17862 18232 17868 18244
rect 17920 18232 17926 18284
rect 19153 18275 19211 18281
rect 19153 18272 19165 18275
rect 18156 18244 19165 18272
rect 18156 18216 18184 18244
rect 19153 18241 19165 18244
rect 19199 18241 19211 18275
rect 19444 18272 19472 18371
rect 20346 18368 20352 18380
rect 20404 18368 20410 18420
rect 20165 18275 20223 18281
rect 20165 18272 20177 18275
rect 19444 18244 20177 18272
rect 19153 18235 19211 18241
rect 20165 18241 20177 18244
rect 20211 18241 20223 18275
rect 20622 18272 20628 18284
rect 20583 18244 20628 18272
rect 20165 18235 20223 18241
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 12894 18204 12900 18216
rect 12855 18176 12900 18204
rect 12894 18164 12900 18176
rect 12952 18164 12958 18216
rect 13909 18207 13967 18213
rect 13909 18173 13921 18207
rect 13955 18204 13967 18207
rect 14366 18204 14372 18216
rect 13955 18176 14372 18204
rect 13955 18173 13967 18176
rect 13909 18167 13967 18173
rect 14366 18164 14372 18176
rect 14424 18164 14430 18216
rect 14826 18204 14832 18216
rect 14787 18176 14832 18204
rect 14826 18164 14832 18176
rect 14884 18164 14890 18216
rect 14918 18164 14924 18216
rect 14976 18204 14982 18216
rect 15013 18207 15071 18213
rect 15013 18204 15025 18207
rect 14976 18176 15025 18204
rect 14976 18164 14982 18176
rect 15013 18173 15025 18176
rect 15059 18173 15071 18207
rect 15013 18167 15071 18173
rect 17678 18164 17684 18216
rect 17736 18204 17742 18216
rect 17957 18207 18015 18213
rect 17957 18204 17969 18207
rect 17736 18176 17969 18204
rect 17736 18164 17742 18176
rect 17957 18173 17969 18176
rect 18003 18204 18015 18207
rect 18046 18204 18052 18216
rect 18003 18176 18052 18204
rect 18003 18173 18015 18176
rect 17957 18167 18015 18173
rect 18046 18164 18052 18176
rect 18104 18164 18110 18216
rect 18138 18164 18144 18216
rect 18196 18204 18202 18216
rect 18196 18176 18289 18204
rect 18196 18164 18202 18176
rect 20346 18164 20352 18216
rect 20404 18204 20410 18216
rect 21100 18204 21128 18235
rect 20404 18176 21128 18204
rect 20404 18164 20410 18176
rect 13262 18136 13268 18148
rect 8435 18108 13268 18136
rect 8435 18105 8447 18108
rect 8389 18099 8447 18105
rect 13262 18096 13268 18108
rect 13320 18096 13326 18148
rect 10042 18068 10048 18080
rect 8036 18040 10048 18068
rect 10042 18028 10048 18040
rect 10100 18028 10106 18080
rect 12066 18028 12072 18080
rect 12124 18068 12130 18080
rect 12621 18071 12679 18077
rect 12621 18068 12633 18071
rect 12124 18040 12633 18068
rect 12124 18028 12130 18040
rect 12621 18037 12633 18040
rect 12667 18037 12679 18071
rect 13446 18068 13452 18080
rect 13407 18040 13452 18068
rect 12621 18031 12679 18037
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 14461 18071 14519 18077
rect 14461 18037 14473 18071
rect 14507 18068 14519 18071
rect 15378 18068 15384 18080
rect 14507 18040 15384 18068
rect 14507 18037 14519 18040
rect 14461 18031 14519 18037
rect 15378 18028 15384 18040
rect 15436 18028 15442 18080
rect 15473 18071 15531 18077
rect 15473 18037 15485 18071
rect 15519 18068 15531 18071
rect 17402 18068 17408 18080
rect 15519 18040 17408 18068
rect 15519 18037 15531 18040
rect 15473 18031 15531 18037
rect 17402 18028 17408 18040
rect 17460 18028 17466 18080
rect 17497 18071 17555 18077
rect 17497 18037 17509 18071
rect 17543 18068 17555 18071
rect 17862 18068 17868 18080
rect 17543 18040 17868 18068
rect 17543 18037 17555 18040
rect 17497 18031 17555 18037
rect 17862 18028 17868 18040
rect 17920 18028 17926 18080
rect 18506 18068 18512 18080
rect 18467 18040 18512 18068
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 19702 18028 19708 18080
rect 19760 18068 19766 18080
rect 19797 18071 19855 18077
rect 19797 18068 19809 18071
rect 19760 18040 19809 18068
rect 19760 18028 19766 18040
rect 19797 18037 19809 18040
rect 19843 18037 19855 18071
rect 19797 18031 19855 18037
rect 20809 18071 20867 18077
rect 20809 18037 20821 18071
rect 20855 18068 20867 18071
rect 20990 18068 20996 18080
rect 20855 18040 20996 18068
rect 20855 18037 20867 18040
rect 20809 18031 20867 18037
rect 20990 18028 20996 18040
rect 21048 18028 21054 18080
rect 21269 18071 21327 18077
rect 21269 18037 21281 18071
rect 21315 18068 21327 18071
rect 21358 18068 21364 18080
rect 21315 18040 21364 18068
rect 21315 18037 21327 18040
rect 21269 18031 21327 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 4433 17867 4491 17873
rect 4433 17833 4445 17867
rect 4479 17864 4491 17867
rect 4706 17864 4712 17876
rect 4479 17836 4712 17864
rect 4479 17833 4491 17836
rect 4433 17827 4491 17833
rect 4706 17824 4712 17836
rect 4764 17824 4770 17876
rect 7742 17824 7748 17876
rect 7800 17864 7806 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7800 17836 7849 17864
rect 7800 17824 7806 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 9582 17824 9588 17876
rect 9640 17864 9646 17876
rect 13633 17867 13691 17873
rect 13633 17864 13645 17867
rect 9640 17836 13645 17864
rect 9640 17824 9646 17836
rect 13633 17833 13645 17836
rect 13679 17864 13691 17867
rect 14550 17864 14556 17876
rect 13679 17836 14556 17864
rect 13679 17833 13691 17836
rect 13633 17827 13691 17833
rect 14550 17824 14556 17836
rect 14608 17824 14614 17876
rect 15102 17864 15108 17876
rect 15063 17836 15108 17864
rect 15102 17824 15108 17836
rect 15160 17824 15166 17876
rect 19337 17867 19395 17873
rect 19337 17864 19349 17867
rect 15212 17836 19349 17864
rect 1949 17799 2007 17805
rect 1949 17765 1961 17799
rect 1995 17765 2007 17799
rect 1949 17759 2007 17765
rect 1673 17663 1731 17669
rect 1673 17629 1685 17663
rect 1719 17660 1731 17663
rect 1964 17660 1992 17759
rect 3234 17756 3240 17808
rect 3292 17796 3298 17808
rect 3421 17799 3479 17805
rect 3421 17796 3433 17799
rect 3292 17768 3433 17796
rect 3292 17756 3298 17768
rect 3421 17765 3433 17768
rect 3467 17796 3479 17799
rect 5994 17796 6000 17808
rect 3467 17768 6000 17796
rect 3467 17765 3479 17768
rect 3421 17759 3479 17765
rect 5994 17756 6000 17768
rect 6052 17756 6058 17808
rect 10321 17799 10379 17805
rect 10321 17765 10333 17799
rect 10367 17765 10379 17799
rect 10321 17759 10379 17765
rect 2774 17728 2780 17740
rect 2148 17700 2780 17728
rect 2148 17669 2176 17700
rect 2774 17688 2780 17700
rect 2832 17688 2838 17740
rect 3326 17688 3332 17740
rect 3384 17728 3390 17740
rect 4985 17731 5043 17737
rect 4985 17728 4997 17731
rect 3384 17700 4997 17728
rect 3384 17688 3390 17700
rect 4985 17697 4997 17700
rect 5031 17697 5043 17731
rect 10336 17728 10364 17759
rect 13814 17756 13820 17808
rect 13872 17796 13878 17808
rect 15212 17796 15240 17836
rect 19337 17833 19349 17836
rect 19383 17833 19395 17867
rect 19337 17827 19395 17833
rect 13872 17768 15240 17796
rect 15488 17768 15792 17796
rect 13872 17756 13878 17768
rect 10410 17728 10416 17740
rect 10323 17700 10416 17728
rect 4985 17691 5043 17697
rect 10410 17688 10416 17700
rect 10468 17728 10474 17740
rect 12805 17731 12863 17737
rect 12805 17728 12817 17731
rect 10468 17700 10732 17728
rect 10468 17688 10474 17700
rect 1719 17632 1992 17660
rect 2133 17663 2191 17669
rect 1719 17629 1731 17632
rect 1673 17623 1731 17629
rect 2133 17629 2145 17663
rect 2179 17629 2191 17663
rect 2133 17623 2191 17629
rect 2593 17663 2651 17669
rect 2593 17629 2605 17663
rect 2639 17660 2651 17663
rect 3053 17663 3111 17669
rect 2639 17632 2774 17660
rect 2639 17629 2651 17632
rect 2593 17623 2651 17629
rect 1486 17524 1492 17536
rect 1447 17496 1492 17524
rect 1486 17484 1492 17496
rect 1544 17484 1550 17536
rect 2038 17484 2044 17536
rect 2096 17524 2102 17536
rect 2409 17527 2467 17533
rect 2409 17524 2421 17527
rect 2096 17496 2421 17524
rect 2096 17484 2102 17496
rect 2409 17493 2421 17496
rect 2455 17493 2467 17527
rect 2746 17524 2774 17632
rect 3053 17629 3065 17663
rect 3099 17660 3111 17663
rect 4246 17660 4252 17672
rect 3099 17632 4252 17660
rect 3099 17629 3111 17632
rect 3053 17623 3111 17629
rect 4246 17620 4252 17632
rect 4304 17620 4310 17672
rect 7190 17660 7196 17672
rect 7151 17632 7196 17660
rect 7190 17620 7196 17632
rect 7248 17620 7254 17672
rect 8021 17663 8079 17669
rect 8021 17629 8033 17663
rect 8067 17660 8079 17663
rect 8386 17660 8392 17672
rect 8067 17632 8392 17660
rect 8067 17629 8079 17632
rect 8021 17623 8079 17629
rect 8386 17620 8392 17632
rect 8444 17620 8450 17672
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17660 8999 17663
rect 9490 17660 9496 17672
rect 8987 17632 9496 17660
rect 8987 17629 8999 17632
rect 8941 17623 8999 17629
rect 9490 17620 9496 17632
rect 9548 17660 9554 17672
rect 10597 17663 10655 17669
rect 10597 17660 10609 17663
rect 9548 17632 10609 17660
rect 9548 17620 9554 17632
rect 10597 17629 10609 17632
rect 10643 17629 10655 17663
rect 10704 17660 10732 17700
rect 12406 17700 12817 17728
rect 10864 17663 10922 17669
rect 10864 17660 10876 17663
rect 10704 17632 10876 17660
rect 10597 17623 10655 17629
rect 10864 17629 10876 17632
rect 10910 17660 10922 17663
rect 12406 17660 12434 17700
rect 12805 17697 12817 17700
rect 12851 17697 12863 17731
rect 12805 17691 12863 17697
rect 14277 17731 14335 17737
rect 14277 17697 14289 17731
rect 14323 17728 14335 17731
rect 14366 17728 14372 17740
rect 14323 17700 14372 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 14366 17688 14372 17700
rect 14424 17688 14430 17740
rect 15488 17728 15516 17768
rect 15304 17700 15516 17728
rect 10910 17632 12434 17660
rect 14384 17656 14412 17688
rect 15304 17660 15332 17700
rect 15562 17688 15568 17740
rect 15620 17728 15626 17740
rect 15657 17731 15715 17737
rect 15657 17728 15669 17731
rect 15620 17700 15669 17728
rect 15620 17688 15626 17700
rect 15657 17697 15669 17700
rect 15703 17697 15715 17731
rect 15764 17728 15792 17768
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 15764 17700 16681 17728
rect 15657 17691 15715 17697
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 14568 17656 15332 17660
rect 14384 17632 15332 17656
rect 10910 17629 10922 17632
rect 10864 17623 10922 17629
rect 14384 17628 14596 17632
rect 15378 17620 15384 17672
rect 15436 17660 15442 17672
rect 15473 17663 15531 17669
rect 15473 17660 15485 17663
rect 15436 17632 15485 17660
rect 15436 17620 15442 17632
rect 15473 17629 15485 17632
rect 15519 17629 15531 17663
rect 18874 17660 18880 17672
rect 18835 17632 18880 17660
rect 15473 17623 15531 17629
rect 18874 17620 18880 17632
rect 18932 17620 18938 17672
rect 3142 17552 3148 17604
rect 3200 17592 3206 17604
rect 3789 17595 3847 17601
rect 3789 17592 3801 17595
rect 3200 17564 3801 17592
rect 3200 17552 3206 17564
rect 3789 17561 3801 17564
rect 3835 17561 3847 17595
rect 3789 17555 3847 17561
rect 4801 17595 4859 17601
rect 4801 17561 4813 17595
rect 4847 17592 4859 17595
rect 6730 17592 6736 17604
rect 4847 17564 6736 17592
rect 4847 17561 4859 17564
rect 4801 17555 4859 17561
rect 6730 17552 6736 17564
rect 6788 17552 6794 17604
rect 6914 17592 6920 17604
rect 6972 17601 6978 17604
rect 6884 17564 6920 17592
rect 6914 17552 6920 17564
rect 6972 17555 6984 17601
rect 6972 17552 6978 17555
rect 8110 17552 8116 17604
rect 8168 17592 8174 17604
rect 9208 17595 9266 17601
rect 9208 17592 9220 17595
rect 8168 17564 9220 17592
rect 8168 17552 8174 17564
rect 9208 17561 9220 17564
rect 9254 17592 9266 17595
rect 12158 17592 12164 17604
rect 9254 17564 12164 17592
rect 9254 17561 9266 17564
rect 9208 17555 9266 17561
rect 12158 17552 12164 17564
rect 12216 17552 12222 17604
rect 12713 17595 12771 17601
rect 12713 17561 12725 17595
rect 12759 17592 12771 17595
rect 16206 17592 16212 17604
rect 12759 17564 16212 17592
rect 12759 17561 12771 17564
rect 12713 17555 12771 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 16298 17552 16304 17604
rect 16356 17592 16362 17604
rect 16577 17595 16635 17601
rect 16577 17592 16589 17595
rect 16356 17564 16589 17592
rect 16356 17552 16362 17564
rect 16577 17561 16589 17564
rect 16623 17561 16635 17595
rect 16577 17555 16635 17561
rect 18506 17552 18512 17604
rect 18564 17592 18570 17604
rect 18610 17595 18668 17601
rect 18610 17592 18622 17595
rect 18564 17564 18622 17592
rect 18564 17552 18570 17564
rect 18610 17561 18622 17564
rect 18656 17561 18668 17595
rect 19352 17592 19380 17827
rect 19518 17824 19524 17876
rect 19576 17864 19582 17876
rect 19705 17867 19763 17873
rect 19705 17864 19717 17867
rect 19576 17836 19717 17864
rect 19576 17824 19582 17836
rect 19705 17833 19717 17836
rect 19751 17833 19763 17867
rect 20346 17864 20352 17876
rect 20307 17836 20352 17864
rect 19705 17827 19763 17833
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 19702 17688 19708 17740
rect 19760 17728 19766 17740
rect 19760 17700 20668 17728
rect 19760 17688 19766 17700
rect 19886 17660 19892 17672
rect 19847 17632 19892 17660
rect 19886 17620 19892 17632
rect 19944 17620 19950 17672
rect 20640 17669 20668 17700
rect 20165 17663 20223 17669
rect 20165 17629 20177 17663
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20625 17663 20683 17669
rect 20625 17629 20637 17663
rect 20671 17629 20683 17663
rect 20625 17623 20683 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 20180 17592 20208 17623
rect 19352 17564 20208 17592
rect 18610 17555 18668 17561
rect 20346 17552 20352 17604
rect 20404 17592 20410 17604
rect 21100 17592 21128 17623
rect 20404 17564 21128 17592
rect 20404 17552 20410 17564
rect 2869 17527 2927 17533
rect 2869 17524 2881 17527
rect 2746 17496 2881 17524
rect 2409 17487 2467 17493
rect 2869 17493 2881 17496
rect 2915 17493 2927 17527
rect 2869 17487 2927 17493
rect 4893 17527 4951 17533
rect 4893 17493 4905 17527
rect 4939 17524 4951 17527
rect 4982 17524 4988 17536
rect 4939 17496 4988 17524
rect 4939 17493 4951 17496
rect 4893 17487 4951 17493
rect 4982 17484 4988 17496
rect 5040 17484 5046 17536
rect 5534 17524 5540 17536
rect 5495 17496 5540 17524
rect 5534 17484 5540 17496
rect 5592 17484 5598 17536
rect 5813 17527 5871 17533
rect 5813 17493 5825 17527
rect 5859 17524 5871 17527
rect 5902 17524 5908 17536
rect 5859 17496 5908 17524
rect 5859 17493 5871 17496
rect 5813 17487 5871 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 7466 17524 7472 17536
rect 7427 17496 7472 17524
rect 7466 17484 7472 17496
rect 7524 17484 7530 17536
rect 11974 17524 11980 17536
rect 11935 17496 11980 17524
rect 11974 17484 11980 17496
rect 12032 17484 12038 17536
rect 12250 17524 12256 17536
rect 12211 17496 12256 17524
rect 12250 17484 12256 17496
rect 12308 17484 12314 17536
rect 12618 17524 12624 17536
rect 12579 17496 12624 17524
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 14366 17524 14372 17536
rect 14327 17496 14372 17524
rect 14366 17484 14372 17496
rect 14424 17484 14430 17536
rect 14461 17527 14519 17533
rect 14461 17493 14473 17527
rect 14507 17524 14519 17527
rect 14550 17524 14556 17536
rect 14507 17496 14556 17524
rect 14507 17493 14519 17496
rect 14461 17487 14519 17493
rect 14550 17484 14556 17496
rect 14608 17484 14614 17536
rect 14829 17527 14887 17533
rect 14829 17493 14841 17527
rect 14875 17524 14887 17527
rect 15102 17524 15108 17536
rect 14875 17496 15108 17524
rect 14875 17493 14887 17496
rect 14829 17487 14887 17493
rect 15102 17484 15108 17496
rect 15160 17484 15166 17536
rect 15562 17524 15568 17536
rect 15523 17496 15568 17524
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 16114 17524 16120 17536
rect 16075 17496 16120 17524
rect 16114 17484 16120 17496
rect 16172 17484 16178 17536
rect 16390 17484 16396 17536
rect 16448 17524 16454 17536
rect 16485 17527 16543 17533
rect 16485 17524 16497 17527
rect 16448 17496 16497 17524
rect 16448 17484 16454 17496
rect 16485 17493 16497 17496
rect 16531 17493 16543 17527
rect 17494 17524 17500 17536
rect 17455 17496 17500 17524
rect 16485 17487 16543 17493
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 20809 17527 20867 17533
rect 20809 17493 20821 17527
rect 20855 17524 20867 17527
rect 21082 17524 21088 17536
rect 20855 17496 21088 17524
rect 20855 17493 20867 17496
rect 20809 17487 20867 17493
rect 21082 17484 21088 17496
rect 21140 17484 21146 17536
rect 21266 17524 21272 17536
rect 21227 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 2409 17323 2467 17329
rect 2409 17289 2421 17323
rect 2455 17289 2467 17323
rect 3878 17320 3884 17332
rect 3839 17292 3884 17320
rect 2409 17283 2467 17289
rect 2424 17252 2452 17283
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 4982 17320 4988 17332
rect 4943 17292 4988 17320
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 5721 17323 5779 17329
rect 5721 17289 5733 17323
rect 5767 17320 5779 17323
rect 5994 17320 6000 17332
rect 5767 17292 6000 17320
rect 5767 17289 5779 17292
rect 5721 17283 5779 17289
rect 5994 17280 6000 17292
rect 6052 17320 6058 17332
rect 6365 17323 6423 17329
rect 6365 17320 6377 17323
rect 6052 17292 6377 17320
rect 6052 17280 6058 17292
rect 6365 17289 6377 17292
rect 6411 17289 6423 17323
rect 6365 17283 6423 17289
rect 6730 17280 6736 17332
rect 6788 17320 6794 17332
rect 6917 17323 6975 17329
rect 6917 17320 6929 17323
rect 6788 17292 6929 17320
rect 6788 17280 6794 17292
rect 6917 17289 6929 17292
rect 6963 17289 6975 17323
rect 8205 17323 8263 17329
rect 8205 17320 8217 17323
rect 6917 17283 6975 17289
rect 7024 17292 8217 17320
rect 1688 17224 2452 17252
rect 3421 17255 3479 17261
rect 1688 17193 1716 17224
rect 3421 17221 3433 17255
rect 3467 17252 3479 17255
rect 4890 17252 4896 17264
rect 3467 17224 4896 17252
rect 3467 17221 3479 17224
rect 3421 17215 3479 17221
rect 4890 17212 4896 17224
rect 4948 17212 4954 17264
rect 5534 17212 5540 17264
rect 5592 17252 5598 17264
rect 5629 17255 5687 17261
rect 5629 17252 5641 17255
rect 5592 17224 5641 17252
rect 5592 17212 5598 17224
rect 5629 17221 5641 17224
rect 5675 17252 5687 17255
rect 6086 17252 6092 17264
rect 5675 17224 6092 17252
rect 5675 17221 5687 17224
rect 5629 17215 5687 17221
rect 6086 17212 6092 17224
rect 6144 17212 6150 17264
rect 1673 17187 1731 17193
rect 1673 17153 1685 17187
rect 1719 17153 1731 17187
rect 1673 17147 1731 17153
rect 2133 17187 2191 17193
rect 2133 17153 2145 17187
rect 2179 17153 2191 17187
rect 2590 17184 2596 17196
rect 2551 17156 2596 17184
rect 2133 17147 2191 17153
rect 2148 17116 2176 17147
rect 2590 17144 2596 17156
rect 2648 17144 2654 17196
rect 2958 17144 2964 17196
rect 3016 17184 3022 17196
rect 3513 17187 3571 17193
rect 3513 17184 3525 17187
rect 3016 17156 3525 17184
rect 3016 17144 3022 17156
rect 3513 17153 3525 17156
rect 3559 17153 3571 17187
rect 3513 17147 3571 17153
rect 4617 17187 4675 17193
rect 4617 17153 4629 17187
rect 4663 17184 4675 17187
rect 6546 17184 6552 17196
rect 4663 17156 6552 17184
rect 4663 17153 4675 17156
rect 4617 17147 4675 17153
rect 6546 17144 6552 17156
rect 6604 17184 6610 17196
rect 7024 17184 7052 17292
rect 8205 17289 8217 17292
rect 8251 17289 8263 17323
rect 8205 17283 8263 17289
rect 8665 17323 8723 17329
rect 8665 17289 8677 17323
rect 8711 17289 8723 17323
rect 8665 17283 8723 17289
rect 9125 17323 9183 17329
rect 9125 17289 9137 17323
rect 9171 17320 9183 17323
rect 9306 17320 9312 17332
rect 9171 17292 9312 17320
rect 9171 17289 9183 17292
rect 9125 17283 9183 17289
rect 8680 17252 8708 17283
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 10781 17323 10839 17329
rect 10781 17289 10793 17323
rect 10827 17320 10839 17323
rect 11977 17323 12035 17329
rect 11977 17320 11989 17323
rect 10827 17292 11989 17320
rect 10827 17289 10839 17292
rect 10781 17283 10839 17289
rect 11977 17289 11989 17292
rect 12023 17289 12035 17323
rect 11977 17283 12035 17289
rect 12345 17323 12403 17329
rect 12345 17289 12357 17323
rect 12391 17320 12403 17323
rect 12894 17320 12900 17332
rect 12391 17292 12900 17320
rect 12391 17289 12403 17292
rect 12345 17283 12403 17289
rect 12894 17280 12900 17292
rect 12952 17280 12958 17332
rect 14366 17320 14372 17332
rect 14327 17292 14372 17320
rect 14366 17280 14372 17292
rect 14424 17280 14430 17332
rect 14737 17323 14795 17329
rect 14737 17289 14749 17323
rect 14783 17320 14795 17323
rect 14918 17320 14924 17332
rect 14783 17292 14924 17320
rect 14783 17289 14795 17292
rect 14737 17283 14795 17289
rect 14918 17280 14924 17292
rect 14976 17280 14982 17332
rect 15102 17320 15108 17332
rect 15063 17292 15108 17320
rect 15102 17280 15108 17292
rect 15160 17280 15166 17332
rect 15197 17323 15255 17329
rect 15197 17289 15209 17323
rect 15243 17320 15255 17323
rect 16114 17320 16120 17332
rect 15243 17292 16120 17320
rect 15243 17289 15255 17292
rect 15197 17283 15255 17289
rect 16114 17280 16120 17292
rect 16172 17280 16178 17332
rect 16390 17280 16396 17332
rect 16448 17320 16454 17332
rect 16669 17323 16727 17329
rect 16669 17320 16681 17323
rect 16448 17292 16681 17320
rect 16448 17280 16454 17292
rect 16669 17289 16681 17292
rect 16715 17289 16727 17323
rect 17954 17320 17960 17332
rect 16669 17283 16727 17289
rect 16776 17292 17960 17320
rect 12618 17252 12624 17264
rect 8680 17224 12624 17252
rect 12618 17212 12624 17224
rect 12676 17212 12682 17264
rect 12912 17224 14136 17252
rect 7282 17184 7288 17196
rect 6604 17156 7052 17184
rect 7243 17156 7288 17184
rect 6604 17144 6610 17156
rect 7282 17144 7288 17156
rect 7340 17144 7346 17196
rect 8297 17187 8355 17193
rect 8297 17184 8309 17187
rect 7392 17156 8309 17184
rect 7392 17128 7420 17156
rect 8297 17153 8309 17156
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 9493 17187 9551 17193
rect 9493 17153 9505 17187
rect 9539 17184 9551 17187
rect 10502 17184 10508 17196
rect 9539 17156 10508 17184
rect 9539 17153 9551 17156
rect 9493 17147 9551 17153
rect 10502 17144 10508 17156
rect 10560 17144 10566 17196
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17184 11759 17187
rect 12342 17184 12348 17196
rect 11747 17156 12348 17184
rect 11747 17153 11759 17156
rect 11701 17147 11759 17153
rect 12342 17144 12348 17156
rect 12400 17184 12406 17196
rect 12437 17187 12495 17193
rect 12437 17184 12449 17187
rect 12400 17156 12449 17184
rect 12400 17144 12406 17156
rect 12437 17153 12449 17156
rect 12483 17184 12495 17187
rect 12912 17184 12940 17224
rect 12483 17156 12940 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 13262 17144 13268 17196
rect 13320 17184 13326 17196
rect 13357 17187 13415 17193
rect 13357 17184 13369 17187
rect 13320 17156 13369 17184
rect 13320 17144 13326 17156
rect 13357 17153 13369 17156
rect 13403 17184 13415 17187
rect 14001 17187 14059 17193
rect 14001 17184 14013 17187
rect 13403 17156 14013 17184
rect 13403 17153 13415 17156
rect 13357 17147 13415 17153
rect 14001 17153 14013 17156
rect 14047 17153 14059 17187
rect 14108 17184 14136 17224
rect 16776 17184 16804 17292
rect 17954 17280 17960 17292
rect 18012 17280 18018 17332
rect 18138 17320 18144 17332
rect 18099 17292 18144 17320
rect 18138 17280 18144 17292
rect 18196 17280 18202 17332
rect 20073 17323 20131 17329
rect 19168 17292 19932 17320
rect 17402 17212 17408 17264
rect 17460 17252 17466 17264
rect 19168 17252 19196 17292
rect 17460 17224 19196 17252
rect 19276 17255 19334 17261
rect 17460 17212 17466 17224
rect 19276 17221 19288 17255
rect 19322 17252 19334 17255
rect 19794 17252 19800 17264
rect 19322 17224 19800 17252
rect 19322 17221 19334 17224
rect 19276 17215 19334 17221
rect 19794 17212 19800 17224
rect 19852 17212 19858 17264
rect 14108 17156 16804 17184
rect 17037 17187 17095 17193
rect 14001 17147 14059 17153
rect 17037 17153 17049 17187
rect 17083 17184 17095 17187
rect 17770 17184 17776 17196
rect 17083 17156 17776 17184
rect 17083 17153 17095 17156
rect 17037 17147 17095 17153
rect 3234 17116 3240 17128
rect 2148 17088 3240 17116
rect 3234 17076 3240 17088
rect 3292 17076 3298 17128
rect 3329 17119 3387 17125
rect 3329 17085 3341 17119
rect 3375 17085 3387 17119
rect 3329 17079 3387 17085
rect 4433 17119 4491 17125
rect 4433 17085 4445 17119
rect 4479 17085 4491 17119
rect 4433 17079 4491 17085
rect 4525 17119 4583 17125
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4571 17088 5304 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 1486 17048 1492 17060
rect 1447 17020 1492 17048
rect 1486 17008 1492 17020
rect 1544 17008 1550 17060
rect 2866 17008 2872 17060
rect 2924 17048 2930 17060
rect 3344 17048 3372 17079
rect 4448 17048 4476 17079
rect 5276 17057 5304 17088
rect 5810 17076 5816 17128
rect 5868 17116 5874 17128
rect 7374 17116 7380 17128
rect 5868 17088 5913 17116
rect 7335 17088 7380 17116
rect 5868 17076 5874 17088
rect 7374 17076 7380 17088
rect 7432 17076 7438 17128
rect 7469 17119 7527 17125
rect 7469 17085 7481 17119
rect 7515 17085 7527 17119
rect 8110 17116 8116 17128
rect 8071 17088 8116 17116
rect 7469 17079 7527 17085
rect 5261 17051 5319 17057
rect 2924 17020 4752 17048
rect 2924 17008 2930 17020
rect 1946 16980 1952 16992
rect 1907 16952 1952 16980
rect 1946 16940 1952 16952
rect 2004 16940 2010 16992
rect 4724 16980 4752 17020
rect 5261 17017 5273 17051
rect 5307 17017 5319 17051
rect 5261 17011 5319 17017
rect 5902 17008 5908 17060
rect 5960 17048 5966 17060
rect 7484 17048 7512 17079
rect 8110 17076 8116 17088
rect 8168 17076 8174 17128
rect 8570 17076 8576 17128
rect 8628 17116 8634 17128
rect 9582 17116 9588 17128
rect 8628 17088 9588 17116
rect 8628 17076 8634 17088
rect 9582 17076 9588 17088
rect 9640 17076 9646 17128
rect 9677 17119 9735 17125
rect 9677 17085 9689 17119
rect 9723 17085 9735 17119
rect 9677 17079 9735 17085
rect 5960 17020 7512 17048
rect 5960 17008 5966 17020
rect 8662 17008 8668 17060
rect 8720 17048 8726 17060
rect 9692 17048 9720 17079
rect 10410 17076 10416 17128
rect 10468 17116 10474 17128
rect 10597 17119 10655 17125
rect 10597 17116 10609 17119
rect 10468 17088 10609 17116
rect 10468 17076 10474 17088
rect 10597 17085 10609 17088
rect 10643 17085 10655 17119
rect 10597 17079 10655 17085
rect 10689 17119 10747 17125
rect 10689 17085 10701 17119
rect 10735 17116 10747 17119
rect 11054 17116 11060 17128
rect 10735 17088 11060 17116
rect 10735 17085 10747 17088
rect 10689 17079 10747 17085
rect 11054 17076 11060 17088
rect 11112 17076 11118 17128
rect 12158 17076 12164 17128
rect 12216 17116 12222 17128
rect 12621 17119 12679 17125
rect 12621 17116 12633 17119
rect 12216 17088 12633 17116
rect 12216 17076 12222 17088
rect 12621 17085 12633 17088
rect 12667 17085 12679 17119
rect 12621 17079 12679 17085
rect 13630 17076 13636 17128
rect 13688 17116 13694 17128
rect 13817 17119 13875 17125
rect 13817 17116 13829 17119
rect 13688 17088 13829 17116
rect 13688 17076 13694 17088
rect 13817 17085 13829 17088
rect 13863 17085 13875 17119
rect 13817 17079 13875 17085
rect 13909 17119 13967 17125
rect 13909 17085 13921 17119
rect 13955 17085 13967 17119
rect 14016 17116 14044 17147
rect 17770 17144 17776 17156
rect 17828 17144 17834 17196
rect 18874 17184 18880 17196
rect 17880 17156 18880 17184
rect 14642 17116 14648 17128
rect 14016 17088 14648 17116
rect 13909 17079 13967 17085
rect 12526 17048 12532 17060
rect 8720 17020 9720 17048
rect 9784 17020 12532 17048
rect 8720 17008 8726 17020
rect 4798 16980 4804 16992
rect 4711 16952 4804 16980
rect 4798 16940 4804 16952
rect 4856 16980 4862 16992
rect 5920 16980 5948 17008
rect 4856 16952 5948 16980
rect 4856 16940 4862 16952
rect 6086 16940 6092 16992
rect 6144 16980 6150 16992
rect 9784 16980 9812 17020
rect 12526 17008 12532 17020
rect 12584 17008 12590 17060
rect 13924 17048 13952 17079
rect 14642 17076 14648 17088
rect 14700 17076 14706 17128
rect 15381 17119 15439 17125
rect 15381 17085 15393 17119
rect 15427 17116 15439 17119
rect 15470 17116 15476 17128
rect 15427 17088 15476 17116
rect 15427 17085 15439 17088
rect 15381 17079 15439 17085
rect 15470 17076 15476 17088
rect 15528 17076 15534 17128
rect 17126 17116 17132 17128
rect 17087 17088 17132 17116
rect 17126 17076 17132 17088
rect 17184 17076 17190 17128
rect 17218 17076 17224 17128
rect 17276 17116 17282 17128
rect 17276 17088 17321 17116
rect 17276 17076 17282 17088
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 17880 17116 17908 17156
rect 18874 17144 18880 17156
rect 18932 17184 18938 17196
rect 19904 17193 19932 17292
rect 20073 17289 20085 17323
rect 20119 17320 20131 17323
rect 20622 17320 20628 17332
rect 20119 17292 20628 17320
rect 20119 17289 20131 17292
rect 20073 17283 20131 17289
rect 20622 17280 20628 17292
rect 20680 17280 20686 17332
rect 19521 17187 19579 17193
rect 19521 17184 19533 17187
rect 18932 17156 19533 17184
rect 18932 17144 18938 17156
rect 19521 17153 19533 17156
rect 19567 17153 19579 17187
rect 19521 17147 19579 17153
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17184 20683 17187
rect 20806 17184 20812 17196
rect 20671 17156 20812 17184
rect 20671 17153 20683 17156
rect 20625 17147 20683 17153
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 21082 17184 21088 17196
rect 21043 17156 21088 17184
rect 21082 17144 21088 17156
rect 21140 17144 21146 17196
rect 17552 17088 17908 17116
rect 17552 17076 17558 17088
rect 15102 17048 15108 17060
rect 13924 17020 15108 17048
rect 15102 17008 15108 17020
rect 15160 17048 15166 17060
rect 17954 17048 17960 17060
rect 15160 17020 17960 17048
rect 15160 17008 15166 17020
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 11146 16980 11152 16992
rect 6144 16952 9812 16980
rect 11107 16952 11152 16980
rect 6144 16940 6150 16952
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 13814 16980 13820 16992
rect 11848 16952 13820 16980
rect 11848 16940 11854 16952
rect 13814 16940 13820 16952
rect 13872 16940 13878 16992
rect 17126 16940 17132 16992
rect 17184 16980 17190 16992
rect 17681 16983 17739 16989
rect 17681 16980 17693 16983
rect 17184 16952 17693 16980
rect 17184 16940 17190 16952
rect 17681 16949 17693 16952
rect 17727 16949 17739 16983
rect 17681 16943 17739 16949
rect 20809 16983 20867 16989
rect 20809 16949 20821 16983
rect 20855 16980 20867 16983
rect 21082 16980 21088 16992
rect 20855 16952 21088 16980
rect 20855 16949 20867 16952
rect 20809 16943 20867 16949
rect 21082 16940 21088 16952
rect 21140 16940 21146 16992
rect 21266 16980 21272 16992
rect 21227 16952 21272 16980
rect 21266 16940 21272 16952
rect 21324 16940 21330 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 2774 16736 2780 16788
rect 2832 16776 2838 16788
rect 5810 16776 5816 16788
rect 2832 16748 5396 16776
rect 5771 16748 5816 16776
rect 2832 16736 2838 16748
rect 2498 16668 2504 16720
rect 2556 16708 2562 16720
rect 5368 16708 5396 16748
rect 5810 16736 5816 16748
rect 5868 16736 5874 16788
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 8570 16776 8576 16788
rect 7340 16748 8248 16776
rect 8531 16748 8576 16776
rect 7340 16736 7346 16748
rect 7650 16708 7656 16720
rect 2556 16680 3004 16708
rect 5368 16680 7656 16708
rect 2556 16668 2562 16680
rect 2866 16640 2872 16652
rect 2827 16612 2872 16640
rect 2866 16600 2872 16612
rect 2924 16600 2930 16652
rect 2976 16649 3004 16680
rect 7650 16668 7656 16680
rect 7708 16668 7714 16720
rect 8220 16717 8248 16748
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 8662 16736 8668 16788
rect 8720 16776 8726 16788
rect 8941 16779 8999 16785
rect 8941 16776 8953 16779
rect 8720 16748 8953 16776
rect 8720 16736 8726 16748
rect 8941 16745 8953 16748
rect 8987 16745 8999 16779
rect 8941 16739 8999 16745
rect 9416 16748 10364 16776
rect 8205 16711 8263 16717
rect 8205 16677 8217 16711
rect 8251 16708 8263 16711
rect 9416 16708 9444 16748
rect 8251 16680 9444 16708
rect 10336 16708 10364 16748
rect 10502 16736 10508 16788
rect 10560 16776 10566 16788
rect 10597 16779 10655 16785
rect 10597 16776 10609 16779
rect 10560 16748 10609 16776
rect 10560 16736 10566 16748
rect 10597 16745 10609 16748
rect 10643 16776 10655 16779
rect 12618 16776 12624 16788
rect 10643 16748 12624 16776
rect 10643 16745 10655 16748
rect 10597 16739 10655 16745
rect 12618 16736 12624 16748
rect 12676 16776 12682 16788
rect 13725 16779 13783 16785
rect 13725 16776 13737 16779
rect 12676 16748 13737 16776
rect 12676 16736 12682 16748
rect 10686 16708 10692 16720
rect 10336 16680 10692 16708
rect 8251 16677 8263 16680
rect 8205 16671 8263 16677
rect 10686 16668 10692 16680
rect 10744 16668 10750 16720
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16609 3019 16643
rect 2961 16603 3019 16609
rect 3234 16600 3240 16652
rect 3292 16640 3298 16652
rect 3789 16643 3847 16649
rect 3789 16640 3801 16643
rect 3292 16612 3801 16640
rect 3292 16600 3298 16612
rect 3789 16609 3801 16612
rect 3835 16609 3847 16643
rect 3789 16603 3847 16609
rect 4338 16600 4344 16652
rect 4396 16640 4402 16652
rect 4433 16643 4491 16649
rect 4433 16640 4445 16643
rect 4396 16612 4445 16640
rect 4396 16600 4402 16612
rect 4433 16609 4445 16612
rect 4479 16609 4491 16643
rect 4433 16603 4491 16609
rect 5626 16600 5632 16652
rect 5684 16640 5690 16652
rect 7285 16643 7343 16649
rect 5684 16612 7236 16640
rect 5684 16600 5690 16612
rect 1670 16572 1676 16584
rect 1631 16544 1676 16572
rect 1670 16532 1676 16544
rect 1728 16532 1734 16584
rect 1946 16572 1952 16584
rect 1907 16544 1952 16572
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 3053 16575 3111 16581
rect 3053 16541 3065 16575
rect 3099 16572 3111 16575
rect 3142 16572 3148 16584
rect 3099 16544 3148 16572
rect 3099 16541 3111 16544
rect 3053 16535 3111 16541
rect 3142 16532 3148 16544
rect 3200 16532 3206 16584
rect 5810 16532 5816 16584
rect 5868 16572 5874 16584
rect 6089 16575 6147 16581
rect 6089 16572 6101 16575
rect 5868 16544 6101 16572
rect 5868 16532 5874 16544
rect 6089 16541 6101 16544
rect 6135 16541 6147 16575
rect 6089 16535 6147 16541
rect 6733 16575 6791 16581
rect 6733 16541 6745 16575
rect 6779 16572 6791 16575
rect 6914 16572 6920 16584
rect 6779 16544 6920 16572
rect 6779 16541 6791 16544
rect 6733 16535 6791 16541
rect 6914 16532 6920 16544
rect 6972 16532 6978 16584
rect 7208 16572 7236 16612
rect 7285 16609 7297 16643
rect 7331 16640 7343 16643
rect 8662 16640 8668 16652
rect 7331 16612 8668 16640
rect 7331 16609 7343 16612
rect 7285 16603 7343 16609
rect 8662 16600 8668 16612
rect 8720 16600 8726 16652
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16640 10379 16643
rect 10962 16640 10968 16652
rect 10367 16612 10968 16640
rect 10367 16609 10379 16612
rect 10321 16603 10379 16609
rect 7377 16575 7435 16581
rect 7377 16572 7389 16575
rect 7208 16544 7389 16572
rect 7377 16541 7389 16544
rect 7423 16541 7435 16575
rect 7377 16535 7435 16541
rect 9490 16532 9496 16584
rect 9548 16572 9554 16584
rect 10336 16572 10364 16603
rect 10962 16600 10968 16612
rect 11020 16600 11026 16652
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 11974 16640 11980 16652
rect 11563 16612 11980 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12250 16640 12256 16652
rect 12084 16612 12256 16640
rect 9548 16544 10364 16572
rect 9548 16532 9554 16544
rect 11146 16532 11152 16584
rect 11204 16572 11210 16584
rect 11701 16575 11759 16581
rect 11701 16572 11713 16575
rect 11204 16544 11713 16572
rect 11204 16532 11210 16544
rect 11701 16541 11713 16544
rect 11747 16541 11759 16575
rect 11701 16535 11759 16541
rect 4700 16507 4758 16513
rect 4700 16473 4712 16507
rect 4746 16504 4758 16507
rect 5718 16504 5724 16516
rect 4746 16476 5724 16504
rect 4746 16473 4758 16476
rect 4700 16467 4758 16473
rect 5718 16464 5724 16476
rect 5776 16464 5782 16516
rect 10076 16507 10134 16513
rect 10076 16473 10088 16507
rect 10122 16504 10134 16507
rect 10318 16504 10324 16516
rect 10122 16476 10324 16504
rect 10122 16473 10134 16476
rect 10076 16467 10134 16473
rect 10318 16464 10324 16476
rect 10376 16464 10382 16516
rect 11609 16507 11667 16513
rect 11609 16473 11621 16507
rect 11655 16504 11667 16507
rect 12084 16504 12112 16612
rect 12250 16600 12256 16612
rect 12308 16600 12314 16652
rect 12894 16600 12900 16652
rect 12952 16640 12958 16652
rect 13265 16643 13323 16649
rect 13265 16640 13277 16643
rect 12952 16612 13277 16640
rect 12952 16600 12958 16612
rect 13265 16609 13277 16612
rect 13311 16609 13323 16643
rect 13556 16640 13584 16748
rect 13725 16745 13737 16748
rect 13771 16745 13783 16779
rect 13725 16739 13783 16745
rect 14829 16779 14887 16785
rect 14829 16745 14841 16779
rect 14875 16776 14887 16779
rect 15562 16776 15568 16788
rect 14875 16748 15568 16776
rect 14875 16745 14887 16748
rect 14829 16739 14887 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 16298 16736 16304 16788
rect 16356 16776 16362 16788
rect 16393 16779 16451 16785
rect 16393 16776 16405 16779
rect 16356 16748 16405 16776
rect 16356 16736 16362 16748
rect 16393 16745 16405 16748
rect 16439 16745 16451 16779
rect 16393 16739 16451 16745
rect 17770 16736 17776 16788
rect 17828 16776 17834 16788
rect 18417 16779 18475 16785
rect 18417 16776 18429 16779
rect 17828 16748 18429 16776
rect 17828 16736 17834 16748
rect 18417 16745 18429 16748
rect 18463 16745 18475 16779
rect 20346 16776 20352 16788
rect 20307 16748 20352 16776
rect 18417 16739 18475 16745
rect 20346 16736 20352 16748
rect 20404 16736 20410 16788
rect 20806 16776 20812 16788
rect 20767 16748 20812 16776
rect 20806 16736 20812 16748
rect 20864 16736 20870 16788
rect 13630 16668 13636 16720
rect 13688 16708 13694 16720
rect 16022 16708 16028 16720
rect 13688 16680 15884 16708
rect 15983 16680 16028 16708
rect 13688 16668 13694 16680
rect 14277 16643 14335 16649
rect 13556 16612 14228 16640
rect 13265 16603 13323 16609
rect 14200 16572 14228 16612
rect 14277 16609 14289 16643
rect 14323 16640 14335 16643
rect 14458 16640 14464 16652
rect 14323 16612 14464 16640
rect 14323 16609 14335 16612
rect 14277 16603 14335 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 15102 16640 15108 16652
rect 15063 16612 15108 16640
rect 15102 16600 15108 16612
rect 15160 16600 15166 16652
rect 15856 16640 15884 16680
rect 16022 16668 16028 16680
rect 16080 16668 16086 16720
rect 16206 16668 16212 16720
rect 16264 16708 16270 16720
rect 17405 16711 17463 16717
rect 17405 16708 17417 16711
rect 16264 16680 17417 16708
rect 16264 16668 16270 16680
rect 17405 16677 17417 16680
rect 17451 16677 17463 16711
rect 17405 16671 17463 16677
rect 17586 16668 17592 16720
rect 17644 16708 17650 16720
rect 17644 16680 18000 16708
rect 17644 16668 17650 16680
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 15856 16612 16957 16640
rect 16945 16609 16957 16612
rect 16991 16640 17003 16643
rect 17218 16640 17224 16652
rect 16991 16612 17224 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17218 16600 17224 16612
rect 17276 16600 17282 16652
rect 17862 16640 17868 16652
rect 17823 16612 17868 16640
rect 17862 16600 17868 16612
rect 17920 16600 17926 16652
rect 17972 16649 18000 16680
rect 17957 16643 18015 16649
rect 17957 16609 17969 16643
rect 18003 16609 18015 16643
rect 20346 16640 20352 16652
rect 17957 16603 18015 16609
rect 18064 16612 20352 16640
rect 14369 16575 14427 16581
rect 14369 16572 14381 16575
rect 14200 16544 14381 16572
rect 14369 16541 14381 16544
rect 14415 16541 14427 16575
rect 14369 16535 14427 16541
rect 16761 16575 16819 16581
rect 16761 16541 16773 16575
rect 16807 16572 16819 16575
rect 17586 16572 17592 16584
rect 16807 16544 17592 16572
rect 16807 16541 16819 16544
rect 16761 16535 16819 16541
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 17678 16532 17684 16584
rect 17736 16572 17742 16584
rect 18064 16572 18092 16612
rect 20346 16600 20352 16612
rect 20404 16600 20410 16652
rect 17736 16544 18092 16572
rect 17736 16532 17742 16544
rect 18506 16532 18512 16584
rect 18564 16572 18570 16584
rect 19245 16575 19303 16581
rect 19245 16572 19257 16575
rect 18564 16544 19257 16572
rect 18564 16532 18570 16544
rect 19245 16541 19257 16544
rect 19291 16541 19303 16575
rect 19245 16535 19303 16541
rect 19794 16532 19800 16584
rect 19852 16572 19858 16584
rect 19889 16575 19947 16581
rect 19889 16572 19901 16575
rect 19852 16544 19901 16572
rect 19852 16532 19858 16544
rect 19889 16541 19901 16544
rect 19935 16541 19947 16575
rect 20162 16572 20168 16584
rect 20123 16544 20168 16572
rect 19889 16535 19947 16541
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20625 16575 20683 16581
rect 20625 16541 20637 16575
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 20640 16504 20668 16535
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20772 16544 21097 16572
rect 20772 16532 20778 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 11655 16476 12112 16504
rect 12820 16476 20668 16504
rect 11655 16473 11667 16476
rect 11609 16467 11667 16473
rect 1486 16436 1492 16448
rect 1447 16408 1492 16436
rect 1486 16396 1492 16408
rect 1544 16396 1550 16448
rect 2130 16436 2136 16448
rect 2091 16408 2136 16436
rect 2130 16396 2136 16408
rect 2188 16396 2194 16448
rect 3418 16436 3424 16448
rect 3379 16408 3424 16436
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 7469 16439 7527 16445
rect 7469 16436 7481 16439
rect 7156 16408 7481 16436
rect 7156 16396 7162 16408
rect 7469 16405 7481 16408
rect 7515 16405 7527 16439
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7469 16399 7527 16405
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 12069 16439 12127 16445
rect 12069 16405 12081 16439
rect 12115 16436 12127 16439
rect 12820 16436 12848 16476
rect 12115 16408 12848 16436
rect 12115 16405 12127 16408
rect 12069 16399 12127 16405
rect 12894 16396 12900 16448
rect 12952 16436 12958 16448
rect 14461 16439 14519 16445
rect 14461 16436 14473 16439
rect 12952 16408 14473 16436
rect 12952 16396 12958 16408
rect 14461 16405 14473 16408
rect 14507 16436 14519 16439
rect 15010 16436 15016 16448
rect 14507 16408 15016 16436
rect 14507 16405 14519 16408
rect 14461 16399 14519 16405
rect 15010 16396 15016 16408
rect 15068 16396 15074 16448
rect 16853 16439 16911 16445
rect 16853 16405 16865 16439
rect 16899 16436 16911 16439
rect 17678 16436 17684 16448
rect 16899 16408 17684 16436
rect 16899 16405 16911 16408
rect 16853 16399 16911 16405
rect 17678 16396 17684 16408
rect 17736 16396 17742 16448
rect 17773 16439 17831 16445
rect 17773 16405 17785 16439
rect 17819 16436 17831 16439
rect 17954 16436 17960 16448
rect 17819 16408 17960 16436
rect 17819 16405 17831 16408
rect 17773 16399 17831 16405
rect 17954 16396 17960 16408
rect 18012 16436 18018 16448
rect 18785 16439 18843 16445
rect 18785 16436 18797 16439
rect 18012 16408 18797 16436
rect 18012 16396 18018 16408
rect 18785 16405 18797 16408
rect 18831 16405 18843 16439
rect 21266 16436 21272 16448
rect 21227 16408 21272 16436
rect 18785 16399 18843 16405
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 1949 16235 2007 16241
rect 1949 16201 1961 16235
rect 1995 16201 2007 16235
rect 2590 16232 2596 16244
rect 2551 16204 2596 16232
rect 1949 16195 2007 16201
rect 1673 16099 1731 16105
rect 1673 16065 1685 16099
rect 1719 16096 1731 16099
rect 1964 16096 1992 16195
rect 2590 16192 2596 16204
rect 2648 16192 2654 16244
rect 3326 16192 3332 16244
rect 3384 16232 3390 16244
rect 8021 16235 8079 16241
rect 8021 16232 8033 16235
rect 3384 16204 8033 16232
rect 3384 16192 3390 16204
rect 8021 16201 8033 16204
rect 8067 16201 8079 16235
rect 8021 16195 8079 16201
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 11517 16235 11575 16241
rect 11517 16232 11529 16235
rect 11112 16204 11529 16232
rect 11112 16192 11118 16204
rect 11517 16201 11529 16204
rect 11563 16201 11575 16235
rect 18322 16232 18328 16244
rect 11517 16195 11575 16201
rect 14660 16204 18328 16232
rect 2682 16124 2688 16176
rect 2740 16164 2746 16176
rect 3973 16167 4031 16173
rect 3973 16164 3985 16167
rect 2740 16136 3985 16164
rect 2740 16124 2746 16136
rect 3973 16133 3985 16136
rect 4019 16133 4031 16167
rect 7558 16164 7564 16176
rect 3973 16127 4031 16133
rect 4908 16136 7564 16164
rect 1719 16068 1992 16096
rect 2133 16099 2191 16105
rect 1719 16065 1731 16068
rect 1673 16059 1731 16065
rect 2133 16065 2145 16099
rect 2179 16065 2191 16099
rect 2133 16059 2191 16065
rect 2409 16099 2467 16105
rect 2409 16065 2421 16099
rect 2455 16096 2467 16099
rect 4798 16096 4804 16108
rect 2455 16068 4804 16096
rect 2455 16065 2467 16068
rect 2409 16059 2467 16065
rect 2148 16028 2176 16059
rect 4798 16056 4804 16068
rect 4856 16056 4862 16108
rect 2148 16000 2774 16028
rect 2746 15960 2774 16000
rect 2866 15988 2872 16040
rect 2924 16028 2930 16040
rect 3237 16031 3295 16037
rect 3237 16028 3249 16031
rect 2924 16000 3249 16028
rect 2924 15988 2930 16000
rect 3237 15997 3249 16000
rect 3283 15997 3295 16031
rect 3237 15991 3295 15997
rect 3697 16031 3755 16037
rect 3697 15997 3709 16031
rect 3743 16028 3755 16031
rect 3970 16028 3976 16040
rect 3743 16000 3976 16028
rect 3743 15997 3755 16000
rect 3697 15991 3755 15997
rect 3970 15988 3976 16000
rect 4028 15988 4034 16040
rect 2961 15963 3019 15969
rect 2961 15960 2973 15963
rect 2746 15932 2973 15960
rect 2961 15929 2973 15932
rect 3007 15960 3019 15963
rect 4908 15960 4936 16136
rect 7558 16124 7564 16136
rect 7616 16124 7622 16176
rect 8389 16099 8447 16105
rect 8389 16096 8401 16099
rect 6196 16068 8401 16096
rect 4985 16031 5043 16037
rect 4985 15997 4997 16031
rect 5031 16028 5043 16031
rect 5074 16028 5080 16040
rect 5031 16000 5080 16028
rect 5031 15997 5043 16000
rect 4985 15991 5043 15997
rect 5074 15988 5080 16000
rect 5132 16028 5138 16040
rect 6196 16028 6224 16068
rect 8389 16065 8401 16068
rect 8435 16065 8447 16099
rect 9122 16096 9128 16108
rect 9083 16068 9128 16096
rect 8389 16059 8447 16065
rect 9122 16056 9128 16068
rect 9180 16056 9186 16108
rect 11054 16056 11060 16108
rect 11112 16096 11118 16108
rect 11882 16096 11888 16108
rect 11112 16068 11888 16096
rect 11112 16056 11118 16068
rect 11882 16056 11888 16068
rect 11940 16056 11946 16108
rect 14550 16096 14556 16108
rect 14511 16068 14556 16096
rect 14550 16056 14556 16068
rect 14608 16056 14614 16108
rect 5132 16000 6224 16028
rect 5132 15988 5138 16000
rect 6730 15988 6736 16040
rect 6788 16028 6794 16040
rect 7285 16031 7343 16037
rect 7285 16028 7297 16031
rect 6788 16000 7297 16028
rect 6788 15988 6794 16000
rect 7285 15997 7297 16000
rect 7331 15997 7343 16031
rect 7285 15991 7343 15997
rect 7745 16031 7803 16037
rect 7745 15997 7757 16031
rect 7791 16028 7803 16031
rect 8018 16028 8024 16040
rect 7791 16000 8024 16028
rect 7791 15997 7803 16000
rect 7745 15991 7803 15997
rect 8018 15988 8024 16000
rect 8076 15988 8082 16040
rect 8202 15988 8208 16040
rect 8260 16028 8266 16040
rect 10229 16031 10287 16037
rect 10229 16028 10241 16031
rect 8260 16000 10241 16028
rect 8260 15988 8266 16000
rect 10229 15997 10241 16000
rect 10275 15997 10287 16031
rect 11977 16031 12035 16037
rect 11977 16028 11989 16031
rect 10229 15991 10287 15997
rect 10704 16000 11989 16028
rect 5534 15960 5540 15972
rect 3007 15932 4936 15960
rect 5495 15932 5540 15960
rect 3007 15929 3019 15932
rect 2961 15923 3019 15929
rect 5534 15920 5540 15932
rect 5592 15920 5598 15972
rect 6457 15963 6515 15969
rect 6457 15929 6469 15963
rect 6503 15960 6515 15963
rect 7374 15960 7380 15972
rect 6503 15932 7380 15960
rect 6503 15929 6515 15932
rect 6457 15923 6515 15929
rect 7374 15920 7380 15932
rect 7432 15920 7438 15972
rect 10704 15904 10732 16000
rect 11977 15997 11989 16000
rect 12023 15997 12035 16031
rect 12158 16028 12164 16040
rect 12119 16000 12164 16028
rect 11977 15991 12035 15997
rect 12158 15988 12164 16000
rect 12216 15988 12222 16040
rect 13814 15988 13820 16040
rect 13872 16028 13878 16040
rect 14660 16037 14688 16204
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 19429 16235 19487 16241
rect 19429 16201 19441 16235
rect 19475 16232 19487 16235
rect 19610 16232 19616 16244
rect 19475 16204 19616 16232
rect 19475 16201 19487 16204
rect 19429 16195 19487 16201
rect 19610 16192 19616 16204
rect 19668 16192 19674 16244
rect 20162 16232 20168 16244
rect 20123 16204 20168 16232
rect 20162 16192 20168 16204
rect 20220 16192 20226 16244
rect 17221 16167 17279 16173
rect 17221 16133 17233 16167
rect 17267 16164 17279 16167
rect 18598 16164 18604 16176
rect 17267 16136 18604 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 18598 16124 18604 16136
rect 18656 16124 18662 16176
rect 15194 16096 15200 16108
rect 15155 16068 15200 16096
rect 15194 16056 15200 16068
rect 15252 16056 15258 16108
rect 17494 16096 17500 16108
rect 17455 16068 17500 16096
rect 17494 16056 17500 16068
rect 17552 16056 17558 16108
rect 17764 16099 17822 16105
rect 17764 16065 17776 16099
rect 17810 16096 17822 16099
rect 18046 16096 18052 16108
rect 17810 16068 18052 16096
rect 17810 16065 17822 16068
rect 17764 16059 17822 16065
rect 18046 16056 18052 16068
rect 18104 16056 18110 16108
rect 18230 16056 18236 16108
rect 18288 16096 18294 16108
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 18288 16068 19993 16096
rect 18288 16056 18294 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 20625 16059 20683 16065
rect 20824 16068 21097 16096
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 13872 16000 14657 16028
rect 13872 15988 13878 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 14737 16031 14795 16037
rect 14737 15997 14749 16031
rect 14783 15997 14795 16031
rect 14737 15991 14795 15997
rect 12802 15920 12808 15972
rect 12860 15960 12866 15972
rect 14752 15960 14780 15991
rect 19058 15988 19064 16040
rect 19116 16028 19122 16040
rect 20640 16028 20668 16059
rect 19116 16000 20668 16028
rect 19116 15988 19122 16000
rect 12860 15932 14780 15960
rect 12860 15920 12866 15932
rect 15010 15920 15016 15972
rect 15068 15960 15074 15972
rect 20824 15969 20852 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 20809 15963 20867 15969
rect 15068 15932 17540 15960
rect 15068 15920 15074 15932
rect 1486 15892 1492 15904
rect 1447 15864 1492 15892
rect 1486 15852 1492 15864
rect 1544 15852 1550 15904
rect 4154 15852 4160 15904
rect 4212 15892 4218 15904
rect 4341 15895 4399 15901
rect 4341 15892 4353 15895
rect 4212 15864 4353 15892
rect 4212 15852 4218 15864
rect 4341 15861 4353 15864
rect 4387 15861 4399 15895
rect 4341 15855 4399 15861
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5813 15895 5871 15901
rect 5813 15892 5825 15895
rect 5040 15864 5825 15892
rect 5040 15852 5046 15864
rect 5813 15861 5825 15864
rect 5859 15861 5871 15895
rect 5813 15855 5871 15861
rect 7009 15895 7067 15901
rect 7009 15861 7021 15895
rect 7055 15892 7067 15895
rect 7098 15892 7104 15904
rect 7055 15864 7104 15892
rect 7055 15861 7067 15864
rect 7009 15855 7067 15861
rect 7098 15852 7104 15864
rect 7156 15852 7162 15904
rect 8478 15852 8484 15904
rect 8536 15892 8542 15904
rect 8757 15895 8815 15901
rect 8757 15892 8769 15895
rect 8536 15864 8769 15892
rect 8536 15852 8542 15864
rect 8757 15861 8769 15864
rect 8803 15861 8815 15895
rect 9490 15892 9496 15904
rect 9451 15864 9496 15892
rect 8757 15855 8815 15861
rect 9490 15852 9496 15864
rect 9548 15852 9554 15904
rect 9858 15892 9864 15904
rect 9819 15864 9864 15892
rect 9858 15852 9864 15864
rect 9916 15852 9922 15904
rect 10686 15892 10692 15904
rect 10647 15864 10692 15892
rect 10686 15852 10692 15864
rect 10744 15852 10750 15904
rect 11054 15892 11060 15904
rect 11015 15864 11060 15892
rect 11054 15852 11060 15864
rect 11112 15852 11118 15904
rect 13814 15892 13820 15904
rect 13775 15864 13820 15892
rect 13814 15852 13820 15864
rect 13872 15852 13878 15904
rect 14185 15895 14243 15901
rect 14185 15861 14197 15895
rect 14231 15892 14243 15895
rect 14458 15892 14464 15904
rect 14231 15864 14464 15892
rect 14231 15861 14243 15864
rect 14185 15855 14243 15861
rect 14458 15852 14464 15864
rect 14516 15852 14522 15904
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 15841 15895 15899 15901
rect 15841 15892 15853 15895
rect 15804 15864 15853 15892
rect 15804 15852 15810 15864
rect 15841 15861 15853 15864
rect 15887 15861 15899 15895
rect 16206 15892 16212 15904
rect 16167 15864 16212 15892
rect 15841 15855 15899 15861
rect 16206 15852 16212 15864
rect 16264 15852 16270 15904
rect 16853 15895 16911 15901
rect 16853 15861 16865 15895
rect 16899 15892 16911 15895
rect 17402 15892 17408 15904
rect 16899 15864 17408 15892
rect 16899 15861 16911 15864
rect 16853 15855 16911 15861
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 17512 15892 17540 15932
rect 20809 15929 20821 15963
rect 20855 15929 20867 15963
rect 20809 15923 20867 15929
rect 18414 15892 18420 15904
rect 17512 15864 18420 15892
rect 18414 15852 18420 15864
rect 18472 15852 18478 15904
rect 18506 15852 18512 15904
rect 18564 15892 18570 15904
rect 18877 15895 18935 15901
rect 18877 15892 18889 15895
rect 18564 15864 18889 15892
rect 18564 15852 18570 15864
rect 18877 15861 18889 15864
rect 18923 15861 18935 15895
rect 21266 15892 21272 15904
rect 21227 15864 21272 15892
rect 18877 15855 18935 15861
rect 21266 15852 21272 15864
rect 21324 15852 21330 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1670 15648 1676 15700
rect 1728 15688 1734 15700
rect 2409 15691 2467 15697
rect 2409 15688 2421 15691
rect 1728 15660 2421 15688
rect 1728 15648 1734 15660
rect 2409 15657 2421 15660
rect 2455 15657 2467 15691
rect 3329 15691 3387 15697
rect 3329 15688 3341 15691
rect 2409 15651 2467 15657
rect 2746 15660 3341 15688
rect 2038 15552 2044 15564
rect 1688 15524 2044 15552
rect 1688 15493 1716 15524
rect 2038 15512 2044 15524
rect 2096 15512 2102 15564
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 1949 15487 2007 15493
rect 1949 15453 1961 15487
rect 1995 15484 2007 15487
rect 2498 15484 2504 15496
rect 1995 15456 2504 15484
rect 1995 15453 2007 15456
rect 1949 15447 2007 15453
rect 2498 15444 2504 15456
rect 2556 15444 2562 15496
rect 2593 15487 2651 15493
rect 2593 15453 2605 15487
rect 2639 15484 2651 15487
rect 2746 15484 2774 15660
rect 3329 15657 3341 15660
rect 3375 15688 3387 15691
rect 5258 15688 5264 15700
rect 3375 15660 5264 15688
rect 3375 15657 3387 15660
rect 3329 15651 3387 15657
rect 5258 15648 5264 15660
rect 5316 15648 5322 15700
rect 7282 15648 7288 15700
rect 7340 15688 7346 15700
rect 7561 15691 7619 15697
rect 7561 15688 7573 15691
rect 7340 15660 7573 15688
rect 7340 15648 7346 15660
rect 7561 15657 7573 15660
rect 7607 15688 7619 15691
rect 9674 15688 9680 15700
rect 7607 15660 9680 15688
rect 7607 15657 7619 15660
rect 7561 15651 7619 15657
rect 9674 15648 9680 15660
rect 9732 15648 9738 15700
rect 10318 15688 10324 15700
rect 10279 15660 10324 15688
rect 10318 15648 10324 15660
rect 10376 15648 10382 15700
rect 12802 15688 12808 15700
rect 11440 15660 12664 15688
rect 12763 15660 12808 15688
rect 8662 15580 8668 15632
rect 8720 15620 8726 15632
rect 11440 15620 11468 15660
rect 8720 15592 11468 15620
rect 12636 15620 12664 15660
rect 12802 15648 12808 15660
rect 12860 15648 12866 15700
rect 17678 15688 17684 15700
rect 15600 15660 17684 15688
rect 15600 15620 15628 15660
rect 17678 15648 17684 15660
rect 17736 15688 17742 15700
rect 18785 15691 18843 15697
rect 18785 15688 18797 15691
rect 17736 15660 18797 15688
rect 17736 15648 17742 15660
rect 18785 15657 18797 15660
rect 18831 15688 18843 15691
rect 19889 15691 19947 15697
rect 18831 15660 19334 15688
rect 18831 15657 18843 15660
rect 18785 15651 18843 15657
rect 12636 15592 15628 15620
rect 16945 15623 17003 15629
rect 8720 15580 8726 15592
rect 16945 15589 16957 15623
rect 16991 15620 17003 15623
rect 18322 15620 18328 15632
rect 16991 15592 18328 15620
rect 16991 15589 17003 15592
rect 16945 15583 17003 15589
rect 18322 15580 18328 15592
rect 18380 15580 18386 15632
rect 18414 15580 18420 15632
rect 18472 15620 18478 15632
rect 18472 15592 18517 15620
rect 18472 15580 18478 15592
rect 11054 15552 11060 15564
rect 9140 15524 11060 15552
rect 2639 15456 2774 15484
rect 3789 15487 3847 15493
rect 2639 15453 2651 15456
rect 2593 15447 2651 15453
rect 3789 15453 3801 15487
rect 3835 15484 3847 15487
rect 4338 15484 4344 15496
rect 3835 15456 4344 15484
rect 3835 15453 3847 15456
rect 3789 15447 3847 15453
rect 4338 15444 4344 15456
rect 4396 15444 4402 15496
rect 7190 15484 7196 15496
rect 6932 15456 7196 15484
rect 6932 15428 6960 15456
rect 7190 15444 7196 15456
rect 7248 15484 7254 15496
rect 7285 15487 7343 15493
rect 7285 15484 7297 15487
rect 7248 15456 7297 15484
rect 7248 15444 7254 15456
rect 7285 15453 7297 15456
rect 7331 15453 7343 15487
rect 7926 15484 7932 15496
rect 7887 15456 7932 15484
rect 7285 15447 7343 15453
rect 7926 15444 7932 15456
rect 7984 15444 7990 15496
rect 4034 15419 4092 15425
rect 4034 15416 4046 15419
rect 2608 15388 4046 15416
rect 2608 15360 2636 15388
rect 4034 15385 4046 15388
rect 4080 15385 4092 15419
rect 4034 15379 4092 15385
rect 5537 15419 5595 15425
rect 5537 15385 5549 15419
rect 5583 15416 5595 15419
rect 5583 15388 6868 15416
rect 5583 15385 5595 15388
rect 5537 15379 5595 15385
rect 1486 15348 1492 15360
rect 1447 15320 1492 15348
rect 1486 15308 1492 15320
rect 1544 15308 1550 15360
rect 2130 15348 2136 15360
rect 2091 15320 2136 15348
rect 2130 15308 2136 15320
rect 2188 15308 2194 15360
rect 2590 15308 2596 15360
rect 2648 15308 2654 15360
rect 2961 15351 3019 15357
rect 2961 15317 2973 15351
rect 3007 15348 3019 15351
rect 3142 15348 3148 15360
rect 3007 15320 3148 15348
rect 3007 15317 3019 15320
rect 2961 15311 3019 15317
rect 3142 15308 3148 15320
rect 3200 15308 3206 15360
rect 5166 15348 5172 15360
rect 5127 15320 5172 15348
rect 5166 15308 5172 15320
rect 5224 15308 5230 15360
rect 5902 15348 5908 15360
rect 5863 15320 5908 15348
rect 5902 15308 5908 15320
rect 5960 15308 5966 15360
rect 6840 15348 6868 15388
rect 6914 15376 6920 15428
rect 6972 15376 6978 15428
rect 7006 15376 7012 15428
rect 7064 15425 7070 15428
rect 7064 15416 7076 15425
rect 9140 15416 9168 15524
rect 11054 15512 11060 15524
rect 11112 15512 11118 15564
rect 14182 15552 14188 15564
rect 14143 15524 14188 15552
rect 14182 15512 14188 15524
rect 14240 15512 14246 15564
rect 14550 15512 14556 15564
rect 14608 15552 14614 15564
rect 15105 15555 15163 15561
rect 15105 15552 15117 15555
rect 14608 15524 15117 15552
rect 14608 15512 14614 15524
rect 15105 15521 15117 15524
rect 15151 15521 15163 15555
rect 15105 15515 15163 15521
rect 19150 15512 19156 15564
rect 19208 15552 19214 15564
rect 19306 15552 19334 15660
rect 19889 15657 19901 15691
rect 19935 15688 19947 15691
rect 20714 15688 20720 15700
rect 19935 15660 20720 15688
rect 19935 15657 19947 15660
rect 19889 15651 19947 15657
rect 20714 15648 20720 15660
rect 20772 15648 20778 15700
rect 19208 15524 19748 15552
rect 19208 15512 19214 15524
rect 9582 15444 9588 15496
rect 9640 15484 9646 15496
rect 9677 15487 9735 15493
rect 9677 15484 9689 15487
rect 9640 15456 9689 15484
rect 9640 15444 9646 15456
rect 9677 15453 9689 15456
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 10962 15444 10968 15496
rect 11020 15484 11026 15496
rect 11425 15487 11483 15493
rect 11425 15484 11437 15487
rect 11020 15456 11437 15484
rect 11020 15444 11026 15456
rect 11425 15453 11437 15456
rect 11471 15453 11483 15487
rect 11425 15447 11483 15453
rect 11692 15487 11750 15493
rect 11692 15453 11704 15487
rect 11738 15484 11750 15487
rect 12066 15484 12072 15496
rect 11738 15456 12072 15484
rect 11738 15453 11750 15456
rect 11692 15447 11750 15453
rect 12066 15444 12072 15456
rect 12124 15444 12130 15496
rect 14458 15484 14464 15496
rect 14419 15456 14464 15484
rect 14458 15444 14464 15456
rect 14516 15444 14522 15496
rect 15565 15487 15623 15493
rect 15565 15453 15577 15487
rect 15611 15484 15623 15487
rect 17494 15484 17500 15496
rect 15611 15456 17500 15484
rect 15611 15453 15623 15456
rect 15565 15447 15623 15453
rect 17494 15444 17500 15456
rect 17552 15444 17558 15496
rect 17954 15444 17960 15496
rect 18012 15484 18018 15496
rect 18049 15487 18107 15493
rect 18049 15484 18061 15487
rect 18012 15456 18061 15484
rect 18012 15444 18018 15456
rect 18049 15453 18061 15456
rect 18095 15484 18107 15487
rect 19058 15484 19064 15496
rect 18095 15456 19064 15484
rect 18095 15453 18107 15456
rect 18049 15447 18107 15453
rect 19058 15444 19064 15456
rect 19116 15444 19122 15496
rect 19720 15493 19748 15524
rect 19705 15487 19763 15493
rect 19705 15453 19717 15487
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20622 15484 20628 15496
rect 20583 15456 20628 15484
rect 20165 15447 20223 15453
rect 9306 15416 9312 15428
rect 7064 15388 7109 15416
rect 8404 15388 9168 15416
rect 9267 15388 9312 15416
rect 7064 15379 7076 15388
rect 7064 15376 7070 15379
rect 8404 15348 8432 15388
rect 9306 15376 9312 15388
rect 9364 15376 9370 15428
rect 15654 15416 15660 15428
rect 14844 15388 15660 15416
rect 8570 15348 8576 15360
rect 6840 15320 8432 15348
rect 8531 15320 8576 15348
rect 8570 15308 8576 15320
rect 8628 15308 8634 15360
rect 8662 15308 8668 15360
rect 8720 15348 8726 15360
rect 8941 15351 8999 15357
rect 8941 15348 8953 15351
rect 8720 15320 8953 15348
rect 8720 15308 8726 15320
rect 8941 15317 8953 15320
rect 8987 15317 8999 15351
rect 10594 15348 10600 15360
rect 10555 15320 10600 15348
rect 8941 15311 8999 15317
rect 10594 15308 10600 15320
rect 10652 15308 10658 15360
rect 13354 15308 13360 15360
rect 13412 15348 13418 15360
rect 14844 15357 14872 15388
rect 15654 15376 15660 15388
rect 15712 15376 15718 15428
rect 15832 15419 15890 15425
rect 15832 15385 15844 15419
rect 15878 15416 15890 15419
rect 17034 15416 17040 15428
rect 15878 15388 17040 15416
rect 15878 15385 15890 15388
rect 15832 15379 15890 15385
rect 17034 15376 17040 15388
rect 17092 15376 17098 15428
rect 17405 15419 17463 15425
rect 17405 15385 17417 15419
rect 17451 15416 17463 15419
rect 18138 15416 18144 15428
rect 17451 15388 18144 15416
rect 17451 15385 17463 15388
rect 17405 15379 17463 15385
rect 18138 15376 18144 15388
rect 18196 15376 18202 15428
rect 18414 15376 18420 15428
rect 18472 15416 18478 15428
rect 20180 15416 20208 15447
rect 20622 15444 20628 15456
rect 20680 15444 20686 15496
rect 21082 15484 21088 15496
rect 21043 15456 21088 15484
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 18472 15388 20208 15416
rect 18472 15376 18478 15388
rect 14369 15351 14427 15357
rect 14369 15348 14381 15351
rect 13412 15320 14381 15348
rect 13412 15308 13418 15320
rect 14369 15317 14381 15320
rect 14415 15317 14427 15351
rect 14369 15311 14427 15317
rect 14829 15351 14887 15357
rect 14829 15317 14841 15351
rect 14875 15317 14887 15351
rect 14829 15311 14887 15317
rect 15010 15308 15016 15360
rect 15068 15348 15074 15360
rect 17681 15351 17739 15357
rect 17681 15348 17693 15351
rect 15068 15320 17693 15348
rect 15068 15308 15074 15320
rect 17681 15317 17693 15320
rect 17727 15317 17739 15351
rect 19426 15348 19432 15360
rect 19387 15320 19432 15348
rect 17681 15311 17739 15317
rect 19426 15308 19432 15320
rect 19484 15308 19490 15360
rect 20349 15351 20407 15357
rect 20349 15317 20361 15351
rect 20395 15348 20407 15351
rect 20714 15348 20720 15360
rect 20395 15320 20720 15348
rect 20395 15317 20407 15320
rect 20349 15311 20407 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 20809 15351 20867 15357
rect 20809 15317 20821 15351
rect 20855 15348 20867 15351
rect 21082 15348 21088 15360
rect 20855 15320 21088 15348
rect 20855 15317 20867 15320
rect 20809 15311 20867 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 5718 15104 5724 15156
rect 5776 15144 5782 15156
rect 5813 15147 5871 15153
rect 5813 15144 5825 15147
rect 5776 15116 5825 15144
rect 5776 15104 5782 15116
rect 5813 15113 5825 15116
rect 5859 15113 5871 15147
rect 5813 15107 5871 15113
rect 9309 15147 9367 15153
rect 9309 15113 9321 15147
rect 9355 15144 9367 15147
rect 9490 15144 9496 15156
rect 9355 15116 9496 15144
rect 9355 15113 9367 15116
rect 9309 15107 9367 15113
rect 9490 15104 9496 15116
rect 9548 15104 9554 15156
rect 13357 15147 13415 15153
rect 13357 15113 13369 15147
rect 13403 15144 13415 15147
rect 15013 15147 15071 15153
rect 13403 15116 13860 15144
rect 13403 15113 13415 15116
rect 13357 15107 13415 15113
rect 3142 15036 3148 15088
rect 3200 15076 3206 15088
rect 8196 15079 8254 15085
rect 3200 15048 7420 15076
rect 3200 15036 3206 15048
rect 1673 15011 1731 15017
rect 1673 14977 1685 15011
rect 1719 15008 1731 15011
rect 1946 15008 1952 15020
rect 1719 14980 1952 15008
rect 1719 14977 1731 14980
rect 1673 14971 1731 14977
rect 1946 14968 1952 14980
rect 2004 14968 2010 15020
rect 2130 15008 2136 15020
rect 2091 14980 2136 15008
rect 2130 14968 2136 14980
rect 2188 14968 2194 15020
rect 3717 15011 3775 15017
rect 3717 14977 3729 15011
rect 3763 15008 3775 15011
rect 4062 15008 4068 15020
rect 3763 14980 4068 15008
rect 3763 14977 3775 14980
rect 3717 14971 3775 14977
rect 4062 14968 4068 14980
rect 4120 14968 4126 15020
rect 4246 14968 4252 15020
rect 4304 15008 4310 15020
rect 5166 15008 5172 15020
rect 4304 14980 5172 15008
rect 4304 14968 4310 14980
rect 5166 14968 5172 14980
rect 5224 14968 5230 15020
rect 5994 14968 6000 15020
rect 6052 15008 6058 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 6052 14980 6745 15008
rect 6052 14968 6058 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 7282 15008 7288 15020
rect 6871 14980 7288 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 7282 14968 7288 14980
rect 7340 14968 7346 15020
rect 7392 15008 7420 15048
rect 8196 15045 8208 15079
rect 8242 15076 8254 15079
rect 8570 15076 8576 15088
rect 8242 15048 8576 15076
rect 8242 15045 8254 15048
rect 8196 15039 8254 15045
rect 8570 15036 8576 15048
rect 8628 15036 8634 15088
rect 13832 15076 13860 15116
rect 15013 15113 15025 15147
rect 15059 15144 15071 15147
rect 15194 15144 15200 15156
rect 15059 15116 15200 15144
rect 15059 15113 15071 15116
rect 15013 15107 15071 15113
rect 15194 15104 15200 15116
rect 15252 15104 15258 15156
rect 15654 15144 15660 15156
rect 15615 15116 15660 15144
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 18046 15144 18052 15156
rect 16071 15116 17908 15144
rect 18007 15116 18052 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 13900 15079 13958 15085
rect 13900 15076 13912 15079
rect 11992 15048 13584 15076
rect 13832 15048 13912 15076
rect 9214 15008 9220 15020
rect 7392 14980 9220 15008
rect 9214 14968 9220 14980
rect 9272 14968 9278 15020
rect 10686 14968 10692 15020
rect 10744 15017 10750 15020
rect 11992 15017 12020 15048
rect 10744 15008 10756 15017
rect 11977 15011 12035 15017
rect 10744 14980 10789 15008
rect 10744 14971 10756 14980
rect 11977 14977 11989 15011
rect 12023 14977 12035 15011
rect 11977 14971 12035 14977
rect 12244 15011 12302 15017
rect 12244 14977 12256 15011
rect 12290 15008 12302 15011
rect 12802 15008 12808 15020
rect 12290 14980 12808 15008
rect 12290 14977 12302 14980
rect 12244 14971 12302 14977
rect 10744 14968 10750 14971
rect 12802 14968 12808 14980
rect 12860 14968 12866 15020
rect 13556 15008 13584 15048
rect 13900 15045 13912 15048
rect 13946 15076 13958 15079
rect 14182 15076 14188 15088
rect 13946 15048 14188 15076
rect 13946 15045 13958 15048
rect 13900 15039 13958 15045
rect 14182 15036 14188 15048
rect 14240 15076 14246 15088
rect 14366 15076 14372 15088
rect 14240 15048 14372 15076
rect 14240 15036 14246 15048
rect 14366 15036 14372 15048
rect 14424 15036 14430 15088
rect 17494 15076 17500 15088
rect 16684 15048 17500 15076
rect 13630 15008 13636 15020
rect 13556 14980 13636 15008
rect 13630 14968 13636 14980
rect 13688 15008 13694 15020
rect 13688 14980 13733 15008
rect 13688 14968 13694 14980
rect 16574 14968 16580 15020
rect 16632 15008 16638 15020
rect 16684 15017 16712 15048
rect 17494 15036 17500 15048
rect 17552 15036 17558 15088
rect 17880 15076 17908 15116
rect 18046 15104 18052 15116
rect 18104 15104 18110 15156
rect 19426 15104 19432 15156
rect 19484 15144 19490 15156
rect 19705 15147 19763 15153
rect 19705 15144 19717 15147
rect 19484 15116 19717 15144
rect 19484 15104 19490 15116
rect 19705 15113 19717 15116
rect 19751 15113 19763 15147
rect 19705 15107 19763 15113
rect 20533 15147 20591 15153
rect 20533 15113 20545 15147
rect 20579 15144 20591 15147
rect 20622 15144 20628 15156
rect 20579 15116 20628 15144
rect 20579 15113 20591 15116
rect 20533 15107 20591 15113
rect 20622 15104 20628 15116
rect 20680 15104 20686 15156
rect 18230 15076 18236 15088
rect 17880 15048 18236 15076
rect 18230 15036 18236 15048
rect 18288 15036 18294 15088
rect 16942 15017 16948 15020
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 16632 14980 16681 15008
rect 16632 14968 16638 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 16669 14971 16727 14977
rect 16936 14971 16948 15017
rect 17000 15008 17006 15020
rect 18693 15011 18751 15017
rect 17000 14980 17036 15008
rect 16942 14968 16948 14971
rect 17000 14968 17006 14980
rect 18693 14977 18705 15011
rect 18739 15008 18751 15011
rect 18782 15008 18788 15020
rect 18739 14980 18788 15008
rect 18739 14977 18751 14980
rect 18693 14971 18751 14977
rect 18782 14968 18788 14980
rect 18840 14968 18846 15020
rect 19702 15008 19708 15020
rect 18984 14980 19708 15008
rect 3973 14943 4031 14949
rect 3973 14909 3985 14943
rect 4019 14940 4031 14943
rect 4338 14940 4344 14952
rect 4019 14912 4344 14940
rect 4019 14909 4031 14912
rect 3973 14903 4031 14909
rect 4338 14900 4344 14912
rect 4396 14900 4402 14952
rect 4798 14900 4804 14952
rect 4856 14940 4862 14952
rect 7009 14943 7067 14949
rect 4856 14912 6408 14940
rect 4856 14900 4862 14912
rect 4249 14875 4307 14881
rect 4249 14841 4261 14875
rect 4295 14872 4307 14875
rect 5350 14872 5356 14884
rect 4295 14844 5356 14872
rect 4295 14841 4307 14844
rect 4249 14835 4307 14841
rect 5350 14832 5356 14844
rect 5408 14832 5414 14884
rect 6380 14881 6408 14912
rect 7009 14909 7021 14943
rect 7055 14940 7067 14943
rect 7834 14940 7840 14952
rect 7055 14912 7840 14940
rect 7055 14909 7067 14912
rect 7009 14903 7067 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 7929 14943 7987 14949
rect 7929 14909 7941 14943
rect 7975 14909 7987 14943
rect 7929 14903 7987 14909
rect 6365 14875 6423 14881
rect 6365 14841 6377 14875
rect 6411 14841 6423 14875
rect 6365 14835 6423 14841
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 1670 14764 1676 14816
rect 1728 14804 1734 14816
rect 1949 14807 2007 14813
rect 1949 14804 1961 14807
rect 1728 14776 1961 14804
rect 1728 14764 1734 14776
rect 1949 14773 1961 14776
rect 1995 14773 2007 14807
rect 2590 14804 2596 14816
rect 2551 14776 2596 14804
rect 1949 14767 2007 14773
rect 2590 14764 2596 14776
rect 2648 14764 2654 14816
rect 4522 14764 4528 14816
rect 4580 14804 4586 14816
rect 4617 14807 4675 14813
rect 4617 14804 4629 14807
rect 4580 14776 4629 14804
rect 4580 14764 4586 14776
rect 4617 14773 4629 14776
rect 4663 14773 4675 14807
rect 4617 14767 4675 14773
rect 7469 14807 7527 14813
rect 7469 14773 7481 14807
rect 7515 14804 7527 14807
rect 7558 14804 7564 14816
rect 7515 14776 7564 14804
rect 7515 14773 7527 14776
rect 7469 14767 7527 14773
rect 7558 14764 7564 14776
rect 7616 14764 7622 14816
rect 7944 14804 7972 14903
rect 10962 14900 10968 14952
rect 11020 14940 11026 14952
rect 11020 14912 11113 14940
rect 11020 14900 11026 14912
rect 15194 14900 15200 14952
rect 15252 14940 15258 14952
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 15252 14912 15393 14940
rect 15252 14900 15258 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15562 14940 15568 14952
rect 15523 14912 15568 14940
rect 15381 14903 15439 14909
rect 15562 14900 15568 14912
rect 15620 14900 15626 14952
rect 18506 14940 18512 14952
rect 18467 14912 18512 14940
rect 18506 14900 18512 14912
rect 18564 14900 18570 14952
rect 18601 14943 18659 14949
rect 18601 14909 18613 14943
rect 18647 14940 18659 14943
rect 18874 14940 18880 14952
rect 18647 14912 18880 14940
rect 18647 14909 18659 14912
rect 18601 14903 18659 14909
rect 18874 14900 18880 14912
rect 18932 14900 18938 14952
rect 9140 14844 10088 14872
rect 9140 14816 9168 14844
rect 9122 14804 9128 14816
rect 7944 14776 9128 14804
rect 9122 14764 9128 14776
rect 9180 14764 9186 14816
rect 9582 14804 9588 14816
rect 9543 14776 9588 14804
rect 9582 14764 9588 14776
rect 9640 14764 9646 14816
rect 10060 14804 10088 14844
rect 10980 14804 11008 14900
rect 18984 14872 19012 14980
rect 19702 14968 19708 14980
rect 19760 14968 19766 15020
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 19518 14900 19524 14952
rect 19576 14940 19582 14952
rect 19797 14943 19855 14949
rect 19797 14940 19809 14943
rect 19576 14912 19809 14940
rect 19576 14900 19582 14912
rect 19797 14909 19809 14912
rect 19843 14909 19855 14943
rect 19797 14903 19855 14909
rect 19886 14900 19892 14952
rect 19944 14940 19950 14952
rect 19944 14912 19989 14940
rect 19944 14900 19950 14912
rect 18340 14844 19012 14872
rect 19061 14875 19119 14881
rect 10060 14776 11008 14804
rect 13630 14764 13636 14816
rect 13688 14804 13694 14816
rect 14274 14804 14280 14816
rect 13688 14776 14280 14804
rect 13688 14764 13694 14776
rect 14274 14764 14280 14776
rect 14332 14764 14338 14816
rect 17034 14764 17040 14816
rect 17092 14804 17098 14816
rect 18340 14804 18368 14844
rect 19061 14841 19073 14875
rect 19107 14872 19119 14875
rect 20364 14872 20392 14971
rect 20714 14968 20720 15020
rect 20772 15008 20778 15020
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20772 14980 21097 15008
rect 20772 14968 20778 14980
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 19107 14844 20392 14872
rect 19107 14841 19119 14844
rect 19061 14835 19119 14841
rect 17092 14776 18368 14804
rect 17092 14764 17098 14776
rect 18414 14764 18420 14816
rect 18472 14804 18478 14816
rect 19337 14807 19395 14813
rect 19337 14804 19349 14807
rect 18472 14776 19349 14804
rect 18472 14764 18478 14776
rect 19337 14773 19349 14776
rect 19383 14773 19395 14807
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 19337 14767 19395 14773
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1946 14600 1952 14612
rect 1907 14572 1952 14600
rect 1946 14560 1952 14572
rect 2004 14560 2010 14612
rect 2498 14560 2504 14612
rect 2556 14600 2562 14612
rect 2685 14603 2743 14609
rect 2685 14600 2697 14603
rect 2556 14572 2697 14600
rect 2556 14560 2562 14572
rect 2685 14569 2697 14572
rect 2731 14569 2743 14603
rect 6914 14600 6920 14612
rect 2685 14563 2743 14569
rect 6564 14572 6920 14600
rect 1210 14492 1216 14544
rect 1268 14532 1274 14544
rect 6181 14535 6239 14541
rect 6181 14532 6193 14535
rect 1268 14504 6193 14532
rect 1268 14492 1274 14504
rect 6181 14501 6193 14504
rect 6227 14501 6239 14535
rect 6181 14495 6239 14501
rect 3142 14464 3148 14476
rect 2148 14436 3148 14464
rect 1670 14396 1676 14408
rect 1631 14368 1676 14396
rect 1670 14356 1676 14368
rect 1728 14356 1734 14408
rect 2148 14405 2176 14436
rect 3142 14424 3148 14436
rect 3200 14424 3206 14476
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14464 3387 14467
rect 4246 14464 4252 14476
rect 3375 14436 4252 14464
rect 3375 14433 3387 14436
rect 3329 14427 3387 14433
rect 4246 14424 4252 14436
rect 4304 14424 4310 14476
rect 4341 14467 4399 14473
rect 4341 14433 4353 14467
rect 4387 14433 4399 14467
rect 4341 14427 4399 14433
rect 2133 14399 2191 14405
rect 2133 14365 2145 14399
rect 2179 14365 2191 14399
rect 2133 14359 2191 14365
rect 2590 14356 2596 14408
rect 2648 14396 2654 14408
rect 4356 14396 4384 14427
rect 4430 14424 4436 14476
rect 4488 14464 4494 14476
rect 6564 14473 6592 14572
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 7926 14600 7932 14612
rect 7887 14572 7932 14600
rect 7926 14560 7932 14572
rect 7984 14560 7990 14612
rect 8110 14560 8116 14612
rect 8168 14600 8174 14612
rect 12161 14603 12219 14609
rect 8168 14572 10088 14600
rect 8168 14560 8174 14572
rect 10060 14532 10088 14572
rect 12161 14569 12173 14603
rect 12207 14600 12219 14603
rect 13354 14600 13360 14612
rect 12207 14572 13360 14600
rect 12207 14569 12219 14572
rect 12161 14563 12219 14569
rect 13354 14560 13360 14572
rect 13412 14560 13418 14612
rect 14829 14603 14887 14609
rect 14829 14569 14841 14603
rect 14875 14600 14887 14603
rect 15562 14600 15568 14612
rect 14875 14572 15568 14600
rect 14875 14569 14887 14572
rect 14829 14563 14887 14569
rect 15562 14560 15568 14572
rect 15620 14560 15626 14612
rect 15672 14572 16712 14600
rect 15672 14532 15700 14572
rect 10060 14504 15700 14532
rect 16684 14532 16712 14572
rect 16942 14560 16948 14612
rect 17000 14600 17006 14612
rect 17129 14603 17187 14609
rect 17129 14600 17141 14603
rect 17000 14572 17141 14600
rect 17000 14560 17006 14572
rect 17129 14569 17141 14572
rect 17175 14600 17187 14603
rect 17954 14600 17960 14612
rect 17175 14572 17960 14600
rect 17175 14569 17187 14572
rect 17129 14563 17187 14569
rect 17954 14560 17960 14572
rect 18012 14560 18018 14612
rect 18506 14600 18512 14612
rect 18432 14572 18512 14600
rect 17218 14532 17224 14544
rect 16684 14504 17224 14532
rect 17218 14492 17224 14504
rect 17276 14492 17282 14544
rect 17310 14492 17316 14544
rect 17368 14532 17374 14544
rect 17405 14535 17463 14541
rect 17405 14532 17417 14535
rect 17368 14504 17417 14532
rect 17368 14492 17374 14504
rect 17405 14501 17417 14504
rect 17451 14501 17463 14535
rect 17405 14495 17463 14501
rect 17678 14492 17684 14544
rect 17736 14532 17742 14544
rect 17773 14535 17831 14541
rect 17773 14532 17785 14535
rect 17736 14504 17785 14532
rect 17736 14492 17742 14504
rect 17773 14501 17785 14504
rect 17819 14501 17831 14535
rect 17773 14495 17831 14501
rect 6549 14467 6607 14473
rect 6549 14464 6561 14467
rect 4488 14436 6561 14464
rect 4488 14424 4494 14436
rect 6549 14433 6561 14436
rect 6595 14433 6607 14467
rect 6549 14427 6607 14433
rect 8294 14424 8300 14476
rect 8352 14464 8358 14476
rect 11609 14467 11667 14473
rect 8352 14436 9260 14464
rect 8352 14424 8358 14436
rect 2648 14368 4384 14396
rect 2648 14356 2654 14368
rect 4706 14356 4712 14408
rect 4764 14396 4770 14408
rect 9122 14396 9128 14408
rect 4764 14368 6960 14396
rect 9083 14368 9128 14396
rect 4764 14356 4770 14368
rect 3878 14288 3884 14340
rect 3936 14328 3942 14340
rect 4249 14331 4307 14337
rect 4249 14328 4261 14331
rect 3936 14300 4261 14328
rect 3936 14288 3942 14300
rect 4249 14297 4261 14300
rect 4295 14297 4307 14331
rect 4249 14291 4307 14297
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 6822 14337 6828 14340
rect 5169 14331 5227 14337
rect 5169 14328 5181 14331
rect 4672 14300 5181 14328
rect 4672 14288 4678 14300
rect 5169 14297 5181 14300
rect 5215 14297 5227 14331
rect 6816 14328 6828 14337
rect 6783 14300 6828 14328
rect 5169 14291 5227 14297
rect 6816 14291 6828 14300
rect 6822 14288 6828 14291
rect 6880 14288 6886 14340
rect 6932 14328 6960 14368
rect 9122 14356 9128 14368
rect 9180 14356 9186 14408
rect 9232 14396 9260 14436
rect 11609 14433 11621 14467
rect 11655 14464 11667 14467
rect 12802 14464 12808 14476
rect 11655 14436 12808 14464
rect 11655 14433 11667 14436
rect 11609 14427 11667 14433
rect 12802 14424 12808 14436
rect 12860 14424 12866 14476
rect 14277 14467 14335 14473
rect 14277 14433 14289 14467
rect 14323 14464 14335 14467
rect 14366 14464 14372 14476
rect 14323 14436 14372 14464
rect 14323 14433 14335 14436
rect 14277 14427 14335 14433
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 18432 14473 18460 14572
rect 18506 14560 18512 14572
rect 18564 14560 18570 14612
rect 18874 14600 18880 14612
rect 18835 14572 18880 14600
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 19518 14600 19524 14612
rect 19479 14572 19524 14600
rect 19518 14560 19524 14572
rect 19576 14560 19582 14612
rect 19058 14492 19064 14544
rect 19116 14532 19122 14544
rect 19116 14504 20024 14532
rect 19116 14492 19122 14504
rect 18233 14467 18291 14473
rect 18233 14464 18245 14467
rect 18104 14436 18245 14464
rect 18104 14424 18110 14436
rect 18233 14433 18245 14436
rect 18279 14433 18291 14467
rect 18233 14427 18291 14433
rect 18417 14467 18475 14473
rect 18417 14433 18429 14467
rect 18463 14433 18475 14467
rect 18874 14464 18880 14476
rect 18417 14427 18475 14433
rect 18625 14436 18880 14464
rect 10502 14396 10508 14408
rect 9232 14368 10508 14396
rect 10502 14356 10508 14368
rect 10560 14356 10566 14408
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14396 11207 14399
rect 11790 14396 11796 14408
rect 11195 14368 11796 14396
rect 11195 14365 11207 14368
rect 11149 14359 11207 14365
rect 11790 14356 11796 14368
rect 11848 14396 11854 14408
rect 12066 14396 12072 14408
rect 11848 14368 12072 14396
rect 11848 14356 11854 14368
rect 12066 14356 12072 14368
rect 12124 14356 12130 14408
rect 13725 14399 13783 14405
rect 13725 14365 13737 14399
rect 13771 14396 13783 14399
rect 15654 14396 15660 14408
rect 13771 14368 15660 14396
rect 13771 14365 13783 14368
rect 13725 14359 13783 14365
rect 15654 14356 15660 14368
rect 15712 14356 15718 14408
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 16574 14396 16580 14408
rect 15795 14368 16580 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 16574 14356 16580 14368
rect 16632 14396 16638 14408
rect 16942 14396 16948 14408
rect 16632 14368 16948 14396
rect 16632 14356 16638 14368
rect 16942 14356 16948 14368
rect 17000 14356 17006 14408
rect 9392 14331 9450 14337
rect 6932 14300 8340 14328
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 3050 14260 3056 14272
rect 3011 14232 3056 14260
rect 3050 14220 3056 14232
rect 3108 14220 3114 14272
rect 3145 14263 3203 14269
rect 3145 14229 3157 14263
rect 3191 14260 3203 14263
rect 3789 14263 3847 14269
rect 3789 14260 3801 14263
rect 3191 14232 3801 14260
rect 3191 14229 3203 14232
rect 3145 14223 3203 14229
rect 3789 14229 3801 14232
rect 3835 14229 3847 14263
rect 4154 14260 4160 14272
rect 4115 14232 4160 14260
rect 3789 14223 3847 14229
rect 4154 14220 4160 14232
rect 4212 14220 4218 14272
rect 4798 14260 4804 14272
rect 4759 14232 4804 14260
rect 4798 14220 4804 14232
rect 4856 14220 4862 14272
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 5721 14263 5779 14269
rect 5721 14260 5733 14263
rect 5132 14232 5733 14260
rect 5132 14220 5138 14232
rect 5721 14229 5733 14232
rect 5767 14229 5779 14263
rect 5721 14223 5779 14229
rect 6638 14220 6644 14272
rect 6696 14260 6702 14272
rect 8110 14260 8116 14272
rect 6696 14232 8116 14260
rect 6696 14220 6702 14232
rect 8110 14220 8116 14232
rect 8168 14260 8174 14272
rect 8205 14263 8263 14269
rect 8205 14260 8217 14263
rect 8168 14232 8217 14260
rect 8168 14220 8174 14232
rect 8205 14229 8217 14232
rect 8251 14229 8263 14263
rect 8312 14260 8340 14300
rect 9392 14297 9404 14331
rect 9438 14328 9450 14331
rect 9490 14328 9496 14340
rect 9438 14300 9496 14328
rect 9438 14297 9450 14300
rect 9392 14291 9450 14297
rect 9490 14288 9496 14300
rect 9548 14288 9554 14340
rect 11882 14328 11888 14340
rect 9600 14300 11888 14328
rect 9600 14260 9628 14300
rect 11882 14288 11888 14300
rect 11940 14288 11946 14340
rect 12250 14288 12256 14340
rect 12308 14328 12314 14340
rect 14461 14331 14519 14337
rect 14461 14328 14473 14331
rect 12308 14300 14473 14328
rect 12308 14288 12314 14300
rect 14461 14297 14473 14300
rect 14507 14297 14519 14331
rect 14461 14291 14519 14297
rect 16016 14331 16074 14337
rect 16016 14297 16028 14331
rect 16062 14328 16074 14331
rect 17126 14328 17132 14340
rect 16062 14300 17132 14328
rect 16062 14297 16074 14300
rect 16016 14291 16074 14297
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 18509 14331 18567 14337
rect 18509 14297 18521 14331
rect 18555 14328 18567 14331
rect 18625 14328 18653 14436
rect 18874 14424 18880 14436
rect 18932 14424 18938 14476
rect 19996 14473 20024 14504
rect 19981 14467 20039 14473
rect 19981 14433 19993 14467
rect 20027 14433 20039 14467
rect 19981 14427 20039 14433
rect 20165 14467 20223 14473
rect 20165 14433 20177 14467
rect 20211 14464 20223 14467
rect 20530 14464 20536 14476
rect 20211 14436 20536 14464
rect 20211 14433 20223 14436
rect 20165 14427 20223 14433
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 19334 14396 19340 14408
rect 18748 14368 19340 14396
rect 18748 14356 18754 14368
rect 19334 14356 19340 14368
rect 19392 14356 19398 14408
rect 19610 14356 19616 14408
rect 19668 14396 19674 14408
rect 20625 14399 20683 14405
rect 20625 14396 20637 14399
rect 19668 14368 20637 14396
rect 19668 14356 19674 14368
rect 20625 14365 20637 14368
rect 20671 14365 20683 14399
rect 21082 14396 21088 14408
rect 21043 14368 21088 14396
rect 20625 14359 20683 14365
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 18555 14300 18653 14328
rect 18555 14297 18567 14300
rect 18509 14291 18567 14297
rect 19794 14288 19800 14340
rect 19852 14328 19858 14340
rect 19889 14331 19947 14337
rect 19889 14328 19901 14331
rect 19852 14300 19901 14328
rect 19852 14288 19858 14300
rect 19889 14297 19901 14300
rect 19935 14328 19947 14331
rect 20070 14328 20076 14340
rect 19935 14300 20076 14328
rect 19935 14297 19947 14300
rect 19889 14291 19947 14297
rect 20070 14288 20076 14300
rect 20128 14288 20134 14340
rect 21174 14328 21180 14340
rect 20180 14300 21180 14328
rect 8312 14232 9628 14260
rect 8205 14223 8263 14229
rect 9766 14220 9772 14272
rect 9824 14260 9830 14272
rect 10505 14263 10563 14269
rect 10505 14260 10517 14263
rect 9824 14232 10517 14260
rect 9824 14220 9830 14232
rect 10505 14229 10517 14232
rect 10551 14260 10563 14263
rect 10686 14260 10692 14272
rect 10551 14232 10692 14260
rect 10551 14229 10563 14232
rect 10505 14223 10563 14229
rect 10686 14220 10692 14232
rect 10744 14220 10750 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11701 14263 11759 14269
rect 11701 14260 11713 14263
rect 11296 14232 11713 14260
rect 11296 14220 11302 14232
rect 11701 14229 11713 14232
rect 11747 14229 11759 14263
rect 13354 14260 13360 14272
rect 13315 14232 13360 14260
rect 11701 14223 11759 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 14366 14260 14372 14272
rect 14327 14232 14372 14260
rect 14366 14220 14372 14232
rect 14424 14220 14430 14272
rect 15470 14260 15476 14272
rect 15431 14232 15476 14260
rect 15470 14220 15476 14232
rect 15528 14220 15534 14272
rect 17310 14220 17316 14272
rect 17368 14260 17374 14272
rect 20180 14260 20208 14300
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 17368 14232 20208 14260
rect 20809 14263 20867 14269
rect 17368 14220 17374 14232
rect 20809 14229 20821 14263
rect 20855 14260 20867 14263
rect 21082 14260 21088 14272
rect 20855 14232 21088 14260
rect 20855 14229 20867 14232
rect 20809 14223 20867 14229
rect 21082 14220 21088 14232
rect 21140 14220 21146 14272
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 3050 14016 3056 14068
rect 3108 14056 3114 14068
rect 3145 14059 3203 14065
rect 3145 14056 3157 14059
rect 3108 14028 3157 14056
rect 3108 14016 3114 14028
rect 3145 14025 3157 14028
rect 3191 14025 3203 14059
rect 3145 14019 3203 14025
rect 4709 14059 4767 14065
rect 4709 14025 4721 14059
rect 4755 14056 4767 14059
rect 5994 14056 6000 14068
rect 4755 14028 5396 14056
rect 5955 14028 6000 14056
rect 4755 14025 4767 14028
rect 4709 14019 4767 14025
rect 1670 13920 1676 13932
rect 1631 13892 1676 13920
rect 1670 13880 1676 13892
rect 1728 13880 1734 13932
rect 2774 13880 2780 13932
rect 2832 13920 2838 13932
rect 3605 13923 3663 13929
rect 2832 13892 2877 13920
rect 2832 13880 2838 13892
rect 3605 13889 3617 13923
rect 3651 13920 3663 13923
rect 4617 13923 4675 13929
rect 3651 13892 4384 13920
rect 3651 13889 3663 13892
rect 3605 13883 3663 13889
rect 2130 13852 2136 13864
rect 2091 13824 2136 13852
rect 2130 13812 2136 13824
rect 2188 13812 2194 13864
rect 2590 13852 2596 13864
rect 2551 13824 2596 13852
rect 2590 13812 2596 13824
rect 2648 13812 2654 13864
rect 2685 13855 2743 13861
rect 2685 13821 2697 13855
rect 2731 13852 2743 13855
rect 3050 13852 3056 13864
rect 2731 13824 3056 13852
rect 2731 13821 2743 13824
rect 2685 13815 2743 13821
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 3418 13852 3424 13864
rect 3379 13824 3424 13852
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 1486 13784 1492 13796
rect 1447 13756 1492 13784
rect 1486 13744 1492 13756
rect 1544 13744 1550 13796
rect 4356 13784 4384 13892
rect 4617 13889 4629 13923
rect 4663 13920 4675 13923
rect 4706 13920 4712 13932
rect 4663 13892 4712 13920
rect 4663 13889 4675 13892
rect 4617 13883 4675 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 4801 13855 4859 13861
rect 4801 13821 4813 13855
rect 4847 13821 4859 13855
rect 4801 13815 4859 13821
rect 4816 13784 4844 13815
rect 4356 13756 4844 13784
rect 4724 13728 4752 13756
rect 3142 13676 3148 13728
rect 3200 13716 3206 13728
rect 4062 13716 4068 13728
rect 3200 13688 4068 13716
rect 3200 13676 3206 13688
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4246 13716 4252 13728
rect 4207 13688 4252 13716
rect 4246 13676 4252 13688
rect 4304 13676 4310 13728
rect 4706 13676 4712 13728
rect 4764 13676 4770 13728
rect 4890 13676 4896 13728
rect 4948 13716 4954 13728
rect 5368 13716 5396 14028
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6638 14016 6644 14068
rect 6696 14056 6702 14068
rect 7469 14059 7527 14065
rect 7469 14056 7481 14059
rect 6696 14028 7481 14056
rect 6696 14016 6702 14028
rect 7469 14025 7481 14028
rect 7515 14025 7527 14059
rect 7469 14019 7527 14025
rect 8205 14059 8263 14065
rect 8205 14025 8217 14059
rect 8251 14056 8263 14059
rect 8294 14056 8300 14068
rect 8251 14028 8300 14056
rect 8251 14025 8263 14028
rect 8205 14019 8263 14025
rect 8294 14016 8300 14028
rect 8352 14016 8358 14068
rect 8386 14016 8392 14068
rect 8444 14056 8450 14068
rect 8573 14059 8631 14065
rect 8573 14056 8585 14059
rect 8444 14028 8585 14056
rect 8444 14016 8450 14028
rect 8573 14025 8585 14028
rect 8619 14025 8631 14059
rect 11793 14059 11851 14065
rect 11793 14056 11805 14059
rect 8573 14019 8631 14025
rect 8680 14028 11805 14056
rect 5537 13923 5595 13929
rect 5537 13889 5549 13923
rect 5583 13889 5595 13923
rect 5537 13883 5595 13889
rect 5629 13923 5687 13929
rect 5629 13889 5641 13923
rect 5675 13920 5687 13923
rect 5994 13920 6000 13932
rect 5675 13892 6000 13920
rect 5675 13889 5687 13892
rect 5629 13883 5687 13889
rect 5445 13855 5503 13861
rect 5445 13821 5457 13855
rect 5491 13821 5503 13855
rect 5552 13852 5580 13883
rect 5994 13880 6000 13892
rect 6052 13880 6058 13932
rect 6638 13920 6644 13932
rect 6288 13892 6644 13920
rect 6288 13852 6316 13892
rect 6638 13880 6644 13892
rect 6696 13880 6702 13932
rect 8680 13920 8708 14028
rect 11793 14025 11805 14028
rect 11839 14025 11851 14059
rect 11793 14019 11851 14025
rect 11882 14016 11888 14068
rect 11940 14056 11946 14068
rect 12250 14056 12256 14068
rect 11940 14028 11985 14056
rect 12211 14028 12256 14056
rect 11940 14016 11946 14028
rect 12250 14016 12256 14028
rect 12308 14016 12314 14068
rect 14366 14016 14372 14068
rect 14424 14056 14430 14068
rect 14461 14059 14519 14065
rect 14461 14056 14473 14059
rect 14424 14028 14473 14056
rect 14424 14016 14430 14028
rect 14461 14025 14473 14028
rect 14507 14025 14519 14059
rect 14461 14019 14519 14025
rect 16853 14059 16911 14065
rect 16853 14025 16865 14059
rect 16899 14056 16911 14059
rect 17034 14056 17040 14068
rect 16899 14028 17040 14056
rect 16899 14025 16911 14028
rect 16853 14019 16911 14025
rect 17034 14016 17040 14028
rect 17092 14016 17098 14068
rect 17589 14059 17647 14065
rect 17589 14025 17601 14059
rect 17635 14056 17647 14059
rect 17862 14056 17868 14068
rect 17635 14028 17868 14056
rect 17635 14025 17647 14028
rect 17589 14019 17647 14025
rect 17862 14016 17868 14028
rect 17920 14016 17926 14068
rect 18414 14056 18420 14068
rect 18375 14028 18420 14056
rect 18414 14016 18420 14028
rect 18472 14016 18478 14068
rect 18782 14056 18788 14068
rect 18743 14028 18788 14056
rect 18782 14016 18788 14028
rect 18840 14016 18846 14068
rect 19061 14059 19119 14065
rect 19061 14025 19073 14059
rect 19107 14025 19119 14059
rect 19061 14019 19119 14025
rect 19521 14059 19579 14065
rect 19521 14025 19533 14059
rect 19567 14056 19579 14059
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 19567 14028 20085 14056
rect 19567 14025 19579 14028
rect 19521 14019 19579 14025
rect 20073 14025 20085 14028
rect 20119 14025 20131 14059
rect 20073 14019 20131 14025
rect 11057 13991 11115 13997
rect 11057 13988 11069 13991
rect 6932 13892 8708 13920
rect 8864 13960 11069 13988
rect 6454 13852 6460 13864
rect 5552 13824 6316 13852
rect 6415 13824 6460 13852
rect 5445 13815 5503 13821
rect 5451 13784 5479 13815
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6730 13852 6736 13864
rect 6691 13824 6736 13852
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 5902 13784 5908 13796
rect 5451 13756 5908 13784
rect 5902 13744 5908 13756
rect 5960 13784 5966 13796
rect 6822 13784 6828 13796
rect 5960 13756 6828 13784
rect 5960 13744 5966 13756
rect 6822 13744 6828 13756
rect 6880 13744 6886 13796
rect 6932 13716 6960 13892
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13821 7251 13855
rect 7193 13815 7251 13821
rect 7377 13855 7435 13861
rect 7377 13821 7389 13855
rect 7423 13852 7435 13855
rect 7650 13852 7656 13864
rect 7423 13824 7656 13852
rect 7423 13821 7435 13824
rect 7377 13815 7435 13821
rect 7098 13744 7104 13796
rect 7156 13784 7162 13796
rect 7208 13784 7236 13815
rect 7650 13812 7656 13824
rect 7708 13852 7714 13864
rect 8294 13852 8300 13864
rect 7708 13824 8300 13852
rect 7708 13812 7714 13824
rect 8294 13812 8300 13824
rect 8352 13812 8358 13864
rect 7156 13756 7236 13784
rect 7156 13744 7162 13756
rect 8110 13744 8116 13796
rect 8168 13784 8174 13796
rect 8864 13784 8892 13960
rect 11057 13957 11069 13960
rect 11103 13988 11115 13991
rect 11238 13988 11244 14000
rect 11103 13960 11244 13988
rect 11103 13957 11115 13960
rect 11057 13951 11115 13957
rect 11238 13948 11244 13960
rect 11296 13948 11302 14000
rect 14918 13988 14924 14000
rect 11716 13960 12434 13988
rect 14879 13960 14924 13988
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9950 13920 9956 13932
rect 8996 13892 9041 13920
rect 9911 13892 9956 13920
rect 8996 13880 9002 13892
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 10042 13880 10048 13932
rect 10100 13920 10106 13932
rect 10597 13923 10655 13929
rect 10597 13920 10609 13923
rect 10100 13892 10609 13920
rect 10100 13880 10106 13892
rect 10597 13889 10609 13892
rect 10643 13920 10655 13923
rect 10643 13892 11652 13920
rect 10643 13889 10655 13892
rect 10597 13883 10655 13889
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9125 13855 9183 13861
rect 9125 13821 9137 13855
rect 9171 13852 9183 13855
rect 9582 13852 9588 13864
rect 9171 13824 9588 13852
rect 9171 13821 9183 13824
rect 9125 13815 9183 13821
rect 8168 13756 8892 13784
rect 9048 13784 9076 13815
rect 9582 13812 9588 13824
rect 9640 13812 9646 13864
rect 10137 13855 10195 13861
rect 10137 13821 10149 13855
rect 10183 13821 10195 13855
rect 10137 13815 10195 13821
rect 9214 13784 9220 13796
rect 9048 13756 9220 13784
rect 8168 13744 8174 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9490 13744 9496 13796
rect 9548 13784 9554 13796
rect 10152 13784 10180 13815
rect 9548 13756 10180 13784
rect 11624 13784 11652 13892
rect 11716 13861 11744 13960
rect 12406 13920 12434 13960
rect 14918 13948 14924 13960
rect 14976 13948 14982 14000
rect 17221 13991 17279 13997
rect 15304 13960 17080 13988
rect 12802 13920 12808 13932
rect 12406 13892 12808 13920
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13920 14243 13923
rect 14458 13920 14464 13932
rect 14231 13892 14464 13920
rect 14231 13889 14243 13892
rect 14185 13883 14243 13889
rect 14458 13880 14464 13892
rect 14516 13880 14522 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13920 14887 13923
rect 15304 13920 15332 13960
rect 14875 13892 15332 13920
rect 14875 13889 14887 13892
rect 14829 13883 14887 13889
rect 15378 13880 15384 13932
rect 15436 13920 15442 13932
rect 16298 13920 16304 13932
rect 15436 13892 16304 13920
rect 15436 13880 15442 13892
rect 16298 13880 16304 13892
rect 16356 13880 16362 13932
rect 17052 13920 17080 13960
rect 17221 13957 17233 13991
rect 17267 13988 17279 13991
rect 17267 13960 18460 13988
rect 17267 13957 17279 13960
rect 17221 13951 17279 13957
rect 18432 13920 18460 13960
rect 18506 13948 18512 14000
rect 18564 13988 18570 14000
rect 19076 13988 19104 14019
rect 20346 14016 20352 14068
rect 20404 14056 20410 14068
rect 20533 14059 20591 14065
rect 20533 14056 20545 14059
rect 20404 14028 20545 14056
rect 20404 14016 20410 14028
rect 20533 14025 20545 14028
rect 20579 14025 20591 14059
rect 21266 14056 21272 14068
rect 21227 14028 21272 14056
rect 20533 14019 20591 14025
rect 21266 14016 21272 14028
rect 21324 14016 21330 14068
rect 18564 13960 19104 13988
rect 18564 13948 18570 13960
rect 19334 13948 19340 14000
rect 19392 13988 19398 14000
rect 20438 13988 20444 14000
rect 19392 13960 20444 13988
rect 19392 13948 19398 13960
rect 20438 13948 20444 13960
rect 20496 13948 20502 14000
rect 18690 13920 18696 13932
rect 17052 13892 17172 13920
rect 18432 13892 18696 13920
rect 11701 13855 11759 13861
rect 11701 13821 11713 13855
rect 11747 13821 11759 13855
rect 12526 13852 12532 13864
rect 11701 13815 11759 13821
rect 11808 13824 12434 13852
rect 12487 13824 12532 13852
rect 11808 13784 11836 13824
rect 11624 13756 11836 13784
rect 12406 13796 12434 13824
rect 12526 13812 12532 13824
rect 12584 13812 12590 13864
rect 12406 13756 12440 13796
rect 9548 13744 9554 13756
rect 12434 13744 12440 13756
rect 12492 13744 12498 13796
rect 12820 13784 12848 13880
rect 13078 13852 13084 13864
rect 13039 13824 13084 13852
rect 13078 13812 13084 13824
rect 13136 13812 13142 13864
rect 13449 13855 13507 13861
rect 13449 13821 13461 13855
rect 13495 13852 13507 13855
rect 13538 13852 13544 13864
rect 13495 13824 13544 13852
rect 13495 13821 13507 13824
rect 13449 13815 13507 13821
rect 13538 13812 13544 13824
rect 13596 13812 13602 13864
rect 13817 13855 13875 13861
rect 13817 13821 13829 13855
rect 13863 13852 13875 13855
rect 14734 13852 14740 13864
rect 13863 13824 14740 13852
rect 13863 13821 13875 13824
rect 13817 13815 13875 13821
rect 14734 13812 14740 13824
rect 14792 13812 14798 13864
rect 15013 13855 15071 13861
rect 15013 13821 15025 13855
rect 15059 13821 15071 13855
rect 15013 13815 15071 13821
rect 16025 13855 16083 13861
rect 16025 13821 16037 13855
rect 16071 13852 16083 13855
rect 17144 13852 17172 13892
rect 18690 13880 18696 13892
rect 18748 13880 18754 13932
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13920 19487 13923
rect 19518 13920 19524 13932
rect 19475 13892 19524 13920
rect 19475 13889 19487 13892
rect 19429 13883 19487 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 21082 13920 21088 13932
rect 21043 13892 21088 13920
rect 21082 13880 21088 13892
rect 21140 13880 21146 13932
rect 17494 13852 17500 13864
rect 16071 13824 17080 13852
rect 17144 13824 17500 13852
rect 16071 13821 16083 13824
rect 16025 13815 16083 13821
rect 15028 13784 15056 13815
rect 12820 13756 15056 13784
rect 17052 13784 17080 13824
rect 17494 13812 17500 13824
rect 17552 13812 17558 13864
rect 18046 13812 18052 13864
rect 18104 13852 18110 13864
rect 18141 13855 18199 13861
rect 18141 13852 18153 13855
rect 18104 13824 18153 13852
rect 18104 13812 18110 13824
rect 18141 13821 18153 13824
rect 18187 13821 18199 13855
rect 18322 13852 18328 13864
rect 18283 13824 18328 13852
rect 18141 13815 18199 13821
rect 18322 13812 18328 13824
rect 18380 13812 18386 13864
rect 19613 13855 19671 13861
rect 19613 13821 19625 13855
rect 19659 13821 19671 13855
rect 19613 13815 19671 13821
rect 17126 13784 17132 13796
rect 17052 13756 17132 13784
rect 17126 13744 17132 13756
rect 17184 13744 17190 13796
rect 17954 13744 17960 13796
rect 18012 13784 18018 13796
rect 19628 13784 19656 13815
rect 20622 13812 20628 13864
rect 20680 13852 20686 13864
rect 20680 13824 20725 13852
rect 20680 13812 20686 13824
rect 19794 13784 19800 13796
rect 18012 13756 19800 13784
rect 18012 13744 18018 13756
rect 19794 13744 19800 13756
rect 19852 13744 19858 13796
rect 4948 13688 6960 13716
rect 4948 13676 4954 13688
rect 7742 13676 7748 13728
rect 7800 13716 7806 13728
rect 7837 13719 7895 13725
rect 7837 13716 7849 13719
rect 7800 13688 7849 13716
rect 7800 13676 7806 13688
rect 7837 13685 7849 13688
rect 7883 13685 7895 13719
rect 9582 13716 9588 13728
rect 9543 13688 9588 13716
rect 7837 13679 7895 13685
rect 9582 13676 9588 13688
rect 9640 13676 9646 13728
rect 12710 13676 12716 13728
rect 12768 13716 12774 13728
rect 17310 13716 17316 13728
rect 12768 13688 17316 13716
rect 12768 13676 12774 13688
rect 17310 13676 17316 13688
rect 17368 13676 17374 13728
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2774 13472 2780 13524
rect 2832 13512 2838 13524
rect 3053 13515 3111 13521
rect 3053 13512 3065 13515
rect 2832 13484 3065 13512
rect 2832 13472 2838 13484
rect 3053 13481 3065 13484
rect 3099 13481 3111 13515
rect 3053 13475 3111 13481
rect 3418 13472 3424 13524
rect 3476 13472 3482 13524
rect 3789 13515 3847 13521
rect 3789 13481 3801 13515
rect 3835 13512 3847 13515
rect 3878 13512 3884 13524
rect 3835 13484 3884 13512
rect 3835 13481 3847 13484
rect 3789 13475 3847 13481
rect 3878 13472 3884 13484
rect 3936 13472 3942 13524
rect 4062 13472 4068 13524
rect 4120 13512 4126 13524
rect 4985 13515 5043 13521
rect 4120 13484 4384 13512
rect 4120 13472 4126 13484
rect 2222 13404 2228 13456
rect 2280 13444 2286 13456
rect 2406 13444 2412 13456
rect 2280 13416 2412 13444
rect 2280 13404 2286 13416
rect 2406 13404 2412 13416
rect 2464 13404 2470 13456
rect 2038 13336 2044 13388
rect 2096 13376 2102 13388
rect 2501 13379 2559 13385
rect 2501 13376 2513 13379
rect 2096 13348 2513 13376
rect 2096 13336 2102 13348
rect 2501 13345 2513 13348
rect 2547 13376 2559 13379
rect 3142 13376 3148 13388
rect 2547 13348 3148 13376
rect 2547 13345 2559 13348
rect 2501 13339 2559 13345
rect 3142 13336 3148 13348
rect 3200 13336 3206 13388
rect 3436 13320 3464 13472
rect 4246 13444 4252 13456
rect 4172 13416 4252 13444
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13277 1731 13311
rect 1673 13271 1731 13277
rect 1688 13240 1716 13271
rect 2130 13268 2136 13320
rect 2188 13308 2194 13320
rect 2685 13311 2743 13317
rect 2685 13308 2697 13311
rect 2188 13280 2697 13308
rect 2188 13268 2194 13280
rect 2685 13277 2697 13280
rect 2731 13277 2743 13311
rect 2685 13271 2743 13277
rect 3418 13268 3424 13320
rect 3476 13268 3482 13320
rect 4172 13317 4200 13416
rect 4246 13404 4252 13416
rect 4304 13404 4310 13456
rect 4356 13385 4384 13484
rect 4985 13481 4997 13515
rect 5031 13512 5043 13515
rect 5258 13512 5264 13524
rect 5031 13484 5264 13512
rect 5031 13481 5043 13484
rect 4985 13475 5043 13481
rect 5258 13472 5264 13484
rect 5316 13472 5322 13524
rect 7282 13512 7288 13524
rect 7243 13484 7288 13512
rect 7282 13472 7288 13484
rect 7340 13472 7346 13524
rect 9214 13512 9220 13524
rect 9175 13484 9220 13512
rect 9214 13472 9220 13484
rect 9272 13472 9278 13524
rect 9950 13472 9956 13524
rect 10008 13512 10014 13524
rect 10413 13515 10471 13521
rect 10413 13512 10425 13515
rect 10008 13484 10425 13512
rect 10008 13472 10014 13484
rect 10413 13481 10425 13484
rect 10459 13481 10471 13515
rect 10413 13475 10471 13481
rect 12342 13472 12348 13524
rect 12400 13512 12406 13524
rect 12894 13512 12900 13524
rect 12400 13484 12900 13512
rect 12400 13472 12406 13484
rect 12894 13472 12900 13484
rect 12952 13472 12958 13524
rect 16942 13512 16948 13524
rect 16903 13484 16948 13512
rect 16942 13472 16948 13484
rect 17000 13472 17006 13524
rect 17862 13472 17868 13524
rect 17920 13472 17926 13524
rect 18322 13472 18328 13524
rect 18380 13512 18386 13524
rect 18417 13515 18475 13521
rect 18417 13512 18429 13515
rect 18380 13484 18429 13512
rect 18380 13472 18386 13484
rect 18417 13481 18429 13484
rect 18463 13481 18475 13515
rect 21634 13512 21640 13524
rect 18417 13475 18475 13481
rect 18524 13484 21640 13512
rect 6822 13404 6828 13456
rect 6880 13444 6886 13456
rect 17880 13444 17908 13472
rect 18524 13444 18552 13484
rect 21634 13472 21640 13484
rect 21692 13472 21698 13524
rect 6880 13416 7880 13444
rect 6880 13404 6886 13416
rect 4341 13379 4399 13385
rect 4341 13345 4353 13379
rect 4387 13345 4399 13379
rect 7742 13376 7748 13388
rect 7703 13348 7748 13376
rect 4341 13339 4399 13345
rect 7742 13336 7748 13348
rect 7800 13336 7806 13388
rect 7852 13385 7880 13416
rect 17779 13416 18552 13444
rect 18877 13447 18935 13453
rect 7837 13379 7895 13385
rect 7837 13345 7849 13379
rect 7883 13345 7895 13379
rect 7837 13339 7895 13345
rect 9582 13336 9588 13388
rect 9640 13376 9646 13388
rect 9677 13379 9735 13385
rect 9677 13376 9689 13379
rect 9640 13348 9689 13376
rect 9640 13336 9646 13348
rect 9677 13345 9689 13348
rect 9723 13345 9735 13379
rect 9677 13339 9735 13345
rect 9766 13336 9772 13388
rect 9824 13376 9830 13388
rect 12250 13376 12256 13388
rect 9824 13348 9869 13376
rect 12211 13348 12256 13376
rect 9824 13336 9830 13348
rect 12250 13336 12256 13348
rect 12308 13336 12314 13388
rect 13078 13336 13084 13388
rect 13136 13376 13142 13388
rect 13136 13348 15608 13376
rect 13136 13336 13142 13348
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13277 4215 13311
rect 7009 13311 7067 13317
rect 4157 13271 4215 13277
rect 4264 13280 6960 13308
rect 2222 13240 2228 13252
rect 1688 13212 2228 13240
rect 2222 13200 2228 13212
rect 2280 13200 2286 13252
rect 4264 13240 4292 13280
rect 2424 13212 4292 13240
rect 1486 13172 1492 13184
rect 1447 13144 1492 13172
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 1854 13132 1860 13184
rect 1912 13172 1918 13184
rect 1949 13175 2007 13181
rect 1949 13172 1961 13175
rect 1912 13144 1961 13172
rect 1912 13132 1918 13144
rect 1949 13141 1961 13144
rect 1995 13172 2007 13175
rect 2424 13172 2452 13212
rect 4338 13200 4344 13252
rect 4396 13240 4402 13252
rect 5261 13243 5319 13249
rect 5261 13240 5273 13243
rect 4396 13212 5273 13240
rect 4396 13200 4402 13212
rect 5261 13209 5273 13212
rect 5307 13209 5319 13243
rect 6932 13240 6960 13280
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 8294 13308 8300 13320
rect 7055 13280 8300 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 8294 13268 8300 13280
rect 8352 13268 8358 13320
rect 11241 13311 11299 13317
rect 11241 13277 11253 13311
rect 11287 13308 11299 13311
rect 11882 13308 11888 13320
rect 11287 13280 11888 13308
rect 11287 13277 11299 13280
rect 11241 13271 11299 13277
rect 11882 13268 11888 13280
rect 11940 13268 11946 13320
rect 12986 13268 12992 13320
rect 13044 13308 13050 13320
rect 13354 13308 13360 13320
rect 13044 13280 13360 13308
rect 13044 13268 13050 13280
rect 13354 13268 13360 13280
rect 13412 13268 13418 13320
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14093 13311 14151 13317
rect 14093 13308 14105 13311
rect 13872 13280 14105 13308
rect 13872 13268 13878 13280
rect 14093 13277 14105 13280
rect 14139 13277 14151 13311
rect 14093 13271 14151 13277
rect 15580 13252 15608 13348
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17779 13376 17807 13416
rect 18877 13413 18889 13447
rect 18923 13444 18935 13447
rect 18923 13416 20392 13444
rect 18923 13413 18935 13416
rect 18877 13407 18935 13413
rect 17000 13348 17807 13376
rect 17865 13379 17923 13385
rect 17000 13336 17006 13348
rect 17865 13345 17877 13379
rect 17911 13376 17923 13379
rect 17954 13376 17960 13388
rect 17911 13348 17960 13376
rect 17911 13345 17923 13348
rect 17865 13339 17923 13345
rect 17954 13336 17960 13348
rect 18012 13336 18018 13388
rect 19794 13376 19800 13388
rect 19755 13348 19800 13376
rect 19794 13336 19800 13348
rect 19852 13336 19858 13388
rect 20364 13376 20392 13416
rect 20438 13404 20444 13456
rect 20496 13444 20502 13456
rect 20533 13447 20591 13453
rect 20533 13444 20545 13447
rect 20496 13416 20545 13444
rect 20496 13404 20502 13416
rect 20533 13413 20545 13416
rect 20579 13444 20591 13447
rect 20622 13444 20628 13456
rect 20579 13416 20628 13444
rect 20579 13413 20591 13416
rect 20533 13407 20591 13413
rect 20622 13404 20628 13416
rect 20680 13404 20686 13456
rect 20898 13376 20904 13388
rect 20364 13348 20904 13376
rect 20898 13336 20904 13348
rect 20956 13336 20962 13388
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 18322 13308 18328 13320
rect 17460 13280 18328 13308
rect 17460 13268 17466 13280
rect 18322 13268 18328 13280
rect 18380 13268 18386 13320
rect 18690 13308 18696 13320
rect 18651 13280 18696 13308
rect 18690 13268 18696 13280
rect 18748 13268 18754 13320
rect 20990 13268 20996 13320
rect 21048 13308 21054 13320
rect 21085 13311 21143 13317
rect 21085 13308 21097 13311
rect 21048 13280 21097 13308
rect 21048 13268 21054 13280
rect 21085 13277 21097 13280
rect 21131 13277 21143 13311
rect 21085 13271 21143 13277
rect 7190 13240 7196 13252
rect 6932 13212 7196 13240
rect 5261 13203 5319 13209
rect 7190 13200 7196 13212
rect 7248 13240 7254 13252
rect 7466 13240 7472 13252
rect 7248 13212 7472 13240
rect 7248 13200 7254 13212
rect 7466 13200 7472 13212
rect 7524 13200 7530 13252
rect 9858 13200 9864 13252
rect 9916 13240 9922 13252
rect 15013 13243 15071 13249
rect 15013 13240 15025 13243
rect 9916 13212 15025 13240
rect 9916 13200 9922 13212
rect 15013 13209 15025 13212
rect 15059 13240 15071 13243
rect 15194 13240 15200 13252
rect 15059 13212 15200 13240
rect 15059 13209 15071 13212
rect 15013 13203 15071 13209
rect 15194 13200 15200 13212
rect 15252 13200 15258 13252
rect 15562 13200 15568 13252
rect 15620 13240 15626 13252
rect 15657 13243 15715 13249
rect 15657 13240 15669 13243
rect 15620 13212 15669 13240
rect 15620 13200 15626 13212
rect 15657 13209 15669 13212
rect 15703 13209 15715 13243
rect 15657 13203 15715 13209
rect 15930 13200 15936 13252
rect 15988 13240 15994 13252
rect 18049 13243 18107 13249
rect 18049 13240 18061 13243
rect 15988 13212 18061 13240
rect 15988 13200 15994 13212
rect 18049 13209 18061 13212
rect 18095 13209 18107 13243
rect 18049 13203 18107 13209
rect 19613 13243 19671 13249
rect 19613 13209 19625 13243
rect 19659 13240 19671 13243
rect 20254 13240 20260 13252
rect 19659 13212 20260 13240
rect 19659 13209 19671 13212
rect 19613 13203 19671 13209
rect 20254 13200 20260 13212
rect 20312 13200 20318 13252
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 20404 13212 20449 13240
rect 20404 13200 20410 13212
rect 2590 13172 2596 13184
rect 1995 13144 2452 13172
rect 2551 13144 2596 13172
rect 1995 13141 2007 13144
rect 1949 13135 2007 13141
rect 2590 13132 2596 13144
rect 2648 13132 2654 13184
rect 3326 13172 3332 13184
rect 3287 13144 3332 13172
rect 3326 13132 3332 13144
rect 3384 13132 3390 13184
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4304 13144 4349 13172
rect 4304 13132 4310 13144
rect 7282 13132 7288 13184
rect 7340 13172 7346 13184
rect 7653 13175 7711 13181
rect 7653 13172 7665 13175
rect 7340 13144 7665 13172
rect 7340 13132 7346 13144
rect 7653 13141 7665 13144
rect 7699 13141 7711 13175
rect 7653 13135 7711 13141
rect 7742 13132 7748 13184
rect 7800 13172 7806 13184
rect 8297 13175 8355 13181
rect 8297 13172 8309 13175
rect 7800 13144 8309 13172
rect 7800 13132 7806 13144
rect 8297 13141 8309 13144
rect 8343 13141 8355 13175
rect 8297 13135 8355 13141
rect 9585 13175 9643 13181
rect 9585 13141 9597 13175
rect 9631 13172 9643 13175
rect 10042 13172 10048 13184
rect 9631 13144 10048 13172
rect 9631 13141 9643 13144
rect 9585 13135 9643 13141
rect 10042 13132 10048 13144
rect 10100 13132 10106 13184
rect 10778 13172 10784 13184
rect 10739 13144 10784 13172
rect 10778 13132 10784 13144
rect 10836 13132 10842 13184
rect 11238 13132 11244 13184
rect 11296 13172 11302 13184
rect 11517 13175 11575 13181
rect 11517 13172 11529 13175
rect 11296 13144 11529 13172
rect 11296 13132 11302 13144
rect 11517 13141 11529 13144
rect 11563 13141 11575 13175
rect 11517 13135 11575 13141
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 11885 13175 11943 13181
rect 11885 13172 11897 13175
rect 11756 13144 11897 13172
rect 11756 13132 11762 13144
rect 11885 13141 11897 13144
rect 11931 13141 11943 13175
rect 12710 13172 12716 13184
rect 12671 13144 12716 13172
rect 11885 13135 11943 13141
rect 12710 13132 12716 13144
rect 12768 13132 12774 13184
rect 13262 13172 13268 13184
rect 13223 13144 13268 13172
rect 13262 13132 13268 13144
rect 13320 13132 13326 13184
rect 13354 13132 13360 13184
rect 13412 13172 13418 13184
rect 13633 13175 13691 13181
rect 13633 13172 13645 13175
rect 13412 13144 13645 13172
rect 13412 13132 13418 13144
rect 13633 13141 13645 13144
rect 13679 13141 13691 13175
rect 13633 13135 13691 13141
rect 14737 13175 14795 13181
rect 14737 13141 14749 13175
rect 14783 13172 14795 13175
rect 14918 13172 14924 13184
rect 14783 13144 14924 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 14918 13132 14924 13144
rect 14976 13132 14982 13184
rect 17402 13132 17408 13184
rect 17460 13172 17466 13184
rect 17957 13175 18015 13181
rect 17957 13172 17969 13175
rect 17460 13144 17969 13172
rect 17460 13132 17466 13144
rect 17957 13141 17969 13144
rect 18003 13141 18015 13175
rect 17957 13135 18015 13141
rect 18874 13132 18880 13184
rect 18932 13172 18938 13184
rect 19245 13175 19303 13181
rect 19245 13172 19257 13175
rect 18932 13144 19257 13172
rect 18932 13132 18938 13144
rect 19245 13141 19257 13144
rect 19291 13141 19303 13175
rect 19245 13135 19303 13141
rect 19702 13132 19708 13184
rect 19760 13172 19766 13184
rect 21266 13172 21272 13184
rect 19760 13144 19805 13172
rect 21227 13144 21272 13172
rect 19760 13132 19766 13144
rect 21266 13132 21272 13144
rect 21324 13132 21330 13184
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 2498 12968 2504 12980
rect 2459 12940 2504 12968
rect 2498 12928 2504 12940
rect 2556 12928 2562 12980
rect 2590 12928 2596 12980
rect 2648 12968 2654 12980
rect 2869 12971 2927 12977
rect 2869 12968 2881 12971
rect 2648 12940 2881 12968
rect 2648 12928 2654 12940
rect 2869 12937 2881 12940
rect 2915 12937 2927 12971
rect 2869 12931 2927 12937
rect 3881 12971 3939 12977
rect 3881 12937 3893 12971
rect 3927 12968 3939 12971
rect 4062 12968 4068 12980
rect 3927 12940 4068 12968
rect 3927 12937 3939 12940
rect 3881 12931 3939 12937
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 4157 12971 4215 12977
rect 4157 12937 4169 12971
rect 4203 12968 4215 12971
rect 4246 12968 4252 12980
rect 4203 12940 4252 12968
rect 4203 12937 4215 12940
rect 4157 12931 4215 12937
rect 4246 12928 4252 12940
rect 4304 12928 4310 12980
rect 4430 12928 4436 12980
rect 4488 12968 4494 12980
rect 4617 12971 4675 12977
rect 4617 12968 4629 12971
rect 4488 12940 4629 12968
rect 4488 12928 4494 12940
rect 4617 12937 4629 12940
rect 4663 12968 4675 12971
rect 5258 12968 5264 12980
rect 4663 12940 5264 12968
rect 4663 12937 4675 12940
rect 4617 12931 4675 12937
rect 5258 12928 5264 12940
rect 5316 12928 5322 12980
rect 5994 12928 6000 12980
rect 6052 12968 6058 12980
rect 6365 12971 6423 12977
rect 6365 12968 6377 12971
rect 6052 12940 6377 12968
rect 6052 12928 6058 12940
rect 6365 12937 6377 12940
rect 6411 12937 6423 12971
rect 6365 12931 6423 12937
rect 6733 12971 6791 12977
rect 6733 12937 6745 12971
rect 6779 12968 6791 12971
rect 7742 12968 7748 12980
rect 6779 12940 7748 12968
rect 6779 12937 6791 12940
rect 6733 12931 6791 12937
rect 7742 12928 7748 12940
rect 7800 12928 7806 12980
rect 10042 12968 10048 12980
rect 10003 12940 10048 12968
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10410 12968 10416 12980
rect 10371 12940 10416 12968
rect 10410 12928 10416 12940
rect 10468 12928 10474 12980
rect 10502 12928 10508 12980
rect 10560 12968 10566 12980
rect 11054 12968 11060 12980
rect 10560 12940 10605 12968
rect 11015 12940 11060 12968
rect 10560 12928 10566 12940
rect 11054 12928 11060 12940
rect 11112 12968 11118 12980
rect 11977 12971 12035 12977
rect 11977 12968 11989 12971
rect 11112 12940 11989 12968
rect 11112 12928 11118 12940
rect 11977 12937 11989 12940
rect 12023 12937 12035 12971
rect 15930 12968 15936 12980
rect 15891 12940 15936 12968
rect 11977 12931 12035 12937
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 16942 12968 16948 12980
rect 16903 12940 16948 12968
rect 16942 12928 16948 12940
rect 17000 12928 17006 12980
rect 17034 12928 17040 12980
rect 17092 12968 17098 12980
rect 17402 12968 17408 12980
rect 17092 12940 17264 12968
rect 17363 12940 17408 12968
rect 17092 12928 17098 12940
rect 3326 12900 3332 12912
rect 1688 12872 3332 12900
rect 1578 12792 1584 12844
rect 1636 12832 1642 12844
rect 1688 12841 1716 12872
rect 3326 12860 3332 12872
rect 3384 12860 3390 12912
rect 4522 12900 4528 12912
rect 4483 12872 4528 12900
rect 4522 12860 4528 12872
rect 4580 12860 4586 12912
rect 7374 12900 7380 12912
rect 7335 12872 7380 12900
rect 7374 12860 7380 12872
rect 7432 12860 7438 12912
rect 7837 12903 7895 12909
rect 7837 12869 7849 12903
rect 7883 12900 7895 12903
rect 8294 12900 8300 12912
rect 7883 12872 8300 12900
rect 7883 12869 7895 12872
rect 7837 12863 7895 12869
rect 8294 12860 8300 12872
rect 8352 12900 8358 12912
rect 12989 12903 13047 12909
rect 12989 12900 13001 12903
rect 8352 12872 13001 12900
rect 8352 12860 8358 12872
rect 12989 12869 13001 12872
rect 13035 12900 13047 12903
rect 13078 12900 13084 12912
rect 13035 12872 13084 12900
rect 13035 12869 13047 12872
rect 12989 12863 13047 12869
rect 13078 12860 13084 12872
rect 13136 12860 13142 12912
rect 15470 12900 15476 12912
rect 15431 12872 15476 12900
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 1673 12835 1731 12841
rect 1673 12832 1685 12835
rect 1636 12804 1685 12832
rect 1636 12792 1642 12804
rect 1673 12801 1685 12804
rect 1719 12801 1731 12835
rect 1673 12795 1731 12801
rect 1854 12792 1860 12844
rect 1912 12832 1918 12844
rect 2409 12835 2467 12841
rect 2409 12832 2421 12835
rect 1912 12804 2421 12832
rect 1912 12792 1918 12804
rect 2409 12801 2421 12804
rect 2455 12801 2467 12835
rect 2409 12795 2467 12801
rect 3513 12835 3571 12841
rect 3513 12801 3525 12835
rect 3559 12832 3571 12835
rect 4062 12832 4068 12844
rect 3559 12804 4068 12832
rect 3559 12801 3571 12804
rect 3513 12795 3571 12801
rect 4062 12792 4068 12804
rect 4120 12792 4126 12844
rect 7926 12792 7932 12844
rect 7984 12832 7990 12844
rect 12342 12832 12348 12844
rect 7984 12804 12348 12832
rect 7984 12792 7990 12804
rect 12342 12792 12348 12804
rect 12400 12792 12406 12844
rect 15194 12792 15200 12844
rect 15252 12832 15258 12844
rect 15565 12835 15623 12841
rect 15565 12832 15577 12835
rect 15252 12804 15577 12832
rect 15252 12792 15258 12804
rect 15565 12801 15577 12804
rect 15611 12801 15623 12835
rect 17037 12835 17095 12841
rect 17037 12832 17049 12835
rect 15565 12795 15623 12801
rect 16224 12804 17049 12832
rect 2314 12764 2320 12776
rect 2275 12736 2320 12764
rect 2314 12724 2320 12736
rect 2372 12724 2378 12776
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3237 12767 3295 12773
rect 3237 12764 3249 12767
rect 3200 12736 3249 12764
rect 3200 12724 3206 12736
rect 3237 12733 3249 12736
rect 3283 12733 3295 12767
rect 3237 12727 3295 12733
rect 3421 12767 3479 12773
rect 3421 12733 3433 12767
rect 3467 12764 3479 12767
rect 4430 12764 4436 12776
rect 3467 12736 4436 12764
rect 3467 12733 3479 12736
rect 3421 12727 3479 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 4801 12767 4859 12773
rect 4801 12733 4813 12767
rect 4847 12764 4859 12767
rect 5258 12764 5264 12776
rect 4847 12736 5264 12764
rect 4847 12733 4859 12736
rect 4801 12727 4859 12733
rect 5258 12724 5264 12736
rect 5316 12764 5322 12776
rect 5721 12767 5779 12773
rect 5721 12764 5733 12767
rect 5316 12736 5733 12764
rect 5316 12724 5322 12736
rect 5721 12733 5733 12736
rect 5767 12733 5779 12767
rect 5994 12764 6000 12776
rect 5955 12736 6000 12764
rect 5721 12727 5779 12733
rect 5994 12724 6000 12736
rect 6052 12724 6058 12776
rect 6822 12764 6828 12776
rect 6783 12736 6828 12764
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 7009 12767 7067 12773
rect 7009 12733 7021 12767
rect 7055 12764 7067 12767
rect 7098 12764 7104 12776
rect 7055 12736 7104 12764
rect 7055 12733 7067 12736
rect 7009 12727 7067 12733
rect 7098 12724 7104 12736
rect 7156 12724 7162 12776
rect 7650 12724 7656 12776
rect 7708 12764 7714 12776
rect 7708 12736 8524 12764
rect 7708 12724 7714 12736
rect 1857 12699 1915 12705
rect 1857 12665 1869 12699
rect 1903 12696 1915 12699
rect 8386 12696 8392 12708
rect 1903 12668 8392 12696
rect 1903 12665 1915 12668
rect 1857 12659 1915 12665
rect 8386 12656 8392 12668
rect 8444 12656 8450 12708
rect 8496 12696 8524 12736
rect 9214 12724 9220 12776
rect 9272 12764 9278 12776
rect 9490 12764 9496 12776
rect 9272 12736 9496 12764
rect 9272 12724 9278 12736
rect 9490 12724 9496 12736
rect 9548 12764 9554 12776
rect 10597 12767 10655 12773
rect 10597 12764 10609 12767
rect 9548 12736 10609 12764
rect 9548 12724 9554 12736
rect 10597 12733 10609 12736
rect 10643 12733 10655 12767
rect 11790 12764 11796 12776
rect 11751 12736 11796 12764
rect 10597 12727 10655 12733
rect 11790 12724 11796 12736
rect 11848 12724 11854 12776
rect 11885 12767 11943 12773
rect 11885 12733 11897 12767
rect 11931 12733 11943 12767
rect 15378 12764 15384 12776
rect 15339 12736 15384 12764
rect 11885 12727 11943 12733
rect 9398 12696 9404 12708
rect 8496 12668 9404 12696
rect 9398 12656 9404 12668
rect 9456 12656 9462 12708
rect 10134 12656 10140 12708
rect 10192 12696 10198 12708
rect 11900 12696 11928 12727
rect 15378 12724 15384 12736
rect 15436 12724 15442 12776
rect 10192 12668 11928 12696
rect 10192 12656 10198 12668
rect 11974 12656 11980 12708
rect 12032 12696 12038 12708
rect 12032 12668 14412 12696
rect 12032 12656 12038 12668
rect 1946 12588 1952 12640
rect 2004 12628 2010 12640
rect 5902 12628 5908 12640
rect 2004 12600 5908 12628
rect 2004 12588 2010 12600
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 8478 12588 8484 12640
rect 8536 12628 8542 12640
rect 9122 12628 9128 12640
rect 8536 12600 9128 12628
rect 8536 12588 8542 12600
rect 9122 12588 9128 12600
rect 9180 12588 9186 12640
rect 12345 12631 12403 12637
rect 12345 12597 12357 12631
rect 12391 12628 12403 12631
rect 12526 12628 12532 12640
rect 12391 12600 12532 12628
rect 12391 12597 12403 12600
rect 12345 12591 12403 12597
rect 12526 12588 12532 12600
rect 12584 12588 12590 12640
rect 12713 12631 12771 12637
rect 12713 12597 12725 12631
rect 12759 12628 12771 12631
rect 13630 12628 13636 12640
rect 12759 12600 13636 12628
rect 12759 12597 12771 12600
rect 12713 12591 12771 12597
rect 13630 12588 13636 12600
rect 13688 12588 13694 12640
rect 14274 12628 14280 12640
rect 14235 12600 14280 12628
rect 14274 12588 14280 12600
rect 14332 12588 14338 12640
rect 14384 12628 14412 12668
rect 16224 12637 16252 12804
rect 17037 12801 17049 12804
rect 17083 12801 17095 12835
rect 17236 12832 17264 12940
rect 17402 12928 17408 12940
rect 17460 12928 17466 12980
rect 17494 12928 17500 12980
rect 17552 12968 17558 12980
rect 18141 12971 18199 12977
rect 18141 12968 18153 12971
rect 17552 12940 18153 12968
rect 17552 12928 17558 12940
rect 18141 12937 18153 12940
rect 18187 12968 18199 12971
rect 19334 12968 19340 12980
rect 18187 12940 19340 12968
rect 18187 12937 18199 12940
rect 18141 12931 18199 12937
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 19429 12971 19487 12977
rect 19429 12937 19441 12971
rect 19475 12968 19487 12971
rect 19702 12968 19708 12980
rect 19475 12940 19708 12968
rect 19475 12937 19487 12940
rect 19429 12931 19487 12937
rect 19702 12928 19708 12940
rect 19760 12928 19766 12980
rect 20254 12928 20260 12980
rect 20312 12968 20318 12980
rect 20441 12971 20499 12977
rect 20441 12968 20453 12971
rect 20312 12940 20453 12968
rect 20312 12928 20318 12940
rect 20441 12937 20453 12940
rect 20487 12937 20499 12971
rect 20441 12931 20499 12937
rect 18049 12903 18107 12909
rect 18049 12869 18061 12903
rect 18095 12900 18107 12903
rect 20806 12900 20812 12912
rect 18095 12872 20812 12900
rect 18095 12869 18107 12872
rect 18049 12863 18107 12869
rect 20806 12860 20812 12872
rect 20864 12860 20870 12912
rect 20901 12903 20959 12909
rect 20901 12869 20913 12903
rect 20947 12900 20959 12903
rect 20990 12900 20996 12912
rect 20947 12872 20996 12900
rect 20947 12869 20959 12872
rect 20901 12863 20959 12869
rect 20990 12860 20996 12872
rect 21048 12860 21054 12912
rect 17862 12832 17868 12844
rect 17236 12804 17868 12832
rect 17037 12795 17095 12801
rect 17862 12792 17868 12804
rect 17920 12792 17926 12844
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 16853 12767 16911 12773
rect 16853 12733 16865 12767
rect 16899 12764 16911 12767
rect 17126 12764 17132 12776
rect 16899 12736 17132 12764
rect 16899 12733 16911 12736
rect 16853 12727 16911 12733
rect 17126 12724 17132 12736
rect 17184 12764 17190 12776
rect 17770 12764 17776 12776
rect 17184 12736 17776 12764
rect 17184 12724 17190 12736
rect 17770 12724 17776 12736
rect 17828 12724 17834 12776
rect 18230 12724 18236 12776
rect 18288 12764 18294 12776
rect 18288 12736 18333 12764
rect 18288 12724 18294 12736
rect 16390 12656 16396 12708
rect 16448 12696 16454 12708
rect 18984 12696 19012 12795
rect 19334 12792 19340 12844
rect 19392 12832 19398 12844
rect 19797 12835 19855 12841
rect 19797 12832 19809 12835
rect 19392 12804 19809 12832
rect 19392 12792 19398 12804
rect 19797 12801 19809 12804
rect 19843 12832 19855 12835
rect 20254 12832 20260 12844
rect 19843 12804 20260 12832
rect 19843 12801 19855 12804
rect 19797 12795 19855 12801
rect 20254 12792 20260 12804
rect 20312 12792 20318 12844
rect 19886 12764 19892 12776
rect 19847 12736 19892 12764
rect 19886 12724 19892 12736
rect 19944 12724 19950 12776
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 20346 12764 20352 12776
rect 20119 12736 20352 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 16448 12668 19012 12696
rect 19153 12699 19211 12705
rect 16448 12656 16454 12668
rect 19153 12665 19165 12699
rect 19199 12696 19211 12699
rect 19610 12696 19616 12708
rect 19199 12668 19616 12696
rect 19199 12665 19211 12668
rect 19153 12659 19211 12665
rect 19610 12656 19616 12668
rect 19668 12656 19674 12708
rect 16209 12631 16267 12637
rect 16209 12628 16221 12631
rect 14384 12600 16221 12628
rect 16209 12597 16221 12600
rect 16255 12597 16267 12631
rect 16209 12591 16267 12597
rect 17310 12588 17316 12640
rect 17368 12628 17374 12640
rect 17681 12631 17739 12637
rect 17681 12628 17693 12631
rect 17368 12600 17693 12628
rect 17368 12588 17374 12600
rect 17681 12597 17693 12600
rect 17727 12597 17739 12631
rect 17681 12591 17739 12597
rect 17770 12588 17776 12640
rect 17828 12628 17834 12640
rect 20088 12628 20116 12727
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 20438 12724 20444 12776
rect 20496 12764 20502 12776
rect 20993 12767 21051 12773
rect 20993 12764 21005 12767
rect 20496 12736 21005 12764
rect 20496 12724 20502 12736
rect 20993 12733 21005 12736
rect 21039 12733 21051 12767
rect 20993 12727 21051 12733
rect 17828 12600 20116 12628
rect 17828 12588 17834 12600
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 4430 12384 4436 12436
rect 4488 12424 4494 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 4488 12396 4721 12424
rect 4488 12384 4494 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 7009 12427 7067 12433
rect 7009 12424 7021 12427
rect 5224 12396 7021 12424
rect 5224 12384 5230 12396
rect 7009 12393 7021 12396
rect 7055 12424 7067 12427
rect 7282 12424 7288 12436
rect 7055 12396 7288 12424
rect 7055 12393 7067 12396
rect 7009 12387 7067 12393
rect 7282 12384 7288 12396
rect 7340 12384 7346 12436
rect 7377 12427 7435 12433
rect 7377 12393 7389 12427
rect 7423 12424 7435 12427
rect 8573 12427 8631 12433
rect 7423 12396 7503 12424
rect 7423 12393 7435 12396
rect 7377 12387 7435 12393
rect 4062 12316 4068 12368
rect 4120 12356 4126 12368
rect 5721 12359 5779 12365
rect 5721 12356 5733 12359
rect 4120 12328 5733 12356
rect 4120 12316 4126 12328
rect 5721 12325 5733 12328
rect 5767 12325 5779 12359
rect 5721 12319 5779 12325
rect 5902 12316 5908 12368
rect 5960 12356 5966 12368
rect 6638 12356 6644 12368
rect 5960 12328 6644 12356
rect 5960 12316 5966 12328
rect 6638 12316 6644 12328
rect 6696 12316 6702 12368
rect 4706 12248 4712 12300
rect 4764 12288 4770 12300
rect 5258 12288 5264 12300
rect 4764 12260 5264 12288
rect 4764 12248 4770 12260
rect 5258 12248 5264 12260
rect 5316 12248 5322 12300
rect 5626 12248 5632 12300
rect 5684 12288 5690 12300
rect 5994 12288 6000 12300
rect 5684 12260 6000 12288
rect 5684 12248 5690 12260
rect 5994 12248 6000 12260
rect 6052 12288 6058 12300
rect 6273 12291 6331 12297
rect 6273 12288 6285 12291
rect 6052 12260 6285 12288
rect 6052 12248 6058 12260
rect 6273 12257 6285 12260
rect 6319 12257 6331 12291
rect 6273 12251 6331 12257
rect 7190 12248 7196 12300
rect 7248 12288 7254 12300
rect 7475 12288 7503 12396
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 12342 12424 12348 12436
rect 8619 12396 12348 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 12342 12384 12348 12396
rect 12400 12384 12406 12436
rect 13078 12384 13084 12436
rect 13136 12424 13142 12436
rect 13725 12427 13783 12433
rect 13725 12424 13737 12427
rect 13136 12396 13737 12424
rect 13136 12384 13142 12396
rect 13725 12393 13737 12396
rect 13771 12424 13783 12427
rect 13814 12424 13820 12436
rect 13771 12396 13820 12424
rect 13771 12393 13783 12396
rect 13725 12387 13783 12393
rect 13814 12384 13820 12396
rect 13872 12384 13878 12436
rect 16209 12427 16267 12433
rect 16209 12393 16221 12427
rect 16255 12424 16267 12427
rect 16298 12424 16304 12436
rect 16255 12396 16304 12424
rect 16255 12393 16267 12396
rect 16209 12387 16267 12393
rect 16298 12384 16304 12396
rect 16356 12384 16362 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17678 12424 17684 12436
rect 17000 12396 17684 12424
rect 17000 12384 17006 12396
rect 17678 12384 17684 12396
rect 17736 12424 17742 12436
rect 20990 12424 20996 12436
rect 17736 12396 20996 12424
rect 17736 12384 17742 12396
rect 20990 12384 20996 12396
rect 21048 12384 21054 12436
rect 7742 12316 7748 12368
rect 7800 12316 7806 12368
rect 8846 12316 8852 12368
rect 8904 12356 8910 12368
rect 8904 12328 9168 12356
rect 8904 12316 8910 12328
rect 7248 12260 7503 12288
rect 7248 12248 7254 12260
rect 3421 12223 3479 12229
rect 1596 12192 3280 12220
rect 1596 12164 1624 12192
rect 1578 12152 1584 12164
rect 1539 12124 1584 12152
rect 1578 12112 1584 12124
rect 1636 12112 1642 12164
rect 1762 12152 1768 12164
rect 1723 12124 1768 12152
rect 1762 12112 1768 12124
rect 1820 12112 1826 12164
rect 2314 12112 2320 12164
rect 2372 12152 2378 12164
rect 3154 12155 3212 12161
rect 3154 12152 3166 12155
rect 2372 12124 3166 12152
rect 2372 12112 2378 12124
rect 3154 12121 3166 12124
rect 3200 12121 3212 12155
rect 3252 12152 3280 12192
rect 3421 12189 3433 12223
rect 3467 12220 3479 12223
rect 4338 12220 4344 12232
rect 3467 12192 4344 12220
rect 3467 12189 3479 12192
rect 3421 12183 3479 12189
rect 4338 12180 4344 12192
rect 4396 12180 4402 12232
rect 5718 12180 5724 12232
rect 5776 12220 5782 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5776 12192 6101 12220
rect 5776 12180 5782 12192
rect 6089 12189 6101 12192
rect 6135 12220 6147 12223
rect 7650 12220 7656 12232
rect 6135 12192 7656 12220
rect 6135 12189 6147 12192
rect 6089 12183 6147 12189
rect 7650 12180 7656 12192
rect 7708 12180 7714 12232
rect 7760 12229 7788 12316
rect 9140 12297 9168 12328
rect 9214 12316 9220 12368
rect 9272 12356 9278 12368
rect 9272 12328 10272 12356
rect 9272 12316 9278 12328
rect 7929 12291 7987 12297
rect 7929 12257 7941 12291
rect 7975 12257 7987 12291
rect 7929 12251 7987 12257
rect 9125 12291 9183 12297
rect 9125 12257 9137 12291
rect 9171 12257 9183 12291
rect 9125 12251 9183 12257
rect 7745 12223 7803 12229
rect 7745 12189 7757 12223
rect 7791 12189 7803 12223
rect 7745 12183 7803 12189
rect 7834 12180 7840 12232
rect 7892 12220 7898 12232
rect 7944 12220 7972 12251
rect 9398 12248 9404 12300
rect 9456 12288 9462 12300
rect 9766 12288 9772 12300
rect 9456 12260 9772 12288
rect 9456 12248 9462 12260
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 10134 12288 10140 12300
rect 10095 12260 10140 12288
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10244 12297 10272 12328
rect 14366 12316 14372 12368
rect 14424 12356 14430 12368
rect 14826 12356 14832 12368
rect 14424 12328 14832 12356
rect 14424 12316 14430 12328
rect 14826 12316 14832 12328
rect 14884 12316 14890 12368
rect 19429 12359 19487 12365
rect 19429 12325 19441 12359
rect 19475 12325 19487 12359
rect 20530 12356 20536 12368
rect 19429 12319 19487 12325
rect 19996 12328 20536 12356
rect 10229 12291 10287 12297
rect 10229 12257 10241 12291
rect 10275 12257 10287 12291
rect 18230 12288 18236 12300
rect 18143 12260 18236 12288
rect 10229 12251 10287 12257
rect 7892 12192 7972 12220
rect 7892 12180 7898 12192
rect 8478 12180 8484 12232
rect 8536 12220 8542 12232
rect 10689 12223 10747 12229
rect 10689 12220 10701 12223
rect 8536 12192 10701 12220
rect 8536 12180 8542 12192
rect 10689 12189 10701 12192
rect 10735 12189 10747 12223
rect 10689 12183 10747 12189
rect 12345 12223 12403 12229
rect 12345 12189 12357 12223
rect 12391 12220 12403 12223
rect 14274 12220 14280 12232
rect 12391 12192 14280 12220
rect 12391 12189 12403 12192
rect 12345 12183 12403 12189
rect 14274 12180 14280 12192
rect 14332 12220 14338 12232
rect 14829 12223 14887 12229
rect 14829 12220 14841 12223
rect 14332 12192 14841 12220
rect 14332 12180 14338 12192
rect 14829 12189 14841 12192
rect 14875 12189 14887 12223
rect 14829 12183 14887 12189
rect 14918 12180 14924 12232
rect 14976 12220 14982 12232
rect 15085 12223 15143 12229
rect 15085 12220 15097 12223
rect 14976 12192 15097 12220
rect 14976 12180 14982 12192
rect 15085 12189 15097 12192
rect 15131 12189 15143 12223
rect 17862 12220 17868 12232
rect 17823 12192 17868 12220
rect 15085 12183 15143 12189
rect 17862 12180 17868 12192
rect 17920 12180 17926 12232
rect 3789 12155 3847 12161
rect 3789 12152 3801 12155
rect 3252 12124 3801 12152
rect 3154 12115 3212 12121
rect 3789 12121 3801 12124
rect 3835 12121 3847 12155
rect 3789 12115 3847 12121
rect 4433 12155 4491 12161
rect 4433 12121 4445 12155
rect 4479 12152 4491 12155
rect 4522 12152 4528 12164
rect 4479 12124 4528 12152
rect 4479 12121 4491 12124
rect 4433 12115 4491 12121
rect 2038 12084 2044 12096
rect 1999 12056 2044 12084
rect 2038 12044 2044 12056
rect 2096 12044 2102 12096
rect 3160 12084 3188 12115
rect 4522 12112 4528 12124
rect 4580 12152 4586 12164
rect 10134 12152 10140 12164
rect 4580 12124 10140 12152
rect 4580 12112 4586 12124
rect 10134 12112 10140 12124
rect 10192 12112 10198 12164
rect 10956 12155 11014 12161
rect 10956 12121 10968 12155
rect 11002 12152 11014 12155
rect 11790 12152 11796 12164
rect 11002 12124 11796 12152
rect 11002 12121 11014 12124
rect 10956 12115 11014 12121
rect 11790 12112 11796 12124
rect 11848 12112 11854 12164
rect 12612 12155 12670 12161
rect 12612 12121 12624 12155
rect 12658 12121 12670 12155
rect 12612 12115 12670 12121
rect 17620 12155 17678 12161
rect 17620 12121 17632 12155
rect 17666 12152 17678 12155
rect 18156 12152 18184 12260
rect 18230 12248 18236 12260
rect 18288 12288 18294 12300
rect 18693 12291 18751 12297
rect 18693 12288 18705 12291
rect 18288 12260 18705 12288
rect 18288 12248 18294 12260
rect 18693 12257 18705 12260
rect 18739 12257 18751 12291
rect 19444 12288 19472 12319
rect 19518 12288 19524 12300
rect 19444 12260 19524 12288
rect 18693 12251 18751 12257
rect 19518 12248 19524 12260
rect 19576 12248 19582 12300
rect 19996 12220 20024 12328
rect 20530 12316 20536 12328
rect 20588 12316 20594 12368
rect 20073 12291 20131 12297
rect 20073 12257 20085 12291
rect 20119 12288 20131 12291
rect 20438 12288 20444 12300
rect 20119 12260 20444 12288
rect 20119 12257 20131 12260
rect 20073 12251 20131 12257
rect 20438 12248 20444 12260
rect 20496 12248 20502 12300
rect 20622 12220 20628 12232
rect 19306 12192 20024 12220
rect 20583 12192 20628 12220
rect 17666 12124 18184 12152
rect 17666 12121 17678 12124
rect 17620 12115 17678 12121
rect 3418 12084 3424 12096
rect 3160 12056 3424 12084
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 4614 12044 4620 12096
rect 4672 12084 4678 12096
rect 4982 12084 4988 12096
rect 4672 12056 4988 12084
rect 4672 12044 4678 12056
rect 4982 12044 4988 12056
rect 5040 12084 5046 12096
rect 5077 12087 5135 12093
rect 5077 12084 5089 12087
rect 5040 12056 5089 12084
rect 5040 12044 5046 12056
rect 5077 12053 5089 12056
rect 5123 12053 5135 12087
rect 5077 12047 5135 12053
rect 5169 12087 5227 12093
rect 5169 12053 5181 12087
rect 5215 12084 5227 12087
rect 5810 12084 5816 12096
rect 5215 12056 5816 12084
rect 5215 12053 5227 12056
rect 5169 12047 5227 12053
rect 5810 12044 5816 12056
rect 5868 12044 5874 12096
rect 6181 12087 6239 12093
rect 6181 12053 6193 12087
rect 6227 12084 6239 12087
rect 6914 12084 6920 12096
rect 6227 12056 6920 12084
rect 6227 12053 6239 12056
rect 6181 12047 6239 12053
rect 6914 12044 6920 12056
rect 6972 12044 6978 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 7837 12087 7895 12093
rect 7837 12084 7849 12087
rect 7340 12056 7849 12084
rect 7340 12044 7346 12056
rect 7837 12053 7849 12056
rect 7883 12084 7895 12087
rect 8754 12084 8760 12096
rect 7883 12056 8760 12084
rect 7883 12053 7895 12056
rect 7837 12047 7895 12053
rect 8754 12044 8760 12056
rect 8812 12044 8818 12096
rect 8938 12044 8944 12096
rect 8996 12084 9002 12096
rect 9677 12087 9735 12093
rect 9677 12084 9689 12087
rect 8996 12056 9689 12084
rect 8996 12044 9002 12056
rect 9677 12053 9689 12056
rect 9723 12053 9735 12087
rect 9677 12047 9735 12053
rect 9766 12044 9772 12096
rect 9824 12084 9830 12096
rect 10045 12087 10103 12093
rect 10045 12084 10057 12087
rect 9824 12056 10057 12084
rect 9824 12044 9830 12056
rect 10045 12053 10057 12056
rect 10091 12053 10103 12087
rect 10045 12047 10103 12053
rect 12069 12087 12127 12093
rect 12069 12053 12081 12087
rect 12115 12084 12127 12087
rect 12158 12084 12164 12096
rect 12115 12056 12164 12084
rect 12115 12053 12127 12056
rect 12069 12047 12127 12053
rect 12158 12044 12164 12056
rect 12216 12084 12222 12096
rect 12636 12084 12664 12115
rect 18414 12112 18420 12164
rect 18472 12152 18478 12164
rect 18601 12155 18659 12161
rect 18601 12152 18613 12155
rect 18472 12124 18613 12152
rect 18472 12112 18478 12124
rect 18601 12121 18613 12124
rect 18647 12152 18659 12155
rect 19306 12152 19334 12192
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 18647 12124 19334 12152
rect 19797 12155 19855 12161
rect 18647 12121 18659 12124
rect 18601 12115 18659 12121
rect 19797 12121 19809 12155
rect 19843 12152 19855 12155
rect 20530 12152 20536 12164
rect 19843 12124 20536 12152
rect 19843 12121 19855 12124
rect 19797 12115 19855 12121
rect 14182 12084 14188 12096
rect 12216 12056 14188 12084
rect 12216 12044 12222 12056
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14277 12087 14335 12093
rect 14277 12053 14289 12087
rect 14323 12084 14335 12087
rect 14458 12084 14464 12096
rect 14323 12056 14464 12084
rect 14323 12053 14335 12056
rect 14277 12047 14335 12053
rect 14458 12044 14464 12056
rect 14516 12044 14522 12096
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 16485 12087 16543 12093
rect 16485 12084 16497 12087
rect 14792 12056 16497 12084
rect 14792 12044 14798 12056
rect 16485 12053 16497 12056
rect 16531 12084 16543 12087
rect 17218 12084 17224 12096
rect 16531 12056 17224 12084
rect 16531 12053 16543 12056
rect 16485 12047 16543 12053
rect 17218 12044 17224 12056
rect 17276 12044 17282 12096
rect 17402 12044 17408 12096
rect 17460 12084 17466 12096
rect 18141 12087 18199 12093
rect 18141 12084 18153 12087
rect 17460 12056 18153 12084
rect 17460 12044 17466 12056
rect 18141 12053 18153 12056
rect 18187 12053 18199 12087
rect 18141 12047 18199 12053
rect 18509 12087 18567 12093
rect 18509 12053 18521 12087
rect 18555 12084 18567 12087
rect 19812 12084 19840 12115
rect 20530 12112 20536 12124
rect 20588 12112 20594 12164
rect 18555 12056 19840 12084
rect 19889 12087 19947 12093
rect 18555 12053 18567 12056
rect 18509 12047 18567 12053
rect 19889 12053 19901 12087
rect 19935 12084 19947 12087
rect 19978 12084 19984 12096
rect 19935 12056 19984 12084
rect 19935 12053 19947 12056
rect 19889 12047 19947 12053
rect 19978 12044 19984 12056
rect 20036 12044 20042 12096
rect 21266 12084 21272 12096
rect 21227 12056 21272 12084
rect 21266 12044 21272 12056
rect 21324 12044 21330 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 3050 11880 3056 11892
rect 3011 11852 3056 11880
rect 3050 11840 3056 11852
rect 3108 11840 3114 11892
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 5166 11880 5172 11892
rect 4304 11852 5172 11880
rect 4304 11840 4310 11852
rect 5166 11840 5172 11852
rect 5224 11840 5230 11892
rect 5626 11880 5632 11892
rect 5587 11852 5632 11880
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6457 11883 6515 11889
rect 6457 11849 6469 11883
rect 6503 11880 6515 11883
rect 6638 11880 6644 11892
rect 6503 11852 6644 11880
rect 6503 11849 6515 11852
rect 6457 11843 6515 11849
rect 6638 11840 6644 11852
rect 6696 11840 6702 11892
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 7193 11883 7251 11889
rect 7193 11880 7205 11883
rect 6788 11852 7205 11880
rect 6788 11840 6794 11852
rect 7193 11849 7205 11852
rect 7239 11849 7251 11883
rect 7193 11843 7251 11849
rect 7926 11840 7932 11892
rect 7984 11880 7990 11892
rect 8110 11880 8116 11892
rect 7984 11852 8116 11880
rect 7984 11840 7990 11852
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 8662 11840 8668 11892
rect 8720 11880 8726 11892
rect 9033 11883 9091 11889
rect 9033 11880 9045 11883
rect 8720 11852 9045 11880
rect 8720 11840 8726 11852
rect 9033 11849 9045 11852
rect 9079 11849 9091 11883
rect 9033 11843 9091 11849
rect 9493 11883 9551 11889
rect 9493 11849 9505 11883
rect 9539 11880 9551 11883
rect 9674 11880 9680 11892
rect 9539 11852 9680 11880
rect 9539 11849 9551 11852
rect 9493 11843 9551 11849
rect 9674 11840 9680 11852
rect 9732 11840 9738 11892
rect 11974 11880 11980 11892
rect 10152 11852 11980 11880
rect 1857 11815 1915 11821
rect 1857 11781 1869 11815
rect 1903 11812 1915 11815
rect 1903 11784 8616 11812
rect 1903 11781 1915 11784
rect 1857 11775 1915 11781
rect 1578 11704 1584 11756
rect 1636 11744 1642 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1636 11716 1685 11744
rect 1636 11704 1642 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 2682 11744 2688 11756
rect 2643 11716 2688 11744
rect 1673 11707 1731 11713
rect 2682 11704 2688 11716
rect 2740 11704 2746 11756
rect 3326 11744 3332 11756
rect 3287 11716 3332 11744
rect 3326 11704 3332 11716
rect 3384 11744 3390 11756
rect 3789 11747 3847 11753
rect 3789 11744 3801 11747
rect 3384 11716 3801 11744
rect 3384 11704 3390 11716
rect 3789 11713 3801 11716
rect 3835 11713 3847 11747
rect 3789 11707 3847 11713
rect 4249 11747 4307 11753
rect 4249 11713 4261 11747
rect 4295 11744 4307 11747
rect 4338 11744 4344 11756
rect 4295 11716 4344 11744
rect 4295 11713 4307 11716
rect 4249 11707 4307 11713
rect 4338 11704 4344 11716
rect 4396 11704 4402 11756
rect 4516 11747 4574 11753
rect 4516 11713 4528 11747
rect 4562 11744 4574 11747
rect 4982 11744 4988 11756
rect 4562 11716 4988 11744
rect 4562 11713 4574 11716
rect 4516 11707 4574 11713
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 7006 11704 7012 11756
rect 7064 11744 7070 11756
rect 7561 11747 7619 11753
rect 7561 11744 7573 11747
rect 7064 11716 7573 11744
rect 7064 11704 7070 11716
rect 7561 11713 7573 11716
rect 7607 11713 7619 11747
rect 7561 11707 7619 11713
rect 7653 11747 7711 11753
rect 7653 11713 7665 11747
rect 7699 11744 7711 11747
rect 7699 11716 8340 11744
rect 7699 11713 7711 11716
rect 7653 11707 7711 11713
rect 2038 11636 2044 11688
rect 2096 11676 2102 11688
rect 2409 11679 2467 11685
rect 2409 11676 2421 11679
rect 2096 11648 2421 11676
rect 2096 11636 2102 11648
rect 2409 11645 2421 11648
rect 2455 11645 2467 11679
rect 2409 11639 2467 11645
rect 2498 11636 2504 11688
rect 2556 11676 2562 11688
rect 2593 11679 2651 11685
rect 2593 11676 2605 11679
rect 2556 11648 2605 11676
rect 2556 11636 2562 11648
rect 2593 11645 2605 11648
rect 2639 11645 2651 11679
rect 2593 11639 2651 11645
rect 5810 11636 5816 11688
rect 5868 11676 5874 11688
rect 5905 11679 5963 11685
rect 5905 11676 5917 11679
rect 5868 11648 5917 11676
rect 5868 11636 5874 11648
rect 5905 11645 5917 11648
rect 5951 11645 5963 11679
rect 6914 11676 6920 11688
rect 6875 11648 6920 11676
rect 5905 11639 5963 11645
rect 6914 11636 6920 11648
rect 6972 11636 6978 11688
rect 7098 11636 7104 11688
rect 7156 11676 7162 11688
rect 7745 11679 7803 11685
rect 7745 11676 7757 11679
rect 7156 11648 7757 11676
rect 7156 11636 7162 11648
rect 7745 11645 7757 11648
rect 7791 11676 7803 11679
rect 7834 11676 7840 11688
rect 7791 11648 7840 11676
rect 7791 11645 7803 11648
rect 7745 11639 7803 11645
rect 7834 11636 7840 11648
rect 7892 11636 7898 11688
rect 8110 11608 8116 11620
rect 5828 11580 8116 11608
rect 3513 11543 3571 11549
rect 3513 11509 3525 11543
rect 3559 11540 3571 11543
rect 5828 11540 5856 11580
rect 8110 11568 8116 11580
rect 8168 11568 8174 11620
rect 8312 11617 8340 11716
rect 8588 11688 8616 11784
rect 8754 11772 8760 11824
rect 8812 11812 8818 11824
rect 10152 11812 10180 11852
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12713 11883 12771 11889
rect 12713 11849 12725 11883
rect 12759 11880 12771 11883
rect 13357 11883 13415 11889
rect 13357 11880 13369 11883
rect 12759 11852 13369 11880
rect 12759 11849 12771 11852
rect 12713 11843 12771 11849
rect 13357 11849 13369 11852
rect 13403 11849 13415 11883
rect 13357 11843 13415 11849
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11849 14151 11883
rect 14458 11880 14464 11892
rect 14419 11852 14464 11880
rect 14093 11843 14151 11849
rect 11790 11812 11796 11824
rect 8812 11784 10180 11812
rect 10244 11784 11796 11812
rect 8812 11772 8818 11784
rect 9401 11747 9459 11753
rect 9401 11713 9413 11747
rect 9447 11744 9459 11747
rect 9766 11744 9772 11756
rect 9447 11716 9772 11744
rect 9447 11713 9459 11716
rect 9401 11707 9459 11713
rect 9766 11704 9772 11716
rect 9824 11704 9830 11756
rect 8570 11636 8576 11688
rect 8628 11636 8634 11688
rect 9030 11636 9036 11688
rect 9088 11676 9094 11688
rect 10244 11685 10272 11784
rect 11790 11772 11796 11784
rect 11848 11772 11854 11824
rect 12345 11815 12403 11821
rect 12345 11781 12357 11815
rect 12391 11812 12403 11815
rect 14108 11812 14136 11843
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 15565 11883 15623 11889
rect 15565 11849 15577 11883
rect 15611 11880 15623 11883
rect 16945 11883 17003 11889
rect 16945 11880 16957 11883
rect 15611 11852 16957 11880
rect 15611 11849 15623 11852
rect 15565 11843 15623 11849
rect 16945 11849 16957 11852
rect 16991 11849 17003 11883
rect 17310 11880 17316 11892
rect 17271 11852 17316 11880
rect 16945 11843 17003 11849
rect 17310 11840 17316 11852
rect 17368 11840 17374 11892
rect 17402 11840 17408 11892
rect 17460 11880 17466 11892
rect 17460 11852 17505 11880
rect 17460 11840 17466 11852
rect 17586 11840 17592 11892
rect 17644 11880 17650 11892
rect 19978 11880 19984 11892
rect 17644 11852 19984 11880
rect 17644 11840 17650 11852
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20898 11840 20904 11892
rect 20956 11880 20962 11892
rect 20993 11883 21051 11889
rect 20993 11880 21005 11883
rect 20956 11852 21005 11880
rect 20956 11840 20962 11852
rect 20993 11849 21005 11852
rect 21039 11849 21051 11883
rect 20993 11843 21051 11849
rect 21085 11883 21143 11889
rect 21085 11849 21097 11883
rect 21131 11880 21143 11883
rect 21174 11880 21180 11892
rect 21131 11852 21180 11880
rect 21131 11849 21143 11852
rect 21085 11843 21143 11849
rect 21174 11840 21180 11852
rect 21232 11840 21238 11892
rect 12391 11784 14136 11812
rect 12391 11781 12403 11784
rect 12345 11775 12403 11781
rect 14182 11772 14188 11824
rect 14240 11812 14246 11824
rect 16301 11815 16359 11821
rect 14240 11784 15700 11812
rect 14240 11772 14246 11784
rect 10410 11744 10416 11756
rect 10371 11716 10416 11744
rect 10410 11704 10416 11716
rect 10468 11704 10474 11756
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 13188 11716 15485 11744
rect 9585 11679 9643 11685
rect 9585 11676 9597 11679
rect 9088 11648 9597 11676
rect 9088 11636 9094 11648
rect 9585 11645 9597 11648
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 10229 11679 10287 11685
rect 10229 11645 10241 11679
rect 10275 11645 10287 11679
rect 10229 11639 10287 11645
rect 10321 11679 10379 11685
rect 10321 11645 10333 11679
rect 10367 11676 10379 11679
rect 10502 11676 10508 11688
rect 10367 11648 10508 11676
rect 10367 11645 10379 11648
rect 10321 11639 10379 11645
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 12158 11676 12164 11688
rect 12119 11648 12164 11676
rect 12158 11636 12164 11648
rect 12216 11636 12222 11688
rect 12253 11679 12311 11685
rect 12253 11645 12265 11679
rect 12299 11676 12311 11679
rect 12526 11676 12532 11688
rect 12299 11648 12532 11676
rect 12299 11645 12311 11648
rect 12253 11639 12311 11645
rect 12526 11636 12532 11648
rect 12584 11636 12590 11688
rect 13078 11676 13084 11688
rect 13039 11648 13084 11676
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 8297 11611 8355 11617
rect 8297 11577 8309 11611
rect 8343 11608 8355 11611
rect 9858 11608 9864 11620
rect 8343 11580 9864 11608
rect 8343 11577 8355 11580
rect 8297 11571 8355 11577
rect 9858 11568 9864 11580
rect 9916 11568 9922 11620
rect 10781 11611 10839 11617
rect 10781 11577 10793 11611
rect 10827 11608 10839 11611
rect 13188 11608 13216 11716
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 13265 11679 13323 11685
rect 13265 11645 13277 11679
rect 13311 11645 13323 11679
rect 13265 11639 13323 11645
rect 10827 11580 13216 11608
rect 13280 11608 13308 11639
rect 14366 11636 14372 11688
rect 14424 11676 14430 11688
rect 14553 11679 14611 11685
rect 14553 11676 14565 11679
rect 14424 11648 14565 11676
rect 14424 11636 14430 11648
rect 14553 11645 14565 11648
rect 14599 11645 14611 11679
rect 14734 11676 14740 11688
rect 14695 11648 14740 11676
rect 14553 11639 14611 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 15672 11685 15700 11784
rect 16301 11781 16313 11815
rect 16347 11812 16359 11815
rect 20254 11812 20260 11824
rect 16347 11784 20260 11812
rect 16347 11781 16359 11784
rect 16301 11775 16359 11781
rect 20254 11772 20260 11784
rect 20312 11772 20318 11824
rect 18325 11747 18383 11753
rect 18325 11713 18337 11747
rect 18371 11744 18383 11747
rect 18598 11744 18604 11756
rect 18371 11716 18604 11744
rect 18371 11713 18383 11716
rect 18325 11707 18383 11713
rect 18598 11704 18604 11716
rect 18656 11704 18662 11756
rect 19058 11744 19064 11756
rect 19019 11716 19064 11744
rect 19058 11704 19064 11716
rect 19116 11704 19122 11756
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11713 20131 11747
rect 20073 11707 20131 11713
rect 15657 11679 15715 11685
rect 15657 11645 15669 11679
rect 15703 11645 15715 11679
rect 15657 11639 15715 11645
rect 17218 11636 17224 11688
rect 17276 11676 17282 11688
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 17276 11648 17509 11676
rect 17276 11636 17282 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 17770 11636 17776 11688
rect 17828 11676 17834 11688
rect 20088 11676 20116 11707
rect 17828 11648 20116 11676
rect 17828 11636 17834 11648
rect 20622 11636 20628 11688
rect 20680 11676 20686 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 20680 11648 21189 11676
rect 20680 11636 20686 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 15105 11611 15163 11617
rect 15105 11608 15117 11611
rect 13280 11580 15117 11608
rect 10827 11577 10839 11580
rect 10781 11571 10839 11577
rect 15105 11577 15117 11580
rect 15151 11577 15163 11611
rect 15105 11571 15163 11577
rect 18785 11611 18843 11617
rect 18785 11577 18797 11611
rect 18831 11608 18843 11611
rect 20070 11608 20076 11620
rect 18831 11580 20076 11608
rect 18831 11577 18843 11580
rect 18785 11571 18843 11577
rect 20070 11568 20076 11580
rect 20128 11568 20134 11620
rect 3559 11512 5856 11540
rect 3559 11509 3571 11512
rect 3513 11503 3571 11509
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 7926 11540 7932 11552
rect 5960 11512 7932 11540
rect 5960 11500 5966 11512
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8018 11500 8024 11552
rect 8076 11540 8082 11552
rect 8573 11543 8631 11549
rect 8573 11540 8585 11543
rect 8076 11512 8585 11540
rect 8076 11500 8082 11512
rect 8573 11509 8585 11512
rect 8619 11509 8631 11543
rect 8573 11503 8631 11509
rect 11149 11543 11207 11549
rect 11149 11509 11161 11543
rect 11195 11540 11207 11543
rect 11238 11540 11244 11552
rect 11195 11512 11244 11540
rect 11195 11509 11207 11512
rect 11149 11503 11207 11509
rect 11238 11500 11244 11512
rect 11296 11500 11302 11552
rect 11701 11543 11759 11549
rect 11701 11509 11713 11543
rect 11747 11540 11759 11543
rect 13630 11540 13636 11552
rect 11747 11512 13636 11540
rect 11747 11509 11759 11512
rect 11701 11503 11759 11509
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 13725 11543 13783 11549
rect 13725 11509 13737 11543
rect 13771 11540 13783 11543
rect 16390 11540 16396 11552
rect 13771 11512 16396 11540
rect 13771 11509 13783 11512
rect 13725 11503 13783 11509
rect 16390 11500 16396 11512
rect 16448 11500 16454 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18322 11540 18328 11552
rect 18104 11512 18328 11540
rect 18104 11500 18110 11512
rect 18322 11500 18328 11512
rect 18380 11500 18386 11552
rect 19518 11500 19524 11552
rect 19576 11540 19582 11552
rect 19705 11543 19763 11549
rect 19705 11540 19717 11543
rect 19576 11512 19717 11540
rect 19576 11500 19582 11512
rect 19705 11509 19717 11512
rect 19751 11509 19763 11543
rect 19705 11503 19763 11509
rect 20254 11500 20260 11552
rect 20312 11540 20318 11552
rect 20625 11543 20683 11549
rect 20625 11540 20637 11543
rect 20312 11512 20637 11540
rect 20312 11500 20318 11512
rect 20625 11509 20637 11512
rect 20671 11509 20683 11543
rect 20625 11503 20683 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 1670 11336 1676 11348
rect 1631 11308 1676 11336
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 2498 11336 2504 11348
rect 2459 11308 2504 11336
rect 2498 11296 2504 11308
rect 2556 11296 2562 11348
rect 9490 11336 9496 11348
rect 2746 11308 9496 11336
rect 2133 11271 2191 11277
rect 2133 11237 2145 11271
rect 2179 11268 2191 11271
rect 2746 11268 2774 11308
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 9766 11336 9772 11348
rect 9727 11308 9772 11336
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 10134 11296 10140 11348
rect 10192 11336 10198 11348
rect 10229 11339 10287 11345
rect 10229 11336 10241 11339
rect 10192 11308 10241 11336
rect 10192 11296 10198 11308
rect 10229 11305 10241 11308
rect 10275 11305 10287 11339
rect 11054 11336 11060 11348
rect 11015 11308 11060 11336
rect 10229 11299 10287 11305
rect 11054 11296 11060 11308
rect 11112 11296 11118 11348
rect 12253 11339 12311 11345
rect 12253 11305 12265 11339
rect 12299 11336 12311 11339
rect 12986 11336 12992 11348
rect 12299 11308 12992 11336
rect 12299 11305 12311 11308
rect 12253 11299 12311 11305
rect 12986 11296 12992 11308
rect 13044 11296 13050 11348
rect 13630 11296 13636 11348
rect 13688 11336 13694 11348
rect 20622 11336 20628 11348
rect 13688 11308 20300 11336
rect 20583 11308 20628 11336
rect 13688 11296 13694 11308
rect 2179 11240 2774 11268
rect 2179 11237 2191 11240
rect 2133 11231 2191 11237
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 4801 11271 4859 11277
rect 4801 11268 4813 11271
rect 3936 11240 4813 11268
rect 3936 11228 3942 11240
rect 4801 11237 4813 11240
rect 4847 11237 4859 11271
rect 4801 11231 4859 11237
rect 5905 11271 5963 11277
rect 5905 11237 5917 11271
rect 5951 11237 5963 11271
rect 5905 11231 5963 11237
rect 7101 11271 7159 11277
rect 7101 11237 7113 11271
rect 7147 11237 7159 11271
rect 7101 11231 7159 11237
rect 2958 11200 2964 11212
rect 2884 11172 2964 11200
rect 1486 11132 1492 11144
rect 1447 11104 1492 11132
rect 1486 11092 1492 11104
rect 1544 11092 1550 11144
rect 1946 11132 1952 11144
rect 1907 11104 1952 11132
rect 1946 11092 1952 11104
rect 2004 11092 2010 11144
rect 2884 11141 2912 11172
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3145 11203 3203 11209
rect 3145 11169 3157 11203
rect 3191 11200 3203 11203
rect 3418 11200 3424 11212
rect 3191 11172 3424 11200
rect 3191 11169 3203 11172
rect 3145 11163 3203 11169
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 5353 11203 5411 11209
rect 5353 11200 5365 11203
rect 3896 11172 5365 11200
rect 2869 11135 2927 11141
rect 2869 11101 2881 11135
rect 2915 11101 2927 11135
rect 2869 11095 2927 11101
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 3896 11141 3924 11172
rect 5353 11169 5365 11172
rect 5399 11169 5411 11203
rect 5353 11163 5411 11169
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3844 11104 3893 11132
rect 3844 11092 3850 11104
rect 3881 11101 3893 11104
rect 3927 11101 3939 11135
rect 3881 11095 3939 11101
rect 4525 11135 4583 11141
rect 4525 11101 4537 11135
rect 4571 11132 4583 11135
rect 4982 11132 4988 11144
rect 4571 11104 4988 11132
rect 4571 11101 4583 11104
rect 4525 11095 4583 11101
rect 4982 11092 4988 11104
rect 5040 11092 5046 11144
rect 5169 11135 5227 11141
rect 5169 11101 5181 11135
rect 5215 11132 5227 11135
rect 5920 11132 5948 11231
rect 5994 11160 6000 11212
rect 6052 11200 6058 11212
rect 6457 11203 6515 11209
rect 6457 11200 6469 11203
rect 6052 11172 6469 11200
rect 6052 11160 6058 11172
rect 6457 11169 6469 11172
rect 6503 11200 6515 11203
rect 7116 11200 7144 11231
rect 11790 11228 11796 11280
rect 11848 11268 11854 11280
rect 14734 11268 14740 11280
rect 11848 11240 14740 11268
rect 11848 11228 11854 11240
rect 14734 11228 14740 11240
rect 14792 11228 14798 11280
rect 16669 11271 16727 11277
rect 16669 11237 16681 11271
rect 16715 11268 16727 11271
rect 17126 11268 17132 11280
rect 16715 11240 17132 11268
rect 16715 11237 16727 11240
rect 16669 11231 16727 11237
rect 17126 11228 17132 11240
rect 17184 11268 17190 11280
rect 17770 11268 17776 11280
rect 17184 11240 17776 11268
rect 17184 11228 17190 11240
rect 17770 11228 17776 11240
rect 17828 11228 17834 11280
rect 8478 11200 8484 11212
rect 6503 11172 7144 11200
rect 8439 11172 8484 11200
rect 6503 11169 6515 11172
rect 6457 11163 6515 11169
rect 8478 11160 8484 11172
rect 8536 11160 8542 11212
rect 9214 11200 9220 11212
rect 9175 11172 9220 11200
rect 9214 11160 9220 11172
rect 9272 11160 9278 11212
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10042 11200 10048 11212
rect 9916 11172 10048 11200
rect 9916 11160 9922 11172
rect 10042 11160 10048 11172
rect 10100 11160 10106 11212
rect 15841 11203 15899 11209
rect 15841 11169 15853 11203
rect 15887 11200 15899 11203
rect 17862 11200 17868 11212
rect 15887 11172 17868 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 17862 11160 17868 11172
rect 17920 11160 17926 11212
rect 18230 11200 18236 11212
rect 18191 11172 18236 11200
rect 18230 11160 18236 11172
rect 18288 11160 18294 11212
rect 5215 11104 5948 11132
rect 6196 11104 6868 11132
rect 5215 11101 5227 11104
rect 5169 11095 5227 11101
rect 2130 11024 2136 11076
rect 2188 11064 2194 11076
rect 2961 11067 3019 11073
rect 2961 11064 2973 11067
rect 2188 11036 2973 11064
rect 2188 11024 2194 11036
rect 2961 11033 2973 11036
rect 3007 11064 3019 11067
rect 3007 11036 5396 11064
rect 3007 11033 3019 11036
rect 2961 11027 3019 11033
rect 5258 10996 5264 11008
rect 5219 10968 5264 10996
rect 5258 10956 5264 10968
rect 5316 10956 5322 11008
rect 5368 10996 5396 11036
rect 5534 10996 5540 11008
rect 5368 10968 5540 10996
rect 5534 10956 5540 10968
rect 5592 10956 5598 11008
rect 5902 10956 5908 11008
rect 5960 10996 5966 11008
rect 6196 10996 6224 11104
rect 6273 11067 6331 11073
rect 6273 11033 6285 11067
rect 6319 11064 6331 11067
rect 6730 11064 6736 11076
rect 6319 11036 6736 11064
rect 6319 11033 6331 11036
rect 6273 11027 6331 11033
rect 6730 11024 6736 11036
rect 6788 11024 6794 11076
rect 5960 10968 6224 10996
rect 6365 10999 6423 11005
rect 5960 10956 5966 10968
rect 6365 10965 6377 10999
rect 6411 10996 6423 10999
rect 6638 10996 6644 11008
rect 6411 10968 6644 10996
rect 6411 10965 6423 10968
rect 6365 10959 6423 10965
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 6840 10996 6868 11104
rect 7098 11092 7104 11144
rect 7156 11132 7162 11144
rect 9398 11132 9404 11144
rect 7156 11104 8340 11132
rect 9359 11104 9404 11132
rect 7156 11092 7162 11104
rect 7282 11024 7288 11076
rect 7340 11064 7346 11076
rect 8214 11067 8272 11073
rect 8214 11064 8226 11067
rect 7340 11036 8226 11064
rect 7340 11024 7346 11036
rect 8214 11033 8226 11036
rect 8260 11033 8272 11067
rect 8312 11064 8340 11104
rect 9398 11092 9404 11104
rect 9456 11092 9462 11144
rect 15585 11135 15643 11141
rect 15585 11101 15597 11135
rect 15631 11132 15643 11135
rect 15746 11132 15752 11144
rect 15631 11104 15752 11132
rect 15631 11101 15643 11104
rect 15585 11095 15643 11101
rect 15746 11092 15752 11104
rect 15804 11092 15810 11144
rect 17034 11092 17040 11144
rect 17092 11132 17098 11144
rect 17313 11135 17371 11141
rect 17313 11132 17325 11135
rect 17092 11104 17325 11132
rect 17092 11092 17098 11104
rect 17313 11101 17325 11104
rect 17359 11101 17371 11135
rect 17880 11132 17908 11160
rect 19518 11141 19524 11144
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 17880 11104 19257 11132
rect 17313 11095 17371 11101
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19512 11132 19524 11141
rect 19479 11104 19524 11132
rect 19245 11095 19303 11101
rect 19512 11095 19524 11104
rect 9309 11067 9367 11073
rect 9309 11064 9321 11067
rect 8312 11036 9321 11064
rect 8214 11027 8272 11033
rect 9309 11033 9321 11036
rect 9355 11033 9367 11067
rect 9309 11027 9367 11033
rect 9858 11024 9864 11076
rect 9916 11064 9922 11076
rect 10597 11067 10655 11073
rect 10597 11064 10609 11067
rect 9916 11036 10609 11064
rect 9916 11024 9922 11036
rect 10597 11033 10609 11036
rect 10643 11033 10655 11067
rect 11974 11064 11980 11076
rect 10597 11027 10655 11033
rect 11348 11036 11980 11064
rect 11146 10996 11152 11008
rect 6840 10968 11152 10996
rect 11146 10956 11152 10968
rect 11204 10996 11210 11008
rect 11348 11005 11376 11036
rect 11974 11024 11980 11036
rect 12032 11024 12038 11076
rect 13538 11064 13544 11076
rect 13499 11036 13544 11064
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14185 11067 14243 11073
rect 14185 11033 14197 11067
rect 14231 11064 14243 11067
rect 14366 11064 14372 11076
rect 14231 11036 14372 11064
rect 14231 11033 14243 11036
rect 14185 11027 14243 11033
rect 14366 11024 14372 11036
rect 14424 11064 14430 11076
rect 15102 11064 15108 11076
rect 14424 11036 15108 11064
rect 14424 11024 14430 11036
rect 15102 11024 15108 11036
rect 15160 11024 15166 11076
rect 15930 11024 15936 11076
rect 15988 11064 15994 11076
rect 16117 11067 16175 11073
rect 16117 11064 16129 11067
rect 15988 11036 16129 11064
rect 15988 11024 15994 11036
rect 16117 11033 16129 11036
rect 16163 11033 16175 11067
rect 17328 11064 17356 11095
rect 19518 11092 19524 11095
rect 19576 11092 19582 11144
rect 20272 11132 20300 11308
rect 20622 11296 20628 11308
rect 20680 11296 20686 11348
rect 21174 11336 21180 11348
rect 21135 11308 21180 11336
rect 21174 11296 21180 11308
rect 21232 11296 21238 11348
rect 21269 11135 21327 11141
rect 21269 11132 21281 11135
rect 20272 11104 21281 11132
rect 21269 11101 21281 11104
rect 21315 11132 21327 11135
rect 21358 11132 21364 11144
rect 21315 11104 21364 11132
rect 21315 11101 21327 11104
rect 21269 11095 21327 11101
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 18049 11067 18107 11073
rect 17328 11036 18000 11064
rect 16117 11027 16175 11033
rect 11333 10999 11391 11005
rect 11333 10996 11345 10999
rect 11204 10968 11345 10996
rect 11204 10956 11210 10968
rect 11333 10965 11345 10968
rect 11379 10965 11391 10999
rect 11333 10959 11391 10965
rect 11698 10956 11704 11008
rect 11756 10996 11762 11008
rect 12894 10996 12900 11008
rect 11756 10968 12900 10996
rect 11756 10956 11762 10968
rect 12894 10956 12900 10968
rect 12952 10956 12958 11008
rect 13814 10956 13820 11008
rect 13872 10996 13878 11008
rect 14461 10999 14519 11005
rect 14461 10996 14473 10999
rect 13872 10968 14473 10996
rect 13872 10956 13878 10968
rect 14461 10965 14473 10968
rect 14507 10996 14519 10999
rect 16390 10996 16396 11008
rect 14507 10968 16396 10996
rect 14507 10965 14519 10968
rect 14461 10959 14519 10965
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 16942 10996 16948 11008
rect 16903 10968 16948 10996
rect 16942 10956 16948 10968
rect 17000 10956 17006 11008
rect 17678 10996 17684 11008
rect 17639 10968 17684 10996
rect 17678 10956 17684 10968
rect 17736 10956 17742 11008
rect 17972 10996 18000 11036
rect 18049 11033 18061 11067
rect 18095 11064 18107 11067
rect 18693 11067 18751 11073
rect 18693 11064 18705 11067
rect 18095 11036 18705 11064
rect 18095 11033 18107 11036
rect 18049 11027 18107 11033
rect 18693 11033 18705 11036
rect 18739 11033 18751 11067
rect 18693 11027 18751 11033
rect 18141 10999 18199 11005
rect 18141 10996 18153 10999
rect 17972 10968 18153 10996
rect 18141 10965 18153 10968
rect 18187 10965 18199 10999
rect 18141 10959 18199 10965
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 1578 10752 1584 10804
rect 1636 10792 1642 10804
rect 2133 10795 2191 10801
rect 2133 10792 2145 10795
rect 1636 10764 2145 10792
rect 1636 10752 1642 10764
rect 2133 10761 2145 10764
rect 2179 10761 2191 10795
rect 2133 10755 2191 10761
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2682 10792 2688 10804
rect 2547 10764 2688 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2682 10752 2688 10764
rect 2740 10752 2746 10804
rect 2869 10795 2927 10801
rect 2869 10761 2881 10795
rect 2915 10792 2927 10795
rect 3050 10792 3056 10804
rect 2915 10764 3056 10792
rect 2915 10761 2927 10764
rect 2869 10755 2927 10761
rect 3050 10752 3056 10764
rect 3108 10792 3114 10804
rect 3602 10792 3608 10804
rect 3108 10764 3608 10792
rect 3108 10752 3114 10764
rect 3602 10752 3608 10764
rect 3660 10752 3666 10804
rect 3786 10792 3792 10804
rect 3747 10764 3792 10792
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 4706 10752 4712 10804
rect 4764 10792 4770 10804
rect 5902 10792 5908 10804
rect 4764 10764 5908 10792
rect 4764 10752 4770 10764
rect 5902 10752 5908 10764
rect 5960 10752 5966 10804
rect 6730 10792 6736 10804
rect 6691 10764 6736 10792
rect 6730 10752 6736 10764
rect 6788 10752 6794 10804
rect 6914 10752 6920 10804
rect 6972 10792 6978 10804
rect 7101 10795 7159 10801
rect 7101 10792 7113 10795
rect 6972 10764 7113 10792
rect 6972 10752 6978 10764
rect 7101 10761 7113 10764
rect 7147 10761 7159 10795
rect 7101 10755 7159 10761
rect 7193 10795 7251 10801
rect 7193 10761 7205 10795
rect 7239 10792 7251 10795
rect 7466 10792 7472 10804
rect 7239 10764 7472 10792
rect 7239 10761 7251 10764
rect 7193 10755 7251 10761
rect 7466 10752 7472 10764
rect 7524 10752 7530 10804
rect 7650 10752 7656 10804
rect 7708 10792 7714 10804
rect 7708 10764 8524 10792
rect 7708 10752 7714 10764
rect 4430 10724 4436 10736
rect 2746 10696 4436 10724
rect 1670 10656 1676 10668
rect 1631 10628 1676 10656
rect 1670 10616 1676 10628
rect 1728 10656 1734 10668
rect 2746 10656 2774 10696
rect 4430 10684 4436 10696
rect 4488 10684 4494 10736
rect 4924 10727 4982 10733
rect 4924 10693 4936 10727
rect 4970 10724 4982 10727
rect 8389 10727 8447 10733
rect 8389 10724 8401 10727
rect 4970 10696 8401 10724
rect 4970 10693 4982 10696
rect 4924 10687 4982 10693
rect 8389 10693 8401 10696
rect 8435 10693 8447 10727
rect 8496 10724 8524 10764
rect 8570 10752 8576 10804
rect 8628 10792 8634 10804
rect 11698 10792 11704 10804
rect 8628 10764 11704 10792
rect 8628 10752 8634 10764
rect 11698 10752 11704 10764
rect 11756 10752 11762 10804
rect 11885 10795 11943 10801
rect 11885 10761 11897 10795
rect 11931 10792 11943 10795
rect 11974 10792 11980 10804
rect 11931 10764 11980 10792
rect 11931 10761 11943 10764
rect 11885 10755 11943 10761
rect 11974 10752 11980 10764
rect 12032 10752 12038 10804
rect 12253 10795 12311 10801
rect 12253 10761 12265 10795
rect 12299 10792 12311 10795
rect 14829 10795 14887 10801
rect 14829 10792 14841 10795
rect 12299 10764 14841 10792
rect 12299 10761 12311 10764
rect 12253 10755 12311 10761
rect 14829 10761 14841 10764
rect 14875 10761 14887 10795
rect 14829 10755 14887 10761
rect 17037 10795 17095 10801
rect 17037 10761 17049 10795
rect 17083 10792 17095 10795
rect 17678 10792 17684 10804
rect 17083 10764 17684 10792
rect 17083 10761 17095 10764
rect 17037 10755 17095 10761
rect 17678 10752 17684 10764
rect 17736 10752 17742 10804
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 18966 10792 18972 10804
rect 18840 10764 18972 10792
rect 18840 10752 18846 10764
rect 18966 10752 18972 10764
rect 19024 10752 19030 10804
rect 9493 10727 9551 10733
rect 9493 10724 9505 10727
rect 8496 10696 9505 10724
rect 8389 10687 8447 10693
rect 9493 10693 9505 10696
rect 9539 10693 9551 10727
rect 9493 10687 9551 10693
rect 10134 10684 10140 10736
rect 10192 10724 10198 10736
rect 10192 10696 12020 10724
rect 10192 10684 10198 10696
rect 1728 10628 2774 10656
rect 2961 10659 3019 10665
rect 1728 10616 1734 10628
rect 2961 10625 2973 10659
rect 3007 10656 3019 10659
rect 3326 10656 3332 10668
rect 3007 10628 3332 10656
rect 3007 10625 3019 10628
rect 2961 10619 3019 10625
rect 3326 10616 3332 10628
rect 3384 10616 3390 10668
rect 5074 10616 5080 10668
rect 5132 10656 5138 10668
rect 5629 10659 5687 10665
rect 5629 10656 5641 10659
rect 5132 10628 5641 10656
rect 5132 10616 5138 10628
rect 5629 10625 5641 10628
rect 5675 10625 5687 10659
rect 5629 10619 5687 10625
rect 5994 10616 6000 10668
rect 6052 10656 6058 10668
rect 7745 10659 7803 10665
rect 7745 10656 7757 10659
rect 6052 10628 7757 10656
rect 6052 10616 6058 10628
rect 7745 10625 7757 10628
rect 7791 10625 7803 10659
rect 7745 10619 7803 10625
rect 9766 10616 9772 10668
rect 9824 10656 9830 10668
rect 10781 10659 10839 10665
rect 10781 10656 10793 10659
rect 9824 10628 10793 10656
rect 9824 10616 9830 10628
rect 10781 10625 10793 10628
rect 10827 10625 10839 10659
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 10781 10619 10839 10625
rect 10879 10628 11805 10656
rect 3145 10591 3203 10597
rect 3145 10557 3157 10591
rect 3191 10588 3203 10591
rect 3418 10588 3424 10600
rect 3191 10560 3424 10588
rect 3191 10557 3203 10560
rect 3145 10551 3203 10557
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 5166 10588 5172 10600
rect 5127 10560 5172 10588
rect 5166 10548 5172 10560
rect 5224 10548 5230 10600
rect 7282 10588 7288 10600
rect 7243 10560 7288 10588
rect 7282 10548 7288 10560
rect 7340 10548 7346 10600
rect 7374 10548 7380 10600
rect 7432 10588 7438 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 7432 10560 9137 10588
rect 7432 10548 7438 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9125 10551 9183 10557
rect 9398 10548 9404 10600
rect 9456 10588 9462 10600
rect 9953 10591 10011 10597
rect 9953 10588 9965 10591
rect 9456 10560 9965 10588
rect 9456 10548 9462 10560
rect 9953 10557 9965 10560
rect 9999 10557 10011 10591
rect 9953 10551 10011 10557
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10505 10591 10563 10597
rect 10505 10588 10517 10591
rect 10376 10560 10517 10588
rect 10376 10548 10382 10560
rect 10505 10557 10517 10560
rect 10551 10557 10563 10591
rect 10686 10588 10692 10600
rect 10647 10560 10692 10588
rect 10505 10551 10563 10557
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 1857 10523 1915 10529
rect 1857 10489 1869 10523
rect 1903 10520 1915 10523
rect 2498 10520 2504 10532
rect 1903 10492 2504 10520
rect 1903 10489 1915 10492
rect 1857 10483 1915 10489
rect 2498 10480 2504 10492
rect 2556 10480 2562 10532
rect 6457 10523 6515 10529
rect 2746 10492 3924 10520
rect 2222 10412 2228 10464
rect 2280 10452 2286 10464
rect 2746 10452 2774 10492
rect 2280 10424 2774 10452
rect 3896 10452 3924 10492
rect 6457 10489 6469 10523
rect 6503 10520 6515 10523
rect 7466 10520 7472 10532
rect 6503 10492 7472 10520
rect 6503 10489 6515 10492
rect 6457 10483 6515 10489
rect 7466 10480 7472 10492
rect 7524 10480 7530 10532
rect 8478 10480 8484 10532
rect 8536 10520 8542 10532
rect 10879 10520 10907 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 11146 10548 11152 10600
rect 11204 10588 11210 10600
rect 11609 10591 11667 10597
rect 11609 10588 11621 10591
rect 11204 10560 11621 10588
rect 11204 10548 11210 10560
rect 11609 10557 11621 10560
rect 11655 10557 11667 10591
rect 11992 10588 12020 10696
rect 12066 10684 12072 10736
rect 12124 10724 12130 10736
rect 12710 10724 12716 10736
rect 12124 10696 12716 10724
rect 12124 10684 12130 10696
rect 12710 10684 12716 10696
rect 12768 10684 12774 10736
rect 17948 10727 18006 10733
rect 17948 10693 17960 10727
rect 17994 10724 18006 10727
rect 18230 10724 18236 10736
rect 17994 10696 18236 10724
rect 17994 10693 18006 10696
rect 17948 10687 18006 10693
rect 18230 10684 18236 10696
rect 18288 10684 18294 10736
rect 19518 10724 19524 10736
rect 19306 10696 19524 10724
rect 13078 10656 13084 10668
rect 13039 10628 13084 10656
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 15286 10656 15292 10668
rect 14783 10628 15292 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 15286 10616 15292 10628
rect 15344 10616 15350 10668
rect 16298 10656 16304 10668
rect 15396 10628 16304 10656
rect 15013 10591 15071 10597
rect 11992 10560 14964 10588
rect 11609 10551 11667 10557
rect 12802 10520 12808 10532
rect 8536 10492 10907 10520
rect 12763 10492 12808 10520
rect 8536 10480 8542 10492
rect 12802 10480 12808 10492
rect 12860 10480 12866 10532
rect 14093 10523 14151 10529
rect 14093 10489 14105 10523
rect 14139 10520 14151 10523
rect 14274 10520 14280 10532
rect 14139 10492 14280 10520
rect 14139 10489 14151 10492
rect 14093 10483 14151 10489
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 14936 10520 14964 10560
rect 15013 10557 15025 10591
rect 15059 10588 15071 10591
rect 15396 10588 15424 10628
rect 16298 10616 16304 10628
rect 16356 10616 16362 10668
rect 19306 10656 19334 10696
rect 19518 10684 19524 10696
rect 19576 10684 19582 10736
rect 21116 10727 21174 10733
rect 21116 10693 21128 10727
rect 21162 10724 21174 10727
rect 21266 10724 21272 10736
rect 21162 10696 21272 10724
rect 21162 10693 21174 10696
rect 21116 10687 21174 10693
rect 21266 10684 21272 10696
rect 21324 10684 21330 10736
rect 17236 10628 19334 10656
rect 15654 10588 15660 10600
rect 15059 10560 15424 10588
rect 15615 10560 15660 10588
rect 15059 10557 15071 10560
rect 15013 10551 15071 10557
rect 15654 10548 15660 10560
rect 15712 10548 15718 10600
rect 17126 10588 17132 10600
rect 17087 10560 17132 10588
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17034 10520 17040 10532
rect 14936 10492 17040 10520
rect 17034 10480 17040 10492
rect 17092 10520 17098 10532
rect 17236 10520 17264 10628
rect 17313 10591 17371 10597
rect 17313 10557 17325 10591
rect 17359 10557 17371 10591
rect 17678 10588 17684 10600
rect 17639 10560 17684 10588
rect 17313 10551 17371 10557
rect 17092 10492 17264 10520
rect 17092 10480 17098 10492
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 3896 10424 5457 10452
rect 2280 10412 2286 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 5902 10452 5908 10464
rect 5863 10424 5908 10452
rect 5445 10415 5503 10421
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 8849 10455 8907 10461
rect 8849 10421 8861 10455
rect 8895 10452 8907 10455
rect 9214 10452 9220 10464
rect 8895 10424 9220 10452
rect 8895 10421 8907 10424
rect 8849 10415 8907 10421
rect 9214 10412 9220 10424
rect 9272 10412 9278 10464
rect 11054 10412 11060 10464
rect 11112 10452 11118 10464
rect 11149 10455 11207 10461
rect 11149 10452 11161 10455
rect 11112 10424 11161 10452
rect 11112 10412 11118 10424
rect 11149 10421 11161 10424
rect 11195 10421 11207 10455
rect 11149 10415 11207 10421
rect 13725 10455 13783 10461
rect 13725 10421 13737 10455
rect 13771 10452 13783 10455
rect 13814 10452 13820 10464
rect 13771 10424 13820 10452
rect 13771 10421 13783 10424
rect 13725 10415 13783 10421
rect 13814 10412 13820 10424
rect 13872 10412 13878 10464
rect 14366 10452 14372 10464
rect 14327 10424 14372 10452
rect 14366 10412 14372 10424
rect 14424 10412 14430 10464
rect 15838 10412 15844 10464
rect 15896 10452 15902 10464
rect 15933 10455 15991 10461
rect 15933 10452 15945 10455
rect 15896 10424 15945 10452
rect 15896 10412 15902 10424
rect 15933 10421 15945 10424
rect 15979 10421 15991 10455
rect 15933 10415 15991 10421
rect 16669 10455 16727 10461
rect 16669 10421 16681 10455
rect 16715 10452 16727 10455
rect 16942 10452 16948 10464
rect 16715 10424 16948 10452
rect 16715 10421 16727 10424
rect 16669 10415 16727 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 17328 10452 17356 10551
rect 17678 10548 17684 10560
rect 17736 10548 17742 10600
rect 19705 10591 19763 10597
rect 19705 10557 19717 10591
rect 19751 10588 19763 10591
rect 20346 10588 20352 10600
rect 19751 10560 20352 10588
rect 19751 10557 19763 10560
rect 19705 10551 19763 10557
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 21358 10588 21364 10600
rect 21319 10560 21364 10588
rect 21358 10548 21364 10560
rect 21416 10548 21422 10600
rect 19058 10452 19064 10464
rect 17328 10424 19064 10452
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 19886 10412 19892 10464
rect 19944 10452 19950 10464
rect 19981 10455 20039 10461
rect 19981 10452 19993 10455
rect 19944 10424 19993 10452
rect 19944 10412 19950 10424
rect 19981 10421 19993 10424
rect 20027 10421 20039 10455
rect 19981 10415 20039 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 2133 10251 2191 10257
rect 2133 10248 2145 10251
rect 1544 10220 2145 10248
rect 1544 10208 1550 10220
rect 2133 10217 2145 10220
rect 2179 10217 2191 10251
rect 4706 10248 4712 10260
rect 2133 10211 2191 10217
rect 2746 10220 4712 10248
rect 1946 10140 1952 10192
rect 2004 10180 2010 10192
rect 2746 10180 2774 10220
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 4893 10251 4951 10257
rect 4893 10217 4905 10251
rect 4939 10248 4951 10251
rect 5074 10248 5080 10260
rect 4939 10220 5080 10248
rect 4939 10217 4951 10220
rect 4893 10211 4951 10217
rect 5074 10208 5080 10220
rect 5132 10208 5138 10260
rect 5258 10208 5264 10260
rect 5316 10248 5322 10260
rect 5445 10251 5503 10257
rect 5445 10248 5457 10251
rect 5316 10220 5457 10248
rect 5316 10208 5322 10220
rect 5445 10217 5457 10220
rect 5491 10217 5503 10251
rect 5445 10211 5503 10217
rect 6457 10251 6515 10257
rect 6457 10217 6469 10251
rect 6503 10248 6515 10251
rect 6638 10248 6644 10260
rect 6503 10220 6644 10248
rect 6503 10217 6515 10220
rect 6457 10211 6515 10217
rect 6638 10208 6644 10220
rect 6696 10208 6702 10260
rect 8662 10248 8668 10260
rect 6748 10220 8668 10248
rect 2004 10152 2774 10180
rect 3053 10183 3111 10189
rect 2004 10140 2010 10152
rect 3053 10149 3065 10183
rect 3099 10180 3111 10183
rect 4338 10180 4344 10192
rect 3099 10152 4344 10180
rect 3099 10149 3111 10152
rect 3053 10143 3111 10149
rect 4338 10140 4344 10152
rect 4396 10140 4402 10192
rect 6748 10180 6776 10220
rect 8662 10208 8668 10220
rect 8720 10208 8726 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 9766 10248 9772 10260
rect 9272 10220 9444 10248
rect 9727 10220 9772 10248
rect 9272 10208 9278 10220
rect 5276 10152 6776 10180
rect 5276 10124 5304 10152
rect 8110 10140 8116 10192
rect 8168 10180 8174 10192
rect 9416 10180 9444 10220
rect 9766 10208 9772 10220
rect 9824 10208 9830 10260
rect 11422 10248 11428 10260
rect 9876 10220 11008 10248
rect 11383 10220 11428 10248
rect 9876 10180 9904 10220
rect 8168 10152 9352 10180
rect 9416 10152 9904 10180
rect 10980 10180 11008 10220
rect 11422 10208 11428 10220
rect 11480 10208 11486 10260
rect 14274 10208 14280 10260
rect 14332 10248 14338 10260
rect 14332 10220 15516 10248
rect 14332 10208 14338 10220
rect 12066 10180 12072 10192
rect 10980 10152 12072 10180
rect 8168 10140 8174 10152
rect 1854 10112 1860 10124
rect 1815 10084 1860 10112
rect 1854 10072 1860 10084
rect 1912 10072 1918 10124
rect 3878 10112 3884 10124
rect 2746 10084 3884 10112
rect 2317 10047 2375 10053
rect 2317 10013 2329 10047
rect 2363 10044 2375 10047
rect 2746 10044 2774 10084
rect 3878 10072 3884 10084
rect 3936 10072 3942 10124
rect 5258 10072 5264 10124
rect 5316 10072 5322 10124
rect 5994 10112 6000 10124
rect 5955 10084 6000 10112
rect 5994 10072 6000 10084
rect 6052 10072 6058 10124
rect 6638 10072 6644 10124
rect 6696 10112 6702 10124
rect 7009 10115 7067 10121
rect 7009 10112 7021 10115
rect 6696 10084 7021 10112
rect 6696 10072 6702 10084
rect 7009 10081 7021 10084
rect 7055 10112 7067 10115
rect 7282 10112 7288 10124
rect 7055 10084 7288 10112
rect 7055 10081 7067 10084
rect 7009 10075 7067 10081
rect 7282 10072 7288 10084
rect 7340 10112 7346 10124
rect 9324 10121 9352 10152
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 13725 10183 13783 10189
rect 13725 10149 13737 10183
rect 13771 10149 13783 10183
rect 15488 10180 15516 10220
rect 17126 10208 17132 10260
rect 17184 10248 17190 10260
rect 17773 10251 17831 10257
rect 17773 10248 17785 10251
rect 17184 10220 17785 10248
rect 17184 10208 17190 10220
rect 17773 10217 17785 10220
rect 17819 10217 17831 10251
rect 17773 10211 17831 10217
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 19058 10248 19064 10260
rect 18012 10220 19064 10248
rect 18012 10208 18018 10220
rect 19058 10208 19064 10220
rect 19116 10208 19122 10260
rect 19518 10248 19524 10260
rect 19479 10220 19524 10248
rect 19518 10208 19524 10220
rect 19576 10208 19582 10260
rect 18598 10180 18604 10192
rect 15488 10152 18604 10180
rect 13725 10143 13783 10149
rect 8021 10115 8079 10121
rect 8021 10112 8033 10115
rect 7340 10084 8033 10112
rect 7340 10072 7346 10084
rect 8021 10081 8033 10084
rect 8067 10081 8079 10115
rect 8021 10075 8079 10081
rect 9217 10115 9275 10121
rect 9217 10081 9229 10115
rect 9263 10081 9275 10115
rect 9217 10075 9275 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 2363 10016 2774 10044
rect 2869 10047 2927 10053
rect 2363 10013 2375 10016
rect 2317 10007 2375 10013
rect 2869 10013 2881 10047
rect 2915 10013 2927 10047
rect 2869 10007 2927 10013
rect 1670 9976 1676 9988
rect 1631 9948 1676 9976
rect 1670 9936 1676 9948
rect 1728 9976 1734 9988
rect 2774 9976 2780 9988
rect 1728 9948 2780 9976
rect 1728 9936 1734 9948
rect 2774 9936 2780 9948
rect 2832 9936 2838 9988
rect 2884 9976 2912 10007
rect 3418 10004 3424 10056
rect 3476 10044 3482 10056
rect 3789 10047 3847 10053
rect 3789 10044 3801 10047
rect 3476 10016 3801 10044
rect 3476 10004 3482 10016
rect 3789 10013 3801 10016
rect 3835 10013 3847 10047
rect 4706 10044 4712 10056
rect 4667 10016 4712 10044
rect 3789 10007 3847 10013
rect 4706 10004 4712 10016
rect 4764 10004 4770 10056
rect 5534 10004 5540 10056
rect 5592 10044 5598 10056
rect 6917 10047 6975 10053
rect 6917 10044 6929 10047
rect 5592 10016 6929 10044
rect 5592 10004 5598 10016
rect 6917 10013 6929 10016
rect 6963 10013 6975 10047
rect 6917 10007 6975 10013
rect 3510 9976 3516 9988
rect 2884 9948 3516 9976
rect 3510 9936 3516 9948
rect 3568 9976 3574 9988
rect 5350 9976 5356 9988
rect 3568 9948 5356 9976
rect 3568 9936 3574 9948
rect 5350 9936 5356 9948
rect 5408 9936 5414 9988
rect 5905 9979 5963 9985
rect 5905 9945 5917 9979
rect 5951 9976 5963 9979
rect 5951 9948 7512 9976
rect 5951 9945 5963 9948
rect 5905 9939 5963 9945
rect 3421 9911 3479 9917
rect 3421 9877 3433 9911
rect 3467 9908 3479 9911
rect 4062 9908 4068 9920
rect 3467 9880 4068 9908
rect 3467 9877 3479 9880
rect 3421 9871 3479 9877
rect 4062 9868 4068 9880
rect 4120 9868 4126 9920
rect 4430 9908 4436 9920
rect 4391 9880 4436 9908
rect 4430 9868 4436 9880
rect 4488 9868 4494 9920
rect 5813 9911 5871 9917
rect 5813 9877 5825 9911
rect 5859 9908 5871 9911
rect 6730 9908 6736 9920
rect 5859 9880 6736 9908
rect 5859 9877 5871 9880
rect 5813 9871 5871 9877
rect 6730 9868 6736 9880
rect 6788 9868 6794 9920
rect 6822 9868 6828 9920
rect 6880 9908 6886 9920
rect 7484 9917 7512 9948
rect 8018 9936 8024 9988
rect 8076 9976 8082 9988
rect 8481 9979 8539 9985
rect 8481 9976 8493 9979
rect 8076 9948 8493 9976
rect 8076 9936 8082 9948
rect 8481 9945 8493 9948
rect 8527 9945 8539 9979
rect 8481 9939 8539 9945
rect 8938 9936 8944 9988
rect 8996 9976 9002 9988
rect 9232 9976 9260 10075
rect 9582 10072 9588 10124
rect 9640 10112 9646 10124
rect 9766 10112 9772 10124
rect 9640 10084 9772 10112
rect 9640 10072 9646 10084
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 13740 10056 13768 10143
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 19426 10140 19432 10192
rect 19484 10180 19490 10192
rect 19886 10180 19892 10192
rect 19484 10152 19892 10180
rect 19484 10140 19490 10152
rect 19886 10140 19892 10152
rect 19944 10180 19950 10192
rect 19944 10152 20576 10180
rect 19944 10140 19950 10152
rect 20548 10124 20576 10152
rect 16298 10112 16304 10124
rect 15396 10084 16304 10112
rect 9398 10044 9404 10056
rect 9359 10016 9404 10044
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 10045 10047 10103 10053
rect 10045 10013 10057 10047
rect 10091 10044 10103 10047
rect 10134 10044 10140 10056
rect 10091 10016 10140 10044
rect 10091 10013 10103 10016
rect 10045 10007 10103 10013
rect 10134 10004 10140 10016
rect 10192 10004 10198 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 12345 10047 12403 10053
rect 12345 10044 12357 10047
rect 11756 10016 12357 10044
rect 11756 10004 11762 10016
rect 12345 10013 12357 10016
rect 12391 10013 12403 10047
rect 12612 10047 12670 10053
rect 12612 10044 12624 10047
rect 12345 10007 12403 10013
rect 12544 10016 12624 10044
rect 9582 9976 9588 9988
rect 8996 9948 9588 9976
rect 8996 9936 9002 9948
rect 9582 9936 9588 9948
rect 9640 9976 9646 9988
rect 10290 9979 10348 9985
rect 10290 9976 10302 9979
rect 9640 9948 10302 9976
rect 9640 9936 9646 9948
rect 10290 9945 10302 9948
rect 10336 9945 10348 9979
rect 10290 9939 10348 9945
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 12544 9976 12572 10016
rect 12612 10013 12624 10016
rect 12658 10044 12670 10047
rect 13630 10044 13636 10056
rect 12658 10016 13636 10044
rect 12658 10013 12670 10016
rect 12612 10007 12670 10013
rect 13630 10004 13636 10016
rect 13688 10004 13694 10056
rect 13722 10004 13728 10056
rect 13780 10044 13786 10056
rect 15396 10044 15424 10084
rect 16298 10072 16304 10084
rect 16356 10072 16362 10124
rect 16390 10072 16396 10124
rect 16448 10112 16454 10124
rect 17313 10115 17371 10121
rect 17313 10112 17325 10115
rect 16448 10084 17325 10112
rect 16448 10072 16454 10084
rect 17313 10081 17325 10084
rect 17359 10081 17371 10115
rect 17313 10075 17371 10081
rect 18230 10072 18236 10124
rect 18288 10112 18294 10124
rect 18325 10115 18383 10121
rect 18325 10112 18337 10115
rect 18288 10084 18337 10112
rect 18288 10072 18294 10084
rect 18325 10081 18337 10084
rect 18371 10081 18383 10115
rect 20530 10112 20536 10124
rect 20443 10084 20536 10112
rect 18325 10075 18383 10081
rect 20530 10072 20536 10084
rect 20588 10072 20594 10124
rect 20990 10072 20996 10124
rect 21048 10112 21054 10124
rect 21085 10115 21143 10121
rect 21085 10112 21097 10115
rect 21048 10084 21097 10112
rect 21048 10072 21054 10084
rect 21085 10081 21097 10084
rect 21131 10081 21143 10115
rect 21085 10075 21143 10081
rect 13780 10016 15424 10044
rect 15473 10047 15531 10053
rect 13780 10004 13786 10016
rect 15473 10013 15485 10047
rect 15519 10044 15531 10047
rect 17678 10044 17684 10056
rect 15519 10016 17684 10044
rect 15519 10013 15531 10016
rect 15473 10007 15531 10013
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 18877 10047 18935 10053
rect 18877 10044 18889 10047
rect 18156 10016 18889 10044
rect 18156 9988 18184 10016
rect 18877 10013 18889 10016
rect 18923 10013 18935 10047
rect 18877 10007 18935 10013
rect 18966 10004 18972 10056
rect 19024 10044 19030 10056
rect 19613 10047 19671 10053
rect 19613 10044 19625 10047
rect 19024 10016 19625 10044
rect 19024 10004 19030 10016
rect 19613 10013 19625 10016
rect 19659 10013 19671 10047
rect 20346 10044 20352 10056
rect 20307 10016 20352 10044
rect 19613 10007 19671 10013
rect 20346 10004 20352 10016
rect 20404 10004 20410 10056
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 21269 10047 21327 10053
rect 21269 10044 21281 10047
rect 20772 10016 21281 10044
rect 20772 10004 20778 10016
rect 21269 10013 21281 10016
rect 21315 10013 21327 10047
rect 21269 10007 21327 10013
rect 11204 9948 12572 9976
rect 13924 9948 14228 9976
rect 11204 9936 11210 9948
rect 7469 9911 7527 9917
rect 6880 9880 6925 9908
rect 6880 9868 6886 9880
rect 7469 9877 7481 9911
rect 7515 9877 7527 9911
rect 7834 9908 7840 9920
rect 7795 9880 7840 9908
rect 7469 9871 7527 9877
rect 7834 9868 7840 9880
rect 7892 9868 7898 9920
rect 7926 9868 7932 9920
rect 7984 9908 7990 9920
rect 7984 9880 8029 9908
rect 7984 9868 7990 9880
rect 8386 9868 8392 9920
rect 8444 9908 8450 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 8444 9880 11989 9908
rect 8444 9868 8450 9880
rect 11977 9877 11989 9880
rect 12023 9908 12035 9911
rect 13924 9908 13952 9948
rect 14090 9908 14096 9920
rect 12023 9880 13952 9908
rect 14051 9880 14096 9908
rect 12023 9877 12035 9880
rect 11977 9871 12035 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14200 9908 14228 9948
rect 14274 9936 14280 9988
rect 14332 9976 14338 9988
rect 15206 9979 15264 9985
rect 15206 9976 15218 9979
rect 14332 9948 15218 9976
rect 14332 9936 14338 9948
rect 15206 9945 15218 9948
rect 15252 9945 15264 9979
rect 15838 9976 15844 9988
rect 15206 9939 15264 9945
rect 15304 9948 15844 9976
rect 15304 9908 15332 9948
rect 15838 9936 15844 9948
rect 15896 9936 15902 9988
rect 16850 9936 16856 9988
rect 16908 9976 16914 9988
rect 17129 9979 17187 9985
rect 17129 9976 17141 9979
rect 16908 9948 17141 9976
rect 16908 9936 16914 9948
rect 17129 9945 17141 9948
rect 17175 9945 17187 9979
rect 17129 9939 17187 9945
rect 17221 9979 17279 9985
rect 17221 9945 17233 9979
rect 17267 9976 17279 9979
rect 17586 9976 17592 9988
rect 17267 9948 17592 9976
rect 17267 9945 17279 9948
rect 17221 9939 17279 9945
rect 17586 9936 17592 9948
rect 17644 9936 17650 9988
rect 18138 9976 18144 9988
rect 18099 9948 18144 9976
rect 18138 9936 18144 9948
rect 18196 9936 18202 9988
rect 19150 9936 19156 9988
rect 19208 9976 19214 9988
rect 20441 9979 20499 9985
rect 20441 9976 20453 9979
rect 19208 9948 20453 9976
rect 19208 9936 19214 9948
rect 20441 9945 20453 9948
rect 20487 9945 20499 9979
rect 20441 9939 20499 9945
rect 14200 9880 15332 9908
rect 15378 9868 15384 9920
rect 15436 9908 15442 9920
rect 15749 9911 15807 9917
rect 15749 9908 15761 9911
rect 15436 9880 15761 9908
rect 15436 9868 15442 9880
rect 15749 9877 15761 9880
rect 15795 9877 15807 9911
rect 16114 9908 16120 9920
rect 16075 9880 16120 9908
rect 15749 9871 15807 9877
rect 16114 9868 16120 9880
rect 16172 9868 16178 9920
rect 16209 9911 16267 9917
rect 16209 9877 16221 9911
rect 16255 9908 16267 9911
rect 16761 9911 16819 9917
rect 16761 9908 16773 9911
rect 16255 9880 16773 9908
rect 16255 9877 16267 9880
rect 16209 9871 16267 9877
rect 16761 9877 16773 9880
rect 16807 9877 16819 9911
rect 16761 9871 16819 9877
rect 17770 9868 17776 9920
rect 17828 9908 17834 9920
rect 18233 9911 18291 9917
rect 18233 9908 18245 9911
rect 17828 9880 18245 9908
rect 17828 9868 17834 9880
rect 18233 9877 18245 9880
rect 18279 9877 18291 9911
rect 18233 9871 18291 9877
rect 19702 9868 19708 9920
rect 19760 9908 19766 9920
rect 19981 9911 20039 9917
rect 19981 9908 19993 9911
rect 19760 9880 19993 9908
rect 19760 9868 19766 9880
rect 19981 9877 19993 9880
rect 20027 9877 20039 9911
rect 19981 9871 20039 9877
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 2866 9704 2872 9716
rect 1964 9676 2872 9704
rect 1578 9568 1584 9580
rect 1539 9540 1584 9568
rect 1578 9528 1584 9540
rect 1636 9568 1642 9580
rect 1964 9568 1992 9676
rect 2866 9664 2872 9676
rect 2924 9664 2930 9716
rect 3050 9704 3056 9716
rect 2976 9676 3056 9704
rect 2222 9596 2228 9648
rect 2280 9596 2286 9648
rect 2976 9636 3004 9676
rect 3050 9664 3056 9676
rect 3108 9664 3114 9716
rect 3326 9664 3332 9716
rect 3384 9704 3390 9716
rect 6822 9704 6828 9716
rect 3384 9676 6828 9704
rect 3384 9664 3390 9676
rect 6822 9664 6828 9676
rect 6880 9664 6886 9716
rect 8665 9707 8723 9713
rect 8665 9673 8677 9707
rect 8711 9673 8723 9707
rect 8938 9704 8944 9716
rect 8899 9676 8944 9704
rect 8665 9667 8723 9673
rect 2746 9608 3004 9636
rect 4240 9639 4298 9645
rect 1636 9540 1992 9568
rect 2041 9571 2099 9577
rect 1636 9528 1642 9540
rect 2041 9537 2053 9571
rect 2087 9568 2099 9571
rect 2240 9568 2268 9596
rect 2746 9580 2774 9608
rect 4240 9605 4252 9639
rect 4286 9636 4298 9639
rect 4430 9636 4436 9648
rect 4286 9608 4436 9636
rect 4286 9605 4298 9608
rect 4240 9599 4298 9605
rect 4430 9596 4436 9608
rect 4488 9596 4494 9648
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 8205 9639 8263 9645
rect 8205 9636 8217 9639
rect 6972 9608 8217 9636
rect 6972 9596 6978 9608
rect 8205 9605 8217 9608
rect 8251 9605 8263 9639
rect 8680 9636 8708 9667
rect 8938 9664 8944 9676
rect 8996 9664 9002 9716
rect 10594 9664 10600 9716
rect 10652 9704 10658 9716
rect 10870 9704 10876 9716
rect 10652 9676 10876 9704
rect 10652 9664 10658 9676
rect 10870 9664 10876 9676
rect 10928 9664 10934 9716
rect 14093 9707 14151 9713
rect 14093 9673 14105 9707
rect 14139 9704 14151 9707
rect 14274 9704 14280 9716
rect 14139 9676 14280 9704
rect 14139 9673 14151 9676
rect 14093 9667 14151 9673
rect 14274 9664 14280 9676
rect 14332 9664 14338 9716
rect 14366 9664 14372 9716
rect 14424 9704 14430 9716
rect 14737 9707 14795 9713
rect 14737 9704 14749 9707
rect 14424 9676 14749 9704
rect 14424 9664 14430 9676
rect 14737 9673 14749 9676
rect 14783 9673 14795 9707
rect 14737 9667 14795 9673
rect 15654 9664 15660 9716
rect 15712 9704 15718 9716
rect 15749 9707 15807 9713
rect 15749 9704 15761 9707
rect 15712 9676 15761 9704
rect 15712 9664 15718 9676
rect 15749 9673 15761 9676
rect 15795 9673 15807 9707
rect 15749 9667 15807 9673
rect 15838 9664 15844 9716
rect 15896 9704 15902 9716
rect 18141 9707 18199 9713
rect 15896 9676 18092 9704
rect 15896 9664 15902 9676
rect 14645 9639 14703 9645
rect 8680 9608 14320 9636
rect 8205 9599 8263 9605
rect 2087 9540 2268 9568
rect 2308 9571 2366 9577
rect 2087 9537 2099 9540
rect 2041 9531 2099 9537
rect 2308 9537 2320 9571
rect 2354 9568 2366 9571
rect 2590 9568 2596 9580
rect 2354 9540 2596 9568
rect 2354 9537 2366 9540
rect 2308 9531 2366 9537
rect 2590 9528 2596 9540
rect 2648 9528 2654 9580
rect 2682 9528 2688 9580
rect 2740 9540 2774 9580
rect 3973 9571 4031 9577
rect 2740 9528 2746 9540
rect 3973 9537 3985 9571
rect 4019 9568 4031 9571
rect 4614 9568 4620 9580
rect 4019 9540 4620 9568
rect 4019 9537 4031 9540
rect 3973 9531 4031 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 5902 9568 5908 9580
rect 5132 9540 5908 9568
rect 5132 9528 5138 9540
rect 5902 9528 5908 9540
rect 5960 9568 5966 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 5960 9540 6377 9568
rect 5960 9528 5966 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6365 9531 6423 9537
rect 7006 9528 7012 9580
rect 7064 9568 7070 9580
rect 7285 9571 7343 9577
rect 7285 9568 7297 9571
rect 7064 9540 7297 9568
rect 7064 9528 7070 9540
rect 7285 9537 7297 9540
rect 7331 9537 7343 9571
rect 7285 9531 7343 9537
rect 7558 9528 7564 9580
rect 7616 9568 7622 9580
rect 8297 9571 8355 9577
rect 8297 9568 8309 9571
rect 7616 9540 8309 9568
rect 7616 9528 7622 9540
rect 8297 9537 8309 9540
rect 8343 9537 8355 9571
rect 8297 9531 8355 9537
rect 10065 9571 10123 9577
rect 10065 9537 10077 9571
rect 10111 9568 10123 9571
rect 10226 9568 10232 9580
rect 10111 9540 10232 9568
rect 10111 9537 10123 9540
rect 10065 9531 10123 9537
rect 10226 9528 10232 9540
rect 10284 9528 10290 9580
rect 10594 9528 10600 9580
rect 10652 9568 10658 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10652 9540 10701 9568
rect 10652 9528 10658 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 11698 9568 11704 9580
rect 11659 9540 11704 9568
rect 10689 9531 10747 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 11974 9577 11980 9580
rect 11968 9531 11980 9577
rect 12032 9568 12038 9580
rect 13449 9571 13507 9577
rect 12032 9540 12068 9568
rect 11974 9528 11980 9531
rect 12032 9528 12038 9540
rect 13449 9537 13461 9571
rect 13495 9568 13507 9571
rect 13722 9568 13728 9580
rect 13495 9540 13728 9568
rect 13495 9537 13507 9540
rect 13449 9531 13507 9537
rect 13722 9528 13728 9540
rect 13780 9528 13786 9580
rect 14292 9568 14320 9608
rect 14645 9605 14657 9639
rect 14691 9636 14703 9639
rect 15378 9636 15384 9648
rect 14691 9608 15384 9636
rect 14691 9605 14703 9608
rect 14645 9599 14703 9605
rect 15378 9596 15384 9608
rect 15436 9596 15442 9648
rect 17678 9636 17684 9648
rect 16776 9608 17684 9636
rect 16776 9580 16804 9608
rect 17678 9596 17684 9608
rect 17736 9596 17742 9648
rect 18064 9636 18092 9676
rect 18141 9673 18153 9707
rect 18187 9704 18199 9707
rect 18230 9704 18236 9716
rect 18187 9676 18236 9704
rect 18187 9673 18199 9676
rect 18141 9667 18199 9673
rect 18230 9664 18236 9676
rect 18288 9664 18294 9716
rect 18782 9704 18788 9716
rect 18616 9676 18788 9704
rect 18616 9636 18644 9676
rect 18782 9664 18788 9676
rect 18840 9704 18846 9716
rect 19150 9704 19156 9716
rect 18840 9676 19156 9704
rect 18840 9664 18846 9676
rect 19150 9664 19156 9676
rect 19208 9664 19214 9716
rect 18064 9608 18644 9636
rect 19245 9639 19303 9645
rect 19245 9605 19257 9639
rect 19291 9636 19303 9639
rect 20254 9636 20260 9648
rect 19291 9608 20260 9636
rect 19291 9605 19303 9608
rect 19245 9599 19303 9605
rect 20254 9596 20260 9608
rect 20312 9596 20318 9648
rect 16114 9568 16120 9580
rect 14292 9540 16120 9568
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 16758 9568 16764 9580
rect 16671 9540 16764 9568
rect 16758 9528 16764 9540
rect 16816 9528 16822 9580
rect 17028 9571 17086 9577
rect 17028 9537 17040 9571
rect 17074 9568 17086 9571
rect 18506 9568 18512 9580
rect 17074 9540 18512 9568
rect 17074 9537 17086 9540
rect 17028 9531 17086 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 19337 9571 19395 9577
rect 19337 9568 19349 9571
rect 18656 9540 18701 9568
rect 18800 9540 19349 9568
rect 18656 9528 18662 9540
rect 4982 9460 4988 9512
rect 5040 9500 5046 9512
rect 5629 9503 5687 9509
rect 5629 9500 5641 9503
rect 5040 9472 5641 9500
rect 5040 9460 5046 9472
rect 5629 9469 5641 9472
rect 5675 9469 5687 9503
rect 7374 9500 7380 9512
rect 7335 9472 7380 9500
rect 5629 9463 5687 9469
rect 7374 9460 7380 9472
rect 7432 9460 7438 9512
rect 7469 9503 7527 9509
rect 7469 9469 7481 9503
rect 7515 9469 7527 9503
rect 7469 9463 7527 9469
rect 8113 9503 8171 9509
rect 8113 9469 8125 9503
rect 8159 9469 8171 9503
rect 10318 9500 10324 9512
rect 10279 9472 10324 9500
rect 8113 9463 8171 9469
rect 6546 9432 6552 9444
rect 6507 9404 6552 9432
rect 6546 9392 6552 9404
rect 6604 9392 6610 9444
rect 6730 9392 6736 9444
rect 6788 9432 6794 9444
rect 6917 9435 6975 9441
rect 6917 9432 6929 9435
rect 6788 9404 6929 9432
rect 6788 9392 6794 9404
rect 6917 9401 6929 9404
rect 6963 9401 6975 9435
rect 6917 9395 6975 9401
rect 1673 9367 1731 9373
rect 1673 9333 1685 9367
rect 1719 9364 1731 9367
rect 3234 9364 3240 9376
rect 1719 9336 3240 9364
rect 1719 9333 1731 9336
rect 1673 9327 1731 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 3418 9364 3424 9376
rect 3379 9336 3424 9364
rect 3418 9324 3424 9336
rect 3476 9324 3482 9376
rect 5350 9364 5356 9376
rect 5311 9336 5356 9364
rect 5350 9324 5356 9336
rect 5408 9324 5414 9376
rect 6638 9324 6644 9376
rect 6696 9364 6702 9376
rect 7484 9364 7512 9463
rect 8128 9432 8156 9463
rect 10318 9460 10324 9472
rect 10376 9460 10382 9512
rect 11146 9500 11152 9512
rect 11072 9472 11152 9500
rect 8128 9404 9444 9432
rect 6696 9336 7512 9364
rect 9416 9364 9444 9404
rect 11072 9364 11100 9472
rect 11146 9460 11152 9472
rect 11204 9460 11210 9512
rect 14090 9460 14096 9512
rect 14148 9500 14154 9512
rect 14274 9500 14280 9512
rect 14148 9472 14280 9500
rect 14148 9460 14154 9472
rect 14274 9460 14280 9472
rect 14332 9500 14338 9512
rect 14461 9503 14519 9509
rect 14461 9500 14473 9503
rect 14332 9472 14473 9500
rect 14332 9460 14338 9472
rect 14461 9469 14473 9472
rect 14507 9469 14519 9503
rect 14461 9463 14519 9469
rect 16025 9503 16083 9509
rect 16025 9469 16037 9503
rect 16071 9500 16083 9503
rect 16390 9500 16396 9512
rect 16071 9472 16396 9500
rect 16071 9469 16083 9472
rect 16025 9463 16083 9469
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 17770 9460 17776 9512
rect 17828 9500 17834 9512
rect 18800 9500 18828 9540
rect 19337 9537 19349 9540
rect 19383 9537 19395 9571
rect 19337 9531 19395 9537
rect 17828 9472 18828 9500
rect 19153 9503 19211 9509
rect 17828 9460 17834 9472
rect 19153 9469 19165 9503
rect 19199 9469 19211 9503
rect 19352 9500 19380 9531
rect 19518 9528 19524 9580
rect 19576 9568 19582 9580
rect 19794 9568 19800 9580
rect 19576 9540 19800 9568
rect 19576 9528 19582 9540
rect 19794 9528 19800 9540
rect 19852 9528 19858 9580
rect 20530 9528 20536 9580
rect 20588 9568 20594 9580
rect 21094 9571 21152 9577
rect 21094 9568 21106 9571
rect 20588 9540 21106 9568
rect 20588 9528 20594 9540
rect 21094 9537 21106 9540
rect 21140 9537 21152 9571
rect 21094 9531 21152 9537
rect 21358 9500 21364 9512
rect 19352 9472 20392 9500
rect 21319 9472 21364 9500
rect 19153 9463 19211 9469
rect 13354 9432 13360 9444
rect 12912 9404 13360 9432
rect 9416 9336 11100 9364
rect 11149 9367 11207 9373
rect 6696 9324 6702 9336
rect 11149 9333 11161 9367
rect 11195 9364 11207 9367
rect 12912 9364 12940 9404
rect 13354 9392 13360 9404
rect 13412 9392 13418 9444
rect 14642 9392 14648 9444
rect 14700 9432 14706 9444
rect 15105 9435 15163 9441
rect 15105 9432 15117 9435
rect 14700 9404 15117 9432
rect 14700 9392 14706 9404
rect 15105 9401 15117 9404
rect 15151 9401 15163 9435
rect 15105 9395 15163 9401
rect 15286 9392 15292 9444
rect 15344 9432 15350 9444
rect 15381 9435 15439 9441
rect 15381 9432 15393 9435
rect 15344 9404 15393 9432
rect 15344 9392 15350 9404
rect 15381 9401 15393 9404
rect 15427 9401 15439 9435
rect 15381 9395 15439 9401
rect 18046 9392 18052 9444
rect 18104 9432 18110 9444
rect 18417 9435 18475 9441
rect 18417 9432 18429 9435
rect 18104 9404 18429 9432
rect 18104 9392 18110 9404
rect 18417 9401 18429 9404
rect 18463 9401 18475 9435
rect 19168 9432 19196 9463
rect 19426 9432 19432 9444
rect 19168 9404 19432 9432
rect 18417 9395 18475 9401
rect 19426 9392 19432 9404
rect 19484 9392 19490 9444
rect 13078 9364 13084 9376
rect 11195 9336 12940 9364
rect 12991 9336 13084 9364
rect 11195 9333 11207 9336
rect 11149 9327 11207 9333
rect 13078 9324 13084 9336
rect 13136 9364 13142 9376
rect 13722 9364 13728 9376
rect 13136 9336 13728 9364
rect 13136 9324 13142 9336
rect 13722 9324 13728 9336
rect 13780 9324 13786 9376
rect 15470 9324 15476 9376
rect 15528 9364 15534 9376
rect 15930 9364 15936 9376
rect 15528 9336 15936 9364
rect 15528 9324 15534 9336
rect 15930 9324 15936 9336
rect 15988 9364 15994 9376
rect 17954 9364 17960 9376
rect 15988 9336 17960 9364
rect 15988 9324 15994 9336
rect 17954 9324 17960 9336
rect 18012 9324 18018 9376
rect 19705 9367 19763 9373
rect 19705 9333 19717 9367
rect 19751 9364 19763 9367
rect 19794 9364 19800 9376
rect 19751 9336 19800 9364
rect 19751 9333 19763 9336
rect 19705 9327 19763 9333
rect 19794 9324 19800 9336
rect 19852 9324 19858 9376
rect 19978 9364 19984 9376
rect 19939 9336 19984 9364
rect 19978 9324 19984 9336
rect 20036 9324 20042 9376
rect 20364 9364 20392 9472
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 20438 9364 20444 9376
rect 20364 9336 20444 9364
rect 20438 9324 20444 9336
rect 20496 9324 20502 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 3053 9163 3111 9169
rect 3053 9129 3065 9163
rect 3099 9160 3111 9163
rect 4706 9160 4712 9172
rect 3099 9132 4712 9160
rect 3099 9129 3111 9132
rect 3053 9123 3111 9129
rect 4706 9120 4712 9132
rect 4764 9120 4770 9172
rect 6638 9160 6644 9172
rect 6599 9132 6644 9160
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7653 9163 7711 9169
rect 7653 9129 7665 9163
rect 7699 9160 7711 9163
rect 7834 9160 7840 9172
rect 7699 9132 7840 9160
rect 7699 9129 7711 9132
rect 7653 9123 7711 9129
rect 7834 9120 7840 9132
rect 7892 9120 7898 9172
rect 10505 9163 10563 9169
rect 10505 9129 10517 9163
rect 10551 9160 10563 9163
rect 10686 9160 10692 9172
rect 10551 9132 10692 9160
rect 10551 9129 10563 9132
rect 10505 9123 10563 9129
rect 10686 9120 10692 9132
rect 10744 9120 10750 9172
rect 11146 9160 11152 9172
rect 11107 9132 11152 9160
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11974 9120 11980 9172
rect 12032 9160 12038 9172
rect 12069 9163 12127 9169
rect 12069 9160 12081 9163
rect 12032 9132 12081 9160
rect 12032 9120 12038 9132
rect 12069 9129 12081 9132
rect 12115 9129 12127 9163
rect 12069 9123 12127 9129
rect 15930 9120 15936 9172
rect 15988 9160 15994 9172
rect 15988 9132 17080 9160
rect 15988 9120 15994 9132
rect 2038 9052 2044 9104
rect 2096 9092 2102 9104
rect 4982 9092 4988 9104
rect 2096 9064 4988 9092
rect 2096 9052 2102 9064
rect 4982 9052 4988 9064
rect 5040 9052 5046 9104
rect 6546 9052 6552 9104
rect 6604 9092 6610 9104
rect 8297 9095 8355 9101
rect 8297 9092 8309 9095
rect 6604 9064 8309 9092
rect 6604 9052 6610 9064
rect 8297 9061 8309 9064
rect 8343 9061 8355 9095
rect 8297 9055 8355 9061
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 12894 9092 12900 9104
rect 10652 9064 12900 9092
rect 10652 9052 10658 9064
rect 12894 9052 12900 9064
rect 12952 9052 12958 9104
rect 2501 9027 2559 9033
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 3418 9024 3424 9036
rect 2547 8996 3424 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 4522 9024 4528 9036
rect 4483 8996 4528 9024
rect 4522 8984 4528 8996
rect 4580 8984 4586 9036
rect 4706 9024 4712 9036
rect 4667 8996 4712 9024
rect 4706 8984 4712 8996
rect 4764 8984 4770 9036
rect 7009 9027 7067 9033
rect 7009 8993 7021 9027
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 3142 8956 3148 8968
rect 1688 8928 3148 8956
rect 1688 8900 1716 8928
rect 3142 8916 3148 8928
rect 3200 8916 3206 8968
rect 4614 8916 4620 8968
rect 4672 8956 4678 8968
rect 5166 8956 5172 8968
rect 4672 8928 5172 8956
rect 4672 8916 4678 8928
rect 5166 8916 5172 8928
rect 5224 8956 5230 8968
rect 5261 8959 5319 8965
rect 5261 8956 5273 8959
rect 5224 8928 5273 8956
rect 5224 8916 5230 8928
rect 5261 8925 5273 8928
rect 5307 8925 5319 8959
rect 5261 8919 5319 8925
rect 5350 8916 5356 8968
rect 5408 8956 5414 8968
rect 5517 8959 5575 8965
rect 5517 8956 5529 8959
rect 5408 8928 5529 8956
rect 5408 8916 5414 8928
rect 5517 8925 5529 8928
rect 5563 8956 5575 8959
rect 7024 8956 7052 8987
rect 9582 8984 9588 9036
rect 9640 9024 9646 9036
rect 9861 9027 9919 9033
rect 9861 9024 9873 9027
rect 9640 8996 9873 9024
rect 9640 8984 9646 8996
rect 9861 8993 9873 8996
rect 9907 8993 9919 9027
rect 9861 8987 9919 8993
rect 9968 8996 11560 9024
rect 5563 8928 7052 8956
rect 5563 8925 5575 8928
rect 5517 8919 5575 8925
rect 7098 8916 7104 8968
rect 7156 8956 7162 8968
rect 7285 8959 7343 8965
rect 7285 8956 7297 8959
rect 7156 8928 7297 8956
rect 7156 8916 7162 8928
rect 7285 8925 7297 8928
rect 7331 8956 7343 8959
rect 7558 8956 7564 8968
rect 7331 8928 7564 8956
rect 7331 8925 7343 8928
rect 7285 8919 7343 8925
rect 7558 8916 7564 8928
rect 7616 8916 7622 8968
rect 1670 8888 1676 8900
rect 1631 8860 1676 8888
rect 1670 8848 1676 8860
rect 1728 8848 1734 8900
rect 1854 8888 1860 8900
rect 1815 8860 1860 8888
rect 1854 8848 1860 8860
rect 1912 8848 1918 8900
rect 2590 8888 2596 8900
rect 2551 8860 2596 8888
rect 2590 8848 2596 8860
rect 2648 8848 2654 8900
rect 3234 8848 3240 8900
rect 3292 8888 3298 8900
rect 9968 8888 9996 8996
rect 10042 8916 10048 8968
rect 10100 8956 10106 8968
rect 10100 8928 10145 8956
rect 10100 8916 10106 8928
rect 11238 8916 11244 8968
rect 11296 8956 11302 8968
rect 11425 8959 11483 8965
rect 11425 8956 11437 8959
rect 11296 8928 11437 8956
rect 11296 8916 11302 8928
rect 11425 8925 11437 8928
rect 11471 8925 11483 8959
rect 11532 8956 11560 8996
rect 12434 8984 12440 9036
rect 12492 9024 12498 9036
rect 13630 9024 13636 9036
rect 12492 8996 13636 9024
rect 12492 8984 12498 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 12986 8956 12992 8968
rect 11532 8928 12992 8956
rect 11425 8919 11483 8925
rect 12986 8916 12992 8928
rect 13044 8956 13050 8968
rect 13446 8956 13452 8968
rect 13044 8928 13452 8956
rect 13044 8916 13050 8928
rect 13446 8916 13452 8928
rect 13504 8916 13510 8968
rect 14185 8959 14243 8965
rect 14185 8925 14197 8959
rect 14231 8956 14243 8959
rect 14274 8956 14280 8968
rect 14231 8928 14280 8956
rect 14231 8925 14243 8928
rect 14185 8919 14243 8925
rect 14274 8916 14280 8928
rect 14332 8916 14338 8968
rect 15470 8956 15476 8968
rect 15431 8928 15476 8956
rect 15470 8916 15476 8928
rect 15528 8916 15534 8968
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 16758 8956 16764 8968
rect 15795 8928 16764 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16758 8916 16764 8928
rect 16816 8916 16822 8968
rect 17052 8956 17080 9132
rect 18506 9120 18512 9172
rect 18564 9160 18570 9172
rect 20993 9163 21051 9169
rect 20993 9160 21005 9163
rect 18564 9132 21005 9160
rect 18564 9120 18570 9132
rect 20993 9129 21005 9132
rect 21039 9129 21051 9163
rect 20993 9123 21051 9129
rect 17129 9095 17187 9101
rect 17129 9061 17141 9095
rect 17175 9092 17187 9095
rect 18874 9092 18880 9104
rect 17175 9064 18880 9092
rect 17175 9061 17187 9064
rect 17129 9055 17187 9061
rect 18874 9052 18880 9064
rect 18932 9052 18938 9104
rect 19337 9095 19395 9101
rect 19337 9061 19349 9095
rect 19383 9061 19395 9095
rect 19337 9055 19395 9061
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 19352 9024 19380 9055
rect 19794 9024 19800 9036
rect 17552 8996 19380 9024
rect 19755 8996 19800 9024
rect 17552 8984 17558 8996
rect 19794 8984 19800 8996
rect 19852 8984 19858 9036
rect 19978 8984 19984 9036
rect 20036 9024 20042 9036
rect 20530 9024 20536 9036
rect 20036 8996 20536 9024
rect 20036 8984 20042 8996
rect 20530 8984 20536 8996
rect 20588 8984 20594 9036
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17052 8928 17417 8956
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 17586 8916 17592 8968
rect 17644 8956 17650 8968
rect 18601 8959 18659 8965
rect 18601 8956 18613 8959
rect 17644 8928 18613 8956
rect 17644 8916 17650 8928
rect 18601 8925 18613 8928
rect 18647 8925 18659 8959
rect 19702 8956 19708 8968
rect 19663 8928 19708 8956
rect 18601 8919 18659 8925
rect 19702 8916 19708 8928
rect 19760 8916 19766 8968
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8925 20407 8959
rect 20349 8919 20407 8925
rect 10137 8891 10195 8897
rect 10137 8888 10149 8891
rect 3292 8860 9996 8888
rect 10060 8860 10149 8888
rect 3292 8848 3298 8860
rect 2682 8820 2688 8832
rect 2643 8792 2688 8820
rect 2682 8780 2688 8792
rect 2740 8780 2746 8832
rect 2774 8780 2780 8832
rect 2832 8820 2838 8832
rect 2958 8820 2964 8832
rect 2832 8792 2964 8820
rect 2832 8780 2838 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3142 8780 3148 8832
rect 3200 8820 3206 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3200 8792 3341 8820
rect 3200 8780 3206 8792
rect 3329 8789 3341 8792
rect 3375 8820 3387 8823
rect 3786 8820 3792 8832
rect 3375 8792 3792 8820
rect 3375 8789 3387 8792
rect 3329 8783 3387 8789
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 3970 8780 3976 8832
rect 4028 8820 4034 8832
rect 4065 8823 4123 8829
rect 4065 8820 4077 8823
rect 4028 8792 4077 8820
rect 4028 8780 4034 8792
rect 4065 8789 4077 8792
rect 4111 8789 4123 8823
rect 4065 8783 4123 8789
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 5718 8820 5724 8832
rect 4479 8792 5724 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 5718 8780 5724 8792
rect 5776 8820 5782 8832
rect 6822 8820 6828 8832
rect 5776 8792 6828 8820
rect 5776 8780 5782 8792
rect 6822 8780 6828 8792
rect 6880 8780 6886 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 6972 8792 7205 8820
rect 6972 8780 6978 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 8021 8823 8079 8829
rect 8021 8789 8033 8823
rect 8067 8820 8079 8823
rect 8110 8820 8116 8832
rect 8067 8792 8116 8820
rect 8067 8789 8079 8792
rect 8021 8783 8079 8789
rect 8110 8780 8116 8792
rect 8168 8780 8174 8832
rect 8570 8780 8576 8832
rect 8628 8820 8634 8832
rect 8941 8823 8999 8829
rect 8941 8820 8953 8823
rect 8628 8792 8953 8820
rect 8628 8780 8634 8792
rect 8941 8789 8953 8792
rect 8987 8789 8999 8823
rect 9398 8820 9404 8832
rect 9359 8792 9404 8820
rect 8941 8783 8999 8789
rect 9398 8780 9404 8792
rect 9456 8820 9462 8832
rect 10060 8820 10088 8860
rect 10137 8857 10149 8860
rect 10183 8857 10195 8891
rect 10137 8851 10195 8857
rect 16016 8891 16074 8897
rect 16016 8857 16028 8891
rect 16062 8888 16074 8891
rect 16390 8888 16396 8900
rect 16062 8860 16396 8888
rect 16062 8857 16074 8860
rect 16016 8851 16074 8857
rect 9456 8792 10088 8820
rect 10152 8820 10180 8851
rect 16390 8848 16396 8860
rect 16448 8848 16454 8900
rect 17770 8848 17776 8900
rect 17828 8888 17834 8900
rect 18782 8888 18788 8900
rect 17828 8860 18788 8888
rect 17828 8848 17834 8860
rect 18782 8848 18788 8860
rect 18840 8848 18846 8900
rect 18874 8848 18880 8900
rect 18932 8888 18938 8900
rect 20364 8888 20392 8919
rect 18932 8860 20392 8888
rect 18932 8848 18938 8860
rect 12158 8820 12164 8832
rect 10152 8792 12164 8820
rect 9456 8780 9462 8792
rect 12158 8780 12164 8792
rect 12216 8780 12222 8832
rect 12710 8820 12716 8832
rect 12671 8792 12716 8820
rect 12710 8780 12716 8792
rect 12768 8780 12774 8832
rect 13081 8823 13139 8829
rect 13081 8789 13093 8823
rect 13127 8820 13139 8823
rect 13446 8820 13452 8832
rect 13127 8792 13452 8820
rect 13127 8789 13139 8792
rect 13081 8783 13139 8789
rect 13446 8780 13452 8792
rect 13504 8780 13510 8832
rect 13630 8820 13636 8832
rect 13591 8792 13636 8820
rect 13630 8780 13636 8792
rect 13688 8780 13694 8832
rect 14826 8820 14832 8832
rect 14787 8792 14832 8820
rect 14826 8780 14832 8792
rect 14884 8780 14890 8832
rect 15286 8820 15292 8832
rect 15247 8792 15292 8820
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 17586 8780 17592 8832
rect 17644 8820 17650 8832
rect 18049 8823 18107 8829
rect 18049 8820 18061 8823
rect 17644 8792 18061 8820
rect 17644 8780 17650 8792
rect 18049 8789 18061 8792
rect 18095 8789 18107 8823
rect 18049 8783 18107 8789
rect 20898 8780 20904 8832
rect 20956 8820 20962 8832
rect 21361 8823 21419 8829
rect 21361 8820 21373 8823
rect 20956 8792 21373 8820
rect 20956 8780 20962 8792
rect 21361 8789 21373 8792
rect 21407 8820 21419 8823
rect 21450 8820 21456 8832
rect 21407 8792 21456 8820
rect 21407 8789 21419 8792
rect 21361 8783 21419 8789
rect 21450 8780 21456 8792
rect 21508 8780 21514 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 1949 8619 2007 8625
rect 1949 8585 1961 8619
rect 1995 8616 2007 8619
rect 2498 8616 2504 8628
rect 1995 8588 2504 8616
rect 1995 8585 2007 8588
rect 1949 8579 2007 8585
rect 2498 8576 2504 8588
rect 2556 8576 2562 8628
rect 2590 8576 2596 8628
rect 2648 8616 2654 8628
rect 3605 8619 3663 8625
rect 3605 8616 3617 8619
rect 2648 8588 3617 8616
rect 2648 8576 2654 8588
rect 3605 8585 3617 8588
rect 3651 8585 3663 8619
rect 3970 8616 3976 8628
rect 3931 8588 3976 8616
rect 3605 8579 3663 8585
rect 3970 8576 3976 8588
rect 4028 8576 4034 8628
rect 4062 8576 4068 8628
rect 4120 8616 4126 8628
rect 4120 8588 4844 8616
rect 4120 8576 4126 8588
rect 2516 8548 2544 8576
rect 2516 8520 3740 8548
rect 1486 8480 1492 8492
rect 1447 8452 1492 8480
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 1946 8480 1952 8492
rect 1719 8452 1952 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 1946 8440 1952 8452
rect 2004 8440 2010 8492
rect 3073 8483 3131 8489
rect 3073 8449 3085 8483
rect 3119 8480 3131 8483
rect 3234 8480 3240 8492
rect 3119 8452 3240 8480
rect 3119 8449 3131 8452
rect 3073 8443 3131 8449
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3712 8480 3740 8520
rect 3786 8508 3792 8560
rect 3844 8548 3850 8560
rect 4816 8548 4844 8588
rect 4890 8576 4896 8628
rect 4948 8616 4954 8628
rect 5261 8619 5319 8625
rect 5261 8616 5273 8619
rect 4948 8588 5273 8616
rect 4948 8576 4954 8588
rect 5261 8585 5273 8588
rect 5307 8585 5319 8619
rect 5261 8579 5319 8585
rect 6549 8619 6607 8625
rect 6549 8585 6561 8619
rect 6595 8616 6607 8619
rect 7098 8616 7104 8628
rect 6595 8588 7104 8616
rect 6595 8585 6607 8588
rect 6549 8579 6607 8585
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7561 8619 7619 8625
rect 7561 8585 7573 8619
rect 7607 8616 7619 8619
rect 7926 8616 7932 8628
rect 7607 8588 7932 8616
rect 7607 8585 7619 8588
rect 7561 8579 7619 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 9033 8619 9091 8625
rect 9033 8585 9045 8619
rect 9079 8616 9091 8619
rect 9766 8616 9772 8628
rect 9079 8588 9772 8616
rect 9079 8585 9091 8588
rect 9033 8579 9091 8585
rect 9766 8576 9772 8588
rect 9824 8576 9830 8628
rect 10042 8576 10048 8628
rect 10100 8616 10106 8628
rect 10137 8619 10195 8625
rect 10137 8616 10149 8619
rect 10100 8588 10149 8616
rect 10100 8576 10106 8588
rect 10137 8585 10149 8588
rect 10183 8585 10195 8619
rect 18506 8616 18512 8628
rect 10137 8579 10195 8585
rect 14568 8588 18512 8616
rect 6914 8548 6920 8560
rect 3844 8520 4292 8548
rect 4816 8520 6920 8548
rect 3844 8508 3850 8520
rect 4264 8480 4292 8520
rect 6914 8508 6920 8520
rect 6972 8508 6978 8560
rect 7193 8551 7251 8557
rect 7193 8517 7205 8551
rect 7239 8548 7251 8551
rect 8665 8551 8723 8557
rect 8665 8548 8677 8551
rect 7239 8520 8677 8548
rect 7239 8517 7251 8520
rect 7193 8511 7251 8517
rect 8665 8517 8677 8520
rect 8711 8548 8723 8551
rect 9674 8548 9680 8560
rect 8711 8520 9680 8548
rect 8711 8517 8723 8520
rect 8665 8511 8723 8517
rect 9674 8508 9680 8520
rect 9732 8508 9738 8560
rect 3712 8452 4200 8480
rect 4264 8452 4844 8480
rect 3329 8415 3387 8421
rect 3329 8381 3341 8415
rect 3375 8412 3387 8415
rect 3418 8412 3424 8424
rect 3375 8384 3424 8412
rect 3375 8381 3387 8384
rect 3329 8375 3387 8381
rect 3418 8372 3424 8384
rect 3476 8412 3482 8424
rect 4062 8412 4068 8424
rect 3476 8384 3924 8412
rect 4023 8384 4068 8412
rect 3476 8372 3482 8384
rect 3050 8236 3056 8288
rect 3108 8276 3114 8288
rect 3326 8276 3332 8288
rect 3108 8248 3332 8276
rect 3108 8236 3114 8248
rect 3326 8236 3332 8248
rect 3384 8236 3390 8288
rect 3896 8276 3924 8384
rect 4062 8372 4068 8384
rect 4120 8372 4126 8424
rect 4172 8421 4200 8452
rect 4157 8415 4215 8421
rect 4157 8381 4169 8415
rect 4203 8381 4215 8415
rect 4157 8375 4215 8381
rect 4430 8372 4436 8424
rect 4488 8412 4494 8424
rect 4617 8415 4675 8421
rect 4617 8412 4629 8415
rect 4488 8384 4629 8412
rect 4488 8372 4494 8384
rect 4617 8381 4629 8384
rect 4663 8381 4675 8415
rect 4816 8412 4844 8452
rect 4890 8440 4896 8492
rect 4948 8480 4954 8492
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4948 8452 5089 8480
rect 4948 8440 4954 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5537 8483 5595 8489
rect 5537 8449 5549 8483
rect 5583 8449 5595 8483
rect 6362 8480 6368 8492
rect 6323 8452 6368 8480
rect 5537 8443 5595 8449
rect 5552 8412 5580 8443
rect 6362 8440 6368 8452
rect 6420 8440 6426 8492
rect 6638 8440 6644 8492
rect 6696 8480 6702 8492
rect 7101 8483 7159 8489
rect 7101 8480 7113 8483
rect 6696 8452 7113 8480
rect 6696 8440 6702 8452
rect 7101 8449 7113 8452
rect 7147 8480 7159 8483
rect 7466 8480 7472 8492
rect 7147 8452 7472 8480
rect 7147 8449 7159 8452
rect 7101 8443 7159 8449
rect 7466 8440 7472 8452
rect 7524 8480 7530 8492
rect 7837 8483 7895 8489
rect 7524 8452 7788 8480
rect 7524 8440 7530 8452
rect 7009 8415 7067 8421
rect 7009 8412 7021 8415
rect 4816 8384 5580 8412
rect 5644 8384 7021 8412
rect 4617 8375 4675 8381
rect 4246 8304 4252 8356
rect 4304 8344 4310 8356
rect 4890 8344 4896 8356
rect 4304 8316 4896 8344
rect 4304 8304 4310 8316
rect 4890 8304 4896 8316
rect 4948 8304 4954 8356
rect 5350 8304 5356 8356
rect 5408 8344 5414 8356
rect 5644 8344 5672 8384
rect 7009 8381 7021 8384
rect 7055 8381 7067 8415
rect 7760 8412 7788 8452
rect 7837 8449 7849 8483
rect 7883 8480 7895 8483
rect 8110 8480 8116 8492
rect 7883 8452 8116 8480
rect 7883 8449 7895 8452
rect 7837 8443 7895 8449
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 9784 8480 9812 8576
rect 14568 8548 14596 8588
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 11072 8520 14596 8548
rect 14636 8551 14694 8557
rect 10042 8480 10048 8492
rect 9784 8452 10048 8480
rect 10042 8440 10048 8452
rect 10100 8440 10106 8492
rect 8297 8415 8355 8421
rect 8297 8412 8309 8415
rect 7009 8375 7067 8381
rect 7116 8384 7328 8412
rect 7760 8384 8309 8412
rect 5408 8316 5672 8344
rect 5721 8347 5779 8353
rect 5408 8304 5414 8316
rect 5721 8313 5733 8347
rect 5767 8344 5779 8347
rect 7116 8344 7144 8384
rect 5767 8316 7144 8344
rect 7300 8344 7328 8384
rect 8297 8381 8309 8384
rect 8343 8412 8355 8415
rect 9582 8412 9588 8424
rect 8343 8384 8800 8412
rect 9543 8384 9588 8412
rect 8343 8381 8355 8384
rect 8297 8375 8355 8381
rect 8662 8344 8668 8356
rect 7300 8316 8668 8344
rect 5767 8313 5779 8316
rect 5721 8307 5779 8313
rect 8662 8304 8668 8316
rect 8720 8304 8726 8356
rect 8772 8344 8800 8384
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 9677 8415 9735 8421
rect 9677 8381 9689 8415
rect 9723 8412 9735 8415
rect 10870 8412 10876 8424
rect 9723 8384 10876 8412
rect 9723 8381 9735 8384
rect 9677 8375 9735 8381
rect 10870 8372 10876 8384
rect 10928 8372 10934 8424
rect 11072 8344 11100 8520
rect 14636 8517 14648 8551
rect 14682 8548 14694 8551
rect 14826 8548 14832 8560
rect 14682 8520 14832 8548
rect 14682 8517 14694 8520
rect 14636 8511 14694 8517
rect 14826 8508 14832 8520
rect 14884 8508 14890 8560
rect 16945 8551 17003 8557
rect 16945 8517 16957 8551
rect 16991 8548 17003 8551
rect 17126 8548 17132 8560
rect 16991 8520 17132 8548
rect 16991 8517 17003 8520
rect 16945 8511 17003 8517
rect 17126 8508 17132 8520
rect 17184 8508 17190 8560
rect 17678 8508 17684 8560
rect 17736 8548 17742 8560
rect 20806 8548 20812 8560
rect 17736 8520 20812 8548
rect 17736 8508 17742 8520
rect 12526 8440 12532 8492
rect 12584 8480 12590 8492
rect 13538 8480 13544 8492
rect 12584 8452 12629 8480
rect 13499 8452 13544 8480
rect 12584 8440 12590 8452
rect 13538 8440 13544 8452
rect 13596 8440 13602 8492
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 14366 8480 14372 8492
rect 13688 8452 14228 8480
rect 14327 8452 14372 8480
rect 13688 8440 13694 8452
rect 11882 8412 11888 8424
rect 11843 8384 11888 8412
rect 11882 8372 11888 8384
rect 11940 8372 11946 8424
rect 12250 8412 12256 8424
rect 12211 8384 12256 8412
rect 12250 8372 12256 8384
rect 12308 8372 12314 8424
rect 12434 8372 12440 8424
rect 12492 8412 12498 8424
rect 12492 8384 12537 8412
rect 12492 8372 12498 8384
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14200 8412 14228 8452
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 14476 8480 14596 8484
rect 16114 8480 16120 8492
rect 14476 8456 15424 8480
rect 14476 8412 14504 8456
rect 14568 8452 15424 8456
rect 16075 8452 16120 8480
rect 13780 8384 13825 8412
rect 14200 8384 14504 8412
rect 15396 8412 15424 8452
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16390 8440 16396 8492
rect 16448 8480 16454 8492
rect 17037 8483 17095 8489
rect 16448 8452 16804 8480
rect 16448 8440 16454 8452
rect 16776 8421 16804 8452
rect 17037 8449 17049 8483
rect 17083 8480 17095 8483
rect 17218 8480 17224 8492
rect 17083 8452 17224 8480
rect 17083 8449 17095 8452
rect 17037 8443 17095 8449
rect 17218 8440 17224 8452
rect 17276 8440 17282 8492
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18690 8480 18696 8492
rect 18095 8452 18696 8480
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 18690 8440 18696 8452
rect 18748 8440 18754 8492
rect 18892 8489 18920 8520
rect 20806 8508 20812 8520
rect 20864 8548 20870 8560
rect 21358 8548 21364 8560
rect 20864 8520 21364 8548
rect 20864 8508 20870 8520
rect 21358 8508 21364 8520
rect 21416 8508 21422 8560
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8449 18935 8483
rect 18877 8443 18935 8449
rect 19144 8483 19202 8489
rect 19144 8449 19156 8483
rect 19190 8480 19202 8483
rect 20530 8480 20536 8492
rect 19190 8452 20208 8480
rect 20491 8452 20536 8480
rect 19190 8449 19202 8452
rect 19144 8443 19202 8449
rect 16761 8415 16819 8421
rect 15396 8384 16436 8412
rect 13780 8372 13786 8384
rect 8772 8316 11100 8344
rect 12802 8304 12808 8356
rect 12860 8344 12866 8356
rect 12897 8347 12955 8353
rect 12897 8344 12909 8347
rect 12860 8316 12909 8344
rect 12860 8304 12866 8316
rect 12897 8313 12909 8316
rect 12943 8313 12955 8347
rect 13538 8344 13544 8356
rect 12897 8307 12955 8313
rect 13004 8316 13544 8344
rect 4614 8276 4620 8288
rect 3896 8248 4620 8276
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 8021 8279 8079 8285
rect 8021 8245 8033 8279
rect 8067 8276 8079 8279
rect 8386 8276 8392 8288
rect 8067 8248 8392 8276
rect 8067 8245 8079 8248
rect 8021 8239 8079 8245
rect 8386 8236 8392 8248
rect 8444 8236 8450 8288
rect 10505 8279 10563 8285
rect 10505 8245 10517 8279
rect 10551 8276 10563 8279
rect 10870 8276 10876 8288
rect 10551 8248 10876 8276
rect 10551 8245 10563 8248
rect 10505 8239 10563 8245
rect 10870 8236 10876 8248
rect 10928 8236 10934 8288
rect 11149 8279 11207 8285
rect 11149 8245 11161 8279
rect 11195 8276 11207 8279
rect 13004 8276 13032 8316
rect 13538 8304 13544 8316
rect 13596 8304 13602 8356
rect 15749 8347 15807 8353
rect 15749 8313 15761 8347
rect 15795 8344 15807 8347
rect 15838 8344 15844 8356
rect 15795 8316 15844 8344
rect 15795 8313 15807 8316
rect 15749 8307 15807 8313
rect 15838 8304 15844 8316
rect 15896 8304 15902 8356
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 16080 8316 16313 8344
rect 16080 8304 16086 8316
rect 16301 8313 16313 8316
rect 16347 8313 16359 8347
rect 16408 8344 16436 8384
rect 16761 8381 16773 8415
rect 16807 8412 16819 8415
rect 16807 8384 17908 8412
rect 16807 8381 16819 8384
rect 16761 8375 16819 8381
rect 17405 8347 17463 8353
rect 16408 8316 16712 8344
rect 16301 8307 16359 8313
rect 13170 8276 13176 8288
rect 11195 8248 13032 8276
rect 13131 8248 13176 8276
rect 11195 8245 11207 8248
rect 11149 8239 11207 8245
rect 13170 8236 13176 8248
rect 13228 8236 13234 8288
rect 16684 8276 16712 8316
rect 17405 8313 17417 8347
rect 17451 8344 17463 8347
rect 17770 8344 17776 8356
rect 17451 8316 17776 8344
rect 17451 8313 17463 8316
rect 17405 8307 17463 8313
rect 17770 8304 17776 8316
rect 17828 8304 17834 8356
rect 17880 8344 17908 8384
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18141 8415 18199 8421
rect 18141 8412 18153 8415
rect 18012 8384 18153 8412
rect 18012 8372 18018 8384
rect 18141 8381 18153 8384
rect 18187 8381 18199 8415
rect 18141 8375 18199 8381
rect 18233 8415 18291 8421
rect 18233 8381 18245 8415
rect 18279 8381 18291 8415
rect 20180 8412 20208 8452
rect 20530 8440 20536 8452
rect 20588 8440 20594 8492
rect 21177 8415 21235 8421
rect 21177 8412 21189 8415
rect 20180 8384 21189 8412
rect 18233 8375 18291 8381
rect 21177 8381 21189 8384
rect 21223 8381 21235 8415
rect 21177 8375 21235 8381
rect 18248 8344 18276 8375
rect 17880 8316 18276 8344
rect 17972 8288 18000 8316
rect 17126 8276 17132 8288
rect 16684 8248 17132 8276
rect 17126 8236 17132 8248
rect 17184 8236 17190 8288
rect 17681 8279 17739 8285
rect 17681 8245 17693 8279
rect 17727 8276 17739 8279
rect 17862 8276 17868 8288
rect 17727 8248 17868 8276
rect 17727 8245 17739 8248
rect 17681 8239 17739 8245
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 17954 8236 17960 8288
rect 18012 8236 18018 8288
rect 20254 8276 20260 8288
rect 20215 8248 20260 8276
rect 20254 8236 20260 8248
rect 20312 8236 20318 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2501 8075 2559 8081
rect 2501 8041 2513 8075
rect 2547 8072 2559 8075
rect 2682 8072 2688 8084
rect 2547 8044 2688 8072
rect 2547 8041 2559 8044
rect 2501 8035 2559 8041
rect 2682 8032 2688 8044
rect 2740 8032 2746 8084
rect 4080 8044 7512 8072
rect 2240 7976 3188 8004
rect 2240 7880 2268 7976
rect 2498 7896 2504 7948
rect 2556 7936 2562 7948
rect 3053 7939 3111 7945
rect 3053 7936 3065 7939
rect 2556 7908 3065 7936
rect 2556 7896 2562 7908
rect 3053 7905 3065 7908
rect 3099 7905 3111 7939
rect 3160 7936 3188 7976
rect 3418 7936 3424 7948
rect 3160 7908 3424 7936
rect 3053 7899 3111 7905
rect 3418 7896 3424 7908
rect 3476 7896 3482 7948
rect 1946 7868 1952 7880
rect 1907 7840 1952 7868
rect 1946 7828 1952 7840
rect 2004 7828 2010 7880
rect 2222 7868 2228 7880
rect 2183 7840 2228 7868
rect 2222 7828 2228 7840
rect 2280 7828 2286 7880
rect 2406 7828 2412 7880
rect 2464 7868 2470 7880
rect 2464 7840 3096 7868
rect 2464 7828 2470 7840
rect 2961 7803 3019 7809
rect 2961 7800 2973 7803
rect 2746 7772 2973 7800
rect 2498 7692 2504 7744
rect 2556 7732 2562 7744
rect 2746 7732 2774 7772
rect 2961 7769 2973 7772
rect 3007 7769 3019 7803
rect 3068 7800 3096 7840
rect 3326 7828 3332 7880
rect 3384 7868 3390 7880
rect 4080 7868 4108 8044
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 4212 7976 4384 8004
rect 4212 7964 4218 7976
rect 4356 7945 4384 7976
rect 4522 7964 4528 8016
rect 4580 8004 4586 8016
rect 7285 8007 7343 8013
rect 7285 8004 7297 8007
rect 4580 7976 7297 8004
rect 4580 7964 4586 7976
rect 7285 7973 7297 7976
rect 7331 7973 7343 8007
rect 7285 7967 7343 7973
rect 4341 7939 4399 7945
rect 4341 7905 4353 7939
rect 4387 7936 4399 7939
rect 4706 7936 4712 7948
rect 4387 7908 4712 7936
rect 4387 7905 4399 7908
rect 4341 7899 4399 7905
rect 4706 7896 4712 7908
rect 4764 7936 4770 7948
rect 5626 7936 5632 7948
rect 4764 7908 5632 7936
rect 4764 7896 4770 7908
rect 5626 7896 5632 7908
rect 5684 7896 5690 7948
rect 7484 7936 7512 8044
rect 7650 8032 7656 8084
rect 7708 8072 7714 8084
rect 8110 8072 8116 8084
rect 7708 8044 8116 8072
rect 7708 8032 7714 8044
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 11241 8075 11299 8081
rect 11241 8041 11253 8075
rect 11287 8072 11299 8075
rect 12250 8072 12256 8084
rect 11287 8044 12256 8072
rect 11287 8041 11299 8044
rect 11241 8035 11299 8041
rect 12250 8032 12256 8044
rect 12308 8032 12314 8084
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12897 8075 12955 8081
rect 12897 8072 12909 8075
rect 12492 8044 12909 8072
rect 12492 8032 12498 8044
rect 12897 8041 12909 8044
rect 12943 8041 12955 8075
rect 20622 8072 20628 8084
rect 12897 8035 12955 8041
rect 14844 8044 20628 8072
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8478 8004 8484 8016
rect 7984 7976 8484 8004
rect 7984 7964 7990 7976
rect 8478 7964 8484 7976
rect 8536 7964 8542 8016
rect 12710 7964 12716 8016
rect 12768 8004 12774 8016
rect 14737 8007 14795 8013
rect 14737 8004 14749 8007
rect 12768 7976 14749 8004
rect 12768 7964 12774 7976
rect 14737 7973 14749 7976
rect 14783 7973 14795 8007
rect 14737 7967 14795 7973
rect 8941 7939 8999 7945
rect 8941 7936 8953 7939
rect 7484 7908 8953 7936
rect 3384 7840 4108 7868
rect 4157 7871 4215 7877
rect 3384 7828 3390 7840
rect 4157 7837 4169 7871
rect 4203 7868 4215 7871
rect 4430 7868 4436 7880
rect 4203 7840 4436 7868
rect 4203 7837 4215 7840
rect 4157 7831 4215 7837
rect 4430 7828 4436 7840
rect 4488 7828 4494 7880
rect 7484 7877 7512 7908
rect 8941 7905 8953 7908
rect 8987 7905 8999 7939
rect 8941 7899 8999 7905
rect 13170 7896 13176 7948
rect 13228 7936 13234 7948
rect 13357 7939 13415 7945
rect 13357 7936 13369 7939
rect 13228 7908 13369 7936
rect 13228 7896 13234 7908
rect 13357 7905 13369 7908
rect 13403 7905 13415 7939
rect 13357 7899 13415 7905
rect 13446 7896 13452 7948
rect 13504 7936 13510 7948
rect 13504 7908 13549 7936
rect 13504 7896 13510 7908
rect 7469 7871 7527 7877
rect 7469 7837 7481 7871
rect 7515 7837 7527 7871
rect 7742 7868 7748 7880
rect 7703 7840 7748 7868
rect 7469 7831 7527 7837
rect 7742 7828 7748 7840
rect 7800 7828 7806 7880
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 9490 7868 9496 7880
rect 8444 7840 9496 7868
rect 8444 7828 8450 7840
rect 9490 7828 9496 7840
rect 9548 7828 9554 7880
rect 9585 7871 9643 7877
rect 9585 7837 9597 7871
rect 9631 7868 9643 7871
rect 10318 7868 10324 7880
rect 9631 7840 10324 7868
rect 9631 7837 9643 7840
rect 9585 7831 9643 7837
rect 10318 7828 10324 7840
rect 10376 7828 10382 7880
rect 12621 7871 12679 7877
rect 12621 7868 12633 7871
rect 11716 7840 12633 7868
rect 11716 7812 11744 7840
rect 12621 7837 12633 7840
rect 12667 7868 12679 7871
rect 14366 7868 14372 7880
rect 12667 7840 14372 7868
rect 12667 7837 12679 7840
rect 12621 7831 12679 7837
rect 14366 7828 14372 7840
rect 14424 7828 14430 7880
rect 3068 7772 4292 7800
rect 2961 7763 3019 7769
rect 4264 7741 4292 7772
rect 4614 7760 4620 7812
rect 4672 7800 4678 7812
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 4672 7772 5273 7800
rect 4672 7760 4678 7772
rect 5261 7769 5273 7772
rect 5307 7800 5319 7803
rect 5902 7800 5908 7812
rect 5307 7772 5908 7800
rect 5307 7769 5319 7772
rect 5261 7763 5319 7769
rect 5902 7760 5908 7772
rect 5960 7760 5966 7812
rect 7009 7803 7067 7809
rect 7009 7769 7021 7803
rect 7055 7800 7067 7803
rect 8294 7800 8300 7812
rect 7055 7772 8300 7800
rect 7055 7769 7067 7772
rect 7009 7763 7067 7769
rect 8294 7760 8300 7772
rect 8352 7800 8358 7812
rect 8478 7800 8484 7812
rect 8352 7772 8484 7800
rect 8352 7760 8358 7772
rect 8478 7760 8484 7772
rect 8536 7760 8542 7812
rect 9852 7803 9910 7809
rect 9852 7769 9864 7803
rect 9898 7800 9910 7803
rect 11238 7800 11244 7812
rect 9898 7772 11244 7800
rect 9898 7769 9910 7772
rect 9852 7763 9910 7769
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 11698 7760 11704 7812
rect 11756 7760 11762 7812
rect 12376 7803 12434 7809
rect 12376 7769 12388 7803
rect 12422 7800 12434 7803
rect 13446 7800 13452 7812
rect 12422 7772 13452 7800
rect 12422 7769 12434 7772
rect 12376 7763 12434 7769
rect 13446 7760 13452 7772
rect 13504 7760 13510 7812
rect 14844 7800 14872 8044
rect 20622 8032 20628 8044
rect 20680 8032 20686 8084
rect 18874 8004 18880 8016
rect 18340 7976 18880 8004
rect 17405 7939 17463 7945
rect 17405 7905 17417 7939
rect 17451 7936 17463 7939
rect 17678 7936 17684 7948
rect 17451 7908 17684 7936
rect 17451 7905 17463 7908
rect 17405 7899 17463 7905
rect 17678 7896 17684 7908
rect 17736 7896 17742 7948
rect 17770 7896 17776 7948
rect 17828 7936 17834 7948
rect 18340 7945 18368 7976
rect 18874 7964 18880 7976
rect 18932 7964 18938 8016
rect 18141 7939 18199 7945
rect 18141 7936 18153 7939
rect 17828 7908 18153 7936
rect 17828 7896 17834 7908
rect 18141 7905 18153 7908
rect 18187 7905 18199 7939
rect 18141 7899 18199 7905
rect 18325 7939 18383 7945
rect 18325 7905 18337 7939
rect 18371 7905 18383 7939
rect 18690 7936 18696 7948
rect 18651 7908 18696 7936
rect 18325 7899 18383 7905
rect 18690 7896 18696 7908
rect 18748 7896 18754 7948
rect 20254 7936 20260 7948
rect 20215 7908 20260 7936
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 14921 7871 14979 7877
rect 14921 7837 14933 7871
rect 14967 7837 14979 7871
rect 14921 7831 14979 7837
rect 15381 7871 15439 7877
rect 15381 7837 15393 7871
rect 15427 7868 15439 7871
rect 15470 7868 15476 7880
rect 15427 7840 15476 7868
rect 15427 7837 15439 7840
rect 15381 7831 15439 7837
rect 14476 7772 14872 7800
rect 14936 7800 14964 7831
rect 15470 7828 15476 7840
rect 15528 7828 15534 7880
rect 15562 7828 15568 7880
rect 15620 7868 15626 7880
rect 15657 7871 15715 7877
rect 15657 7868 15669 7871
rect 15620 7840 15669 7868
rect 15620 7828 15626 7840
rect 15657 7837 15669 7840
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 17862 7828 17868 7880
rect 17920 7868 17926 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17920 7840 18061 7868
rect 17920 7828 17926 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18782 7828 18788 7880
rect 18840 7868 18846 7880
rect 19058 7868 19064 7880
rect 18840 7840 19064 7868
rect 18840 7828 18846 7840
rect 19058 7828 19064 7840
rect 19116 7828 19122 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 14936 7772 17724 7800
rect 2556 7704 2774 7732
rect 2869 7735 2927 7741
rect 2556 7692 2562 7704
rect 2869 7701 2881 7735
rect 2915 7732 2927 7735
rect 3789 7735 3847 7741
rect 3789 7732 3801 7735
rect 2915 7704 3801 7732
rect 2915 7701 2927 7704
rect 2869 7695 2927 7701
rect 3789 7701 3801 7704
rect 3835 7701 3847 7735
rect 3789 7695 3847 7701
rect 4249 7735 4307 7741
rect 4249 7701 4261 7735
rect 4295 7732 4307 7735
rect 4430 7732 4436 7744
rect 4295 7704 4436 7732
rect 4295 7701 4307 7704
rect 4249 7695 4307 7701
rect 4430 7692 4436 7704
rect 4488 7692 4494 7744
rect 4798 7732 4804 7744
rect 4759 7704 4804 7732
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 8386 7732 8392 7744
rect 8347 7704 8392 7732
rect 8386 7692 8392 7704
rect 8444 7692 8450 7744
rect 10962 7732 10968 7744
rect 10923 7704 10968 7732
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 13262 7732 13268 7744
rect 13223 7704 13268 7732
rect 13262 7692 13268 7704
rect 13320 7692 13326 7744
rect 14476 7741 14504 7772
rect 14461 7735 14519 7741
rect 14461 7701 14473 7735
rect 14507 7701 14519 7735
rect 14461 7695 14519 7701
rect 14550 7692 14556 7744
rect 14608 7732 14614 7744
rect 17696 7741 17724 7772
rect 17770 7760 17776 7812
rect 17828 7800 17834 7812
rect 19444 7800 19472 7831
rect 20070 7828 20076 7880
rect 20128 7868 20134 7880
rect 20165 7871 20223 7877
rect 20165 7868 20177 7871
rect 20128 7840 20177 7868
rect 20128 7828 20134 7840
rect 20165 7837 20177 7840
rect 20211 7837 20223 7871
rect 20272 7868 20300 7896
rect 20717 7871 20775 7877
rect 20717 7868 20729 7871
rect 20272 7840 20729 7868
rect 20165 7831 20223 7837
rect 20717 7837 20729 7840
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 17828 7772 19472 7800
rect 17828 7760 17834 7772
rect 15197 7735 15255 7741
rect 15197 7732 15209 7735
rect 14608 7704 15209 7732
rect 14608 7692 14614 7704
rect 15197 7701 15209 7704
rect 15243 7701 15255 7735
rect 15197 7695 15255 7701
rect 17681 7735 17739 7741
rect 17681 7701 17693 7735
rect 17727 7701 17739 7735
rect 17681 7695 17739 7701
rect 19058 7692 19064 7744
rect 19116 7732 19122 7744
rect 19245 7735 19303 7741
rect 19245 7732 19257 7735
rect 19116 7704 19257 7732
rect 19116 7692 19122 7704
rect 19245 7701 19257 7704
rect 19291 7701 19303 7735
rect 19702 7732 19708 7744
rect 19663 7704 19708 7732
rect 19245 7695 19303 7701
rect 19702 7692 19708 7704
rect 19760 7692 19766 7744
rect 19794 7692 19800 7744
rect 19852 7732 19858 7744
rect 20073 7735 20131 7741
rect 20073 7732 20085 7735
rect 19852 7704 20085 7732
rect 19852 7692 19858 7704
rect 20073 7701 20085 7704
rect 20119 7701 20131 7735
rect 21358 7732 21364 7744
rect 21319 7704 21364 7732
rect 20073 7695 20131 7701
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 2498 7528 2504 7540
rect 2459 7500 2504 7528
rect 2498 7488 2504 7500
rect 2556 7488 2562 7540
rect 2866 7528 2872 7540
rect 2827 7500 2872 7528
rect 2866 7488 2872 7500
rect 2924 7488 2930 7540
rect 4338 7488 4344 7540
rect 4396 7528 4402 7540
rect 4525 7531 4583 7537
rect 4525 7528 4537 7531
rect 4396 7500 4537 7528
rect 4396 7488 4402 7500
rect 4525 7497 4537 7500
rect 4571 7497 4583 7531
rect 4525 7491 4583 7497
rect 4617 7531 4675 7537
rect 4617 7497 4629 7531
rect 4663 7528 4675 7531
rect 4798 7528 4804 7540
rect 4663 7500 4804 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 4798 7488 4804 7500
rect 4856 7488 4862 7540
rect 4985 7531 5043 7537
rect 4985 7497 4997 7531
rect 5031 7528 5043 7531
rect 5629 7531 5687 7537
rect 5629 7528 5641 7531
rect 5031 7500 5641 7528
rect 5031 7497 5043 7500
rect 4985 7491 5043 7497
rect 5629 7497 5641 7500
rect 5675 7497 5687 7531
rect 5629 7491 5687 7497
rect 5997 7531 6055 7537
rect 5997 7497 6009 7531
rect 6043 7528 6055 7531
rect 7190 7528 7196 7540
rect 6043 7500 7196 7528
rect 6043 7497 6055 7500
rect 5997 7491 6055 7497
rect 7190 7488 7196 7500
rect 7248 7488 7254 7540
rect 9401 7531 9459 7537
rect 9401 7497 9413 7531
rect 9447 7528 9459 7531
rect 9674 7528 9680 7540
rect 9447 7500 9680 7528
rect 9447 7497 9459 7500
rect 9401 7491 9459 7497
rect 9674 7488 9680 7500
rect 9732 7488 9738 7540
rect 10226 7488 10232 7540
rect 10284 7528 10290 7540
rect 10321 7531 10379 7537
rect 10321 7528 10333 7531
rect 10284 7500 10333 7528
rect 10284 7488 10290 7500
rect 10321 7497 10333 7500
rect 10367 7497 10379 7531
rect 11882 7528 11888 7540
rect 11843 7500 11888 7528
rect 10321 7491 10379 7497
rect 11882 7488 11888 7500
rect 11940 7488 11946 7540
rect 12253 7531 12311 7537
rect 12253 7497 12265 7531
rect 12299 7528 12311 7531
rect 12526 7528 12532 7540
rect 12299 7500 12532 7528
rect 12299 7497 12311 7500
rect 12253 7491 12311 7497
rect 12526 7488 12532 7500
rect 12584 7488 12590 7540
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7528 12863 7531
rect 13262 7528 13268 7540
rect 12851 7500 13268 7528
rect 12851 7497 12863 7500
rect 12805 7491 12863 7497
rect 1854 7460 1860 7472
rect 1815 7432 1860 7460
rect 1854 7420 1860 7432
rect 1912 7420 1918 7472
rect 2774 7420 2780 7472
rect 2832 7460 2838 7472
rect 7466 7460 7472 7472
rect 2832 7432 7472 7460
rect 2832 7420 2838 7432
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 1670 7392 1676 7404
rect 1452 7364 1676 7392
rect 1452 7352 1458 7364
rect 1670 7352 1676 7364
rect 1728 7352 1734 7404
rect 2976 7401 3004 7432
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 8288 7463 8346 7469
rect 8288 7429 8300 7463
rect 8334 7460 8346 7463
rect 8386 7460 8392 7472
rect 8334 7432 8392 7460
rect 8334 7429 8346 7432
rect 8288 7423 8346 7429
rect 8386 7420 8392 7432
rect 8444 7420 8450 7472
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7361 3019 7395
rect 2961 7355 3019 7361
rect 3418 7352 3424 7404
rect 3476 7392 3482 7404
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3476 7364 3709 7392
rect 3476 7352 3482 7364
rect 3697 7361 3709 7364
rect 3743 7392 3755 7395
rect 3878 7392 3884 7404
rect 3743 7364 3884 7392
rect 3743 7361 3755 7364
rect 3697 7355 3755 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 9692 7401 9720 7488
rect 9766 7420 9772 7472
rect 9824 7460 9830 7472
rect 11793 7463 11851 7469
rect 11793 7460 11805 7463
rect 9824 7432 11805 7460
rect 9824 7420 9830 7432
rect 11793 7429 11805 7432
rect 11839 7429 11851 7463
rect 11793 7423 11851 7429
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 12820 7460 12848 7491
rect 13262 7488 13268 7500
rect 13320 7488 13326 7540
rect 16942 7528 16948 7540
rect 15580 7500 16948 7528
rect 12124 7432 12848 7460
rect 12124 7420 12130 7432
rect 13814 7420 13820 7472
rect 13872 7460 13878 7472
rect 14194 7463 14252 7469
rect 14194 7460 14206 7463
rect 13872 7432 14206 7460
rect 13872 7420 13878 7432
rect 14194 7429 14206 7432
rect 14240 7429 14252 7463
rect 14194 7423 14252 7429
rect 6621 7395 6679 7401
rect 6621 7392 6633 7395
rect 5828 7364 6633 7392
rect 3145 7327 3203 7333
rect 3145 7293 3157 7327
rect 3191 7324 3203 7327
rect 3234 7324 3240 7336
rect 3191 7296 3240 7324
rect 3191 7293 3203 7296
rect 3145 7287 3203 7293
rect 3234 7284 3240 7296
rect 3292 7324 3298 7336
rect 4154 7324 4160 7336
rect 3292 7296 4160 7324
rect 3292 7284 3298 7296
rect 4154 7284 4160 7296
rect 4212 7284 4218 7336
rect 4433 7327 4491 7333
rect 4433 7293 4445 7327
rect 4479 7324 4491 7327
rect 5166 7324 5172 7336
rect 4479 7296 5172 7324
rect 4479 7293 4491 7296
rect 4433 7287 4491 7293
rect 5166 7284 5172 7296
rect 5224 7284 5230 7336
rect 5353 7327 5411 7333
rect 5353 7293 5365 7327
rect 5399 7293 5411 7327
rect 5534 7324 5540 7336
rect 5495 7296 5540 7324
rect 5353 7287 5411 7293
rect 2225 7191 2283 7197
rect 2225 7157 2237 7191
rect 2271 7188 2283 7191
rect 2406 7188 2412 7200
rect 2271 7160 2412 7188
rect 2271 7157 2283 7160
rect 2225 7151 2283 7157
rect 2406 7148 2412 7160
rect 2464 7148 2470 7200
rect 2590 7148 2596 7200
rect 2648 7188 2654 7200
rect 3513 7191 3571 7197
rect 3513 7188 3525 7191
rect 2648 7160 3525 7188
rect 2648 7148 2654 7160
rect 3513 7157 3525 7160
rect 3559 7157 3571 7191
rect 5368 7188 5396 7287
rect 5534 7284 5540 7296
rect 5592 7284 5598 7336
rect 5828 7188 5856 7364
rect 6621 7361 6633 7364
rect 6667 7361 6679 7395
rect 6621 7355 6679 7361
rect 9677 7395 9735 7401
rect 9677 7361 9689 7395
rect 9723 7361 9735 7395
rect 9677 7355 9735 7361
rect 14366 7352 14372 7404
rect 14424 7392 14430 7404
rect 14461 7395 14519 7401
rect 14461 7392 14473 7395
rect 14424 7364 14473 7392
rect 14424 7352 14430 7364
rect 14461 7361 14473 7364
rect 14507 7361 14519 7395
rect 14461 7355 14519 7361
rect 15381 7395 15439 7401
rect 15381 7361 15393 7395
rect 15427 7392 15439 7395
rect 15580 7392 15608 7500
rect 16942 7488 16948 7500
rect 17000 7488 17006 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18049 7531 18107 7537
rect 18049 7528 18061 7531
rect 18012 7500 18061 7528
rect 18012 7488 18018 7500
rect 18049 7497 18061 7500
rect 18095 7497 18107 7531
rect 18049 7491 18107 7497
rect 18690 7488 18696 7540
rect 18748 7528 18754 7540
rect 19518 7528 19524 7540
rect 18748 7500 19524 7528
rect 18748 7488 18754 7500
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 21174 7528 21180 7540
rect 21135 7500 21180 7528
rect 21174 7488 21180 7500
rect 21232 7488 21238 7540
rect 17678 7460 17684 7472
rect 16684 7432 17684 7460
rect 15427 7364 15608 7392
rect 15657 7395 15715 7401
rect 15427 7361 15439 7364
rect 15381 7355 15439 7361
rect 15657 7361 15669 7395
rect 15703 7392 15715 7395
rect 16574 7392 16580 7404
rect 15703 7364 16580 7392
rect 15703 7361 15715 7364
rect 15657 7355 15715 7361
rect 16574 7352 16580 7364
rect 16632 7352 16638 7404
rect 16684 7401 16712 7432
rect 17678 7420 17684 7432
rect 17736 7420 17742 7472
rect 18598 7420 18604 7472
rect 18656 7460 18662 7472
rect 20564 7463 20622 7469
rect 18656 7432 20484 7460
rect 18656 7420 18662 7432
rect 16942 7401 16948 7404
rect 16669 7395 16727 7401
rect 16669 7361 16681 7395
rect 16715 7361 16727 7395
rect 16669 7355 16727 7361
rect 16936 7355 16948 7401
rect 17000 7392 17006 7404
rect 19153 7395 19211 7401
rect 17000 7364 17036 7392
rect 16942 7352 16948 7355
rect 17000 7352 17006 7364
rect 19153 7361 19165 7395
rect 19199 7392 19211 7395
rect 19518 7392 19524 7404
rect 19199 7364 19524 7392
rect 19199 7361 19211 7364
rect 19153 7355 19211 7361
rect 19518 7352 19524 7364
rect 19576 7352 19582 7404
rect 20456 7392 20484 7432
rect 20564 7429 20576 7463
rect 20610 7460 20622 7463
rect 21358 7460 21364 7472
rect 20610 7432 21364 7460
rect 20610 7429 20622 7432
rect 20564 7423 20622 7429
rect 21358 7420 21364 7432
rect 21416 7420 21422 7472
rect 21269 7395 21327 7401
rect 21269 7392 21281 7395
rect 20456 7364 21281 7392
rect 21269 7361 21281 7364
rect 21315 7361 21327 7395
rect 21269 7355 21327 7361
rect 5902 7284 5908 7336
rect 5960 7324 5966 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 5960 7296 6377 7324
rect 5960 7284 5966 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 8021 7327 8079 7333
rect 8021 7293 8033 7327
rect 8067 7293 8079 7327
rect 8021 7287 8079 7293
rect 5902 7188 5908 7200
rect 5368 7160 5908 7188
rect 3513 7151 3571 7157
rect 5902 7148 5908 7160
rect 5960 7148 5966 7200
rect 7006 7148 7012 7200
rect 7064 7188 7070 7200
rect 7742 7188 7748 7200
rect 7064 7160 7748 7188
rect 7064 7148 7070 7160
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8036 7188 8064 7287
rect 9122 7284 9128 7336
rect 9180 7324 9186 7336
rect 11057 7327 11115 7333
rect 11057 7324 11069 7327
rect 9180 7296 11069 7324
rect 9180 7284 9186 7296
rect 11057 7293 11069 7296
rect 11103 7293 11115 7327
rect 11057 7287 11115 7293
rect 11701 7327 11759 7333
rect 11701 7293 11713 7327
rect 11747 7293 11759 7327
rect 11701 7287 11759 7293
rect 14921 7327 14979 7333
rect 14921 7293 14933 7327
rect 14967 7293 14979 7327
rect 14921 7287 14979 7293
rect 8294 7188 8300 7200
rect 8036 7160 8300 7188
rect 8294 7148 8300 7160
rect 8352 7148 8358 7200
rect 9766 7148 9772 7200
rect 9824 7188 9830 7200
rect 10597 7191 10655 7197
rect 10597 7188 10609 7191
rect 9824 7160 10609 7188
rect 9824 7148 9830 7160
rect 10597 7157 10609 7160
rect 10643 7157 10655 7191
rect 11072 7188 11100 7287
rect 11716 7256 11744 7287
rect 13081 7259 13139 7265
rect 13081 7256 13093 7259
rect 11716 7228 13093 7256
rect 13081 7225 13093 7228
rect 13127 7256 13139 7259
rect 13446 7256 13452 7268
rect 13127 7228 13452 7256
rect 13127 7225 13139 7228
rect 13081 7219 13139 7225
rect 13446 7216 13452 7228
rect 13504 7216 13510 7268
rect 14936 7256 14964 7287
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 16114 7324 16120 7336
rect 15068 7296 16120 7324
rect 15068 7284 15074 7296
rect 16114 7284 16120 7296
rect 16172 7284 16178 7336
rect 16301 7327 16359 7333
rect 16301 7293 16313 7327
rect 16347 7324 16359 7327
rect 16390 7324 16396 7336
rect 16347 7296 16396 7324
rect 16347 7293 16359 7296
rect 16301 7287 16359 7293
rect 16390 7284 16396 7296
rect 16448 7284 16454 7336
rect 19794 7324 19800 7336
rect 18432 7296 19800 7324
rect 14936 7228 16712 7256
rect 14642 7188 14648 7200
rect 11072 7160 14648 7188
rect 10597 7151 10655 7157
rect 14642 7148 14648 7160
rect 14700 7148 14706 7200
rect 15194 7188 15200 7200
rect 15155 7160 15200 7188
rect 15194 7148 15200 7160
rect 15252 7148 15258 7200
rect 15841 7191 15899 7197
rect 15841 7157 15853 7191
rect 15887 7188 15899 7191
rect 15930 7188 15936 7200
rect 15887 7160 15936 7188
rect 15887 7157 15899 7160
rect 15841 7151 15899 7157
rect 15930 7148 15936 7160
rect 15988 7148 15994 7200
rect 16684 7188 16712 7228
rect 18432 7188 18460 7296
rect 19794 7284 19800 7296
rect 19852 7284 19858 7336
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21174 7324 21180 7336
rect 20864 7296 21180 7324
rect 20864 7284 20870 7296
rect 21174 7284 21180 7296
rect 21232 7284 21238 7336
rect 18509 7259 18567 7265
rect 18509 7225 18521 7259
rect 18555 7256 18567 7259
rect 18555 7228 19932 7256
rect 18555 7225 18567 7228
rect 18509 7219 18567 7225
rect 16684 7160 18460 7188
rect 19429 7191 19487 7197
rect 19429 7157 19441 7191
rect 19475 7188 19487 7191
rect 19518 7188 19524 7200
rect 19475 7160 19524 7188
rect 19475 7157 19487 7160
rect 19429 7151 19487 7157
rect 19518 7148 19524 7160
rect 19576 7148 19582 7200
rect 19904 7188 19932 7228
rect 20806 7188 20812 7200
rect 19904 7160 20812 7188
rect 20806 7148 20812 7160
rect 20864 7148 20870 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 5350 6984 5356 6996
rect 4632 6956 5356 6984
rect 2314 6848 2320 6860
rect 2275 6820 2320 6848
rect 2314 6808 2320 6820
rect 2372 6808 2378 6860
rect 2406 6808 2412 6860
rect 2464 6848 2470 6860
rect 3786 6848 3792 6860
rect 2464 6820 3792 6848
rect 2464 6808 2470 6820
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4632 6848 4660 6956
rect 5350 6944 5356 6956
rect 5408 6944 5414 6996
rect 10686 6944 10692 6996
rect 10744 6984 10750 6996
rect 11057 6987 11115 6993
rect 11057 6984 11069 6987
rect 10744 6956 11069 6984
rect 10744 6944 10750 6956
rect 11057 6953 11069 6956
rect 11103 6984 11115 6987
rect 13078 6984 13084 6996
rect 11103 6956 13084 6984
rect 11103 6953 11115 6956
rect 11057 6947 11115 6953
rect 13078 6944 13084 6956
rect 13136 6944 13142 6996
rect 15654 6984 15660 6996
rect 13648 6956 15660 6984
rect 5626 6876 5632 6928
rect 5684 6916 5690 6928
rect 8941 6919 8999 6925
rect 5684 6888 7144 6916
rect 5684 6876 5690 6888
rect 4172 6820 4660 6848
rect 4172 6792 4200 6820
rect 5718 6808 5724 6860
rect 5776 6848 5782 6860
rect 7006 6848 7012 6860
rect 5776 6820 6316 6848
rect 6967 6820 7012 6848
rect 5776 6808 5782 6820
rect 934 6740 940 6792
rect 992 6780 998 6792
rect 1673 6783 1731 6789
rect 1673 6780 1685 6783
rect 992 6752 1685 6780
rect 992 6740 998 6752
rect 1673 6749 1685 6752
rect 1719 6749 1731 6783
rect 3234 6780 3240 6792
rect 3195 6752 3240 6780
rect 1673 6743 1731 6749
rect 3234 6740 3240 6752
rect 3292 6740 3298 6792
rect 4154 6780 4160 6792
rect 4067 6752 4160 6780
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4614 6780 4620 6792
rect 4575 6752 4620 6780
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 6288 6789 6316 6820
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7116 6848 7144 6888
rect 8941 6885 8953 6919
rect 8987 6885 8999 6919
rect 13648 6916 13676 6956
rect 15654 6944 15660 6956
rect 15712 6944 15718 6996
rect 16942 6984 16948 6996
rect 16903 6956 16948 6984
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17405 6987 17463 6993
rect 17405 6953 17417 6987
rect 17451 6984 17463 6987
rect 17770 6984 17776 6996
rect 17451 6956 17776 6984
rect 17451 6953 17463 6956
rect 17405 6947 17463 6953
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 17862 6944 17868 6996
rect 17920 6984 17926 6996
rect 17920 6956 18368 6984
rect 17920 6944 17926 6956
rect 15470 6916 15476 6928
rect 8941 6879 8999 6885
rect 13464 6888 13676 6916
rect 15212 6888 15476 6916
rect 8481 6851 8539 6857
rect 8481 6848 8493 6851
rect 7116 6820 8493 6848
rect 8481 6817 8493 6820
rect 8527 6848 8539 6851
rect 8956 6848 8984 6879
rect 8527 6820 8984 6848
rect 8527 6817 8539 6820
rect 8481 6811 8539 6817
rect 11238 6808 11244 6860
rect 11296 6848 11302 6860
rect 11333 6851 11391 6857
rect 11333 6848 11345 6851
rect 11296 6820 11345 6848
rect 11296 6808 11302 6820
rect 11333 6817 11345 6820
rect 11379 6817 11391 6851
rect 11333 6811 11391 6817
rect 12437 6851 12495 6857
rect 12437 6817 12449 6851
rect 12483 6848 12495 6851
rect 13464 6848 13492 6888
rect 15010 6848 15016 6860
rect 12483 6820 13492 6848
rect 13556 6820 15016 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 6273 6783 6331 6789
rect 4816 6752 6224 6780
rect 1854 6712 1860 6724
rect 1815 6684 1860 6712
rect 1854 6672 1860 6684
rect 1912 6672 1918 6724
rect 2222 6672 2228 6724
rect 2280 6712 2286 6724
rect 2501 6715 2559 6721
rect 2501 6712 2513 6715
rect 2280 6684 2513 6712
rect 2280 6672 2286 6684
rect 2501 6681 2513 6684
rect 2547 6681 2559 6715
rect 2501 6675 2559 6681
rect 3881 6715 3939 6721
rect 3881 6681 3893 6715
rect 3927 6712 3939 6715
rect 4816 6712 4844 6752
rect 3927 6684 4844 6712
rect 4884 6715 4942 6721
rect 3927 6681 3939 6684
rect 3881 6675 3939 6681
rect 4884 6681 4896 6715
rect 4930 6712 4942 6715
rect 5166 6712 5172 6724
rect 4930 6684 5172 6712
rect 4930 6681 4942 6684
rect 4884 6675 4942 6681
rect 5166 6672 5172 6684
rect 5224 6672 5230 6724
rect 5626 6672 5632 6724
rect 5684 6712 5690 6724
rect 5810 6712 5816 6724
rect 5684 6684 5816 6712
rect 5684 6672 5690 6684
rect 5810 6672 5816 6684
rect 5868 6672 5874 6724
rect 6196 6712 6224 6752
rect 6273 6749 6285 6783
rect 6319 6749 6331 6783
rect 7190 6780 7196 6792
rect 7151 6752 7196 6780
rect 6273 6743 6331 6749
rect 7190 6740 7196 6752
rect 7248 6740 7254 6792
rect 9674 6740 9680 6792
rect 9732 6780 9738 6792
rect 10054 6783 10112 6789
rect 10054 6780 10066 6783
rect 9732 6752 10066 6780
rect 9732 6740 9738 6752
rect 10054 6749 10066 6752
rect 10100 6749 10112 6783
rect 10318 6780 10324 6792
rect 10279 6752 10324 6780
rect 10054 6743 10112 6749
rect 10318 6740 10324 6752
rect 10376 6740 10382 6792
rect 11977 6783 12035 6789
rect 11977 6749 11989 6783
rect 12023 6780 12035 6783
rect 12250 6780 12256 6792
rect 12023 6752 12256 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 13556 6789 13584 6820
rect 15010 6808 15016 6820
rect 15068 6808 15074 6860
rect 15105 6851 15163 6857
rect 15105 6817 15117 6851
rect 15151 6848 15163 6851
rect 15212 6848 15240 6888
rect 15470 6876 15476 6888
rect 15528 6916 15534 6928
rect 17954 6916 17960 6928
rect 15528 6888 17960 6916
rect 15528 6876 15534 6888
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 18046 6876 18052 6928
rect 18104 6916 18110 6928
rect 18104 6888 18149 6916
rect 18104 6876 18110 6888
rect 18340 6848 18368 6956
rect 15151 6820 15240 6848
rect 15304 6820 18276 6848
rect 18340 6820 20208 6848
rect 15151 6817 15163 6820
rect 15105 6811 15163 6817
rect 13081 6783 13139 6789
rect 13081 6780 13093 6783
rect 12400 6752 13093 6780
rect 12400 6740 12406 6752
rect 13081 6749 13093 6752
rect 13127 6749 13139 6783
rect 13081 6743 13139 6749
rect 13541 6783 13599 6789
rect 13541 6749 13553 6783
rect 13587 6749 13599 6783
rect 13541 6743 13599 6749
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 14366 6780 14372 6792
rect 14139 6752 14372 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 15304 6712 15332 6820
rect 18248 6792 18276 6820
rect 15381 6783 15439 6789
rect 15381 6749 15393 6783
rect 15427 6749 15439 6783
rect 15381 6743 15439 6749
rect 6196 6684 15332 6712
rect 15396 6712 15424 6743
rect 15654 6740 15660 6792
rect 15712 6780 15718 6792
rect 15841 6783 15899 6789
rect 15841 6780 15853 6783
rect 15712 6752 15853 6780
rect 15712 6740 15718 6752
rect 15841 6749 15853 6752
rect 15887 6749 15899 6783
rect 16298 6780 16304 6792
rect 16259 6752 16304 6780
rect 15841 6743 15899 6749
rect 16298 6740 16304 6752
rect 16356 6740 16362 6792
rect 16574 6740 16580 6792
rect 16632 6780 16638 6792
rect 17034 6780 17040 6792
rect 16632 6752 17040 6780
rect 16632 6740 16638 6752
rect 17034 6740 17040 6752
rect 17092 6740 17098 6792
rect 17221 6783 17279 6789
rect 17221 6749 17233 6783
rect 17267 6776 17279 6783
rect 17310 6776 17316 6792
rect 17267 6749 17316 6776
rect 17221 6748 17316 6749
rect 17221 6743 17279 6748
rect 17310 6740 17316 6748
rect 17368 6776 17374 6792
rect 17862 6780 17868 6792
rect 17788 6776 17868 6780
rect 17368 6752 17868 6776
rect 17368 6748 17816 6752
rect 17368 6740 17374 6748
rect 17862 6740 17868 6752
rect 17920 6740 17926 6792
rect 18230 6780 18236 6792
rect 18191 6752 18236 6780
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18322 6740 18328 6792
rect 18380 6780 18386 6792
rect 18785 6783 18843 6789
rect 18785 6780 18797 6783
rect 18380 6752 18797 6780
rect 18380 6740 18386 6752
rect 18785 6749 18797 6752
rect 18831 6749 18843 6783
rect 18785 6743 18843 6749
rect 18966 6740 18972 6792
rect 19024 6780 19030 6792
rect 19613 6783 19671 6789
rect 19613 6780 19625 6783
rect 19024 6752 19625 6780
rect 19024 6740 19030 6752
rect 19613 6749 19625 6752
rect 19659 6749 19671 6783
rect 19613 6743 19671 6749
rect 17954 6712 17960 6724
rect 15396 6684 17960 6712
rect 17954 6672 17960 6684
rect 18012 6672 18018 6724
rect 18598 6712 18604 6724
rect 18559 6684 18604 6712
rect 18598 6672 18604 6684
rect 18656 6672 18662 6724
rect 19426 6712 19432 6724
rect 19387 6684 19432 6712
rect 19426 6672 19432 6684
rect 19484 6672 19490 6724
rect 20070 6712 20076 6724
rect 19536 6684 20076 6712
rect 2406 6644 2412 6656
rect 2367 6616 2412 6644
rect 2406 6604 2412 6616
rect 2464 6604 2470 6656
rect 2869 6647 2927 6653
rect 2869 6613 2881 6647
rect 2915 6644 2927 6647
rect 3050 6644 3056 6656
rect 2915 6616 3056 6644
rect 2915 6613 2927 6616
rect 2869 6607 2927 6613
rect 3050 6604 3056 6616
rect 3108 6604 3114 6656
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 3970 6644 3976 6656
rect 3467 6616 3976 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4341 6647 4399 6653
rect 4341 6613 4353 6647
rect 4387 6644 4399 6647
rect 4706 6644 4712 6656
rect 4387 6616 4712 6644
rect 4387 6613 4399 6616
rect 4341 6607 4399 6613
rect 4706 6604 4712 6616
rect 4764 6604 4770 6656
rect 5350 6604 5356 6656
rect 5408 6644 5414 6656
rect 5902 6644 5908 6656
rect 5408 6616 5908 6644
rect 5408 6604 5414 6616
rect 5902 6604 5908 6616
rect 5960 6644 5966 6656
rect 5997 6647 6055 6653
rect 5997 6644 6009 6647
rect 5960 6616 6009 6644
rect 5960 6604 5966 6616
rect 5997 6613 6009 6616
rect 6043 6613 6055 6647
rect 5997 6607 6055 6613
rect 6457 6647 6515 6653
rect 6457 6613 6469 6647
rect 6503 6644 6515 6647
rect 6730 6644 6736 6656
rect 6503 6616 6736 6644
rect 6503 6613 6515 6616
rect 6457 6607 6515 6613
rect 6730 6604 6736 6616
rect 6788 6604 6794 6656
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7374 6604 7380 6656
rect 7432 6644 7438 6656
rect 7561 6647 7619 6653
rect 7561 6644 7573 6647
rect 7432 6616 7573 6644
rect 7432 6604 7438 6616
rect 7561 6613 7573 6616
rect 7607 6613 7619 6647
rect 7561 6607 7619 6613
rect 7742 6604 7748 6656
rect 7800 6644 7806 6656
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 7800 6616 7849 6644
rect 7800 6604 7806 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 8202 6644 8208 6656
rect 8163 6616 8208 6644
rect 7837 6607 7895 6613
rect 8202 6604 8208 6616
rect 8260 6604 8266 6656
rect 8297 6647 8355 6653
rect 8297 6613 8309 6647
rect 8343 6644 8355 6647
rect 8846 6644 8852 6656
rect 8343 6616 8852 6644
rect 8343 6613 8355 6616
rect 8297 6607 8355 6613
rect 8846 6604 8852 6616
rect 8904 6604 8910 6656
rect 9306 6604 9312 6656
rect 9364 6644 9370 6656
rect 10597 6647 10655 6653
rect 10597 6644 10609 6647
rect 9364 6616 10609 6644
rect 9364 6604 9370 6616
rect 10597 6613 10609 6616
rect 10643 6644 10655 6647
rect 10870 6644 10876 6656
rect 10643 6616 10876 6644
rect 10643 6613 10655 6616
rect 10597 6607 10655 6613
rect 10870 6604 10876 6616
rect 10928 6604 10934 6656
rect 12805 6647 12863 6653
rect 12805 6613 12817 6647
rect 12851 6644 12863 6647
rect 12986 6644 12992 6656
rect 12851 6616 12992 6644
rect 12851 6613 12863 6616
rect 12805 6607 12863 6613
rect 12986 6604 12992 6616
rect 13044 6604 13050 6656
rect 13170 6604 13176 6656
rect 13228 6644 13234 6656
rect 13265 6647 13323 6653
rect 13265 6644 13277 6647
rect 13228 6616 13277 6644
rect 13228 6604 13234 6616
rect 13265 6613 13277 6616
rect 13311 6613 13323 6647
rect 13722 6644 13728 6656
rect 13683 6616 13728 6644
rect 13265 6607 13323 6613
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 14734 6644 14740 6656
rect 14695 6616 14740 6644
rect 14734 6604 14740 6616
rect 14792 6604 14798 6656
rect 15565 6647 15623 6653
rect 15565 6613 15577 6647
rect 15611 6644 15623 6647
rect 15746 6644 15752 6656
rect 15611 6616 15752 6644
rect 15611 6613 15623 6616
rect 15565 6607 15623 6613
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 16025 6647 16083 6653
rect 16025 6613 16037 6647
rect 16071 6644 16083 6647
rect 17310 6644 17316 6656
rect 16071 6616 17316 6644
rect 16071 6613 16083 6616
rect 16025 6607 16083 6613
rect 17310 6604 17316 6616
rect 17368 6604 17374 6656
rect 17494 6604 17500 6656
rect 17552 6644 17558 6656
rect 17681 6647 17739 6653
rect 17681 6644 17693 6647
rect 17552 6616 17693 6644
rect 17552 6604 17558 6616
rect 17681 6613 17693 6616
rect 17727 6613 17739 6647
rect 17681 6607 17739 6613
rect 17770 6604 17776 6656
rect 17828 6644 17834 6656
rect 19536 6644 19564 6684
rect 20070 6672 20076 6684
rect 20128 6672 20134 6724
rect 20180 6712 20208 6820
rect 20254 6740 20260 6792
rect 20312 6780 20318 6792
rect 20530 6780 20536 6792
rect 20312 6752 20536 6780
rect 20312 6740 20318 6752
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 20806 6740 20812 6792
rect 20864 6780 20870 6792
rect 21094 6783 21152 6789
rect 21094 6780 21106 6783
rect 20864 6752 21106 6780
rect 20864 6740 20870 6752
rect 21094 6749 21106 6752
rect 21140 6749 21152 6783
rect 21094 6743 21152 6749
rect 21266 6740 21272 6792
rect 21324 6780 21330 6792
rect 21361 6783 21419 6789
rect 21361 6780 21373 6783
rect 21324 6752 21373 6780
rect 21324 6740 21330 6752
rect 21361 6749 21373 6752
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 21818 6712 21824 6724
rect 20180 6684 21824 6712
rect 21818 6672 21824 6684
rect 21876 6672 21882 6724
rect 19978 6644 19984 6656
rect 17828 6616 19564 6644
rect 19939 6616 19984 6644
rect 17828 6604 17834 6616
rect 19978 6604 19984 6616
rect 20036 6604 20042 6656
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 1857 6443 1915 6449
rect 1857 6409 1869 6443
rect 1903 6440 1915 6443
rect 2038 6440 2044 6452
rect 1903 6412 2044 6440
rect 1903 6409 1915 6412
rect 1857 6403 1915 6409
rect 2038 6400 2044 6412
rect 2096 6400 2102 6452
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 2406 6400 2412 6452
rect 2464 6440 2470 6452
rect 2501 6443 2559 6449
rect 2501 6440 2513 6443
rect 2464 6412 2513 6440
rect 2464 6400 2470 6412
rect 2501 6409 2513 6412
rect 2547 6409 2559 6443
rect 2501 6403 2559 6409
rect 2682 6400 2688 6452
rect 2740 6440 2746 6452
rect 2869 6443 2927 6449
rect 2869 6440 2881 6443
rect 2740 6412 2881 6440
rect 2740 6400 2746 6412
rect 2869 6409 2881 6412
rect 2915 6440 2927 6443
rect 2915 6412 4016 6440
rect 2915 6409 2927 6412
rect 2869 6403 2927 6409
rect 1765 6375 1823 6381
rect 1765 6341 1777 6375
rect 1811 6372 1823 6375
rect 2590 6372 2596 6384
rect 1811 6344 2596 6372
rect 1811 6341 1823 6344
rect 1765 6335 1823 6341
rect 2590 6332 2596 6344
rect 2648 6332 2654 6384
rect 2958 6372 2964 6384
rect 2919 6344 2964 6372
rect 2958 6332 2964 6344
rect 3016 6332 3022 6384
rect 3418 6264 3424 6316
rect 3476 6304 3482 6316
rect 3513 6307 3571 6313
rect 3513 6304 3525 6307
rect 3476 6276 3525 6304
rect 3476 6264 3482 6276
rect 3513 6273 3525 6276
rect 3559 6273 3571 6307
rect 3513 6267 3571 6273
rect 1673 6239 1731 6245
rect 1673 6205 1685 6239
rect 1719 6205 1731 6239
rect 1673 6199 1731 6205
rect 3053 6239 3111 6245
rect 3053 6205 3065 6239
rect 3099 6205 3111 6239
rect 3988 6236 4016 6412
rect 4706 6400 4712 6452
rect 4764 6440 4770 6452
rect 5074 6440 5080 6452
rect 4764 6412 5080 6440
rect 4764 6400 4770 6412
rect 5074 6400 5080 6412
rect 5132 6400 5138 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5592 6412 6009 6440
rect 5592 6400 5598 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 5997 6403 6055 6409
rect 6196 6412 6837 6440
rect 6196 6384 6224 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7653 6443 7711 6449
rect 7653 6440 7665 6443
rect 6972 6412 7665 6440
rect 6972 6400 6978 6412
rect 7653 6409 7665 6412
rect 7699 6409 7711 6443
rect 7653 6403 7711 6409
rect 7834 6400 7840 6452
rect 7892 6440 7898 6452
rect 7929 6443 7987 6449
rect 7929 6440 7941 6443
rect 7892 6412 7941 6440
rect 7892 6400 7898 6412
rect 7929 6409 7941 6412
rect 7975 6409 7987 6443
rect 8846 6440 8852 6452
rect 8807 6412 8852 6440
rect 7929 6403 7987 6409
rect 8846 6400 8852 6412
rect 8904 6400 8910 6452
rect 9122 6400 9128 6452
rect 9180 6440 9186 6452
rect 9217 6443 9275 6449
rect 9217 6440 9229 6443
rect 9180 6412 9229 6440
rect 9180 6400 9186 6412
rect 9217 6409 9229 6412
rect 9263 6409 9275 6443
rect 9217 6403 9275 6409
rect 9306 6400 9312 6452
rect 9364 6440 9370 6452
rect 10045 6443 10103 6449
rect 9364 6412 9409 6440
rect 9364 6400 9370 6412
rect 10045 6409 10057 6443
rect 10091 6440 10103 6443
rect 10410 6440 10416 6452
rect 10091 6412 10416 6440
rect 10091 6409 10103 6412
rect 10045 6403 10103 6409
rect 10410 6400 10416 6412
rect 10468 6400 10474 6452
rect 10686 6440 10692 6452
rect 10647 6412 10692 6440
rect 10686 6400 10692 6412
rect 10744 6400 10750 6452
rect 13357 6443 13415 6449
rect 13357 6409 13369 6443
rect 13403 6440 13415 6443
rect 14642 6440 14648 6452
rect 13403 6412 14648 6440
rect 13403 6409 13415 6412
rect 13357 6403 13415 6409
rect 14642 6400 14648 6412
rect 14700 6400 14706 6452
rect 17037 6443 17095 6449
rect 14752 6412 16252 6440
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 4120 6344 6132 6372
rect 4120 6332 4126 6344
rect 4801 6307 4859 6313
rect 4801 6273 4813 6307
rect 4847 6304 4859 6307
rect 4890 6304 4896 6316
rect 4847 6276 4896 6304
rect 4847 6273 4859 6276
rect 4801 6267 4859 6273
rect 4890 6264 4896 6276
rect 4948 6304 4954 6316
rect 5074 6304 5080 6316
rect 4948 6276 5080 6304
rect 4948 6264 4954 6276
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 5534 6304 5540 6316
rect 5495 6276 5540 6304
rect 5534 6264 5540 6276
rect 5592 6264 5598 6316
rect 5629 6307 5687 6313
rect 5629 6273 5641 6307
rect 5675 6273 5687 6307
rect 6104 6304 6132 6344
rect 6178 6332 6184 6384
rect 6236 6332 6242 6384
rect 7742 6372 7748 6384
rect 6288 6344 7748 6372
rect 6288 6304 6316 6344
rect 7742 6332 7748 6344
rect 7800 6332 7806 6384
rect 8570 6372 8576 6384
rect 8128 6344 8576 6372
rect 6104 6276 6316 6304
rect 6380 6276 7144 6304
rect 5629 6267 5687 6273
rect 5258 6236 5264 6248
rect 3988 6208 5264 6236
rect 3053 6199 3111 6205
rect 1688 6168 1716 6199
rect 2590 6168 2596 6180
rect 1688 6140 2596 6168
rect 2590 6128 2596 6140
rect 2648 6168 2654 6180
rect 3068 6168 3096 6199
rect 5258 6196 5264 6208
rect 5316 6196 5322 6248
rect 5445 6239 5503 6245
rect 5445 6205 5457 6239
rect 5491 6205 5503 6239
rect 5644 6236 5672 6267
rect 6086 6236 6092 6248
rect 5644 6208 6092 6236
rect 5445 6199 5503 6205
rect 2648 6140 3096 6168
rect 4525 6171 4583 6177
rect 2648 6128 2654 6140
rect 4525 6137 4537 6171
rect 4571 6168 4583 6171
rect 4571 6140 5120 6168
rect 4571 6137 4583 6140
rect 4525 6131 4583 6137
rect 4154 6100 4160 6112
rect 4115 6072 4160 6100
rect 4154 6060 4160 6072
rect 4212 6060 4218 6112
rect 4982 6100 4988 6112
rect 4943 6072 4988 6100
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5092 6100 5120 6140
rect 5166 6128 5172 6180
rect 5224 6168 5230 6180
rect 5460 6168 5488 6199
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 6270 6196 6276 6248
rect 6328 6236 6334 6248
rect 6380 6236 6408 6276
rect 6328 6208 6408 6236
rect 6328 6196 6334 6208
rect 6638 6196 6644 6248
rect 6696 6236 6702 6248
rect 6917 6239 6975 6245
rect 6917 6236 6929 6239
rect 6696 6208 6929 6236
rect 6696 6196 6702 6208
rect 6917 6205 6929 6208
rect 6963 6205 6975 6239
rect 6917 6199 6975 6205
rect 7009 6239 7067 6245
rect 7009 6205 7021 6239
rect 7055 6205 7067 6239
rect 7116 6236 7144 6276
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7469 6307 7527 6313
rect 7469 6304 7481 6307
rect 7248 6276 7481 6304
rect 7248 6264 7254 6276
rect 7469 6273 7481 6276
rect 7515 6304 7527 6307
rect 8018 6304 8024 6316
rect 7515 6276 8024 6304
rect 7515 6273 7527 6276
rect 7469 6267 7527 6273
rect 8018 6264 8024 6276
rect 8076 6264 8082 6316
rect 8128 6313 8156 6344
rect 8570 6332 8576 6344
rect 8628 6332 8634 6384
rect 9674 6372 9680 6384
rect 9508 6344 9680 6372
rect 8113 6307 8171 6313
rect 8113 6273 8125 6307
rect 8159 6273 8171 6307
rect 8113 6267 8171 6273
rect 8389 6307 8447 6313
rect 8389 6273 8401 6307
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 8404 6236 8432 6267
rect 9508 6245 9536 6344
rect 9674 6332 9680 6344
rect 9732 6372 9738 6384
rect 14752 6372 14780 6412
rect 15470 6372 15476 6384
rect 9732 6344 14780 6372
rect 15120 6344 15476 6372
rect 9732 6332 9738 6344
rect 9766 6264 9772 6316
rect 9824 6304 9830 6316
rect 9861 6307 9919 6313
rect 9861 6304 9873 6307
rect 9824 6276 9873 6304
rect 9824 6264 9830 6276
rect 9861 6273 9873 6276
rect 9907 6273 9919 6307
rect 9861 6267 9919 6273
rect 10686 6264 10692 6316
rect 10744 6304 10750 6316
rect 10781 6307 10839 6313
rect 10781 6304 10793 6307
rect 10744 6276 10793 6304
rect 10744 6264 10750 6276
rect 10781 6273 10793 6276
rect 10827 6273 10839 6307
rect 11882 6304 11888 6316
rect 11843 6276 11888 6304
rect 10781 6267 10839 6273
rect 11882 6264 11888 6276
rect 11940 6264 11946 6316
rect 12158 6264 12164 6316
rect 12216 6304 12222 6316
rect 12621 6307 12679 6313
rect 12216 6276 12434 6304
rect 12216 6264 12222 6276
rect 7116 6208 8432 6236
rect 9493 6239 9551 6245
rect 7009 6199 7067 6205
rect 9493 6205 9505 6239
rect 9539 6205 9551 6239
rect 9493 6199 9551 6205
rect 10597 6239 10655 6245
rect 10597 6205 10609 6239
rect 10643 6236 10655 6239
rect 10962 6236 10968 6248
rect 10643 6208 10968 6236
rect 10643 6205 10655 6208
rect 10597 6199 10655 6205
rect 6822 6168 6828 6180
rect 5224 6140 6828 6168
rect 5224 6128 5230 6140
rect 6822 6128 6828 6140
rect 6880 6168 6886 6180
rect 7024 6168 7052 6199
rect 10962 6196 10968 6208
rect 11020 6196 11026 6248
rect 11974 6236 11980 6248
rect 11935 6208 11980 6236
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12406 6236 12434 6276
rect 12621 6273 12633 6307
rect 12667 6304 12679 6307
rect 12710 6304 12716 6316
rect 12667 6276 12716 6304
rect 12667 6273 12679 6276
rect 12621 6267 12679 6273
rect 12710 6264 12716 6276
rect 12768 6264 12774 6316
rect 13449 6307 13507 6313
rect 13449 6304 13461 6307
rect 12912 6276 13461 6304
rect 12912 6236 12940 6276
rect 13449 6273 13461 6276
rect 13495 6273 13507 6307
rect 14844 6304 15056 6308
rect 15120 6304 15148 6344
rect 15470 6332 15476 6344
rect 15528 6332 15534 6384
rect 13449 6267 13507 6273
rect 14292 6280 15148 6304
rect 14292 6276 14872 6280
rect 15028 6276 15148 6280
rect 15188 6307 15246 6313
rect 13262 6236 13268 6248
rect 12406 6208 12940 6236
rect 13223 6208 13268 6236
rect 12069 6199 12127 6205
rect 8573 6171 8631 6177
rect 6880 6140 7052 6168
rect 7116 6140 7788 6168
rect 6880 6128 6886 6140
rect 5534 6100 5540 6112
rect 5092 6072 5540 6100
rect 5534 6060 5540 6072
rect 5592 6100 5598 6112
rect 6270 6100 6276 6112
rect 5592 6072 6276 6100
rect 5592 6060 5598 6072
rect 6270 6060 6276 6072
rect 6328 6060 6334 6112
rect 6457 6103 6515 6109
rect 6457 6069 6469 6103
rect 6503 6100 6515 6103
rect 6638 6100 6644 6112
rect 6503 6072 6644 6100
rect 6503 6069 6515 6072
rect 6457 6063 6515 6069
rect 6638 6060 6644 6072
rect 6696 6060 6702 6112
rect 6730 6060 6736 6112
rect 6788 6100 6794 6112
rect 7116 6100 7144 6140
rect 6788 6072 7144 6100
rect 7760 6100 7788 6140
rect 8573 6137 8585 6171
rect 8619 6168 8631 6171
rect 10502 6168 10508 6180
rect 8619 6140 10508 6168
rect 8619 6137 8631 6140
rect 8573 6131 8631 6137
rect 10502 6128 10508 6140
rect 10560 6128 10566 6180
rect 10980 6168 11008 6196
rect 12084 6168 12112 6199
rect 13262 6196 13268 6208
rect 13320 6196 13326 6248
rect 14292 6245 14320 6276
rect 15188 6273 15200 6307
rect 15234 6304 15246 6307
rect 16224 6304 16252 6412
rect 17037 6409 17049 6443
rect 17083 6440 17095 6443
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 17083 6412 17693 6440
rect 17083 6409 17095 6412
rect 17037 6403 17095 6409
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 17681 6403 17739 6409
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 19429 6443 19487 6449
rect 19429 6440 19441 6443
rect 18012 6412 19441 6440
rect 18012 6400 18018 6412
rect 19429 6409 19441 6412
rect 19475 6409 19487 6443
rect 19429 6403 19487 6409
rect 19702 6400 19708 6452
rect 19760 6440 19766 6452
rect 19889 6443 19947 6449
rect 19889 6440 19901 6443
rect 19760 6412 19901 6440
rect 19760 6400 19766 6412
rect 19889 6409 19901 6412
rect 19935 6409 19947 6443
rect 19889 6403 19947 6409
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 20809 6443 20867 6449
rect 20809 6440 20821 6443
rect 20680 6412 20821 6440
rect 20680 6400 20686 6412
rect 20809 6409 20821 6412
rect 20855 6409 20867 6443
rect 20809 6403 20867 6409
rect 16390 6332 16396 6384
rect 16448 6372 16454 6384
rect 18049 6375 18107 6381
rect 18049 6372 18061 6375
rect 16448 6344 18061 6372
rect 16448 6332 16454 6344
rect 18049 6341 18061 6344
rect 18095 6341 18107 6375
rect 19978 6372 19984 6384
rect 18049 6335 18107 6341
rect 18156 6344 19984 6372
rect 18156 6304 18184 6344
rect 19978 6332 19984 6344
rect 20036 6332 20042 6384
rect 20070 6332 20076 6384
rect 20128 6372 20134 6384
rect 20714 6372 20720 6384
rect 20128 6344 20720 6372
rect 20128 6332 20134 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 15234 6276 16160 6304
rect 16224 6276 18184 6304
rect 18248 6276 18460 6304
rect 15234 6273 15246 6276
rect 15188 6267 15246 6273
rect 14277 6239 14335 6245
rect 14277 6205 14289 6239
rect 14323 6205 14335 6239
rect 14277 6199 14335 6205
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 14921 6239 14979 6245
rect 14921 6236 14933 6239
rect 14516 6208 14933 6236
rect 14516 6196 14522 6208
rect 14921 6205 14933 6208
rect 14967 6205 14979 6239
rect 16132 6236 16160 6276
rect 16942 6236 16948 6248
rect 16132 6208 16948 6236
rect 14921 6199 14979 6205
rect 16942 6196 16948 6208
rect 17000 6196 17006 6248
rect 17126 6236 17132 6248
rect 17087 6208 17132 6236
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 17221 6239 17279 6245
rect 17221 6205 17233 6239
rect 17267 6205 17279 6239
rect 17221 6199 17279 6205
rect 18141 6239 18199 6245
rect 18141 6205 18153 6239
rect 18187 6236 18199 6239
rect 18248 6236 18276 6276
rect 18187 6208 18276 6236
rect 18325 6239 18383 6245
rect 18187 6205 18199 6208
rect 18141 6199 18199 6205
rect 18325 6205 18337 6239
rect 18371 6205 18383 6239
rect 18432 6236 18460 6276
rect 18506 6264 18512 6316
rect 18564 6304 18570 6316
rect 18877 6307 18935 6313
rect 18877 6304 18889 6307
rect 18564 6276 18889 6304
rect 18564 6264 18570 6276
rect 18877 6273 18889 6276
rect 18923 6273 18935 6307
rect 18877 6267 18935 6273
rect 18966 6264 18972 6316
rect 19024 6304 19030 6316
rect 19061 6307 19119 6313
rect 19061 6304 19073 6307
rect 19024 6276 19073 6304
rect 19024 6264 19030 6276
rect 19061 6273 19073 6276
rect 19107 6273 19119 6307
rect 19794 6304 19800 6316
rect 19755 6276 19800 6304
rect 19061 6267 19119 6273
rect 19794 6264 19800 6276
rect 19852 6264 19858 6316
rect 18690 6236 18696 6248
rect 18432 6208 18696 6236
rect 18325 6199 18383 6205
rect 10980 6140 12112 6168
rect 12158 6128 12164 6180
rect 12216 6168 12222 6180
rect 16298 6168 16304 6180
rect 12216 6140 14964 6168
rect 16211 6140 16304 6168
rect 12216 6128 12222 6140
rect 10594 6100 10600 6112
rect 7760 6072 10600 6100
rect 6788 6060 6794 6072
rect 10594 6060 10600 6072
rect 10652 6060 10658 6112
rect 11146 6100 11152 6112
rect 11107 6072 11152 6100
rect 11146 6060 11152 6072
rect 11204 6060 11210 6112
rect 11238 6060 11244 6112
rect 11296 6100 11302 6112
rect 11517 6103 11575 6109
rect 11517 6100 11529 6103
rect 11296 6072 11529 6100
rect 11296 6060 11302 6072
rect 11517 6069 11529 6072
rect 11563 6069 11575 6103
rect 11517 6063 11575 6069
rect 12805 6103 12863 6109
rect 12805 6069 12817 6103
rect 12851 6100 12863 6103
rect 13630 6100 13636 6112
rect 12851 6072 13636 6100
rect 12851 6069 12863 6072
rect 12805 6063 12863 6069
rect 13630 6060 13636 6072
rect 13688 6060 13694 6112
rect 13814 6100 13820 6112
rect 13775 6072 13820 6100
rect 13814 6060 13820 6072
rect 13872 6060 13878 6112
rect 14936 6100 14964 6140
rect 16298 6128 16304 6140
rect 16356 6168 16362 6180
rect 17236 6168 17264 6199
rect 16356 6140 17264 6168
rect 16356 6128 16362 6140
rect 16390 6100 16396 6112
rect 14936 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16666 6100 16672 6112
rect 16627 6072 16672 6100
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 18138 6100 18144 6112
rect 17000 6072 18144 6100
rect 17000 6060 17006 6072
rect 18138 6060 18144 6072
rect 18196 6100 18202 6112
rect 18340 6100 18368 6199
rect 18690 6196 18696 6208
rect 18748 6196 18754 6248
rect 19518 6196 19524 6248
rect 19576 6236 19582 6248
rect 19981 6239 20039 6245
rect 19981 6236 19993 6239
rect 19576 6208 19993 6236
rect 19576 6196 19582 6208
rect 19981 6205 19993 6208
rect 20027 6205 20039 6239
rect 20898 6236 20904 6248
rect 20859 6208 20904 6236
rect 19981 6199 20039 6205
rect 20898 6196 20904 6208
rect 20956 6196 20962 6248
rect 20993 6239 21051 6245
rect 20993 6205 21005 6239
rect 21039 6205 21051 6239
rect 20993 6199 21051 6205
rect 18874 6128 18880 6180
rect 18932 6168 18938 6180
rect 21008 6168 21036 6199
rect 18932 6140 21036 6168
rect 18932 6128 18938 6140
rect 18196 6072 18368 6100
rect 20441 6103 20499 6109
rect 18196 6060 18202 6072
rect 20441 6069 20453 6103
rect 20487 6100 20499 6103
rect 20622 6100 20628 6112
rect 20487 6072 20628 6100
rect 20487 6069 20499 6072
rect 20441 6063 20499 6069
rect 20622 6060 20628 6072
rect 20680 6060 20686 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1673 5899 1731 5905
rect 1673 5865 1685 5899
rect 1719 5896 1731 5899
rect 2682 5896 2688 5908
rect 1719 5868 2688 5896
rect 1719 5865 1731 5868
rect 1673 5859 1731 5865
rect 2682 5856 2688 5868
rect 2740 5856 2746 5908
rect 3970 5856 3976 5908
rect 4028 5896 4034 5908
rect 5166 5896 5172 5908
rect 4028 5868 4752 5896
rect 5127 5868 5172 5896
rect 4028 5856 4034 5868
rect 4724 5828 4752 5868
rect 5166 5856 5172 5868
rect 5224 5856 5230 5908
rect 6730 5896 6736 5908
rect 5552 5868 6736 5896
rect 5552 5828 5580 5868
rect 6730 5856 6736 5868
rect 6788 5856 6794 5908
rect 7098 5896 7104 5908
rect 7059 5868 7104 5896
rect 7098 5856 7104 5868
rect 7156 5856 7162 5908
rect 8202 5856 8208 5908
rect 8260 5896 8266 5908
rect 9033 5899 9091 5905
rect 9033 5896 9045 5899
rect 8260 5868 9045 5896
rect 8260 5856 8266 5868
rect 9033 5865 9045 5868
rect 9079 5865 9091 5899
rect 9033 5859 9091 5865
rect 9490 5856 9496 5908
rect 9548 5896 9554 5908
rect 12158 5896 12164 5908
rect 9548 5868 12164 5896
rect 9548 5856 9554 5868
rect 12158 5856 12164 5868
rect 12216 5856 12222 5908
rect 13262 5856 13268 5908
rect 13320 5896 13326 5908
rect 13320 5868 15700 5896
rect 13320 5856 13326 5868
rect 4724 5800 5580 5828
rect 5629 5831 5687 5837
rect 5629 5797 5641 5831
rect 5675 5828 5687 5831
rect 5718 5828 5724 5840
rect 5675 5800 5724 5828
rect 5675 5797 5687 5800
rect 5629 5791 5687 5797
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 5994 5788 6000 5840
rect 6052 5828 6058 5840
rect 6089 5831 6147 5837
rect 6089 5828 6101 5831
rect 6052 5800 6101 5828
rect 6052 5788 6058 5800
rect 6089 5797 6101 5800
rect 6135 5797 6147 5831
rect 6089 5791 6147 5797
rect 6914 5788 6920 5840
rect 6972 5828 6978 5840
rect 7377 5831 7435 5837
rect 7377 5828 7389 5831
rect 6972 5800 7389 5828
rect 6972 5788 6978 5800
rect 7377 5797 7389 5800
rect 7423 5797 7435 5831
rect 7377 5791 7435 5797
rect 7466 5788 7472 5840
rect 7524 5828 7530 5840
rect 8297 5831 8355 5837
rect 8297 5828 8309 5831
rect 7524 5800 8309 5828
rect 7524 5788 7530 5800
rect 8297 5797 8309 5800
rect 8343 5797 8355 5831
rect 8297 5791 8355 5797
rect 9674 5788 9680 5840
rect 9732 5788 9738 5840
rect 11974 5828 11980 5840
rect 11935 5800 11980 5828
rect 11974 5788 11980 5800
rect 12032 5788 12038 5840
rect 13725 5831 13783 5837
rect 13725 5797 13737 5831
rect 13771 5828 13783 5831
rect 14366 5828 14372 5840
rect 13771 5800 14372 5828
rect 13771 5797 13783 5800
rect 13725 5791 13783 5797
rect 14366 5788 14372 5800
rect 14424 5828 14430 5840
rect 15105 5831 15163 5837
rect 14424 5800 14688 5828
rect 14424 5788 14430 5800
rect 5258 5720 5264 5772
rect 5316 5760 5322 5772
rect 6457 5763 6515 5769
rect 6457 5760 6469 5763
rect 5316 5732 5580 5760
rect 5316 5720 5322 5732
rect 1578 5692 1584 5704
rect 1539 5664 1584 5692
rect 1578 5652 1584 5664
rect 1636 5652 1642 5704
rect 2041 5695 2099 5701
rect 2041 5661 2053 5695
rect 2087 5692 2099 5695
rect 3789 5695 3847 5701
rect 3789 5692 3801 5695
rect 2087 5664 3801 5692
rect 2087 5661 2099 5664
rect 2041 5655 2099 5661
rect 2976 5636 3004 5664
rect 3789 5661 3801 5664
rect 3835 5692 3847 5695
rect 4614 5692 4620 5704
rect 3835 5664 4620 5692
rect 3835 5661 3847 5664
rect 3789 5655 3847 5661
rect 4614 5652 4620 5664
rect 4672 5652 4678 5704
rect 5442 5692 5448 5704
rect 5403 5664 5448 5692
rect 5442 5652 5448 5664
rect 5500 5652 5506 5704
rect 5552 5692 5580 5732
rect 6012 5732 6469 5760
rect 5902 5692 5908 5704
rect 5552 5664 5908 5692
rect 5902 5652 5908 5664
rect 5960 5652 5966 5704
rect 1854 5584 1860 5636
rect 1912 5624 1918 5636
rect 2314 5633 2320 5636
rect 2286 5627 2320 5633
rect 2286 5624 2298 5627
rect 1912 5596 2298 5624
rect 1912 5584 1918 5596
rect 2286 5593 2298 5596
rect 2372 5624 2378 5636
rect 2372 5596 2434 5624
rect 2286 5587 2320 5593
rect 2314 5584 2320 5587
rect 2372 5584 2378 5596
rect 2958 5584 2964 5636
rect 3016 5584 3022 5636
rect 4056 5627 4114 5633
rect 4056 5593 4068 5627
rect 4102 5624 4114 5627
rect 4154 5624 4160 5636
rect 4102 5596 4160 5624
rect 4102 5593 4114 5596
rect 4056 5587 4114 5593
rect 4154 5584 4160 5596
rect 4212 5584 4218 5636
rect 5350 5584 5356 5636
rect 5408 5624 5414 5636
rect 6012 5624 6040 5732
rect 6457 5729 6469 5732
rect 6503 5729 6515 5763
rect 6638 5760 6644 5772
rect 6599 5732 6644 5760
rect 6457 5723 6515 5729
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 7282 5720 7288 5772
rect 7340 5760 7346 5772
rect 9490 5760 9496 5772
rect 7340 5732 8064 5760
rect 9451 5732 9496 5760
rect 7340 5720 7346 5732
rect 7558 5692 7564 5704
rect 7471 5664 7564 5692
rect 7558 5652 7564 5664
rect 7616 5652 7622 5704
rect 8036 5701 8064 5732
rect 9490 5720 9496 5732
rect 9548 5720 9554 5772
rect 9585 5763 9643 5769
rect 9585 5729 9597 5763
rect 9631 5760 9643 5763
rect 9692 5760 9720 5788
rect 9631 5732 9720 5760
rect 9631 5729 9643 5732
rect 9585 5723 9643 5729
rect 11698 5720 11704 5772
rect 11756 5760 11762 5772
rect 12342 5760 12348 5772
rect 11756 5732 12348 5760
rect 11756 5720 11762 5732
rect 12342 5720 12348 5732
rect 12400 5720 12406 5772
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14660 5769 14688 5800
rect 15105 5797 15117 5831
rect 15151 5797 15163 5831
rect 15105 5791 15163 5797
rect 14553 5763 14611 5769
rect 14553 5760 14565 5763
rect 13872 5732 14565 5760
rect 13872 5720 13878 5732
rect 14553 5729 14565 5732
rect 14599 5729 14611 5763
rect 14553 5723 14611 5729
rect 14645 5763 14703 5769
rect 14645 5729 14657 5763
rect 14691 5729 14703 5763
rect 15120 5760 15148 5791
rect 15672 5769 15700 5868
rect 15838 5856 15844 5908
rect 15896 5896 15902 5908
rect 18874 5896 18880 5908
rect 15896 5868 18552 5896
rect 18835 5868 18880 5896
rect 15896 5856 15902 5868
rect 16224 5769 16252 5868
rect 14645 5723 14703 5729
rect 14844 5732 15148 5760
rect 15657 5763 15715 5769
rect 8021 5695 8079 5701
rect 8021 5661 8033 5695
rect 8067 5692 8079 5695
rect 8110 5692 8116 5704
rect 8067 5664 8116 5692
rect 8067 5661 8079 5664
rect 8021 5655 8079 5661
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8386 5652 8392 5704
rect 8444 5692 8450 5704
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 8444 5664 8493 5692
rect 8444 5652 8450 5664
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 10318 5692 10324 5704
rect 9732 5664 10324 5692
rect 9732 5652 9738 5664
rect 10318 5652 10324 5664
rect 10376 5652 10382 5704
rect 10588 5695 10646 5701
rect 10588 5661 10600 5695
rect 10634 5692 10646 5695
rect 10962 5692 10968 5704
rect 10634 5664 10968 5692
rect 10634 5661 10646 5664
rect 10588 5655 10646 5661
rect 10962 5652 10968 5664
rect 11020 5652 11026 5704
rect 11974 5652 11980 5704
rect 12032 5692 12038 5704
rect 12434 5692 12440 5704
rect 12032 5664 12440 5692
rect 12032 5652 12038 5664
rect 12434 5652 12440 5664
rect 12492 5652 12498 5704
rect 12986 5652 12992 5704
rect 13044 5692 13050 5704
rect 13044 5664 13400 5692
rect 13044 5652 13050 5664
rect 5408 5596 6040 5624
rect 5408 5584 5414 5596
rect 6178 5584 6184 5636
rect 6236 5584 6242 5636
rect 2866 5516 2872 5568
rect 2924 5556 2930 5568
rect 3418 5556 3424 5568
rect 2924 5528 3424 5556
rect 2924 5516 2930 5528
rect 3418 5516 3424 5528
rect 3476 5516 3482 5568
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 6196 5556 6224 5584
rect 6730 5556 6736 5568
rect 4672 5528 6224 5556
rect 6691 5528 6736 5556
rect 4672 5516 4678 5528
rect 6730 5516 6736 5528
rect 6788 5516 6794 5568
rect 6914 5516 6920 5568
rect 6972 5556 6978 5568
rect 7576 5556 7604 5652
rect 12066 5624 12072 5636
rect 7852 5596 12072 5624
rect 7852 5568 7880 5596
rect 12066 5584 12072 5596
rect 12124 5584 12130 5636
rect 12612 5627 12670 5633
rect 12612 5593 12624 5627
rect 12658 5624 12670 5627
rect 12894 5624 12900 5636
rect 12658 5596 12900 5624
rect 12658 5593 12670 5596
rect 12612 5587 12670 5593
rect 12894 5584 12900 5596
rect 12952 5624 12958 5636
rect 13262 5624 13268 5636
rect 12952 5596 13268 5624
rect 12952 5584 12958 5596
rect 13262 5584 13268 5596
rect 13320 5584 13326 5636
rect 13372 5624 13400 5664
rect 14461 5627 14519 5633
rect 13372 5596 14412 5624
rect 7834 5556 7840 5568
rect 6972 5528 7604 5556
rect 7747 5528 7840 5556
rect 6972 5516 6978 5528
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 9398 5556 9404 5568
rect 9359 5528 9404 5556
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 11698 5556 11704 5568
rect 11659 5528 11704 5556
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 14093 5559 14151 5565
rect 14093 5525 14105 5559
rect 14139 5556 14151 5559
rect 14274 5556 14280 5568
rect 14139 5528 14280 5556
rect 14139 5525 14151 5528
rect 14093 5519 14151 5525
rect 14274 5516 14280 5528
rect 14332 5516 14338 5568
rect 14384 5556 14412 5596
rect 14461 5593 14473 5627
rect 14507 5624 14519 5627
rect 14844 5624 14872 5732
rect 15657 5729 15669 5763
rect 15703 5729 15715 5763
rect 15657 5723 15715 5729
rect 16209 5763 16267 5769
rect 16209 5729 16221 5763
rect 16255 5729 16267 5763
rect 16390 5760 16396 5772
rect 16351 5732 16396 5760
rect 16209 5723 16267 5729
rect 16390 5720 16396 5732
rect 16448 5720 16454 5772
rect 18524 5760 18552 5868
rect 18874 5856 18880 5868
rect 18932 5856 18938 5908
rect 20162 5856 20168 5908
rect 20220 5896 20226 5908
rect 20257 5899 20315 5905
rect 20257 5896 20269 5899
rect 20220 5868 20269 5896
rect 20220 5856 20226 5868
rect 20257 5865 20269 5868
rect 20303 5865 20315 5899
rect 20257 5859 20315 5865
rect 20438 5856 20444 5908
rect 20496 5896 20502 5908
rect 21269 5899 21327 5905
rect 21269 5896 21281 5899
rect 20496 5868 21281 5896
rect 20496 5856 20502 5868
rect 21269 5865 21281 5868
rect 21315 5865 21327 5899
rect 21269 5859 21327 5865
rect 18892 5828 18920 5856
rect 19242 5828 19248 5840
rect 18892 5800 19248 5828
rect 19242 5788 19248 5800
rect 19300 5788 19306 5840
rect 20714 5828 20720 5840
rect 19904 5800 20720 5828
rect 19797 5763 19855 5769
rect 19797 5760 19809 5763
rect 18524 5732 19809 5760
rect 19797 5729 19809 5732
rect 19843 5729 19855 5763
rect 19797 5723 19855 5729
rect 15470 5692 15476 5704
rect 15431 5664 15476 5692
rect 15470 5652 15476 5664
rect 15528 5652 15534 5704
rect 17494 5692 17500 5704
rect 17455 5664 17500 5692
rect 17494 5652 17500 5664
rect 17552 5652 17558 5704
rect 17770 5701 17776 5704
rect 17764 5692 17776 5701
rect 17731 5664 17776 5692
rect 17764 5655 17776 5664
rect 17770 5652 17776 5655
rect 17828 5652 17834 5704
rect 19518 5692 19524 5704
rect 17972 5664 19524 5692
rect 17972 5636 18000 5664
rect 19518 5652 19524 5664
rect 19576 5652 19582 5704
rect 19613 5695 19671 5701
rect 19613 5661 19625 5695
rect 19659 5692 19671 5695
rect 19904 5692 19932 5800
rect 20714 5788 20720 5800
rect 20772 5788 20778 5840
rect 20530 5720 20536 5772
rect 20588 5760 20594 5772
rect 20809 5763 20867 5769
rect 20809 5760 20821 5763
rect 20588 5732 20821 5760
rect 20588 5720 20594 5732
rect 20809 5729 20821 5732
rect 20855 5729 20867 5763
rect 20809 5723 20867 5729
rect 20622 5692 20628 5704
rect 19659 5664 19932 5692
rect 20583 5664 20628 5692
rect 19659 5661 19671 5664
rect 19613 5655 19671 5661
rect 20622 5652 20628 5664
rect 20680 5652 20686 5704
rect 14507 5596 14872 5624
rect 14507 5593 14519 5596
rect 14461 5587 14519 5593
rect 15286 5584 15292 5636
rect 15344 5624 15350 5636
rect 16485 5627 16543 5633
rect 16485 5624 16497 5627
rect 15344 5596 16497 5624
rect 15344 5584 15350 5596
rect 16485 5593 16497 5596
rect 16531 5593 16543 5627
rect 17586 5624 17592 5636
rect 16485 5587 16543 5593
rect 16868 5596 17592 5624
rect 16868 5565 16896 5596
rect 17586 5584 17592 5596
rect 17644 5584 17650 5636
rect 17954 5584 17960 5636
rect 18012 5584 18018 5636
rect 18690 5584 18696 5636
rect 18748 5624 18754 5636
rect 20717 5627 20775 5633
rect 20717 5624 20729 5627
rect 18748 5596 20729 5624
rect 18748 5584 18754 5596
rect 20717 5593 20729 5596
rect 20763 5593 20775 5627
rect 20717 5587 20775 5593
rect 15565 5559 15623 5565
rect 15565 5556 15577 5559
rect 14384 5528 15577 5556
rect 15565 5525 15577 5528
rect 15611 5525 15623 5559
rect 15565 5519 15623 5525
rect 16853 5559 16911 5565
rect 16853 5525 16865 5559
rect 16899 5525 16911 5559
rect 16853 5519 16911 5525
rect 17034 5516 17040 5568
rect 17092 5556 17098 5568
rect 17221 5559 17279 5565
rect 17221 5556 17233 5559
rect 17092 5528 17233 5556
rect 17092 5516 17098 5528
rect 17221 5525 17233 5528
rect 17267 5556 17279 5559
rect 17862 5556 17868 5568
rect 17267 5528 17868 5556
rect 17267 5525 17279 5528
rect 17221 5519 17279 5525
rect 17862 5516 17868 5528
rect 17920 5516 17926 5568
rect 18966 5516 18972 5568
rect 19024 5556 19030 5568
rect 19245 5559 19303 5565
rect 19245 5556 19257 5559
rect 19024 5528 19257 5556
rect 19024 5516 19030 5528
rect 19245 5525 19257 5528
rect 19291 5525 19303 5559
rect 19245 5519 19303 5525
rect 19518 5516 19524 5568
rect 19576 5556 19582 5568
rect 19705 5559 19763 5565
rect 19705 5556 19717 5559
rect 19576 5528 19717 5556
rect 19576 5516 19582 5528
rect 19705 5525 19717 5528
rect 19751 5556 19763 5559
rect 20254 5556 20260 5568
rect 19751 5528 20260 5556
rect 19751 5525 19763 5528
rect 19705 5519 19763 5525
rect 20254 5516 20260 5528
rect 20312 5516 20318 5568
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2961 5355 3019 5361
rect 2961 5352 2973 5355
rect 2455 5324 2973 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2961 5321 2973 5324
rect 3007 5321 3019 5355
rect 2961 5315 3019 5321
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3697 5355 3755 5361
rect 3108 5324 3153 5352
rect 3108 5312 3114 5324
rect 3697 5321 3709 5355
rect 3743 5321 3755 5355
rect 3697 5315 3755 5321
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 5902 5352 5908 5364
rect 4111 5324 5908 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 2041 5287 2099 5293
rect 2041 5253 2053 5287
rect 2087 5284 2099 5287
rect 3712 5284 3740 5315
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6457 5355 6515 5361
rect 6457 5321 6469 5355
rect 6503 5352 6515 5355
rect 6730 5352 6736 5364
rect 6503 5324 6736 5352
rect 6503 5321 6515 5324
rect 6457 5315 6515 5321
rect 6730 5312 6736 5324
rect 6788 5312 6794 5364
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 7834 5352 7840 5364
rect 6963 5324 7840 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 5721 5287 5779 5293
rect 5721 5284 5733 5287
rect 2087 5256 3740 5284
rect 3804 5256 5733 5284
rect 2087 5253 2099 5256
rect 2041 5247 2099 5253
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3804 5216 3832 5256
rect 5721 5253 5733 5256
rect 5767 5253 5779 5287
rect 5721 5247 5779 5253
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 6932 5284 6960 5315
rect 7834 5312 7840 5324
rect 7892 5312 7898 5364
rect 10689 5355 10747 5361
rect 10689 5321 10701 5355
rect 10735 5352 10747 5355
rect 11146 5352 11152 5364
rect 10735 5324 11152 5352
rect 10735 5321 10747 5324
rect 10689 5315 10747 5321
rect 11146 5312 11152 5324
rect 11204 5312 11210 5364
rect 13538 5312 13544 5364
rect 13596 5352 13602 5364
rect 13596 5324 15700 5352
rect 13596 5312 13602 5324
rect 5868 5256 6960 5284
rect 5868 5244 5874 5256
rect 8478 5244 8484 5296
rect 8536 5284 8542 5296
rect 9585 5287 9643 5293
rect 9585 5284 9597 5287
rect 8536 5256 9597 5284
rect 8536 5244 8542 5256
rect 9585 5253 9597 5256
rect 9631 5253 9643 5287
rect 9585 5247 9643 5253
rect 10781 5287 10839 5293
rect 10781 5253 10793 5287
rect 10827 5284 10839 5287
rect 11238 5284 11244 5296
rect 10827 5256 11244 5284
rect 10827 5253 10839 5256
rect 10781 5247 10839 5253
rect 11238 5244 11244 5256
rect 11296 5244 11302 5296
rect 12342 5244 12348 5296
rect 12400 5284 12406 5296
rect 12986 5284 12992 5296
rect 12400 5256 12992 5284
rect 12400 5244 12406 5256
rect 12986 5244 12992 5256
rect 13044 5244 13050 5296
rect 14737 5287 14795 5293
rect 14737 5253 14749 5287
rect 14783 5284 14795 5287
rect 15562 5284 15568 5296
rect 14783 5256 15568 5284
rect 14783 5253 14795 5256
rect 14737 5247 14795 5253
rect 15562 5244 15568 5256
rect 15620 5244 15626 5296
rect 15672 5284 15700 5324
rect 16114 5312 16120 5364
rect 16172 5352 16178 5364
rect 16390 5352 16396 5364
rect 16172 5324 16396 5352
rect 16172 5312 16178 5324
rect 16390 5312 16396 5324
rect 16448 5312 16454 5364
rect 16942 5352 16948 5364
rect 16868 5324 16948 5352
rect 15838 5284 15844 5296
rect 15672 5256 15844 5284
rect 3384 5188 3832 5216
rect 3384 5176 3390 5188
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4028 5188 4108 5216
rect 4028 5176 4034 5188
rect 1486 5108 1492 5160
rect 1544 5148 1550 5160
rect 1765 5151 1823 5157
rect 1765 5148 1777 5151
rect 1544 5120 1777 5148
rect 1544 5108 1550 5120
rect 1765 5117 1777 5120
rect 1811 5148 1823 5151
rect 1854 5148 1860 5160
rect 1811 5120 1860 5148
rect 1811 5117 1823 5120
rect 1765 5111 1823 5117
rect 1854 5108 1860 5120
rect 1912 5108 1918 5160
rect 1949 5151 2007 5157
rect 1949 5117 1961 5151
rect 1995 5148 2007 5151
rect 2498 5148 2504 5160
rect 1995 5120 2504 5148
rect 1995 5117 2007 5120
rect 1949 5111 2007 5117
rect 2498 5108 2504 5120
rect 2556 5108 2562 5160
rect 2866 5148 2872 5160
rect 2827 5120 2872 5148
rect 2866 5108 2872 5120
rect 2924 5108 2930 5160
rect 4080 5148 4108 5188
rect 4430 5176 4436 5228
rect 4488 5216 4494 5228
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4488 5188 4721 5216
rect 4488 5176 4494 5188
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4709 5179 4767 5185
rect 5994 5176 6000 5228
rect 6052 5216 6058 5228
rect 6454 5216 6460 5228
rect 6052 5188 6460 5216
rect 6052 5176 6058 5188
rect 6454 5176 6460 5188
rect 6512 5216 6518 5228
rect 6825 5219 6883 5225
rect 6825 5216 6837 5219
rect 6512 5188 6837 5216
rect 6512 5176 6518 5188
rect 6825 5185 6837 5188
rect 6871 5185 6883 5219
rect 6825 5179 6883 5185
rect 7561 5219 7619 5225
rect 7561 5185 7573 5219
rect 7607 5216 7619 5219
rect 9490 5216 9496 5228
rect 7607 5188 9496 5216
rect 7607 5185 7619 5188
rect 7561 5179 7619 5185
rect 9490 5176 9496 5188
rect 9548 5216 9554 5228
rect 9861 5219 9919 5225
rect 9861 5216 9873 5219
rect 9548 5188 9873 5216
rect 9548 5176 9554 5188
rect 9861 5185 9873 5188
rect 9907 5185 9919 5219
rect 11698 5216 11704 5228
rect 9861 5179 9919 5185
rect 10612 5188 11704 5216
rect 10612 5157 10640 5188
rect 11698 5176 11704 5188
rect 11756 5176 11762 5228
rect 15672 5225 15700 5256
rect 15838 5244 15844 5256
rect 15896 5244 15902 5296
rect 15197 5219 15255 5225
rect 15197 5185 15209 5219
rect 15243 5216 15255 5219
rect 15657 5219 15715 5225
rect 15243 5188 15608 5216
rect 15243 5185 15255 5188
rect 15197 5179 15255 5185
rect 4157 5151 4215 5157
rect 4157 5148 4169 5151
rect 4080 5120 4169 5148
rect 4157 5117 4169 5120
rect 4203 5117 4215 5151
rect 4157 5111 4215 5117
rect 4249 5151 4307 5157
rect 4249 5117 4261 5151
rect 4295 5117 4307 5151
rect 7009 5151 7067 5157
rect 7009 5148 7021 5151
rect 4249 5111 4307 5117
rect 6840 5120 7021 5148
rect 2590 5040 2596 5092
rect 2648 5080 2654 5092
rect 4264 5080 4292 5111
rect 6840 5092 6868 5120
rect 7009 5117 7021 5120
rect 7055 5117 7067 5151
rect 7009 5111 7067 5117
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5117 10655 5151
rect 15286 5148 15292 5160
rect 10597 5111 10655 5117
rect 12406 5120 15292 5148
rect 5718 5080 5724 5092
rect 2648 5052 4292 5080
rect 5184 5052 5724 5080
rect 2648 5040 2654 5052
rect 3326 5012 3332 5024
rect 952 4984 3332 5012
rect 952 4888 980 4984
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 5184 5012 5212 5052
rect 5718 5040 5724 5052
rect 5776 5040 5782 5092
rect 6822 5040 6828 5092
rect 6880 5040 6886 5092
rect 9214 5080 9220 5092
rect 8128 5052 9220 5080
rect 5350 5012 5356 5024
rect 3467 4984 5212 5012
rect 5311 4984 5356 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 5350 4972 5356 4984
rect 5408 4972 5414 5024
rect 5813 5015 5871 5021
rect 5813 4981 5825 5015
rect 5859 5012 5871 5015
rect 8128 5012 8156 5052
rect 9214 5040 9220 5052
rect 9272 5040 9278 5092
rect 9398 5040 9404 5092
rect 9456 5080 9462 5092
rect 10045 5083 10103 5089
rect 10045 5080 10057 5083
rect 9456 5052 10057 5080
rect 9456 5040 9462 5052
rect 10045 5049 10057 5052
rect 10091 5080 10103 5083
rect 12406 5080 12434 5120
rect 15286 5108 15292 5120
rect 15344 5108 15350 5160
rect 10091 5052 12434 5080
rect 10091 5049 10103 5052
rect 10045 5043 10103 5049
rect 13078 5040 13084 5092
rect 13136 5080 13142 5092
rect 15473 5083 15531 5089
rect 15473 5080 15485 5083
rect 13136 5052 15485 5080
rect 13136 5040 13142 5052
rect 15473 5049 15485 5052
rect 15519 5049 15531 5083
rect 15580 5080 15608 5188
rect 15657 5185 15669 5219
rect 15703 5185 15715 5219
rect 15930 5216 15936 5228
rect 15891 5188 15936 5216
rect 15657 5179 15715 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16868 5157 16896 5324
rect 16942 5312 16948 5324
rect 17000 5312 17006 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17405 5355 17463 5361
rect 17405 5352 17417 5355
rect 17184 5324 17417 5352
rect 17184 5312 17190 5324
rect 17405 5321 17417 5324
rect 17451 5321 17463 5355
rect 17405 5315 17463 5321
rect 17586 5312 17592 5364
rect 17644 5352 17650 5364
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 17644 5324 18337 5352
rect 17644 5312 17650 5324
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 18690 5352 18696 5364
rect 18651 5324 18696 5352
rect 18325 5315 18383 5321
rect 18690 5312 18696 5324
rect 18748 5312 18754 5364
rect 20349 5355 20407 5361
rect 20349 5321 20361 5355
rect 20395 5352 20407 5355
rect 20530 5352 20536 5364
rect 20395 5324 20536 5352
rect 20395 5321 20407 5324
rect 20349 5315 20407 5321
rect 20530 5312 20536 5324
rect 20588 5312 20594 5364
rect 17034 5284 17040 5296
rect 16995 5256 17040 5284
rect 17034 5244 17040 5256
rect 17092 5244 17098 5296
rect 17494 5244 17500 5296
rect 17552 5284 17558 5296
rect 21174 5284 21180 5296
rect 17552 5256 21180 5284
rect 17552 5244 17558 5256
rect 17770 5176 17776 5228
rect 17828 5216 17834 5228
rect 17954 5216 17960 5228
rect 17828 5188 17960 5216
rect 17828 5176 17834 5188
rect 17954 5176 17960 5188
rect 18012 5176 18018 5228
rect 18233 5219 18291 5225
rect 18233 5185 18245 5219
rect 18279 5216 18291 5219
rect 18874 5216 18880 5228
rect 18279 5188 18880 5216
rect 18279 5185 18291 5188
rect 18233 5179 18291 5185
rect 18874 5176 18880 5188
rect 18932 5176 18938 5228
rect 18984 5225 19012 5256
rect 21174 5244 21180 5256
rect 21232 5244 21238 5296
rect 19242 5225 19248 5228
rect 18969 5219 19027 5225
rect 18969 5185 18981 5219
rect 19015 5185 19027 5219
rect 19236 5216 19248 5225
rect 18969 5179 19027 5185
rect 19076 5188 19248 5216
rect 16853 5151 16911 5157
rect 16853 5117 16865 5151
rect 16899 5117 16911 5151
rect 16853 5111 16911 5117
rect 16942 5108 16948 5160
rect 17000 5148 17006 5160
rect 18141 5151 18199 5157
rect 17000 5120 17045 5148
rect 17000 5108 17006 5120
rect 18141 5117 18153 5151
rect 18187 5148 18199 5151
rect 19076 5148 19104 5188
rect 19236 5179 19248 5188
rect 19242 5176 19248 5179
rect 19300 5176 19306 5228
rect 20530 5176 20536 5228
rect 20588 5216 20594 5228
rect 20625 5219 20683 5225
rect 20625 5216 20637 5219
rect 20588 5188 20637 5216
rect 20588 5176 20594 5188
rect 20625 5185 20637 5188
rect 20671 5185 20683 5219
rect 20625 5179 20683 5185
rect 18187 5120 19104 5148
rect 18187 5117 18199 5120
rect 18141 5111 18199 5117
rect 17954 5080 17960 5092
rect 15580 5052 17960 5080
rect 15473 5043 15531 5049
rect 17954 5040 17960 5052
rect 18012 5040 18018 5092
rect 8294 5012 8300 5024
rect 5859 4984 8156 5012
rect 8255 4984 8300 5012
rect 5859 4981 5871 4984
rect 5813 4975 5871 4981
rect 8294 4972 8300 4984
rect 8352 5012 8358 5024
rect 9582 5012 9588 5024
rect 8352 4984 9588 5012
rect 8352 4972 8358 4984
rect 9582 4972 9588 4984
rect 9640 4972 9646 5024
rect 11149 5015 11207 5021
rect 11149 4981 11161 5015
rect 11195 5012 11207 5015
rect 11238 5012 11244 5024
rect 11195 4984 11244 5012
rect 11195 4981 11207 4984
rect 11149 4975 11207 4981
rect 11238 4972 11244 4984
rect 11296 4972 11302 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12345 5015 12403 5021
rect 12345 5012 12357 5015
rect 11848 4984 12357 5012
rect 11848 4972 11854 4984
rect 12345 4981 12357 4984
rect 12391 4981 12403 5015
rect 12345 4975 12403 4981
rect 12434 4972 12440 5024
rect 12492 5012 12498 5024
rect 12621 5015 12679 5021
rect 12621 5012 12633 5015
rect 12492 4984 12633 5012
rect 12492 4972 12498 4984
rect 12621 4981 12633 4984
rect 12667 4981 12679 5015
rect 12621 4975 12679 4981
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 15013 5015 15071 5021
rect 15013 5012 15025 5015
rect 13596 4984 15025 5012
rect 13596 4972 13602 4984
rect 15013 4981 15025 4984
rect 15059 4981 15071 5015
rect 16114 5012 16120 5024
rect 16075 4984 16120 5012
rect 15013 4975 15071 4981
rect 16114 4972 16120 4984
rect 16172 4972 16178 5024
rect 21266 5012 21272 5024
rect 21227 4984 21272 5012
rect 21266 4972 21272 4984
rect 21324 4972 21330 5024
rect 1104 4922 21896 4944
rect 198 4836 204 4888
rect 256 4876 262 4888
rect 934 4876 940 4888
rect 256 4848 940 4876
rect 256 4836 262 4848
rect 934 4836 940 4848
rect 992 4836 998 4888
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 2498 4808 2504 4820
rect 2459 4780 2504 4808
rect 2498 4768 2504 4780
rect 2556 4768 2562 4820
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 4430 4808 4436 4820
rect 3936 4780 4436 4808
rect 3936 4768 3942 4780
rect 4430 4768 4436 4780
rect 4488 4768 4494 4820
rect 6273 4811 6331 4817
rect 6273 4777 6285 4811
rect 6319 4808 6331 4811
rect 6822 4808 6828 4820
rect 6319 4780 6828 4808
rect 6319 4777 6331 4780
rect 6273 4771 6331 4777
rect 6822 4768 6828 4780
rect 6880 4808 6886 4820
rect 8386 4808 8392 4820
rect 6880 4780 8392 4808
rect 6880 4768 6886 4780
rect 8386 4768 8392 4780
rect 8444 4768 8450 4820
rect 10321 4811 10379 4817
rect 10321 4777 10333 4811
rect 10367 4808 10379 4811
rect 12250 4808 12256 4820
rect 10367 4780 12256 4808
rect 10367 4777 10379 4780
rect 10321 4771 10379 4777
rect 12250 4768 12256 4780
rect 12308 4768 12314 4820
rect 12894 4808 12900 4820
rect 12855 4780 12900 4808
rect 12894 4768 12900 4780
rect 12952 4768 12958 4820
rect 13357 4811 13415 4817
rect 13357 4777 13369 4811
rect 13403 4808 13415 4811
rect 13403 4780 15056 4808
rect 13403 4777 13415 4780
rect 13357 4771 13415 4777
rect 1946 4700 1952 4752
rect 2004 4740 2010 4752
rect 2004 4712 5672 4740
rect 2004 4700 2010 4712
rect 2222 4672 2228 4684
rect 2183 4644 2228 4672
rect 2222 4632 2228 4644
rect 2280 4632 2286 4684
rect 2590 4632 2596 4684
rect 2648 4672 2654 4684
rect 3053 4675 3111 4681
rect 3053 4672 3065 4675
rect 2648 4644 3065 4672
rect 2648 4632 2654 4644
rect 3053 4641 3065 4644
rect 3099 4641 3111 4675
rect 3053 4635 3111 4641
rect 4341 4675 4399 4681
rect 4341 4641 4353 4675
rect 4387 4641 4399 4675
rect 4341 4635 4399 4641
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4672 4491 4675
rect 4798 4672 4804 4684
rect 4479 4644 4804 4672
rect 4479 4641 4491 4644
rect 4433 4635 4491 4641
rect 1949 4607 2007 4613
rect 1949 4573 1961 4607
rect 1995 4604 2007 4607
rect 2130 4604 2136 4616
rect 1995 4576 2136 4604
rect 1995 4573 2007 4576
rect 1949 4567 2007 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 2961 4607 3019 4613
rect 2961 4573 2973 4607
rect 3007 4604 3019 4607
rect 3970 4604 3976 4616
rect 3007 4576 3976 4604
rect 3007 4573 3019 4576
rect 2961 4567 3019 4573
rect 3970 4564 3976 4576
rect 4028 4564 4034 4616
rect 4356 4604 4384 4635
rect 4798 4632 4804 4644
rect 4856 4632 4862 4684
rect 5644 4681 5672 4712
rect 5902 4700 5908 4752
rect 5960 4740 5966 4752
rect 7193 4743 7251 4749
rect 7193 4740 7205 4743
rect 5960 4712 7205 4740
rect 5960 4700 5966 4712
rect 7193 4709 7205 4712
rect 7239 4740 7251 4743
rect 10962 4740 10968 4752
rect 7239 4712 10968 4740
rect 7239 4709 7251 4712
rect 7193 4703 7251 4709
rect 10962 4700 10968 4712
rect 11020 4700 11026 4752
rect 15028 4740 15056 4780
rect 15286 4768 15292 4820
rect 15344 4808 15350 4820
rect 17221 4811 17279 4817
rect 17221 4808 17233 4811
rect 15344 4780 17233 4808
rect 15344 4768 15350 4780
rect 17221 4777 17233 4780
rect 17267 4777 17279 4811
rect 17678 4808 17684 4820
rect 17639 4780 17684 4808
rect 17221 4771 17279 4777
rect 17678 4768 17684 4780
rect 17736 4768 17742 4820
rect 17770 4740 17776 4752
rect 15028 4712 17776 4740
rect 17770 4700 17776 4712
rect 17828 4700 17834 4752
rect 18046 4740 18052 4752
rect 18007 4712 18052 4740
rect 18046 4700 18052 4712
rect 18104 4700 18110 4752
rect 19429 4743 19487 4749
rect 19429 4709 19441 4743
rect 19475 4740 19487 4743
rect 19978 4740 19984 4752
rect 19475 4712 19984 4740
rect 19475 4709 19487 4712
rect 19429 4703 19487 4709
rect 19978 4700 19984 4712
rect 20036 4700 20042 4752
rect 5629 4675 5687 4681
rect 5629 4641 5641 4675
rect 5675 4641 5687 4675
rect 5629 4635 5687 4641
rect 5813 4675 5871 4681
rect 5813 4641 5825 4675
rect 5859 4672 5871 4675
rect 6546 4672 6552 4684
rect 5859 4644 6552 4672
rect 5859 4641 5871 4644
rect 5813 4635 5871 4641
rect 5828 4604 5856 4635
rect 6546 4632 6552 4644
rect 6604 4632 6610 4684
rect 6730 4632 6736 4684
rect 6788 4672 6794 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 6788 4644 7941 4672
rect 6788 4632 6794 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 7929 4635 7987 4641
rect 9214 4632 9220 4684
rect 9272 4672 9278 4684
rect 9401 4675 9459 4681
rect 9401 4672 9413 4675
rect 9272 4644 9413 4672
rect 9272 4632 9278 4644
rect 9401 4641 9413 4644
rect 9447 4641 9459 4675
rect 9582 4672 9588 4684
rect 9543 4644 9588 4672
rect 9401 4635 9459 4641
rect 9582 4632 9588 4644
rect 9640 4632 9646 4684
rect 12986 4632 12992 4684
rect 13044 4672 13050 4684
rect 14090 4672 14096 4684
rect 13044 4644 14096 4672
rect 13044 4632 13050 4644
rect 14090 4632 14096 4644
rect 14148 4632 14154 4684
rect 16114 4632 16120 4684
rect 16172 4672 16178 4684
rect 21174 4672 21180 4684
rect 16172 4644 19288 4672
rect 21135 4644 21180 4672
rect 16172 4632 16178 4644
rect 7006 4604 7012 4616
rect 4356 4576 5856 4604
rect 6967 4576 7012 4604
rect 7006 4564 7012 4576
rect 7064 4564 7070 4616
rect 7469 4607 7527 4613
rect 7469 4573 7481 4607
rect 7515 4604 7527 4607
rect 7558 4604 7564 4616
rect 7515 4576 7564 4604
rect 7515 4573 7527 4576
rect 7469 4567 7527 4573
rect 7558 4564 7564 4576
rect 7616 4564 7622 4616
rect 8573 4607 8631 4613
rect 8573 4573 8585 4607
rect 8619 4604 8631 4607
rect 9122 4604 9128 4616
rect 8619 4576 9128 4604
rect 8619 4573 8631 4576
rect 8573 4567 8631 4573
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 10134 4604 10140 4616
rect 10095 4576 10140 4604
rect 10134 4564 10140 4576
rect 10192 4564 10198 4616
rect 10597 4607 10655 4613
rect 10597 4573 10609 4607
rect 10643 4604 10655 4607
rect 11146 4604 11152 4616
rect 10643 4576 11152 4604
rect 10643 4573 10655 4576
rect 10597 4567 10655 4573
rect 11146 4564 11152 4576
rect 11204 4564 11210 4616
rect 11517 4607 11575 4613
rect 11517 4573 11529 4607
rect 11563 4604 11575 4607
rect 13004 4604 13032 4632
rect 11563 4576 13032 4604
rect 13173 4607 13231 4613
rect 11563 4573 11575 4576
rect 11517 4567 11575 4573
rect 13173 4573 13185 4607
rect 13219 4604 13231 4607
rect 13814 4604 13820 4616
rect 13219 4576 13820 4604
rect 13219 4573 13231 4576
rect 13173 4567 13231 4573
rect 13814 4564 13820 4576
rect 13872 4564 13878 4616
rect 14360 4607 14418 4613
rect 14360 4573 14372 4607
rect 14406 4604 14418 4607
rect 14734 4604 14740 4616
rect 14406 4576 14740 4604
rect 14406 4573 14418 4576
rect 14360 4567 14418 4573
rect 14734 4564 14740 4576
rect 14792 4564 14798 4616
rect 15746 4604 15752 4616
rect 15707 4576 15752 4604
rect 15746 4564 15752 4576
rect 15804 4564 15810 4616
rect 16298 4604 16304 4616
rect 16259 4576 16304 4604
rect 16298 4564 16304 4576
rect 16356 4564 16362 4616
rect 17402 4604 17408 4616
rect 17363 4576 17408 4604
rect 17402 4564 17408 4576
rect 17460 4564 17466 4616
rect 18877 4607 18935 4613
rect 17512 4576 18368 4604
rect 3326 4496 3332 4548
rect 3384 4536 3390 4548
rect 11790 4545 11796 4548
rect 5537 4539 5595 4545
rect 5537 4536 5549 4539
rect 3384 4508 5549 4536
rect 3384 4496 3390 4508
rect 5537 4505 5549 4508
rect 5583 4505 5595 4539
rect 5537 4499 5595 4505
rect 6733 4539 6791 4545
rect 6733 4505 6745 4539
rect 6779 4536 6791 4539
rect 9309 4539 9367 4545
rect 9309 4536 9321 4539
rect 6779 4508 9321 4536
rect 6779 4505 6791 4508
rect 6733 4499 6791 4505
rect 9309 4505 9321 4508
rect 9355 4505 9367 4539
rect 11784 4536 11796 4545
rect 11751 4508 11796 4536
rect 9309 4499 9367 4505
rect 11784 4499 11796 4508
rect 11790 4496 11796 4499
rect 11848 4496 11854 4548
rect 12066 4496 12072 4548
rect 12124 4536 12130 4548
rect 17512 4536 17540 4576
rect 12124 4508 17540 4536
rect 18233 4539 18291 4545
rect 12124 4496 12130 4508
rect 18233 4505 18245 4539
rect 18279 4505 18291 4539
rect 18340 4536 18368 4576
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19058 4604 19064 4616
rect 18923 4576 19064 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 19058 4564 19064 4576
rect 19116 4564 19122 4616
rect 19260 4613 19288 4644
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 19245 4567 19303 4573
rect 20921 4607 20979 4613
rect 20921 4573 20933 4607
rect 20967 4604 20979 4607
rect 21266 4604 21272 4616
rect 20967 4576 21272 4604
rect 20967 4573 20979 4576
rect 20921 4567 20979 4573
rect 21266 4564 21272 4576
rect 21324 4564 21330 4616
rect 18340 4508 19840 4536
rect 18233 4499 18291 4505
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 3234 4468 3240 4480
rect 2915 4440 3240 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 3234 4428 3240 4440
rect 3292 4428 3298 4480
rect 3881 4471 3939 4477
rect 3881 4437 3893 4471
rect 3927 4468 3939 4471
rect 4062 4468 4068 4480
rect 3927 4440 4068 4468
rect 3927 4437 3939 4440
rect 3881 4431 3939 4437
rect 4062 4428 4068 4440
rect 4120 4428 4126 4480
rect 4522 4428 4528 4480
rect 4580 4468 4586 4480
rect 4890 4468 4896 4480
rect 4580 4440 4625 4468
rect 4851 4440 4896 4468
rect 4580 4428 4586 4440
rect 4890 4428 4896 4440
rect 4948 4428 4954 4480
rect 5166 4468 5172 4480
rect 5127 4440 5172 4468
rect 5166 4428 5172 4440
rect 5224 4428 5230 4480
rect 7098 4428 7104 4480
rect 7156 4468 7162 4480
rect 7653 4471 7711 4477
rect 7653 4468 7665 4471
rect 7156 4440 7665 4468
rect 7156 4428 7162 4440
rect 7653 4437 7665 4440
rect 7699 4437 7711 4471
rect 7653 4431 7711 4437
rect 8386 4428 8392 4480
rect 8444 4468 8450 4480
rect 8941 4471 8999 4477
rect 8941 4468 8953 4471
rect 8444 4440 8953 4468
rect 8444 4428 8450 4440
rect 8941 4437 8953 4440
rect 8987 4437 8999 4471
rect 10778 4468 10784 4480
rect 10739 4440 10784 4468
rect 8941 4431 8999 4437
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11241 4471 11299 4477
rect 11241 4437 11253 4471
rect 11287 4468 11299 4471
rect 11882 4468 11888 4480
rect 11287 4440 11888 4468
rect 11287 4437 11299 4440
rect 11241 4431 11299 4437
rect 11882 4428 11888 4440
rect 11940 4428 11946 4480
rect 13725 4471 13783 4477
rect 13725 4437 13737 4471
rect 13771 4468 13783 4471
rect 13814 4468 13820 4480
rect 13771 4440 13820 4468
rect 13771 4437 13783 4440
rect 13725 4431 13783 4437
rect 13814 4428 13820 4440
rect 13872 4468 13878 4480
rect 14366 4468 14372 4480
rect 13872 4440 14372 4468
rect 13872 4428 13878 4440
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 15194 4428 15200 4480
rect 15252 4468 15258 4480
rect 15473 4471 15531 4477
rect 15473 4468 15485 4471
rect 15252 4440 15485 4468
rect 15252 4428 15258 4440
rect 15473 4437 15485 4440
rect 15519 4437 15531 4471
rect 15930 4468 15936 4480
rect 15891 4440 15936 4468
rect 15473 4431 15531 4437
rect 15930 4428 15936 4440
rect 15988 4428 15994 4480
rect 16942 4468 16948 4480
rect 16903 4440 16948 4468
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 18248 4468 18276 4499
rect 18506 4468 18512 4480
rect 18248 4440 18512 4468
rect 18506 4428 18512 4440
rect 18564 4428 18570 4480
rect 18690 4468 18696 4480
rect 18651 4440 18696 4468
rect 18690 4428 18696 4440
rect 18748 4428 18754 4480
rect 19812 4477 19840 4508
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4437 19855 4471
rect 19797 4431 19855 4437
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 1486 4264 1492 4276
rect 1447 4236 1492 4264
rect 1486 4224 1492 4236
rect 1544 4224 1550 4276
rect 3326 4264 3332 4276
rect 3287 4236 3332 4264
rect 3326 4224 3332 4236
rect 3384 4224 3390 4276
rect 4614 4264 4620 4276
rect 3804 4236 4620 4264
rect 1946 4156 1952 4208
rect 2004 4196 2010 4208
rect 3804 4196 3832 4236
rect 4614 4224 4620 4236
rect 4672 4264 4678 4276
rect 6733 4267 6791 4273
rect 6733 4264 6745 4267
rect 4672 4236 6745 4264
rect 4672 4224 4678 4236
rect 6733 4233 6745 4236
rect 6779 4233 6791 4267
rect 6733 4227 6791 4233
rect 8389 4267 8447 4273
rect 8389 4233 8401 4267
rect 8435 4264 8447 4267
rect 8662 4264 8668 4276
rect 8435 4236 8668 4264
rect 8435 4233 8447 4236
rect 8389 4227 8447 4233
rect 8662 4224 8668 4236
rect 8720 4224 8726 4276
rect 10502 4224 10508 4276
rect 10560 4264 10566 4276
rect 10689 4267 10747 4273
rect 10689 4264 10701 4267
rect 10560 4236 10701 4264
rect 10560 4224 10566 4236
rect 10689 4233 10701 4236
rect 10735 4264 10747 4267
rect 10870 4264 10876 4276
rect 10735 4236 10876 4264
rect 10735 4233 10747 4236
rect 10689 4227 10747 4233
rect 10870 4224 10876 4236
rect 10928 4224 10934 4276
rect 11146 4224 11152 4276
rect 11204 4264 11210 4276
rect 11977 4267 12035 4273
rect 11977 4264 11989 4267
rect 11204 4236 11989 4264
rect 11204 4224 11210 4236
rect 11977 4233 11989 4236
rect 12023 4233 12035 4267
rect 11977 4227 12035 4233
rect 14090 4224 14096 4276
rect 14148 4264 14154 4276
rect 18049 4267 18107 4273
rect 14148 4236 14964 4264
rect 14148 4224 14154 4236
rect 2004 4168 3832 4196
rect 2004 4156 2010 4168
rect 3878 4156 3884 4208
rect 3936 4156 3942 4208
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 4798 4196 4804 4208
rect 4488 4168 4804 4196
rect 4488 4156 4494 4168
rect 4798 4156 4804 4168
rect 4856 4156 4862 4208
rect 4985 4199 5043 4205
rect 4985 4165 4997 4199
rect 5031 4196 5043 4199
rect 5166 4196 5172 4208
rect 5031 4168 5172 4196
rect 5031 4165 5043 4168
rect 4985 4159 5043 4165
rect 5166 4156 5172 4168
rect 5224 4156 5230 4208
rect 6638 4196 6644 4208
rect 6599 4168 6644 4196
rect 6638 4156 6644 4168
rect 6696 4156 6702 4208
rect 9582 4196 9588 4208
rect 8680 4168 9588 4196
rect 1578 4088 1584 4140
rect 1636 4128 1642 4140
rect 2590 4128 2596 4140
rect 2648 4137 2654 4140
rect 1636 4100 2596 4128
rect 1636 4088 1642 4100
rect 2590 4088 2596 4100
rect 2648 4091 2660 4137
rect 3896 4128 3924 4156
rect 3712 4100 3924 4128
rect 3973 4131 4031 4137
rect 2648 4088 2654 4091
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 2958 4060 2964 4072
rect 2915 4032 2964 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 2958 4020 2964 4032
rect 3016 4020 3022 4072
rect 3712 4069 3740 4100
rect 3973 4097 3985 4131
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 3697 4063 3755 4069
rect 3697 4029 3709 4063
rect 3743 4029 3755 4063
rect 3878 4060 3884 4072
rect 3839 4032 3884 4060
rect 3697 4023 3755 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 3988 3992 4016 4091
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 5813 4131 5871 4137
rect 5813 4128 5825 4131
rect 5776 4100 5825 4128
rect 5776 4088 5782 4100
rect 5813 4097 5825 4100
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 6086 4088 6092 4140
rect 6144 4128 6150 4140
rect 7377 4131 7435 4137
rect 6144 4100 6500 4128
rect 6144 4088 6150 4100
rect 4890 4020 4896 4072
rect 4948 4060 4954 4072
rect 5077 4063 5135 4069
rect 5077 4060 5089 4063
rect 4948 4032 5089 4060
rect 4948 4020 4954 4032
rect 5077 4029 5089 4032
rect 5123 4029 5135 4063
rect 5077 4023 5135 4029
rect 5166 4020 5172 4072
rect 5224 4060 5230 4072
rect 6472 4060 6500 4100
rect 7377 4097 7389 4131
rect 7423 4128 7435 4131
rect 7742 4128 7748 4140
rect 7423 4100 7748 4128
rect 7423 4097 7435 4100
rect 7377 4091 7435 4097
rect 7742 4088 7748 4100
rect 7800 4088 7806 4140
rect 6546 4060 6552 4072
rect 5224 4032 5269 4060
rect 6472 4032 6552 4060
rect 5224 4020 5230 4032
rect 6546 4020 6552 4032
rect 6604 4020 6610 4072
rect 8478 4060 8484 4072
rect 8439 4032 8484 4060
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 8680 4069 8708 4168
rect 9582 4156 9588 4168
rect 9640 4196 9646 4208
rect 12066 4196 12072 4208
rect 9640 4168 12072 4196
rect 9640 4156 9646 4168
rect 9398 4128 9404 4140
rect 9359 4100 9404 4128
rect 9398 4088 9404 4100
rect 9456 4088 9462 4140
rect 10042 4088 10048 4140
rect 10100 4128 10106 4140
rect 10597 4131 10655 4137
rect 10597 4128 10609 4131
rect 10100 4100 10609 4128
rect 10100 4088 10106 4100
rect 10597 4097 10609 4100
rect 10643 4097 10655 4131
rect 10597 4091 10655 4097
rect 10888 4072 10916 4168
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 14550 4196 14556 4208
rect 14384 4168 14556 4196
rect 11517 4131 11575 4137
rect 11517 4097 11529 4131
rect 11563 4097 11575 4131
rect 11517 4091 11575 4097
rect 12161 4131 12219 4137
rect 12161 4097 12173 4131
rect 12207 4097 12219 4131
rect 12161 4091 12219 4097
rect 8665 4063 8723 4069
rect 8665 4029 8677 4063
rect 8711 4029 8723 4063
rect 9122 4060 9128 4072
rect 9083 4032 9128 4060
rect 8665 4023 8723 4029
rect 9122 4020 9128 4032
rect 9180 4020 9186 4072
rect 9309 4063 9367 4069
rect 9309 4029 9321 4063
rect 9355 4060 9367 4063
rect 9674 4060 9680 4072
rect 9355 4032 9680 4060
rect 9355 4029 9367 4032
rect 9309 4023 9367 4029
rect 9674 4020 9680 4032
rect 9732 4020 9738 4072
rect 10870 4060 10876 4072
rect 10783 4032 10876 4060
rect 10870 4020 10876 4032
rect 10928 4020 10934 4072
rect 4617 3995 4675 4001
rect 4617 3992 4629 3995
rect 3988 3964 4629 3992
rect 4617 3961 4629 3964
rect 4663 3961 4675 3995
rect 4617 3955 4675 3961
rect 5997 3995 6055 4001
rect 5997 3961 6009 3995
rect 6043 3992 6055 3995
rect 9582 3992 9588 4004
rect 6043 3964 9588 3992
rect 6043 3961 6055 3964
rect 5997 3955 6055 3961
rect 9582 3952 9588 3964
rect 9640 3952 9646 4004
rect 9769 3995 9827 4001
rect 9769 3961 9781 3995
rect 9815 3992 9827 3995
rect 11532 3992 11560 4091
rect 12176 4060 12204 4091
rect 12342 4088 12348 4140
rect 12400 4128 12406 4140
rect 12437 4131 12495 4137
rect 12437 4128 12449 4131
rect 12400 4100 12449 4128
rect 12400 4088 12406 4100
rect 12437 4097 12449 4100
rect 12483 4097 12495 4131
rect 13078 4128 13084 4140
rect 13039 4100 13084 4128
rect 12437 4091 12495 4097
rect 13078 4088 13084 4100
rect 13136 4088 13142 4140
rect 13538 4128 13544 4140
rect 13499 4100 13544 4128
rect 13538 4088 13544 4100
rect 13596 4088 13602 4140
rect 14001 4131 14059 4137
rect 14001 4097 14013 4131
rect 14047 4128 14059 4131
rect 14384 4128 14412 4168
rect 14550 4156 14556 4168
rect 14608 4156 14614 4208
rect 14047 4100 14412 4128
rect 14047 4097 14059 4100
rect 14001 4091 14059 4097
rect 14458 4088 14464 4140
rect 14516 4128 14522 4140
rect 14936 4137 14964 4236
rect 16592 4236 17632 4264
rect 15028 4168 15332 4196
rect 14921 4131 14979 4137
rect 14516 4100 14561 4128
rect 14516 4088 14522 4100
rect 14921 4097 14933 4131
rect 14967 4097 14979 4131
rect 14921 4091 14979 4097
rect 14734 4060 14740 4072
rect 12176 4032 14740 4060
rect 14734 4020 14740 4032
rect 14792 4020 14798 4072
rect 15028 4060 15056 4168
rect 15194 4137 15200 4140
rect 15188 4128 15200 4137
rect 15155 4100 15200 4128
rect 15188 4091 15200 4100
rect 15194 4088 15200 4091
rect 15252 4088 15258 4140
rect 15304 4128 15332 4168
rect 16592 4128 16620 4236
rect 17494 4196 17500 4208
rect 16684 4168 17500 4196
rect 16684 4137 16712 4168
rect 17494 4156 17500 4168
rect 17552 4156 17558 4208
rect 16942 4137 16948 4140
rect 15304 4100 16620 4128
rect 16669 4131 16727 4137
rect 16669 4097 16681 4131
rect 16715 4097 16727 4131
rect 16936 4128 16948 4137
rect 16903 4100 16948 4128
rect 16669 4091 16727 4097
rect 16936 4091 16948 4100
rect 16942 4088 16948 4091
rect 17000 4088 17006 4140
rect 17604 4128 17632 4236
rect 18049 4233 18061 4267
rect 18095 4264 18107 4267
rect 18138 4264 18144 4276
rect 18095 4236 18144 4264
rect 18095 4233 18107 4236
rect 18049 4227 18107 4233
rect 18138 4224 18144 4236
rect 18196 4224 18202 4276
rect 18230 4156 18236 4208
rect 18288 4196 18294 4208
rect 20162 4196 20168 4208
rect 18288 4168 20168 4196
rect 18288 4156 18294 4168
rect 20162 4156 20168 4168
rect 20220 4156 20226 4208
rect 18601 4131 18659 4137
rect 18601 4128 18613 4131
rect 17604 4100 18613 4128
rect 18601 4097 18613 4100
rect 18647 4097 18659 4131
rect 18601 4091 18659 4097
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4097 19211 4131
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 19153 4091 19211 4097
rect 20272 4100 20821 4128
rect 19168 4060 19196 4091
rect 14844 4032 15056 4060
rect 17972 4032 19196 4060
rect 12618 3992 12624 4004
rect 9815 3964 11560 3992
rect 12579 3964 12624 3992
rect 9815 3961 9827 3964
rect 9769 3955 9827 3961
rect 12618 3952 12624 3964
rect 12676 3952 12682 4004
rect 13265 3995 13323 4001
rect 13265 3961 13277 3995
rect 13311 3992 13323 3995
rect 14844 3992 14872 4032
rect 13311 3964 14872 3992
rect 16224 3964 16712 3992
rect 13311 3961 13323 3964
rect 13265 3955 13323 3961
rect 4341 3927 4399 3933
rect 4341 3893 4353 3927
rect 4387 3924 4399 3927
rect 5442 3924 5448 3936
rect 4387 3896 5448 3924
rect 4387 3893 4399 3896
rect 4341 3887 4399 3893
rect 5442 3884 5448 3896
rect 5500 3884 5506 3936
rect 6178 3884 6184 3936
rect 6236 3924 6242 3936
rect 6914 3924 6920 3936
rect 6236 3896 6920 3924
rect 6236 3884 6242 3896
rect 6914 3884 6920 3896
rect 6972 3884 6978 3936
rect 7006 3884 7012 3936
rect 7064 3924 7070 3936
rect 7101 3927 7159 3933
rect 7101 3924 7113 3927
rect 7064 3896 7113 3924
rect 7064 3884 7070 3896
rect 7101 3893 7113 3896
rect 7147 3893 7159 3927
rect 7101 3887 7159 3893
rect 7282 3884 7288 3936
rect 7340 3924 7346 3936
rect 7561 3927 7619 3933
rect 7561 3924 7573 3927
rect 7340 3896 7573 3924
rect 7340 3884 7346 3896
rect 7561 3893 7573 3896
rect 7607 3893 7619 3927
rect 7561 3887 7619 3893
rect 8021 3927 8079 3933
rect 8021 3893 8033 3927
rect 8067 3924 8079 3927
rect 8110 3924 8116 3936
rect 8067 3896 8116 3924
rect 8067 3893 8079 3896
rect 8021 3887 8079 3893
rect 8110 3884 8116 3896
rect 8168 3884 8174 3936
rect 8202 3884 8208 3936
rect 8260 3924 8266 3936
rect 10042 3924 10048 3936
rect 8260 3896 10048 3924
rect 8260 3884 8266 3896
rect 10042 3884 10048 3896
rect 10100 3884 10106 3936
rect 10134 3884 10140 3936
rect 10192 3924 10198 3936
rect 10229 3927 10287 3933
rect 10229 3924 10241 3927
rect 10192 3896 10241 3924
rect 10192 3884 10198 3896
rect 10229 3893 10241 3896
rect 10275 3893 10287 3927
rect 11698 3924 11704 3936
rect 11659 3896 11704 3924
rect 10229 3887 10287 3893
rect 11698 3884 11704 3896
rect 11756 3884 11762 3936
rect 13722 3924 13728 3936
rect 13683 3896 13728 3924
rect 13722 3884 13728 3896
rect 13780 3884 13786 3936
rect 14185 3927 14243 3933
rect 14185 3893 14197 3927
rect 14231 3924 14243 3927
rect 14550 3924 14556 3936
rect 14231 3896 14556 3924
rect 14231 3893 14243 3896
rect 14185 3887 14243 3893
rect 14550 3884 14556 3896
rect 14608 3884 14614 3936
rect 14645 3927 14703 3933
rect 14645 3893 14657 3927
rect 14691 3924 14703 3927
rect 16224 3924 16252 3964
rect 14691 3896 16252 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 16298 3884 16304 3936
rect 16356 3924 16362 3936
rect 16684 3924 16712 3964
rect 17972 3924 18000 4032
rect 19610 4020 19616 4072
rect 19668 4060 19674 4072
rect 20272 4060 20300 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 20809 4091 20867 4097
rect 20530 4060 20536 4072
rect 19668 4032 20300 4060
rect 20491 4032 20536 4060
rect 19668 4020 19674 4032
rect 20530 4020 20536 4032
rect 20588 4020 20594 4072
rect 18785 3995 18843 4001
rect 18785 3961 18797 3995
rect 18831 3992 18843 3995
rect 20438 3992 20444 4004
rect 18831 3964 20444 3992
rect 18831 3961 18843 3964
rect 18785 3955 18843 3961
rect 20438 3952 20444 3964
rect 20496 3952 20502 4004
rect 16356 3896 16401 3924
rect 16684 3896 18000 3924
rect 16356 3884 16362 3896
rect 19058 3884 19064 3936
rect 19116 3924 19122 3936
rect 19337 3927 19395 3933
rect 19337 3924 19349 3927
rect 19116 3896 19349 3924
rect 19116 3884 19122 3896
rect 19337 3893 19349 3896
rect 19383 3893 19395 3927
rect 20070 3924 20076 3936
rect 20031 3896 20076 3924
rect 19337 3887 19395 3893
rect 20070 3884 20076 3896
rect 20128 3884 20134 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1026 3680 1032 3732
rect 1084 3720 1090 3732
rect 3050 3720 3056 3732
rect 1084 3692 3056 3720
rect 1084 3680 1090 3692
rect 3050 3680 3056 3692
rect 3108 3680 3114 3732
rect 3878 3680 3884 3732
rect 3936 3720 3942 3732
rect 6549 3723 6607 3729
rect 6549 3720 6561 3723
rect 3936 3692 6561 3720
rect 3936 3680 3942 3692
rect 6549 3689 6561 3692
rect 6595 3689 6607 3723
rect 6549 3683 6607 3689
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 8018 3720 8024 3732
rect 7156 3692 8024 3720
rect 7156 3680 7162 3692
rect 8018 3680 8024 3692
rect 8076 3680 8082 3732
rect 8573 3723 8631 3729
rect 8573 3689 8585 3723
rect 8619 3720 8631 3723
rect 9398 3720 9404 3732
rect 8619 3692 9404 3720
rect 8619 3689 8631 3692
rect 8573 3683 8631 3689
rect 9398 3680 9404 3692
rect 9456 3680 9462 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 12894 3720 12900 3732
rect 9640 3692 12900 3720
rect 9640 3680 9646 3692
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14550 3680 14556 3732
rect 14608 3720 14614 3732
rect 14608 3692 18092 3720
rect 14608 3680 14614 3692
rect 3786 3612 3792 3664
rect 3844 3652 3850 3664
rect 6178 3652 6184 3664
rect 3844 3624 6184 3652
rect 3844 3612 3850 3624
rect 6178 3612 6184 3624
rect 6236 3612 6242 3664
rect 6273 3655 6331 3661
rect 6273 3621 6285 3655
rect 6319 3621 6331 3655
rect 6273 3615 6331 3621
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2225 3587 2283 3593
rect 2225 3553 2237 3587
rect 2271 3584 2283 3587
rect 2314 3584 2320 3596
rect 2271 3556 2320 3584
rect 2271 3553 2283 3556
rect 2225 3547 2283 3553
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 2240 3516 2268 3547
rect 2314 3544 2320 3556
rect 2372 3544 2378 3596
rect 2774 3544 2780 3596
rect 2832 3584 2838 3596
rect 3053 3587 3111 3593
rect 3053 3584 3065 3587
rect 2832 3556 3065 3584
rect 2832 3544 2838 3556
rect 3053 3553 3065 3556
rect 3099 3553 3111 3587
rect 4338 3584 4344 3596
rect 4299 3556 4344 3584
rect 3053 3547 3111 3553
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 4614 3584 4620 3596
rect 4575 3556 4620 3584
rect 4614 3544 4620 3556
rect 4672 3544 4678 3596
rect 5718 3584 5724 3596
rect 5631 3556 5724 3584
rect 5718 3544 5724 3556
rect 5776 3584 5782 3596
rect 6086 3584 6092 3596
rect 5776 3556 6092 3584
rect 5776 3544 5782 3556
rect 6086 3544 6092 3556
rect 6144 3544 6150 3596
rect 624 3488 2268 3516
rect 624 3476 630 3488
rect 3234 3476 3240 3528
rect 3292 3516 3298 3528
rect 3329 3519 3387 3525
rect 3329 3516 3341 3519
rect 3292 3488 3341 3516
rect 3292 3476 3298 3488
rect 3329 3485 3341 3488
rect 3375 3485 3387 3519
rect 5810 3516 5816 3528
rect 5771 3488 5816 3516
rect 3329 3479 3387 3485
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 5994 3516 6000 3528
rect 5951 3488 6000 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6288 3516 6316 3615
rect 6914 3612 6920 3664
rect 6972 3652 6978 3664
rect 6972 3624 7144 3652
rect 6972 3612 6978 3624
rect 7006 3584 7012 3596
rect 6967 3556 7012 3584
rect 7006 3544 7012 3556
rect 7064 3544 7070 3596
rect 7116 3593 7144 3624
rect 7282 3612 7288 3664
rect 7340 3652 7346 3664
rect 7742 3652 7748 3664
rect 7340 3624 7748 3652
rect 7340 3612 7346 3624
rect 7742 3612 7748 3624
rect 7800 3612 7806 3664
rect 8938 3652 8944 3664
rect 7944 3624 8944 3652
rect 7944 3593 7972 3624
rect 8938 3612 8944 3624
rect 8996 3612 9002 3664
rect 10318 3612 10324 3664
rect 10376 3652 10382 3664
rect 11606 3652 11612 3664
rect 10376 3624 11612 3652
rect 10376 3612 10382 3624
rect 11606 3612 11612 3624
rect 11664 3612 11670 3664
rect 13630 3652 13636 3664
rect 13591 3624 13636 3652
rect 13630 3612 13636 3624
rect 13688 3612 13694 3664
rect 13722 3612 13728 3664
rect 13780 3652 13786 3664
rect 13780 3624 17080 3652
rect 13780 3612 13786 3624
rect 7101 3587 7159 3593
rect 7101 3553 7113 3587
rect 7147 3553 7159 3587
rect 7101 3547 7159 3553
rect 7929 3587 7987 3593
rect 7929 3553 7941 3587
rect 7975 3553 7987 3587
rect 8110 3584 8116 3596
rect 8071 3556 8116 3584
rect 7929 3547 7987 3553
rect 8110 3544 8116 3556
rect 8168 3544 8174 3596
rect 10870 3584 10876 3596
rect 10428 3556 10876 3584
rect 6288 3488 6500 3516
rect 4246 3408 4252 3460
rect 4304 3448 4310 3460
rect 4614 3448 4620 3460
rect 4304 3420 4620 3448
rect 4304 3408 4310 3420
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 4982 3448 4988 3460
rect 4943 3420 4988 3448
rect 4982 3408 4988 3420
rect 5040 3408 5046 3460
rect 6472 3448 6500 3488
rect 6546 3476 6552 3528
rect 6604 3516 6610 3528
rect 7650 3516 7656 3528
rect 6604 3488 7656 3516
rect 6604 3476 6610 3488
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8294 3476 8300 3528
rect 8352 3516 8358 3528
rect 10321 3519 10379 3525
rect 10321 3516 10333 3519
rect 8352 3488 10333 3516
rect 8352 3476 8358 3488
rect 10321 3485 10333 3488
rect 10367 3485 10379 3519
rect 10321 3479 10379 3485
rect 6917 3451 6975 3457
rect 6917 3448 6929 3451
rect 6472 3420 6929 3448
rect 6917 3417 6929 3420
rect 6963 3417 6975 3451
rect 6917 3411 6975 3417
rect 8205 3451 8263 3457
rect 8205 3417 8217 3451
rect 8251 3448 8263 3451
rect 8386 3448 8392 3460
rect 8251 3420 8392 3448
rect 8251 3417 8263 3420
rect 8205 3411 8263 3417
rect 8386 3408 8392 3420
rect 8444 3408 8450 3460
rect 8662 3408 8668 3460
rect 8720 3448 8726 3460
rect 9766 3448 9772 3460
rect 8720 3420 9772 3448
rect 8720 3408 8726 3420
rect 9766 3408 9772 3420
rect 9824 3408 9830 3460
rect 10076 3451 10134 3457
rect 10076 3417 10088 3451
rect 10122 3448 10134 3451
rect 10428 3448 10456 3556
rect 10870 3544 10876 3556
rect 10928 3584 10934 3596
rect 11149 3587 11207 3593
rect 11149 3584 11161 3587
rect 10928 3556 11161 3584
rect 10928 3544 10934 3556
rect 11149 3553 11161 3556
rect 11195 3553 11207 3587
rect 14829 3587 14887 3593
rect 11149 3547 11207 3553
rect 11716 3556 14320 3584
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 10652 3488 10732 3516
rect 10652 3476 10658 3488
rect 10122 3420 10456 3448
rect 10122 3417 10134 3420
rect 10076 3411 10134 3417
rect 3326 3340 3332 3392
rect 3384 3380 3390 3392
rect 5077 3383 5135 3389
rect 5077 3380 5089 3383
rect 3384 3352 5089 3380
rect 3384 3340 3390 3352
rect 5077 3349 5089 3352
rect 5123 3380 5135 3383
rect 7926 3380 7932 3392
rect 5123 3352 7932 3380
rect 5123 3349 5135 3352
rect 5077 3343 5135 3349
rect 7926 3340 7932 3352
rect 7984 3380 7990 3392
rect 8110 3380 8116 3392
rect 7984 3352 8116 3380
rect 7984 3340 7990 3352
rect 8110 3340 8116 3352
rect 8168 3340 8174 3392
rect 8938 3380 8944 3392
rect 8899 3352 8944 3380
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 10594 3380 10600 3392
rect 10555 3352 10600 3380
rect 10594 3340 10600 3352
rect 10652 3340 10658 3392
rect 10704 3380 10732 3488
rect 10962 3476 10968 3528
rect 11020 3516 11026 3528
rect 11020 3488 11065 3516
rect 11020 3476 11026 3488
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 11609 3519 11667 3525
rect 11609 3516 11621 3519
rect 11296 3488 11621 3516
rect 11296 3476 11302 3488
rect 11609 3485 11621 3488
rect 11655 3485 11667 3519
rect 11609 3479 11667 3485
rect 10980 3448 11008 3476
rect 11716 3448 11744 3556
rect 12158 3516 12164 3528
rect 12119 3488 12164 3516
rect 12158 3476 12164 3488
rect 12216 3476 12222 3528
rect 12802 3516 12808 3528
rect 12763 3488 12808 3516
rect 12802 3476 12808 3488
rect 12860 3476 12866 3528
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3485 13231 3519
rect 14182 3516 14188 3528
rect 14143 3488 14188 3516
rect 13173 3479 13231 3485
rect 13188 3448 13216 3479
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 14292 3516 14320 3556
rect 14829 3553 14841 3587
rect 14875 3584 14887 3587
rect 15194 3584 15200 3596
rect 14875 3556 15200 3584
rect 14875 3553 14887 3556
rect 14829 3547 14887 3553
rect 15194 3544 15200 3556
rect 15252 3584 15258 3596
rect 16209 3587 16267 3593
rect 16209 3584 16221 3587
rect 15252 3556 16221 3584
rect 15252 3544 15258 3556
rect 16209 3553 16221 3556
rect 16255 3553 16267 3587
rect 16209 3547 16267 3553
rect 15013 3519 15071 3525
rect 15013 3516 15025 3519
rect 14292 3488 15025 3516
rect 15013 3485 15025 3488
rect 15059 3485 15071 3519
rect 15013 3479 15071 3485
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 16945 3519 17003 3525
rect 16945 3516 16957 3519
rect 16080 3488 16957 3516
rect 16080 3476 16086 3488
rect 16945 3485 16957 3488
rect 16991 3485 17003 3519
rect 17052 3516 17080 3624
rect 18064 3525 18092 3692
rect 18690 3680 18696 3732
rect 18748 3720 18754 3732
rect 22278 3720 22284 3732
rect 18748 3692 22284 3720
rect 18748 3680 18754 3692
rect 22278 3680 22284 3692
rect 22336 3680 22342 3732
rect 18233 3655 18291 3661
rect 18233 3621 18245 3655
rect 18279 3652 18291 3655
rect 19518 3652 19524 3664
rect 18279 3624 19524 3652
rect 18279 3621 18291 3624
rect 18233 3615 18291 3621
rect 19518 3612 19524 3624
rect 19576 3612 19582 3664
rect 19429 3587 19487 3593
rect 19429 3553 19441 3587
rect 19475 3584 19487 3587
rect 19794 3584 19800 3596
rect 19475 3556 19800 3584
rect 19475 3553 19487 3556
rect 19429 3547 19487 3553
rect 19794 3544 19800 3556
rect 19852 3544 19858 3596
rect 20809 3587 20867 3593
rect 20809 3553 20821 3587
rect 20855 3584 20867 3587
rect 21634 3584 21640 3596
rect 20855 3556 21640 3584
rect 20855 3553 20867 3556
rect 20809 3547 20867 3553
rect 21634 3544 21640 3556
rect 21692 3544 21698 3596
rect 17497 3519 17555 3525
rect 17497 3516 17509 3519
rect 17052 3488 17509 3516
rect 16945 3479 17003 3485
rect 17497 3485 17509 3488
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 18049 3519 18107 3525
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18601 3519 18659 3525
rect 18601 3485 18613 3519
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 19705 3519 19763 3525
rect 19705 3485 19717 3519
rect 19751 3516 19763 3519
rect 20346 3516 20352 3528
rect 19751 3488 20352 3516
rect 19751 3485 19763 3488
rect 19705 3479 19763 3485
rect 14642 3448 14648 3460
rect 10980 3420 11744 3448
rect 12360 3420 13216 3448
rect 13372 3420 14648 3448
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 10704 3352 11069 3380
rect 11057 3349 11069 3352
rect 11103 3349 11115 3383
rect 11790 3380 11796 3392
rect 11751 3352 11796 3380
rect 11057 3343 11115 3349
rect 11790 3340 11796 3352
rect 11848 3340 11854 3392
rect 12360 3389 12388 3420
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3349 12403 3383
rect 12618 3380 12624 3392
rect 12579 3352 12624 3380
rect 12345 3343 12403 3349
rect 12618 3340 12624 3352
rect 12676 3340 12682 3392
rect 13372 3389 13400 3420
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 15838 3448 15844 3460
rect 14844 3420 15844 3448
rect 13357 3383 13415 3389
rect 13357 3349 13369 3383
rect 13403 3349 13415 3383
rect 13357 3343 13415 3349
rect 14369 3383 14427 3389
rect 14369 3349 14381 3383
rect 14415 3380 14427 3383
rect 14844 3380 14872 3420
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 15930 3408 15936 3460
rect 15988 3448 15994 3460
rect 18616 3448 18644 3479
rect 20346 3476 20352 3488
rect 20404 3476 20410 3528
rect 20533 3519 20591 3525
rect 20533 3485 20545 3519
rect 20579 3485 20591 3519
rect 20533 3479 20591 3485
rect 15988 3420 18644 3448
rect 15988 3408 15994 3420
rect 18966 3408 18972 3460
rect 19024 3448 19030 3460
rect 20548 3448 20576 3479
rect 20622 3448 20628 3460
rect 19024 3420 20628 3448
rect 19024 3408 19030 3420
rect 20622 3408 20628 3420
rect 20680 3408 20686 3460
rect 14415 3352 14872 3380
rect 14921 3383 14979 3389
rect 14415 3349 14427 3352
rect 14369 3343 14427 3349
rect 14921 3349 14933 3383
rect 14967 3380 14979 3383
rect 15102 3380 15108 3392
rect 14967 3352 15108 3380
rect 14967 3349 14979 3352
rect 14921 3343 14979 3349
rect 15102 3340 15108 3352
rect 15160 3340 15166 3392
rect 15378 3380 15384 3392
rect 15339 3352 15384 3380
rect 15378 3340 15384 3352
rect 15436 3340 15442 3392
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 15657 3383 15715 3389
rect 15657 3380 15669 3383
rect 15528 3352 15669 3380
rect 15528 3340 15534 3352
rect 15657 3349 15669 3352
rect 15703 3349 15715 3383
rect 16022 3380 16028 3392
rect 15983 3352 16028 3380
rect 15657 3343 15715 3349
rect 16022 3340 16028 3352
rect 16080 3340 16086 3392
rect 16117 3383 16175 3389
rect 16117 3349 16129 3383
rect 16163 3380 16175 3383
rect 16390 3380 16396 3392
rect 16163 3352 16396 3380
rect 16163 3349 16175 3352
rect 16117 3343 16175 3349
rect 16390 3340 16396 3352
rect 16448 3340 16454 3392
rect 17126 3380 17132 3392
rect 17087 3352 17132 3380
rect 17126 3340 17132 3352
rect 17184 3340 17190 3392
rect 17678 3380 17684 3392
rect 17639 3352 17684 3380
rect 17678 3340 17684 3352
rect 17736 3340 17742 3392
rect 18598 3340 18604 3392
rect 18656 3380 18662 3392
rect 18785 3383 18843 3389
rect 18785 3380 18797 3383
rect 18656 3352 18797 3380
rect 18656 3340 18662 3352
rect 18785 3349 18797 3352
rect 18831 3349 18843 3383
rect 18785 3343 18843 3349
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 2774 3176 2780 3188
rect 2240 3148 2780 3176
rect 1762 3000 1768 3052
rect 1820 3040 1826 3052
rect 2240 3049 2268 3148
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 3970 3176 3976 3188
rect 2875 3148 3832 3176
rect 3931 3148 3976 3176
rect 2875 3117 2903 3148
rect 2860 3111 2918 3117
rect 2860 3077 2872 3111
rect 2906 3077 2918 3111
rect 3804 3108 3832 3148
rect 3970 3136 3976 3148
rect 4028 3136 4034 3188
rect 5721 3179 5779 3185
rect 5721 3145 5733 3179
rect 5767 3176 5779 3179
rect 6914 3176 6920 3188
rect 5767 3148 6920 3176
rect 5767 3145 5779 3148
rect 5721 3139 5779 3145
rect 5166 3108 5172 3120
rect 3804 3080 5172 3108
rect 2860 3071 2918 3077
rect 5166 3068 5172 3080
rect 5224 3108 5230 3120
rect 5736 3108 5764 3139
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 7466 3176 7472 3188
rect 7427 3148 7472 3176
rect 7466 3136 7472 3148
rect 7524 3136 7530 3188
rect 7852 3148 9076 3176
rect 7852 3108 7880 3148
rect 8294 3108 8300 3120
rect 5224 3080 5764 3108
rect 7300 3080 7880 3108
rect 7944 3080 8300 3108
rect 5224 3068 5230 3080
rect 1949 3043 2007 3049
rect 1949 3040 1961 3043
rect 1820 3012 1961 3040
rect 1820 3000 1826 3012
rect 1949 3009 1961 3012
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3009 2283 3043
rect 2225 3003 2283 3009
rect 4608 3043 4666 3049
rect 4608 3009 4620 3043
rect 4654 3040 4666 3043
rect 5718 3040 5724 3052
rect 4654 3012 5724 3040
rect 4654 3009 4666 3012
rect 4608 3003 4666 3009
rect 5718 3000 5724 3012
rect 5776 3000 5782 3052
rect 6914 3040 6920 3052
rect 6875 3012 6920 3040
rect 6914 3000 6920 3012
rect 6972 3000 6978 3052
rect 7098 3000 7104 3052
rect 7156 3040 7162 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 7156 3012 7205 3040
rect 7156 3000 7162 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 2593 2975 2651 2981
rect 2593 2941 2605 2975
rect 2639 2941 2651 2975
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 2593 2935 2651 2941
rect 3896 2944 4353 2972
rect 2608 2836 2636 2935
rect 2958 2836 2964 2848
rect 2608 2808 2964 2836
rect 2958 2796 2964 2808
rect 3016 2836 3022 2848
rect 3896 2836 3924 2944
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 5994 2932 6000 2984
rect 6052 2972 6058 2984
rect 7116 2972 7144 3000
rect 6052 2944 7144 2972
rect 6052 2932 6058 2944
rect 3016 2808 3924 2836
rect 3016 2796 3022 2808
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 7300 2836 7328 3080
rect 7653 3043 7711 3049
rect 7653 3009 7665 3043
rect 7699 3040 7711 3043
rect 7834 3040 7840 3052
rect 7699 3012 7840 3040
rect 7699 3009 7711 3012
rect 7653 3003 7711 3009
rect 7834 3000 7840 3012
rect 7892 3000 7898 3052
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7944 2981 7972 3080
rect 8294 3068 8300 3080
rect 8352 3068 8358 3120
rect 8196 3043 8254 3049
rect 8196 3009 8208 3043
rect 8242 3040 8254 3043
rect 9048 3040 9076 3148
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9309 3179 9367 3185
rect 9309 3176 9321 3179
rect 9180 3148 9321 3176
rect 9180 3136 9186 3148
rect 9309 3145 9321 3148
rect 9355 3145 9367 3179
rect 9674 3176 9680 3188
rect 9635 3148 9680 3176
rect 9309 3139 9367 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 10045 3179 10103 3185
rect 10045 3145 10057 3179
rect 10091 3176 10103 3179
rect 10594 3176 10600 3188
rect 10091 3148 10600 3176
rect 10091 3145 10103 3148
rect 10045 3139 10103 3145
rect 10594 3136 10600 3148
rect 10652 3136 10658 3188
rect 12618 3176 12624 3188
rect 10980 3148 12624 3176
rect 10134 3108 10140 3120
rect 10095 3080 10140 3108
rect 10134 3068 10140 3080
rect 10192 3068 10198 3120
rect 10870 3040 10876 3052
rect 8242 3012 8984 3040
rect 9048 3012 10876 3040
rect 8242 3009 8254 3012
rect 8196 3003 8254 3009
rect 8956 2984 8984 3012
rect 10870 3000 10876 3012
rect 10928 3000 10934 3052
rect 10980 3049 11008 3148
rect 12618 3136 12624 3148
rect 12676 3136 12682 3188
rect 12710 3136 12716 3188
rect 12768 3176 12774 3188
rect 14093 3179 14151 3185
rect 14093 3176 14105 3179
rect 12768 3148 14105 3176
rect 12768 3136 12774 3148
rect 14093 3145 14105 3148
rect 14139 3145 14151 3179
rect 14093 3139 14151 3145
rect 14182 3136 14188 3188
rect 14240 3176 14246 3188
rect 15286 3176 15292 3188
rect 14240 3148 15292 3176
rect 14240 3136 14246 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 15470 3176 15476 3188
rect 15431 3148 15476 3176
rect 15470 3136 15476 3148
rect 15528 3136 15534 3188
rect 16022 3136 16028 3188
rect 16080 3176 16086 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 16080 3148 16129 3176
rect 16080 3136 16086 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 17678 3136 17684 3188
rect 17736 3176 17742 3188
rect 20898 3176 20904 3188
rect 17736 3148 20904 3176
rect 17736 3136 17742 3148
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 11790 3068 11796 3120
rect 11848 3108 11854 3120
rect 11848 3080 13400 3108
rect 11848 3068 11854 3080
rect 10965 3043 11023 3049
rect 10965 3009 10977 3043
rect 11011 3009 11023 3043
rect 10965 3003 11023 3009
rect 11054 3000 11060 3052
rect 11112 3040 11118 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11112 3012 11529 3040
rect 11112 3000 11118 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11756 3012 11989 3040
rect 11756 3000 11762 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 12437 3043 12495 3049
rect 12437 3009 12449 3043
rect 12483 3040 12495 3043
rect 12526 3040 12532 3052
rect 12483 3012 12532 3040
rect 12483 3009 12495 3012
rect 12437 3003 12495 3009
rect 12526 3000 12532 3012
rect 12584 3000 12590 3052
rect 12894 3040 12900 3052
rect 12855 3012 12900 3040
rect 12894 3000 12900 3012
rect 12952 3000 12958 3052
rect 13372 3049 13400 3080
rect 15378 3068 15384 3120
rect 15436 3108 15442 3120
rect 15565 3111 15623 3117
rect 15565 3108 15577 3111
rect 15436 3080 15577 3108
rect 15436 3068 15442 3080
rect 15565 3077 15577 3080
rect 15611 3077 15623 3111
rect 15565 3071 15623 3077
rect 17126 3068 17132 3120
rect 17184 3108 17190 3120
rect 21358 3108 21364 3120
rect 17184 3080 21364 3108
rect 17184 3068 17190 3080
rect 21358 3068 21364 3080
rect 21416 3068 21422 3120
rect 13357 3043 13415 3049
rect 13357 3009 13369 3043
rect 13403 3009 13415 3043
rect 14274 3040 14280 3052
rect 14235 3012 14280 3040
rect 13357 3003 13415 3009
rect 14274 3000 14280 3012
rect 14332 3000 14338 3052
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 7929 2975 7987 2981
rect 7929 2972 7941 2975
rect 7800 2944 7941 2972
rect 7800 2932 7806 2944
rect 7929 2941 7941 2944
rect 7975 2941 7987 2975
rect 7929 2935 7987 2941
rect 8938 2932 8944 2984
rect 8996 2972 9002 2984
rect 10229 2975 10287 2981
rect 10229 2972 10241 2975
rect 8996 2944 10241 2972
rect 8996 2932 9002 2944
rect 10229 2941 10241 2944
rect 10275 2941 10287 2975
rect 12158 2972 12164 2984
rect 10229 2935 10287 2941
rect 10888 2944 12164 2972
rect 7374 2864 7380 2916
rect 7432 2864 7438 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 10318 2904 10324 2916
rect 9732 2876 10324 2904
rect 9732 2864 9738 2876
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 4120 2808 7328 2836
rect 7392 2836 7420 2864
rect 10888 2836 10916 2944
rect 12158 2932 12164 2944
rect 12216 2932 12222 2984
rect 14568 2972 14596 3003
rect 15654 3000 15660 3052
rect 15712 3040 15718 3052
rect 16669 3043 16727 3049
rect 15712 3012 16436 3040
rect 15712 3000 15718 3012
rect 12406 2944 14596 2972
rect 15749 2975 15807 2981
rect 11701 2907 11759 2913
rect 11701 2873 11713 2907
rect 11747 2904 11759 2907
rect 12406 2904 12434 2944
rect 15749 2941 15761 2975
rect 15795 2972 15807 2975
rect 16298 2972 16304 2984
rect 15795 2944 16304 2972
rect 15795 2941 15807 2944
rect 15749 2935 15807 2941
rect 16298 2932 16304 2944
rect 16356 2932 16362 2984
rect 16408 2972 16436 3012
rect 16669 3009 16681 3043
rect 16715 3040 16727 3043
rect 17034 3040 17040 3052
rect 16715 3012 17040 3040
rect 16715 3009 16727 3012
rect 16669 3003 16727 3009
rect 17034 3000 17040 3012
rect 17092 3000 17098 3052
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17405 3043 17463 3049
rect 17405 3040 17417 3043
rect 17368 3012 17417 3040
rect 17368 3000 17374 3012
rect 17405 3009 17417 3012
rect 17451 3009 17463 3043
rect 18046 3040 18052 3052
rect 18007 3012 18052 3040
rect 17405 3003 17463 3009
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18322 3040 18328 3052
rect 18283 3012 18328 3040
rect 18322 3000 18328 3012
rect 18380 3000 18386 3052
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3040 19763 3043
rect 19886 3040 19892 3052
rect 19751 3012 19892 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 19886 3000 19892 3012
rect 19944 3000 19950 3052
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 20070 3040 20076 3052
rect 20027 3012 20076 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 20070 3000 20076 3012
rect 20128 3000 20134 3052
rect 21082 3040 21088 3052
rect 21043 3012 21088 3040
rect 21082 3000 21088 3012
rect 21140 3040 21146 3052
rect 22738 3040 22744 3052
rect 21140 3012 22744 3040
rect 21140 3000 21146 3012
rect 22738 3000 22744 3012
rect 22796 3000 22802 3052
rect 17954 2972 17960 2984
rect 16408 2944 17960 2972
rect 17954 2932 17960 2944
rect 18012 2932 18018 2984
rect 20714 2972 20720 2984
rect 20675 2944 20720 2972
rect 20714 2932 20720 2944
rect 20772 2932 20778 2984
rect 11747 2876 12434 2904
rect 13081 2907 13139 2913
rect 11747 2873 11759 2876
rect 11701 2867 11759 2873
rect 13081 2873 13093 2907
rect 13127 2904 13139 2907
rect 13814 2904 13820 2916
rect 13127 2876 13820 2904
rect 13127 2873 13139 2876
rect 13081 2867 13139 2873
rect 13814 2864 13820 2876
rect 13872 2864 13878 2916
rect 16666 2904 16672 2916
rect 14568 2876 16672 2904
rect 11146 2836 11152 2848
rect 7392 2808 10916 2836
rect 11107 2808 11152 2836
rect 4120 2796 4126 2808
rect 11146 2796 11152 2808
rect 11204 2796 11210 2848
rect 12161 2839 12219 2845
rect 12161 2805 12173 2839
rect 12207 2836 12219 2839
rect 12526 2836 12532 2848
rect 12207 2808 12532 2836
rect 12207 2805 12219 2808
rect 12161 2799 12219 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 12621 2839 12679 2845
rect 12621 2805 12633 2839
rect 12667 2836 12679 2839
rect 12986 2836 12992 2848
rect 12667 2808 12992 2836
rect 12667 2805 12679 2808
rect 12621 2799 12679 2805
rect 12986 2796 12992 2808
rect 13044 2796 13050 2848
rect 13541 2839 13599 2845
rect 13541 2805 13553 2839
rect 13587 2836 13599 2839
rect 14568 2836 14596 2876
rect 16666 2864 16672 2876
rect 16724 2864 16730 2916
rect 14734 2836 14740 2848
rect 13587 2808 14596 2836
rect 14695 2808 14740 2836
rect 13587 2805 13599 2808
rect 13541 2799 13599 2805
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 14826 2796 14832 2848
rect 14884 2836 14890 2848
rect 15105 2839 15163 2845
rect 15105 2836 15117 2839
rect 14884 2808 15117 2836
rect 14884 2796 14890 2808
rect 15105 2805 15117 2808
rect 15151 2805 15163 2839
rect 15105 2799 15163 2805
rect 15930 2796 15936 2848
rect 15988 2836 15994 2848
rect 16853 2839 16911 2845
rect 16853 2836 16865 2839
rect 15988 2808 16865 2836
rect 15988 2796 15994 2808
rect 16853 2805 16865 2808
rect 16899 2805 16911 2839
rect 16853 2799 16911 2805
rect 17310 2796 17316 2848
rect 17368 2836 17374 2848
rect 17589 2839 17647 2845
rect 17589 2836 17601 2839
rect 17368 2808 17601 2836
rect 17368 2796 17374 2808
rect 17589 2805 17601 2808
rect 17635 2805 17647 2839
rect 17589 2799 17647 2805
rect 18230 2796 18236 2848
rect 18288 2836 18294 2848
rect 18509 2839 18567 2845
rect 18509 2836 18521 2839
rect 18288 2808 18521 2836
rect 18288 2796 18294 2808
rect 18509 2805 18521 2808
rect 18555 2805 18567 2839
rect 18509 2799 18567 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 1578 2632 1584 2644
rect 1539 2604 1584 2632
rect 1578 2592 1584 2604
rect 1636 2592 1642 2644
rect 3234 2632 3240 2644
rect 1688 2604 3240 2632
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 1688 2564 1716 2604
rect 3234 2592 3240 2604
rect 3292 2592 3298 2644
rect 3878 2592 3884 2644
rect 3936 2632 3942 2644
rect 6365 2635 6423 2641
rect 3936 2604 5764 2632
rect 3936 2592 3942 2604
rect 1360 2536 1716 2564
rect 1360 2524 1366 2536
rect 2958 2496 2964 2508
rect 2919 2468 2964 2496
rect 2958 2456 2964 2468
rect 3016 2456 3022 2508
rect 5350 2496 5356 2508
rect 3160 2468 5356 2496
rect 2705 2431 2763 2437
rect 2705 2397 2717 2431
rect 2751 2428 2763 2431
rect 3160 2428 3188 2468
rect 5350 2456 5356 2468
rect 5408 2456 5414 2508
rect 5442 2456 5448 2508
rect 5500 2496 5506 2508
rect 5736 2505 5764 2604
rect 6365 2601 6377 2635
rect 6411 2632 6423 2635
rect 6638 2632 6644 2644
rect 6411 2604 6644 2632
rect 6411 2601 6423 2604
rect 6365 2595 6423 2601
rect 6638 2592 6644 2604
rect 6696 2592 6702 2644
rect 8018 2592 8024 2644
rect 8076 2632 8082 2644
rect 8389 2635 8447 2641
rect 8389 2632 8401 2635
rect 8076 2604 8401 2632
rect 8076 2592 8082 2604
rect 8389 2601 8401 2604
rect 8435 2601 8447 2635
rect 9398 2632 9404 2644
rect 9359 2604 9404 2632
rect 8389 2595 8447 2601
rect 9398 2592 9404 2604
rect 9456 2592 9462 2644
rect 9674 2632 9680 2644
rect 9508 2604 9680 2632
rect 9214 2564 9220 2576
rect 8496 2536 9220 2564
rect 5721 2499 5779 2505
rect 5500 2468 5545 2496
rect 5500 2456 5506 2468
rect 5721 2465 5733 2499
rect 5767 2465 5779 2499
rect 7742 2496 7748 2508
rect 7703 2468 7748 2496
rect 5721 2459 5779 2465
rect 7742 2456 7748 2468
rect 7800 2456 7806 2508
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 8021 2499 8079 2505
rect 8021 2496 8033 2499
rect 7984 2468 8033 2496
rect 7984 2456 7990 2468
rect 8021 2465 8033 2468
rect 8067 2465 8079 2499
rect 8021 2459 8079 2465
rect 2751 2400 3188 2428
rect 3237 2431 3295 2437
rect 2751 2397 2763 2400
rect 2705 2391 2763 2397
rect 3237 2397 3249 2431
rect 3283 2397 3295 2431
rect 3237 2391 3295 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 4430 2428 4436 2440
rect 4387 2400 4436 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 3252 2360 3280 2391
rect 4430 2388 4436 2400
rect 4488 2388 4494 2440
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 7478 2431 7536 2437
rect 7478 2428 7490 2431
rect 6788 2400 7490 2428
rect 6788 2388 6794 2400
rect 7478 2397 7490 2400
rect 7524 2397 7536 2431
rect 7478 2391 7536 2397
rect 8496 2360 8524 2536
rect 9214 2524 9220 2536
rect 9272 2524 9278 2576
rect 9508 2496 9536 2604
rect 9674 2592 9680 2604
rect 9732 2592 9738 2644
rect 10042 2632 10048 2644
rect 10003 2604 10048 2632
rect 10042 2592 10048 2604
rect 10100 2592 10106 2644
rect 10410 2592 10416 2644
rect 10468 2632 10474 2644
rect 11747 2635 11805 2641
rect 11747 2632 11759 2635
rect 10468 2604 11759 2632
rect 10468 2592 10474 2604
rect 11747 2601 11759 2604
rect 11793 2601 11805 2635
rect 11747 2595 11805 2601
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 13228 2604 17540 2632
rect 13228 2592 13234 2604
rect 10686 2564 10692 2576
rect 8588 2468 9536 2496
rect 9600 2536 10692 2564
rect 8588 2437 8616 2468
rect 9600 2437 9628 2536
rect 10686 2524 10692 2536
rect 10744 2564 10750 2576
rect 10962 2564 10968 2576
rect 10744 2536 10968 2564
rect 10744 2524 10750 2536
rect 10962 2524 10968 2536
rect 11020 2524 11026 2576
rect 11974 2564 11980 2576
rect 11072 2536 11980 2564
rect 9766 2456 9772 2508
rect 9824 2496 9830 2508
rect 10321 2499 10379 2505
rect 10321 2496 10333 2499
rect 9824 2468 10333 2496
rect 9824 2456 9830 2468
rect 10321 2465 10333 2468
rect 10367 2496 10379 2499
rect 10410 2496 10416 2508
rect 10367 2468 10416 2496
rect 10367 2465 10379 2468
rect 10321 2459 10379 2465
rect 10410 2456 10416 2468
rect 10468 2456 10474 2508
rect 11072 2496 11100 2536
rect 11974 2524 11980 2536
rect 12032 2524 12038 2576
rect 14090 2524 14096 2576
rect 14148 2564 14154 2576
rect 14829 2567 14887 2573
rect 14829 2564 14841 2567
rect 14148 2536 14841 2564
rect 14148 2524 14154 2536
rect 14829 2533 14841 2536
rect 14875 2533 14887 2567
rect 14829 2527 14887 2533
rect 15010 2524 15016 2576
rect 15068 2564 15074 2576
rect 15933 2567 15991 2573
rect 15933 2564 15945 2567
rect 15068 2536 15945 2564
rect 15068 2524 15074 2536
rect 15933 2533 15945 2536
rect 15979 2533 15991 2567
rect 15933 2527 15991 2533
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 17405 2567 17463 2573
rect 17405 2564 17417 2567
rect 16448 2536 17417 2564
rect 16448 2524 16454 2536
rect 17405 2533 17417 2536
rect 17451 2533 17463 2567
rect 17405 2527 17463 2533
rect 10520 2468 11100 2496
rect 8573 2431 8631 2437
rect 8573 2397 8585 2431
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8941 2431 8999 2437
rect 8941 2397 8953 2431
rect 8987 2397 8999 2431
rect 8941 2391 8999 2397
rect 9585 2431 9643 2437
rect 9585 2397 9597 2431
rect 9631 2397 9643 2431
rect 9585 2391 9643 2397
rect 9861 2431 9919 2437
rect 9861 2397 9873 2431
rect 9907 2428 9919 2431
rect 10520 2428 10548 2468
rect 11146 2456 11152 2508
rect 11204 2496 11210 2508
rect 11204 2468 15792 2496
rect 11204 2456 11210 2468
rect 9907 2400 10548 2428
rect 9907 2397 9919 2400
rect 9861 2391 9919 2397
rect 3252 2332 8524 2360
rect 8956 2360 8984 2391
rect 10870 2388 10876 2440
rect 10928 2428 10934 2440
rect 11238 2428 11244 2440
rect 10928 2400 11244 2428
rect 10928 2388 10934 2400
rect 11238 2388 11244 2400
rect 11296 2428 11302 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11296 2400 11529 2428
rect 11296 2388 11302 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12526 2388 12532 2440
rect 12584 2428 12590 2440
rect 12897 2431 12955 2437
rect 12897 2428 12909 2431
rect 12584 2400 12909 2428
rect 12584 2388 12590 2400
rect 12897 2397 12909 2400
rect 12943 2397 12955 2431
rect 12897 2391 12955 2397
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13449 2431 13507 2437
rect 13449 2428 13461 2431
rect 13044 2400 13461 2428
rect 13044 2388 13050 2400
rect 13449 2397 13461 2400
rect 13495 2397 13507 2431
rect 13449 2391 13507 2397
rect 13814 2388 13820 2440
rect 13872 2428 13878 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13872 2400 14105 2428
rect 13872 2388 13878 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14642 2428 14648 2440
rect 14603 2400 14648 2428
rect 14093 2391 14151 2397
rect 14642 2388 14648 2400
rect 14700 2388 14706 2440
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 15764 2437 15792 2468
rect 15838 2456 15844 2508
rect 15896 2496 15902 2508
rect 15896 2468 17356 2496
rect 15896 2456 15902 2468
rect 15197 2431 15255 2437
rect 15197 2428 15209 2431
rect 14792 2400 15209 2428
rect 14792 2388 14798 2400
rect 15197 2397 15209 2400
rect 15243 2397 15255 2431
rect 15197 2391 15255 2397
rect 15749 2431 15807 2437
rect 15749 2397 15761 2431
rect 15795 2397 15807 2431
rect 16666 2428 16672 2440
rect 16627 2400 16672 2428
rect 15749 2391 15807 2397
rect 16666 2388 16672 2400
rect 16724 2388 16730 2440
rect 17221 2431 17279 2437
rect 17221 2397 17233 2431
rect 17267 2397 17279 2431
rect 17221 2391 17279 2397
rect 12618 2360 12624 2372
rect 8956 2332 12624 2360
rect 12618 2320 12624 2332
rect 12676 2320 12682 2372
rect 17236 2360 17264 2391
rect 12728 2332 17264 2360
rect 17328 2360 17356 2468
rect 17512 2428 17540 2604
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 18509 2567 18567 2573
rect 18509 2564 18521 2567
rect 17828 2536 18521 2564
rect 17828 2524 17834 2536
rect 18509 2533 18521 2536
rect 18555 2533 18567 2567
rect 18509 2527 18567 2533
rect 21085 2499 21143 2505
rect 21085 2465 21097 2499
rect 21131 2496 21143 2499
rect 21450 2496 21456 2508
rect 21131 2468 21456 2496
rect 21131 2465 21143 2468
rect 21085 2459 21143 2465
rect 21450 2456 21456 2468
rect 21508 2456 21514 2508
rect 17773 2431 17831 2437
rect 17773 2428 17785 2431
rect 17512 2400 17785 2428
rect 17773 2397 17785 2400
rect 17819 2397 17831 2431
rect 17773 2391 17831 2397
rect 18325 2431 18383 2437
rect 18325 2397 18337 2431
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 18340 2360 18368 2391
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 19981 2431 20039 2437
rect 19981 2428 19993 2431
rect 18564 2400 19993 2428
rect 18564 2388 18570 2400
rect 19981 2397 19993 2400
rect 20027 2397 20039 2431
rect 20254 2428 20260 2440
rect 20215 2400 20260 2428
rect 19981 2391 20039 2397
rect 20254 2388 20260 2400
rect 20312 2388 20318 2440
rect 21266 2388 21272 2440
rect 21324 2428 21330 2440
rect 21361 2431 21419 2437
rect 21361 2428 21373 2431
rect 21324 2400 21373 2428
rect 21324 2388 21330 2400
rect 21361 2397 21373 2400
rect 21407 2397 21419 2431
rect 21361 2391 21419 2397
rect 17328 2332 18368 2360
rect 3418 2292 3424 2304
rect 3379 2264 3424 2292
rect 3418 2252 3424 2264
rect 3476 2252 3482 2304
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 6822 2292 6828 2304
rect 4120 2264 6828 2292
rect 4120 2252 4126 2264
rect 6822 2252 6828 2264
rect 6880 2252 6886 2304
rect 9122 2292 9128 2304
rect 9083 2264 9128 2292
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 10551 2295 10609 2301
rect 10551 2292 10563 2295
rect 9364 2264 10563 2292
rect 9364 2252 9370 2264
rect 10551 2261 10563 2264
rect 10597 2261 10609 2295
rect 10551 2255 10609 2261
rect 10778 2252 10784 2304
rect 10836 2292 10842 2304
rect 12728 2292 12756 2332
rect 10836 2264 12756 2292
rect 10836 2252 10842 2264
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12860 2264 13093 2292
rect 12860 2252 12866 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13081 2255 13139 2261
rect 13262 2252 13268 2304
rect 13320 2292 13326 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13320 2264 13645 2292
rect 13320 2252 13326 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13780 2264 14289 2292
rect 13780 2252 13786 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 14550 2252 14556 2304
rect 14608 2292 14614 2304
rect 15381 2295 15439 2301
rect 15381 2292 15393 2295
rect 14608 2264 15393 2292
rect 14608 2252 14614 2264
rect 15381 2261 15393 2264
rect 15427 2261 15439 2295
rect 15381 2255 15439 2261
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 16853 2295 16911 2301
rect 16853 2292 16865 2295
rect 15528 2264 16865 2292
rect 15528 2252 15534 2264
rect 16853 2261 16865 2264
rect 16899 2261 16911 2295
rect 16853 2255 16911 2261
rect 17218 2252 17224 2304
rect 17276 2292 17282 2304
rect 17957 2295 18015 2301
rect 17957 2292 17969 2295
rect 17276 2264 17969 2292
rect 17276 2252 17282 2264
rect 17957 2261 17969 2264
rect 18003 2261 18015 2295
rect 17957 2255 18015 2261
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
rect 2406 2048 2412 2100
rect 2464 2088 2470 2100
rect 5258 2088 5264 2100
rect 2464 2060 5264 2088
rect 2464 2048 2470 2060
rect 5258 2048 5264 2060
rect 5316 2048 5322 2100
rect 5626 2048 5632 2100
rect 5684 2088 5690 2100
rect 9306 2088 9312 2100
rect 5684 2060 9312 2088
rect 5684 2048 5690 2060
rect 9306 2048 9312 2060
rect 9364 2048 9370 2100
rect 16206 2048 16212 2100
rect 16264 2088 16270 2100
rect 20530 2088 20536 2100
rect 16264 2060 20536 2088
rect 16264 2048 16270 2060
rect 20530 2048 20536 2060
rect 20588 2048 20594 2100
rect 3050 1980 3056 2032
rect 3108 2020 3114 2032
rect 7558 2020 7564 2032
rect 3108 1992 7564 2020
rect 3108 1980 3114 1992
rect 7558 1980 7564 1992
rect 7616 1980 7622 2032
rect 15102 1980 15108 2032
rect 15160 2020 15166 2032
rect 19794 2020 19800 2032
rect 15160 1992 19800 2020
rect 15160 1980 15166 1992
rect 19794 1980 19800 1992
rect 19852 1980 19858 2032
rect 9122 1912 9128 1964
rect 9180 1952 9186 1964
rect 17034 1952 17040 1964
rect 9180 1924 17040 1952
rect 9180 1912 9186 1924
rect 17034 1912 17040 1924
rect 17092 1912 17098 1964
rect 3418 1300 3424 1352
rect 3476 1340 3482 1352
rect 7190 1340 7196 1352
rect 3476 1312 7196 1340
rect 3476 1300 3482 1312
rect 7190 1300 7196 1312
rect 7248 1300 7254 1352
rect 14366 1300 14372 1352
rect 14424 1340 14430 1352
rect 18322 1340 18328 1352
rect 14424 1312 18328 1340
rect 14424 1300 14430 1312
rect 18322 1300 18328 1312
rect 18380 1300 18386 1352
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 1492 20587 1544 20596
rect 1492 20553 1501 20587
rect 1501 20553 1535 20587
rect 1535 20553 1544 20587
rect 1492 20544 1544 20553
rect 2044 20587 2096 20596
rect 2044 20553 2053 20587
rect 2053 20553 2087 20587
rect 2087 20553 2096 20587
rect 2044 20544 2096 20553
rect 2964 20544 3016 20596
rect 2964 20340 3016 20392
rect 2780 20272 2832 20324
rect 3884 20408 3936 20460
rect 9956 20544 10008 20596
rect 17224 20544 17276 20596
rect 19616 20587 19668 20596
rect 19616 20553 19625 20587
rect 19625 20553 19659 20587
rect 19659 20553 19668 20587
rect 19616 20544 19668 20553
rect 20168 20587 20220 20596
rect 20168 20553 20177 20587
rect 20177 20553 20211 20587
rect 20211 20553 20220 20587
rect 20168 20544 20220 20553
rect 4528 20408 4580 20460
rect 5724 20408 5776 20460
rect 10324 20408 10376 20460
rect 18696 20451 18748 20460
rect 18696 20417 18705 20451
rect 18705 20417 18739 20451
rect 18739 20417 18748 20451
rect 18696 20408 18748 20417
rect 18788 20408 18840 20460
rect 19524 20408 19576 20460
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 6552 20340 6604 20392
rect 20444 20340 20496 20392
rect 11244 20272 11296 20324
rect 20720 20315 20772 20324
rect 20720 20281 20729 20315
rect 20729 20281 20763 20315
rect 20763 20281 20772 20315
rect 20720 20272 20772 20281
rect 4988 20204 5040 20256
rect 18052 20204 18104 20256
rect 21364 20204 21416 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 2872 20000 2924 20052
rect 2136 19796 2188 19848
rect 2504 19796 2556 19848
rect 2780 19839 2832 19848
rect 2780 19805 2789 19839
rect 2789 19805 2823 19839
rect 2823 19805 2832 19839
rect 10324 20043 10376 20052
rect 10324 20009 10333 20043
rect 10333 20009 10367 20043
rect 10367 20009 10376 20043
rect 10324 20000 10376 20009
rect 18788 20000 18840 20052
rect 19524 20000 19576 20052
rect 20536 20000 20588 20052
rect 20260 19932 20312 19984
rect 2780 19796 2832 19805
rect 4344 19796 4396 19848
rect 5264 19796 5316 19848
rect 9496 19796 9548 19848
rect 11244 19796 11296 19848
rect 18328 19796 18380 19848
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 18696 19796 18748 19805
rect 19524 19839 19576 19848
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 20076 19796 20128 19848
rect 4804 19728 4856 19780
rect 1492 19703 1544 19712
rect 1492 19669 1501 19703
rect 1501 19669 1535 19703
rect 1535 19669 1544 19703
rect 1492 19660 1544 19669
rect 2044 19703 2096 19712
rect 2044 19669 2053 19703
rect 2053 19669 2087 19703
rect 2087 19669 2096 19703
rect 2044 19660 2096 19669
rect 3148 19660 3200 19712
rect 3332 19660 3384 19712
rect 3884 19660 3936 19712
rect 4068 19660 4120 19712
rect 9404 19728 9456 19780
rect 5724 19660 5776 19712
rect 7748 19660 7800 19712
rect 8392 19660 8444 19712
rect 12624 19660 12676 19712
rect 18328 19660 18380 19712
rect 19616 19728 19668 19780
rect 19524 19660 19576 19712
rect 20720 19703 20772 19712
rect 20720 19669 20729 19703
rect 20729 19669 20763 19703
rect 20763 19669 20772 19703
rect 20720 19660 20772 19669
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 1952 19456 2004 19508
rect 2504 19499 2556 19508
rect 2504 19465 2513 19499
rect 2513 19465 2547 19499
rect 2547 19465 2556 19499
rect 2504 19456 2556 19465
rect 4528 19456 4580 19508
rect 7748 19499 7800 19508
rect 7748 19465 7757 19499
rect 7757 19465 7791 19499
rect 7791 19465 7800 19499
rect 7748 19456 7800 19465
rect 9404 19499 9456 19508
rect 9404 19465 9413 19499
rect 9413 19465 9447 19499
rect 9447 19465 9456 19499
rect 9404 19456 9456 19465
rect 19984 19456 20036 19508
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 2688 19363 2740 19372
rect 2688 19329 2697 19363
rect 2697 19329 2731 19363
rect 2731 19329 2740 19363
rect 2688 19320 2740 19329
rect 3148 19363 3200 19372
rect 3148 19329 3157 19363
rect 3157 19329 3191 19363
rect 3191 19329 3200 19363
rect 3148 19320 3200 19329
rect 4344 19388 4396 19440
rect 3332 19252 3384 19304
rect 7840 19320 7892 19372
rect 8668 19320 8720 19372
rect 12624 19320 12676 19372
rect 13636 19320 13688 19372
rect 18696 19388 18748 19440
rect 20536 19456 20588 19508
rect 20628 19456 20680 19508
rect 14280 19320 14332 19372
rect 14464 19363 14516 19372
rect 14464 19329 14498 19363
rect 14498 19329 14516 19363
rect 14464 19320 14516 19329
rect 17960 19320 18012 19372
rect 20076 19320 20128 19372
rect 20260 19363 20312 19372
rect 20260 19329 20269 19363
rect 20269 19329 20303 19363
rect 20303 19329 20312 19363
rect 20260 19320 20312 19329
rect 20536 19363 20588 19372
rect 20536 19329 20545 19363
rect 20545 19329 20579 19363
rect 20579 19329 20588 19363
rect 20536 19320 20588 19329
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 4896 19116 4948 19168
rect 5264 19116 5316 19168
rect 5816 19159 5868 19168
rect 5816 19125 5825 19159
rect 5825 19125 5859 19159
rect 5859 19125 5868 19159
rect 5816 19116 5868 19125
rect 12900 19116 12952 19168
rect 14372 19116 14424 19168
rect 15108 19116 15160 19168
rect 15568 19159 15620 19168
rect 15568 19125 15577 19159
rect 15577 19125 15611 19159
rect 15611 19125 15620 19159
rect 15568 19116 15620 19125
rect 20352 19116 20404 19168
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1676 18912 1728 18964
rect 2136 18912 2188 18964
rect 2780 18912 2832 18964
rect 8392 18912 8444 18964
rect 13452 18912 13504 18964
rect 4620 18844 4672 18896
rect 19616 18912 19668 18964
rect 20536 18912 20588 18964
rect 1676 18751 1728 18760
rect 1676 18717 1685 18751
rect 1685 18717 1719 18751
rect 1719 18717 1728 18751
rect 1676 18708 1728 18717
rect 2136 18751 2188 18760
rect 2136 18717 2145 18751
rect 2145 18717 2179 18751
rect 2179 18717 2188 18751
rect 2136 18708 2188 18717
rect 8668 18776 8720 18828
rect 4344 18708 4396 18760
rect 5264 18708 5316 18760
rect 5724 18708 5776 18760
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 14280 18708 14332 18760
rect 15568 18708 15620 18760
rect 1308 18640 1360 18692
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 2688 18640 2740 18692
rect 6644 18640 6696 18692
rect 8668 18640 8720 18692
rect 11244 18640 11296 18692
rect 3240 18572 3292 18624
rect 3884 18572 3936 18624
rect 4620 18615 4672 18624
rect 4620 18581 4629 18615
rect 4629 18581 4663 18615
rect 4663 18581 4672 18615
rect 4620 18572 4672 18581
rect 5448 18572 5500 18624
rect 7012 18572 7064 18624
rect 9312 18615 9364 18624
rect 9312 18581 9321 18615
rect 9321 18581 9355 18615
rect 9355 18581 9364 18615
rect 9312 18572 9364 18581
rect 9404 18615 9456 18624
rect 9404 18581 9413 18615
rect 9413 18581 9447 18615
rect 9447 18581 9456 18615
rect 9404 18572 9456 18581
rect 14924 18572 14976 18624
rect 19524 18708 19576 18760
rect 20444 18844 20496 18896
rect 17040 18572 17092 18624
rect 17868 18572 17920 18624
rect 18972 18572 19024 18624
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 1676 18368 1728 18420
rect 3884 18368 3936 18420
rect 9404 18411 9456 18420
rect 9404 18377 9413 18411
rect 9413 18377 9447 18411
rect 9447 18377 9456 18411
rect 9404 18368 9456 18377
rect 3240 18300 3292 18352
rect 6644 18300 6696 18352
rect 13176 18368 13228 18420
rect 13360 18368 13412 18420
rect 20352 18411 20404 18420
rect 2688 18232 2740 18284
rect 3424 18232 3476 18284
rect 3976 18232 4028 18284
rect 3332 18207 3384 18216
rect 3332 18173 3341 18207
rect 3341 18173 3375 18207
rect 3375 18173 3384 18207
rect 3332 18164 3384 18173
rect 3884 18164 3936 18216
rect 4712 18207 4764 18216
rect 4712 18173 4721 18207
rect 4721 18173 4755 18207
rect 4755 18173 4764 18207
rect 4712 18164 4764 18173
rect 4896 18207 4948 18216
rect 4896 18173 4905 18207
rect 4905 18173 4939 18207
rect 4939 18173 4948 18207
rect 4896 18164 4948 18173
rect 2320 18096 2372 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 2780 18028 2832 18080
rect 4252 18071 4304 18080
rect 4252 18037 4261 18071
rect 4261 18037 4295 18071
rect 4295 18037 4304 18071
rect 4252 18028 4304 18037
rect 5264 18071 5316 18080
rect 5264 18037 5273 18071
rect 5273 18037 5307 18071
rect 5307 18037 5316 18071
rect 5264 18028 5316 18037
rect 11980 18275 12032 18284
rect 8668 18164 8720 18216
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 11980 18232 12032 18241
rect 13452 18232 13504 18284
rect 15108 18275 15160 18284
rect 15108 18241 15117 18275
rect 15117 18241 15151 18275
rect 15151 18241 15160 18275
rect 15108 18232 15160 18241
rect 17132 18232 17184 18284
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 20352 18377 20361 18411
rect 20361 18377 20395 18411
rect 20395 18377 20404 18411
rect 20352 18368 20404 18377
rect 20628 18275 20680 18284
rect 20628 18241 20637 18275
rect 20637 18241 20671 18275
rect 20671 18241 20680 18275
rect 20628 18232 20680 18241
rect 12900 18207 12952 18216
rect 12900 18173 12909 18207
rect 12909 18173 12943 18207
rect 12943 18173 12952 18207
rect 12900 18164 12952 18173
rect 14372 18164 14424 18216
rect 14832 18207 14884 18216
rect 14832 18173 14841 18207
rect 14841 18173 14875 18207
rect 14875 18173 14884 18207
rect 14832 18164 14884 18173
rect 14924 18164 14976 18216
rect 17684 18164 17736 18216
rect 18052 18164 18104 18216
rect 18144 18207 18196 18216
rect 18144 18173 18153 18207
rect 18153 18173 18187 18207
rect 18187 18173 18196 18207
rect 18144 18164 18196 18173
rect 20352 18164 20404 18216
rect 13268 18096 13320 18148
rect 10048 18028 10100 18080
rect 12072 18028 12124 18080
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 15384 18028 15436 18080
rect 17408 18028 17460 18080
rect 17868 18028 17920 18080
rect 18512 18071 18564 18080
rect 18512 18037 18521 18071
rect 18521 18037 18555 18071
rect 18555 18037 18564 18071
rect 18512 18028 18564 18037
rect 19708 18028 19760 18080
rect 20996 18028 21048 18080
rect 21364 18028 21416 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 4712 17824 4764 17876
rect 7748 17824 7800 17876
rect 9588 17824 9640 17876
rect 14556 17824 14608 17876
rect 15108 17867 15160 17876
rect 15108 17833 15117 17867
rect 15117 17833 15151 17867
rect 15151 17833 15160 17867
rect 15108 17824 15160 17833
rect 3240 17756 3292 17808
rect 6000 17756 6052 17808
rect 2780 17688 2832 17740
rect 3332 17688 3384 17740
rect 13820 17756 13872 17808
rect 10416 17688 10468 17740
rect 1492 17527 1544 17536
rect 1492 17493 1501 17527
rect 1501 17493 1535 17527
rect 1535 17493 1544 17527
rect 1492 17484 1544 17493
rect 2044 17484 2096 17536
rect 4252 17620 4304 17672
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 8392 17620 8444 17672
rect 9496 17620 9548 17672
rect 14372 17688 14424 17740
rect 15568 17688 15620 17740
rect 15384 17620 15436 17672
rect 18880 17663 18932 17672
rect 18880 17629 18889 17663
rect 18889 17629 18923 17663
rect 18923 17629 18932 17663
rect 18880 17620 18932 17629
rect 3148 17552 3200 17604
rect 6736 17552 6788 17604
rect 6920 17595 6972 17604
rect 6920 17561 6938 17595
rect 6938 17561 6972 17595
rect 6920 17552 6972 17561
rect 8116 17552 8168 17604
rect 12164 17552 12216 17604
rect 16212 17552 16264 17604
rect 16304 17552 16356 17604
rect 18512 17552 18564 17604
rect 19524 17824 19576 17876
rect 20352 17867 20404 17876
rect 20352 17833 20361 17867
rect 20361 17833 20395 17867
rect 20395 17833 20404 17867
rect 20352 17824 20404 17833
rect 19708 17688 19760 17740
rect 19892 17663 19944 17672
rect 19892 17629 19901 17663
rect 19901 17629 19935 17663
rect 19935 17629 19944 17663
rect 19892 17620 19944 17629
rect 20352 17552 20404 17604
rect 4988 17484 5040 17536
rect 5540 17527 5592 17536
rect 5540 17493 5549 17527
rect 5549 17493 5583 17527
rect 5583 17493 5592 17527
rect 5540 17484 5592 17493
rect 5908 17484 5960 17536
rect 7472 17527 7524 17536
rect 7472 17493 7481 17527
rect 7481 17493 7515 17527
rect 7515 17493 7524 17527
rect 7472 17484 7524 17493
rect 11980 17527 12032 17536
rect 11980 17493 11989 17527
rect 11989 17493 12023 17527
rect 12023 17493 12032 17527
rect 11980 17484 12032 17493
rect 12256 17527 12308 17536
rect 12256 17493 12265 17527
rect 12265 17493 12299 17527
rect 12299 17493 12308 17527
rect 12256 17484 12308 17493
rect 12624 17527 12676 17536
rect 12624 17493 12633 17527
rect 12633 17493 12667 17527
rect 12667 17493 12676 17527
rect 12624 17484 12676 17493
rect 14372 17527 14424 17536
rect 14372 17493 14381 17527
rect 14381 17493 14415 17527
rect 14415 17493 14424 17527
rect 14372 17484 14424 17493
rect 14556 17484 14608 17536
rect 15108 17484 15160 17536
rect 15568 17527 15620 17536
rect 15568 17493 15577 17527
rect 15577 17493 15611 17527
rect 15611 17493 15620 17527
rect 15568 17484 15620 17493
rect 16120 17527 16172 17536
rect 16120 17493 16129 17527
rect 16129 17493 16163 17527
rect 16163 17493 16172 17527
rect 16120 17484 16172 17493
rect 16396 17484 16448 17536
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 21088 17484 21140 17536
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 3884 17323 3936 17332
rect 3884 17289 3893 17323
rect 3893 17289 3927 17323
rect 3927 17289 3936 17323
rect 3884 17280 3936 17289
rect 4988 17323 5040 17332
rect 4988 17289 4997 17323
rect 4997 17289 5031 17323
rect 5031 17289 5040 17323
rect 4988 17280 5040 17289
rect 6000 17280 6052 17332
rect 6736 17280 6788 17332
rect 4896 17212 4948 17264
rect 5540 17212 5592 17264
rect 6092 17212 6144 17264
rect 2596 17187 2648 17196
rect 2596 17153 2605 17187
rect 2605 17153 2639 17187
rect 2639 17153 2648 17187
rect 2596 17144 2648 17153
rect 2964 17144 3016 17196
rect 6552 17144 6604 17196
rect 9312 17280 9364 17332
rect 12900 17280 12952 17332
rect 14372 17323 14424 17332
rect 14372 17289 14381 17323
rect 14381 17289 14415 17323
rect 14415 17289 14424 17323
rect 14372 17280 14424 17289
rect 14924 17280 14976 17332
rect 15108 17323 15160 17332
rect 15108 17289 15117 17323
rect 15117 17289 15151 17323
rect 15151 17289 15160 17323
rect 15108 17280 15160 17289
rect 16120 17280 16172 17332
rect 16396 17280 16448 17332
rect 12624 17212 12676 17264
rect 7288 17187 7340 17196
rect 7288 17153 7297 17187
rect 7297 17153 7331 17187
rect 7331 17153 7340 17187
rect 7288 17144 7340 17153
rect 10508 17144 10560 17196
rect 12348 17144 12400 17196
rect 13268 17144 13320 17196
rect 17960 17280 18012 17332
rect 18144 17323 18196 17332
rect 18144 17289 18153 17323
rect 18153 17289 18187 17323
rect 18187 17289 18196 17323
rect 18144 17280 18196 17289
rect 17408 17212 17460 17264
rect 19800 17212 19852 17264
rect 3240 17076 3292 17128
rect 1492 17051 1544 17060
rect 1492 17017 1501 17051
rect 1501 17017 1535 17051
rect 1535 17017 1544 17051
rect 1492 17008 1544 17017
rect 2872 17008 2924 17060
rect 5816 17119 5868 17128
rect 5816 17085 5825 17119
rect 5825 17085 5859 17119
rect 5859 17085 5868 17119
rect 7380 17119 7432 17128
rect 5816 17076 5868 17085
rect 7380 17085 7389 17119
rect 7389 17085 7423 17119
rect 7423 17085 7432 17119
rect 7380 17076 7432 17085
rect 8116 17119 8168 17128
rect 1952 16983 2004 16992
rect 1952 16949 1961 16983
rect 1961 16949 1995 16983
rect 1995 16949 2004 16983
rect 1952 16940 2004 16949
rect 5908 17008 5960 17060
rect 8116 17085 8125 17119
rect 8125 17085 8159 17119
rect 8159 17085 8168 17119
rect 8116 17076 8168 17085
rect 8576 17076 8628 17128
rect 9588 17119 9640 17128
rect 9588 17085 9597 17119
rect 9597 17085 9631 17119
rect 9631 17085 9640 17119
rect 9588 17076 9640 17085
rect 8668 17008 8720 17060
rect 10416 17076 10468 17128
rect 11060 17076 11112 17128
rect 12164 17076 12216 17128
rect 13636 17076 13688 17128
rect 17776 17144 17828 17196
rect 4804 16940 4856 16992
rect 6092 16940 6144 16992
rect 12532 17008 12584 17060
rect 14648 17076 14700 17128
rect 15476 17076 15528 17128
rect 17132 17119 17184 17128
rect 17132 17085 17141 17119
rect 17141 17085 17175 17119
rect 17175 17085 17184 17119
rect 17132 17076 17184 17085
rect 17224 17119 17276 17128
rect 17224 17085 17233 17119
rect 17233 17085 17267 17119
rect 17267 17085 17276 17119
rect 17224 17076 17276 17085
rect 17500 17076 17552 17128
rect 18880 17144 18932 17196
rect 20628 17280 20680 17332
rect 20812 17144 20864 17196
rect 21088 17187 21140 17196
rect 21088 17153 21097 17187
rect 21097 17153 21131 17187
rect 21131 17153 21140 17187
rect 21088 17144 21140 17153
rect 15108 17008 15160 17060
rect 17960 17008 18012 17060
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 11796 16940 11848 16992
rect 13820 16940 13872 16992
rect 17132 16940 17184 16992
rect 21088 16940 21140 16992
rect 21272 16983 21324 16992
rect 21272 16949 21281 16983
rect 21281 16949 21315 16983
rect 21315 16949 21324 16983
rect 21272 16940 21324 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 2780 16736 2832 16788
rect 5816 16779 5868 16788
rect 2504 16668 2556 16720
rect 5816 16745 5825 16779
rect 5825 16745 5859 16779
rect 5859 16745 5868 16779
rect 5816 16736 5868 16745
rect 7288 16736 7340 16788
rect 8576 16779 8628 16788
rect 2872 16643 2924 16652
rect 2872 16609 2881 16643
rect 2881 16609 2915 16643
rect 2915 16609 2924 16643
rect 2872 16600 2924 16609
rect 7656 16668 7708 16720
rect 8576 16745 8585 16779
rect 8585 16745 8619 16779
rect 8619 16745 8628 16779
rect 8576 16736 8628 16745
rect 8668 16736 8720 16788
rect 10508 16736 10560 16788
rect 12624 16736 12676 16788
rect 10692 16668 10744 16720
rect 3240 16600 3292 16652
rect 4344 16600 4396 16652
rect 5632 16600 5684 16652
rect 1676 16575 1728 16584
rect 1676 16541 1685 16575
rect 1685 16541 1719 16575
rect 1719 16541 1728 16575
rect 1676 16532 1728 16541
rect 1952 16575 2004 16584
rect 1952 16541 1961 16575
rect 1961 16541 1995 16575
rect 1995 16541 2004 16575
rect 1952 16532 2004 16541
rect 3148 16532 3200 16584
rect 5816 16532 5868 16584
rect 6920 16532 6972 16584
rect 8668 16600 8720 16652
rect 9496 16532 9548 16584
rect 10968 16600 11020 16652
rect 11980 16600 12032 16652
rect 11152 16532 11204 16584
rect 5724 16464 5776 16516
rect 10324 16464 10376 16516
rect 12256 16600 12308 16652
rect 12900 16600 12952 16652
rect 15568 16736 15620 16788
rect 16304 16736 16356 16788
rect 17776 16736 17828 16788
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 20812 16779 20864 16788
rect 20812 16745 20821 16779
rect 20821 16745 20855 16779
rect 20855 16745 20864 16779
rect 20812 16736 20864 16745
rect 13636 16668 13688 16720
rect 16028 16711 16080 16720
rect 14464 16600 14516 16652
rect 15108 16643 15160 16652
rect 15108 16609 15117 16643
rect 15117 16609 15151 16643
rect 15151 16609 15160 16643
rect 15108 16600 15160 16609
rect 16028 16677 16037 16711
rect 16037 16677 16071 16711
rect 16071 16677 16080 16711
rect 16028 16668 16080 16677
rect 16212 16668 16264 16720
rect 17592 16668 17644 16720
rect 17224 16600 17276 16652
rect 17868 16643 17920 16652
rect 17868 16609 17877 16643
rect 17877 16609 17911 16643
rect 17911 16609 17920 16643
rect 17868 16600 17920 16609
rect 17592 16532 17644 16584
rect 17684 16532 17736 16584
rect 20352 16600 20404 16652
rect 18512 16532 18564 16584
rect 19800 16532 19852 16584
rect 20168 16575 20220 16584
rect 20168 16541 20177 16575
rect 20177 16541 20211 16575
rect 20211 16541 20220 16575
rect 20168 16532 20220 16541
rect 20720 16532 20772 16584
rect 1492 16439 1544 16448
rect 1492 16405 1501 16439
rect 1501 16405 1535 16439
rect 1535 16405 1544 16439
rect 1492 16396 1544 16405
rect 2136 16439 2188 16448
rect 2136 16405 2145 16439
rect 2145 16405 2179 16439
rect 2179 16405 2188 16439
rect 2136 16396 2188 16405
rect 3424 16439 3476 16448
rect 3424 16405 3433 16439
rect 3433 16405 3467 16439
rect 3467 16405 3476 16439
rect 3424 16396 3476 16405
rect 7104 16396 7156 16448
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 12900 16396 12952 16448
rect 15016 16396 15068 16448
rect 17684 16396 17736 16448
rect 17960 16396 18012 16448
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 2596 16235 2648 16244
rect 2596 16201 2605 16235
rect 2605 16201 2639 16235
rect 2639 16201 2648 16235
rect 2596 16192 2648 16201
rect 3332 16192 3384 16244
rect 11060 16192 11112 16244
rect 2688 16124 2740 16176
rect 4804 16056 4856 16108
rect 2872 15988 2924 16040
rect 3976 15988 4028 16040
rect 7564 16124 7616 16176
rect 5080 15988 5132 16040
rect 9128 16099 9180 16108
rect 9128 16065 9137 16099
rect 9137 16065 9171 16099
rect 9171 16065 9180 16099
rect 9128 16056 9180 16065
rect 11060 16056 11112 16108
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 14556 16099 14608 16108
rect 14556 16065 14565 16099
rect 14565 16065 14599 16099
rect 14599 16065 14608 16099
rect 14556 16056 14608 16065
rect 6736 15988 6788 16040
rect 8024 15988 8076 16040
rect 8208 15988 8260 16040
rect 5540 15963 5592 15972
rect 5540 15929 5549 15963
rect 5549 15929 5583 15963
rect 5583 15929 5592 15963
rect 5540 15920 5592 15929
rect 7380 15920 7432 15972
rect 12164 16031 12216 16040
rect 12164 15997 12173 16031
rect 12173 15997 12207 16031
rect 12207 15997 12216 16031
rect 12164 15988 12216 15997
rect 13820 15988 13872 16040
rect 18328 16192 18380 16244
rect 19616 16192 19668 16244
rect 20168 16235 20220 16244
rect 20168 16201 20177 16235
rect 20177 16201 20211 16235
rect 20211 16201 20220 16235
rect 20168 16192 20220 16201
rect 18604 16124 18656 16176
rect 15200 16099 15252 16108
rect 15200 16065 15209 16099
rect 15209 16065 15243 16099
rect 15243 16065 15252 16099
rect 15200 16056 15252 16065
rect 17500 16099 17552 16108
rect 17500 16065 17509 16099
rect 17509 16065 17543 16099
rect 17543 16065 17552 16099
rect 17500 16056 17552 16065
rect 18052 16056 18104 16108
rect 18236 16056 18288 16108
rect 12808 15920 12860 15972
rect 19064 15988 19116 16040
rect 15016 15920 15068 15972
rect 1492 15895 1544 15904
rect 1492 15861 1501 15895
rect 1501 15861 1535 15895
rect 1535 15861 1544 15895
rect 1492 15852 1544 15861
rect 4160 15852 4212 15904
rect 4988 15852 5040 15904
rect 7104 15852 7156 15904
rect 8484 15852 8536 15904
rect 9496 15895 9548 15904
rect 9496 15861 9505 15895
rect 9505 15861 9539 15895
rect 9539 15861 9548 15895
rect 9496 15852 9548 15861
rect 9864 15895 9916 15904
rect 9864 15861 9873 15895
rect 9873 15861 9907 15895
rect 9907 15861 9916 15895
rect 9864 15852 9916 15861
rect 10692 15895 10744 15904
rect 10692 15861 10701 15895
rect 10701 15861 10735 15895
rect 10735 15861 10744 15895
rect 10692 15852 10744 15861
rect 11060 15895 11112 15904
rect 11060 15861 11069 15895
rect 11069 15861 11103 15895
rect 11103 15861 11112 15895
rect 11060 15852 11112 15861
rect 13820 15895 13872 15904
rect 13820 15861 13829 15895
rect 13829 15861 13863 15895
rect 13863 15861 13872 15895
rect 13820 15852 13872 15861
rect 14464 15852 14516 15904
rect 15752 15852 15804 15904
rect 16212 15895 16264 15904
rect 16212 15861 16221 15895
rect 16221 15861 16255 15895
rect 16255 15861 16264 15895
rect 16212 15852 16264 15861
rect 17408 15852 17460 15904
rect 18420 15852 18472 15904
rect 18512 15852 18564 15904
rect 21272 15895 21324 15904
rect 21272 15861 21281 15895
rect 21281 15861 21315 15895
rect 21315 15861 21324 15895
rect 21272 15852 21324 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1676 15648 1728 15700
rect 2044 15512 2096 15564
rect 2504 15444 2556 15496
rect 5264 15648 5316 15700
rect 7288 15648 7340 15700
rect 9680 15648 9732 15700
rect 10324 15691 10376 15700
rect 10324 15657 10333 15691
rect 10333 15657 10367 15691
rect 10367 15657 10376 15691
rect 10324 15648 10376 15657
rect 12808 15691 12860 15700
rect 8668 15580 8720 15632
rect 12808 15657 12817 15691
rect 12817 15657 12851 15691
rect 12851 15657 12860 15691
rect 12808 15648 12860 15657
rect 17684 15648 17736 15700
rect 18328 15580 18380 15632
rect 18420 15623 18472 15632
rect 18420 15589 18429 15623
rect 18429 15589 18463 15623
rect 18463 15589 18472 15623
rect 18420 15580 18472 15589
rect 4344 15444 4396 15496
rect 7196 15444 7248 15496
rect 7932 15487 7984 15496
rect 7932 15453 7941 15487
rect 7941 15453 7975 15487
rect 7975 15453 7984 15487
rect 7932 15444 7984 15453
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 2136 15351 2188 15360
rect 2136 15317 2145 15351
rect 2145 15317 2179 15351
rect 2179 15317 2188 15351
rect 2136 15308 2188 15317
rect 2596 15308 2648 15360
rect 3148 15308 3200 15360
rect 5172 15351 5224 15360
rect 5172 15317 5181 15351
rect 5181 15317 5215 15351
rect 5215 15317 5224 15351
rect 5172 15308 5224 15317
rect 5908 15351 5960 15360
rect 5908 15317 5917 15351
rect 5917 15317 5951 15351
rect 5951 15317 5960 15351
rect 5908 15308 5960 15317
rect 6920 15376 6972 15428
rect 7012 15419 7064 15428
rect 7012 15385 7030 15419
rect 7030 15385 7064 15419
rect 11060 15512 11112 15564
rect 14188 15555 14240 15564
rect 14188 15521 14197 15555
rect 14197 15521 14231 15555
rect 14231 15521 14240 15555
rect 14188 15512 14240 15521
rect 14556 15512 14608 15564
rect 19156 15512 19208 15564
rect 20720 15648 20772 15700
rect 9588 15444 9640 15496
rect 10968 15444 11020 15496
rect 12072 15444 12124 15496
rect 14464 15487 14516 15496
rect 14464 15453 14473 15487
rect 14473 15453 14507 15487
rect 14507 15453 14516 15487
rect 14464 15444 14516 15453
rect 17500 15444 17552 15496
rect 17960 15444 18012 15496
rect 19064 15444 19116 15496
rect 20628 15487 20680 15496
rect 9312 15419 9364 15428
rect 7012 15376 7064 15385
rect 9312 15385 9321 15419
rect 9321 15385 9355 15419
rect 9355 15385 9364 15419
rect 9312 15376 9364 15385
rect 8576 15351 8628 15360
rect 8576 15317 8585 15351
rect 8585 15317 8619 15351
rect 8619 15317 8628 15351
rect 8576 15308 8628 15317
rect 8668 15308 8720 15360
rect 10600 15351 10652 15360
rect 10600 15317 10609 15351
rect 10609 15317 10643 15351
rect 10643 15317 10652 15351
rect 10600 15308 10652 15317
rect 13360 15308 13412 15360
rect 15660 15376 15712 15428
rect 17040 15376 17092 15428
rect 18144 15376 18196 15428
rect 18420 15376 18472 15428
rect 20628 15453 20637 15487
rect 20637 15453 20671 15487
rect 20671 15453 20680 15487
rect 20628 15444 20680 15453
rect 21088 15487 21140 15496
rect 21088 15453 21097 15487
rect 21097 15453 21131 15487
rect 21131 15453 21140 15487
rect 21088 15444 21140 15453
rect 15016 15308 15068 15360
rect 19432 15351 19484 15360
rect 19432 15317 19441 15351
rect 19441 15317 19475 15351
rect 19475 15317 19484 15351
rect 19432 15308 19484 15317
rect 20720 15308 20772 15360
rect 21088 15308 21140 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 5724 15104 5776 15156
rect 9496 15104 9548 15156
rect 3148 15036 3200 15088
rect 1952 14968 2004 15020
rect 2136 15011 2188 15020
rect 2136 14977 2145 15011
rect 2145 14977 2179 15011
rect 2179 14977 2188 15011
rect 2136 14968 2188 14977
rect 4068 14968 4120 15020
rect 4252 14968 4304 15020
rect 5172 15011 5224 15020
rect 5172 14977 5181 15011
rect 5181 14977 5215 15011
rect 5215 14977 5224 15011
rect 5172 14968 5224 14977
rect 6000 14968 6052 15020
rect 7288 14968 7340 15020
rect 8576 15036 8628 15088
rect 15200 15104 15252 15156
rect 15660 15147 15712 15156
rect 15660 15113 15669 15147
rect 15669 15113 15703 15147
rect 15703 15113 15712 15147
rect 15660 15104 15712 15113
rect 18052 15147 18104 15156
rect 9220 14968 9272 15020
rect 10692 15011 10744 15020
rect 10692 14977 10710 15011
rect 10710 14977 10744 15011
rect 10692 14968 10744 14977
rect 12808 14968 12860 15020
rect 14188 15036 14240 15088
rect 14372 15036 14424 15088
rect 13636 15011 13688 15020
rect 13636 14977 13645 15011
rect 13645 14977 13679 15011
rect 13679 14977 13688 15011
rect 13636 14968 13688 14977
rect 16580 14968 16632 15020
rect 17500 15036 17552 15088
rect 18052 15113 18061 15147
rect 18061 15113 18095 15147
rect 18095 15113 18104 15147
rect 18052 15104 18104 15113
rect 19432 15104 19484 15156
rect 20628 15104 20680 15156
rect 18236 15036 18288 15088
rect 16948 15011 17000 15020
rect 16948 14977 16982 15011
rect 16982 14977 17000 15011
rect 16948 14968 17000 14977
rect 18788 14968 18840 15020
rect 4344 14900 4396 14952
rect 4804 14900 4856 14952
rect 5356 14832 5408 14884
rect 7840 14900 7892 14952
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 1676 14764 1728 14816
rect 2596 14807 2648 14816
rect 2596 14773 2605 14807
rect 2605 14773 2639 14807
rect 2639 14773 2648 14807
rect 2596 14764 2648 14773
rect 4528 14764 4580 14816
rect 7564 14764 7616 14816
rect 10968 14943 11020 14952
rect 10968 14909 10977 14943
rect 10977 14909 11011 14943
rect 11011 14909 11020 14943
rect 10968 14900 11020 14909
rect 15200 14900 15252 14952
rect 15568 14943 15620 14952
rect 15568 14909 15577 14943
rect 15577 14909 15611 14943
rect 15611 14909 15620 14943
rect 15568 14900 15620 14909
rect 18512 14943 18564 14952
rect 18512 14909 18521 14943
rect 18521 14909 18555 14943
rect 18555 14909 18564 14943
rect 18512 14900 18564 14909
rect 18880 14900 18932 14952
rect 9128 14764 9180 14816
rect 9588 14807 9640 14816
rect 9588 14773 9597 14807
rect 9597 14773 9631 14807
rect 9631 14773 9640 14807
rect 9588 14764 9640 14773
rect 19708 14968 19760 15020
rect 19524 14900 19576 14952
rect 19892 14943 19944 14952
rect 19892 14909 19901 14943
rect 19901 14909 19935 14943
rect 19935 14909 19944 14943
rect 19892 14900 19944 14909
rect 13636 14764 13688 14816
rect 14280 14764 14332 14816
rect 17040 14764 17092 14816
rect 20720 14968 20772 15020
rect 18420 14764 18472 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1952 14603 2004 14612
rect 1952 14569 1961 14603
rect 1961 14569 1995 14603
rect 1995 14569 2004 14603
rect 1952 14560 2004 14569
rect 2504 14560 2556 14612
rect 1216 14492 1268 14544
rect 1676 14399 1728 14408
rect 1676 14365 1685 14399
rect 1685 14365 1719 14399
rect 1719 14365 1728 14399
rect 1676 14356 1728 14365
rect 3148 14424 3200 14476
rect 4252 14424 4304 14476
rect 2596 14356 2648 14408
rect 4436 14424 4488 14476
rect 6920 14560 6972 14612
rect 7932 14603 7984 14612
rect 7932 14569 7941 14603
rect 7941 14569 7975 14603
rect 7975 14569 7984 14603
rect 7932 14560 7984 14569
rect 8116 14560 8168 14612
rect 13360 14560 13412 14612
rect 15568 14560 15620 14612
rect 16948 14560 17000 14612
rect 17960 14560 18012 14612
rect 17224 14492 17276 14544
rect 17316 14492 17368 14544
rect 17684 14492 17736 14544
rect 8300 14424 8352 14476
rect 4712 14356 4764 14408
rect 9128 14399 9180 14408
rect 3884 14288 3936 14340
rect 4620 14288 4672 14340
rect 6828 14331 6880 14340
rect 6828 14297 6862 14331
rect 6862 14297 6880 14331
rect 6828 14288 6880 14297
rect 9128 14365 9137 14399
rect 9137 14365 9171 14399
rect 9171 14365 9180 14399
rect 9128 14356 9180 14365
rect 12808 14424 12860 14476
rect 14372 14424 14424 14476
rect 18052 14424 18104 14476
rect 18512 14560 18564 14612
rect 18880 14603 18932 14612
rect 18880 14569 18889 14603
rect 18889 14569 18923 14603
rect 18923 14569 18932 14603
rect 18880 14560 18932 14569
rect 19524 14603 19576 14612
rect 19524 14569 19533 14603
rect 19533 14569 19567 14603
rect 19567 14569 19576 14603
rect 19524 14560 19576 14569
rect 19064 14492 19116 14544
rect 10508 14356 10560 14408
rect 11796 14399 11848 14408
rect 11796 14365 11805 14399
rect 11805 14365 11839 14399
rect 11839 14365 11848 14399
rect 11796 14356 11848 14365
rect 12072 14356 12124 14408
rect 15660 14356 15712 14408
rect 16580 14356 16632 14408
rect 16948 14356 17000 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 4160 14263 4212 14272
rect 4160 14229 4169 14263
rect 4169 14229 4203 14263
rect 4203 14229 4212 14263
rect 4160 14220 4212 14229
rect 4804 14263 4856 14272
rect 4804 14229 4813 14263
rect 4813 14229 4847 14263
rect 4847 14229 4856 14263
rect 4804 14220 4856 14229
rect 5080 14220 5132 14272
rect 6644 14220 6696 14272
rect 8116 14220 8168 14272
rect 9496 14288 9548 14340
rect 11888 14288 11940 14340
rect 12256 14288 12308 14340
rect 17132 14288 17184 14340
rect 18880 14424 18932 14476
rect 20536 14424 20588 14476
rect 18696 14356 18748 14408
rect 19340 14356 19392 14408
rect 19616 14356 19668 14408
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 19800 14288 19852 14340
rect 20076 14288 20128 14340
rect 9772 14220 9824 14272
rect 10692 14220 10744 14272
rect 11244 14220 11296 14272
rect 13360 14263 13412 14272
rect 13360 14229 13369 14263
rect 13369 14229 13403 14263
rect 13403 14229 13412 14263
rect 13360 14220 13412 14229
rect 14372 14263 14424 14272
rect 14372 14229 14381 14263
rect 14381 14229 14415 14263
rect 14415 14229 14424 14263
rect 14372 14220 14424 14229
rect 15476 14263 15528 14272
rect 15476 14229 15485 14263
rect 15485 14229 15519 14263
rect 15519 14229 15528 14263
rect 15476 14220 15528 14229
rect 17316 14220 17368 14272
rect 21180 14288 21232 14340
rect 21088 14220 21140 14272
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 3056 14016 3108 14068
rect 6000 14059 6052 14068
rect 1676 13923 1728 13932
rect 1676 13889 1685 13923
rect 1685 13889 1719 13923
rect 1719 13889 1728 13923
rect 1676 13880 1728 13889
rect 2780 13923 2832 13932
rect 2780 13889 2789 13923
rect 2789 13889 2823 13923
rect 2823 13889 2832 13923
rect 2780 13880 2832 13889
rect 2136 13855 2188 13864
rect 2136 13821 2145 13855
rect 2145 13821 2179 13855
rect 2179 13821 2188 13855
rect 2136 13812 2188 13821
rect 2596 13855 2648 13864
rect 2596 13821 2605 13855
rect 2605 13821 2639 13855
rect 2639 13821 2648 13855
rect 2596 13812 2648 13821
rect 3056 13812 3108 13864
rect 3424 13855 3476 13864
rect 3424 13821 3433 13855
rect 3433 13821 3467 13855
rect 3467 13821 3476 13855
rect 3424 13812 3476 13821
rect 1492 13787 1544 13796
rect 1492 13753 1501 13787
rect 1501 13753 1535 13787
rect 1535 13753 1544 13787
rect 1492 13744 1544 13753
rect 4712 13880 4764 13932
rect 3148 13676 3200 13728
rect 4068 13676 4120 13728
rect 4252 13719 4304 13728
rect 4252 13685 4261 13719
rect 4261 13685 4295 13719
rect 4295 13685 4304 13719
rect 4252 13676 4304 13685
rect 4712 13676 4764 13728
rect 4896 13676 4948 13728
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6644 14016 6696 14068
rect 8300 14016 8352 14068
rect 8392 14016 8444 14068
rect 6000 13880 6052 13932
rect 6644 13880 6696 13932
rect 11888 14059 11940 14068
rect 11888 14025 11897 14059
rect 11897 14025 11931 14059
rect 11931 14025 11940 14059
rect 12256 14059 12308 14068
rect 11888 14016 11940 14025
rect 12256 14025 12265 14059
rect 12265 14025 12299 14059
rect 12299 14025 12308 14059
rect 12256 14016 12308 14025
rect 14372 14016 14424 14068
rect 17040 14016 17092 14068
rect 17868 14016 17920 14068
rect 18420 14059 18472 14068
rect 18420 14025 18429 14059
rect 18429 14025 18463 14059
rect 18463 14025 18472 14059
rect 18420 14016 18472 14025
rect 18788 14059 18840 14068
rect 18788 14025 18797 14059
rect 18797 14025 18831 14059
rect 18831 14025 18840 14059
rect 18788 14016 18840 14025
rect 6460 13855 6512 13864
rect 6460 13821 6469 13855
rect 6469 13821 6503 13855
rect 6503 13821 6512 13855
rect 6460 13812 6512 13821
rect 6736 13855 6788 13864
rect 6736 13821 6745 13855
rect 6745 13821 6779 13855
rect 6779 13821 6788 13855
rect 6736 13812 6788 13821
rect 5908 13744 5960 13796
rect 6828 13744 6880 13796
rect 7104 13744 7156 13796
rect 7656 13812 7708 13864
rect 8300 13812 8352 13864
rect 8116 13744 8168 13796
rect 11244 13948 11296 14000
rect 14924 13991 14976 14000
rect 8944 13923 8996 13932
rect 8944 13889 8953 13923
rect 8953 13889 8987 13923
rect 8987 13889 8996 13923
rect 9956 13923 10008 13932
rect 8944 13880 8996 13889
rect 9956 13889 9965 13923
rect 9965 13889 9999 13923
rect 9999 13889 10008 13923
rect 9956 13880 10008 13889
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 9588 13812 9640 13864
rect 9220 13744 9272 13796
rect 9496 13744 9548 13796
rect 14924 13957 14933 13991
rect 14933 13957 14967 13991
rect 14967 13957 14976 13991
rect 14924 13948 14976 13957
rect 12808 13880 12860 13932
rect 14464 13880 14516 13932
rect 15384 13880 15436 13932
rect 16304 13923 16356 13932
rect 16304 13889 16313 13923
rect 16313 13889 16347 13923
rect 16347 13889 16356 13923
rect 16304 13880 16356 13889
rect 18512 13948 18564 14000
rect 20352 14016 20404 14068
rect 21272 14059 21324 14068
rect 21272 14025 21281 14059
rect 21281 14025 21315 14059
rect 21315 14025 21324 14059
rect 21272 14016 21324 14025
rect 19340 13948 19392 14000
rect 20444 13991 20496 14000
rect 20444 13957 20453 13991
rect 20453 13957 20487 13991
rect 20487 13957 20496 13991
rect 20444 13948 20496 13957
rect 12532 13855 12584 13864
rect 12532 13821 12541 13855
rect 12541 13821 12575 13855
rect 12575 13821 12584 13855
rect 12532 13812 12584 13821
rect 12440 13744 12492 13796
rect 13084 13855 13136 13864
rect 13084 13821 13093 13855
rect 13093 13821 13127 13855
rect 13127 13821 13136 13855
rect 13084 13812 13136 13821
rect 13544 13812 13596 13864
rect 14740 13812 14792 13864
rect 18696 13880 18748 13932
rect 19524 13880 19576 13932
rect 21088 13923 21140 13932
rect 21088 13889 21097 13923
rect 21097 13889 21131 13923
rect 21131 13889 21140 13923
rect 21088 13880 21140 13889
rect 17500 13812 17552 13864
rect 18052 13812 18104 13864
rect 18328 13855 18380 13864
rect 18328 13821 18337 13855
rect 18337 13821 18371 13855
rect 18371 13821 18380 13855
rect 18328 13812 18380 13821
rect 17132 13744 17184 13796
rect 17960 13744 18012 13796
rect 20628 13855 20680 13864
rect 20628 13821 20637 13855
rect 20637 13821 20671 13855
rect 20671 13821 20680 13855
rect 20628 13812 20680 13821
rect 19800 13744 19852 13796
rect 7748 13676 7800 13728
rect 9588 13719 9640 13728
rect 9588 13685 9597 13719
rect 9597 13685 9631 13719
rect 9631 13685 9640 13719
rect 9588 13676 9640 13685
rect 12716 13676 12768 13728
rect 17316 13676 17368 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2780 13472 2832 13524
rect 3424 13472 3476 13524
rect 3884 13472 3936 13524
rect 4068 13472 4120 13524
rect 2228 13404 2280 13456
rect 2412 13404 2464 13456
rect 2044 13336 2096 13388
rect 3148 13336 3200 13388
rect 2136 13268 2188 13320
rect 3424 13268 3476 13320
rect 4252 13404 4304 13456
rect 5264 13472 5316 13524
rect 7288 13515 7340 13524
rect 7288 13481 7297 13515
rect 7297 13481 7331 13515
rect 7331 13481 7340 13515
rect 7288 13472 7340 13481
rect 9220 13515 9272 13524
rect 9220 13481 9229 13515
rect 9229 13481 9263 13515
rect 9263 13481 9272 13515
rect 9220 13472 9272 13481
rect 9956 13472 10008 13524
rect 12348 13472 12400 13524
rect 12900 13472 12952 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 17868 13472 17920 13524
rect 18328 13472 18380 13524
rect 6828 13404 6880 13456
rect 21640 13472 21692 13524
rect 7748 13379 7800 13388
rect 7748 13345 7757 13379
rect 7757 13345 7791 13379
rect 7791 13345 7800 13379
rect 7748 13336 7800 13345
rect 9588 13336 9640 13388
rect 9772 13379 9824 13388
rect 9772 13345 9781 13379
rect 9781 13345 9815 13379
rect 9815 13345 9824 13379
rect 12256 13379 12308 13388
rect 9772 13336 9824 13345
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 12256 13336 12308 13345
rect 13084 13336 13136 13388
rect 2228 13200 2280 13252
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 1860 13132 1912 13184
rect 4344 13200 4396 13252
rect 8300 13268 8352 13320
rect 11888 13268 11940 13320
rect 12992 13268 13044 13320
rect 13360 13268 13412 13320
rect 13820 13268 13872 13320
rect 16948 13336 17000 13388
rect 17960 13336 18012 13388
rect 19800 13379 19852 13388
rect 19800 13345 19809 13379
rect 19809 13345 19843 13379
rect 19843 13345 19852 13379
rect 19800 13336 19852 13345
rect 20444 13404 20496 13456
rect 20628 13404 20680 13456
rect 20904 13336 20956 13388
rect 17408 13268 17460 13320
rect 18328 13268 18380 13320
rect 18696 13311 18748 13320
rect 18696 13277 18705 13311
rect 18705 13277 18739 13311
rect 18739 13277 18748 13311
rect 18696 13268 18748 13277
rect 20996 13268 21048 13320
rect 7196 13200 7248 13252
rect 7472 13200 7524 13252
rect 9864 13200 9916 13252
rect 15200 13200 15252 13252
rect 15568 13200 15620 13252
rect 15936 13200 15988 13252
rect 20260 13200 20312 13252
rect 20352 13243 20404 13252
rect 20352 13209 20361 13243
rect 20361 13209 20395 13243
rect 20395 13209 20404 13243
rect 20352 13200 20404 13209
rect 2596 13175 2648 13184
rect 2596 13141 2605 13175
rect 2605 13141 2639 13175
rect 2639 13141 2648 13175
rect 2596 13132 2648 13141
rect 3332 13175 3384 13184
rect 3332 13141 3341 13175
rect 3341 13141 3375 13175
rect 3375 13141 3384 13175
rect 3332 13132 3384 13141
rect 4252 13175 4304 13184
rect 4252 13141 4261 13175
rect 4261 13141 4295 13175
rect 4295 13141 4304 13175
rect 4252 13132 4304 13141
rect 7288 13132 7340 13184
rect 7748 13132 7800 13184
rect 10048 13132 10100 13184
rect 10784 13175 10836 13184
rect 10784 13141 10793 13175
rect 10793 13141 10827 13175
rect 10827 13141 10836 13175
rect 10784 13132 10836 13141
rect 11244 13132 11296 13184
rect 11704 13132 11756 13184
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13268 13175 13320 13184
rect 13268 13141 13277 13175
rect 13277 13141 13311 13175
rect 13311 13141 13320 13175
rect 13268 13132 13320 13141
rect 13360 13132 13412 13184
rect 14924 13132 14976 13184
rect 17408 13132 17460 13184
rect 18880 13132 18932 13184
rect 19708 13175 19760 13184
rect 19708 13141 19717 13175
rect 19717 13141 19751 13175
rect 19751 13141 19760 13175
rect 21272 13175 21324 13184
rect 19708 13132 19760 13141
rect 21272 13141 21281 13175
rect 21281 13141 21315 13175
rect 21315 13141 21324 13175
rect 21272 13132 21324 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 2504 12971 2556 12980
rect 2504 12937 2513 12971
rect 2513 12937 2547 12971
rect 2547 12937 2556 12971
rect 2504 12928 2556 12937
rect 2596 12928 2648 12980
rect 4068 12928 4120 12980
rect 4252 12928 4304 12980
rect 4436 12928 4488 12980
rect 5264 12928 5316 12980
rect 6000 12928 6052 12980
rect 7748 12928 7800 12980
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 10508 12971 10560 12980
rect 10508 12937 10517 12971
rect 10517 12937 10551 12971
rect 10551 12937 10560 12971
rect 11060 12971 11112 12980
rect 10508 12928 10560 12937
rect 11060 12937 11069 12971
rect 11069 12937 11103 12971
rect 11103 12937 11112 12971
rect 11060 12928 11112 12937
rect 15936 12971 15988 12980
rect 15936 12937 15945 12971
rect 15945 12937 15979 12971
rect 15979 12937 15988 12971
rect 15936 12928 15988 12937
rect 16948 12971 17000 12980
rect 16948 12937 16957 12971
rect 16957 12937 16991 12971
rect 16991 12937 17000 12971
rect 16948 12928 17000 12937
rect 17040 12928 17092 12980
rect 17408 12971 17460 12980
rect 1584 12792 1636 12844
rect 3332 12860 3384 12912
rect 4528 12903 4580 12912
rect 4528 12869 4537 12903
rect 4537 12869 4571 12903
rect 4571 12869 4580 12903
rect 4528 12860 4580 12869
rect 7380 12903 7432 12912
rect 7380 12869 7389 12903
rect 7389 12869 7423 12903
rect 7423 12869 7432 12903
rect 7380 12860 7432 12869
rect 8300 12860 8352 12912
rect 13084 12860 13136 12912
rect 15476 12903 15528 12912
rect 15476 12869 15485 12903
rect 15485 12869 15519 12903
rect 15519 12869 15528 12903
rect 15476 12860 15528 12869
rect 1860 12792 1912 12844
rect 4068 12792 4120 12844
rect 7932 12792 7984 12844
rect 12348 12792 12400 12844
rect 15200 12792 15252 12844
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 3148 12724 3200 12776
rect 4436 12724 4488 12776
rect 5264 12724 5316 12776
rect 6000 12767 6052 12776
rect 6000 12733 6009 12767
rect 6009 12733 6043 12767
rect 6043 12733 6052 12767
rect 6000 12724 6052 12733
rect 6828 12767 6880 12776
rect 6828 12733 6837 12767
rect 6837 12733 6871 12767
rect 6871 12733 6880 12767
rect 6828 12724 6880 12733
rect 7104 12724 7156 12776
rect 7656 12724 7708 12776
rect 8392 12656 8444 12708
rect 9220 12724 9272 12776
rect 9496 12724 9548 12776
rect 11796 12767 11848 12776
rect 11796 12733 11805 12767
rect 11805 12733 11839 12767
rect 11839 12733 11848 12767
rect 11796 12724 11848 12733
rect 15384 12767 15436 12776
rect 9404 12656 9456 12708
rect 10140 12656 10192 12708
rect 15384 12733 15393 12767
rect 15393 12733 15427 12767
rect 15427 12733 15436 12767
rect 15384 12724 15436 12733
rect 11980 12656 12032 12708
rect 1952 12588 2004 12640
rect 5908 12588 5960 12640
rect 8484 12588 8536 12640
rect 9128 12631 9180 12640
rect 9128 12597 9137 12631
rect 9137 12597 9171 12631
rect 9171 12597 9180 12631
rect 9128 12588 9180 12597
rect 12532 12588 12584 12640
rect 13636 12588 13688 12640
rect 14280 12631 14332 12640
rect 14280 12597 14289 12631
rect 14289 12597 14323 12631
rect 14323 12597 14332 12631
rect 14280 12588 14332 12597
rect 17408 12937 17417 12971
rect 17417 12937 17451 12971
rect 17451 12937 17460 12971
rect 17408 12928 17460 12937
rect 17500 12928 17552 12980
rect 19340 12928 19392 12980
rect 19708 12928 19760 12980
rect 20260 12928 20312 12980
rect 20812 12903 20864 12912
rect 20812 12869 20821 12903
rect 20821 12869 20855 12903
rect 20855 12869 20864 12903
rect 20812 12860 20864 12869
rect 20996 12860 21048 12912
rect 17868 12792 17920 12844
rect 17132 12724 17184 12776
rect 17776 12724 17828 12776
rect 18236 12767 18288 12776
rect 18236 12733 18245 12767
rect 18245 12733 18279 12767
rect 18279 12733 18288 12767
rect 18236 12724 18288 12733
rect 16396 12656 16448 12708
rect 19340 12792 19392 12844
rect 20260 12792 20312 12844
rect 19892 12767 19944 12776
rect 19892 12733 19901 12767
rect 19901 12733 19935 12767
rect 19935 12733 19944 12767
rect 19892 12724 19944 12733
rect 19616 12656 19668 12708
rect 17316 12588 17368 12640
rect 17776 12588 17828 12640
rect 20352 12724 20404 12776
rect 20444 12724 20496 12776
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 4436 12384 4488 12436
rect 5172 12384 5224 12436
rect 7288 12384 7340 12436
rect 4068 12316 4120 12368
rect 5908 12316 5960 12368
rect 6644 12316 6696 12368
rect 4712 12248 4764 12300
rect 5264 12291 5316 12300
rect 5264 12257 5273 12291
rect 5273 12257 5307 12291
rect 5307 12257 5316 12291
rect 5264 12248 5316 12257
rect 5632 12248 5684 12300
rect 6000 12248 6052 12300
rect 7196 12248 7248 12300
rect 12348 12384 12400 12436
rect 13084 12384 13136 12436
rect 13820 12384 13872 12436
rect 16304 12384 16356 12436
rect 16948 12384 17000 12436
rect 17684 12384 17736 12436
rect 20996 12384 21048 12436
rect 7748 12316 7800 12368
rect 8852 12316 8904 12368
rect 1584 12155 1636 12164
rect 1584 12121 1593 12155
rect 1593 12121 1627 12155
rect 1627 12121 1636 12155
rect 1584 12112 1636 12121
rect 1768 12155 1820 12164
rect 1768 12121 1777 12155
rect 1777 12121 1811 12155
rect 1811 12121 1820 12155
rect 1768 12112 1820 12121
rect 2320 12112 2372 12164
rect 4344 12180 4396 12232
rect 5724 12180 5776 12232
rect 7656 12180 7708 12232
rect 9220 12316 9272 12368
rect 7840 12180 7892 12232
rect 9404 12248 9456 12300
rect 9772 12248 9824 12300
rect 10140 12291 10192 12300
rect 10140 12257 10149 12291
rect 10149 12257 10183 12291
rect 10183 12257 10192 12291
rect 10140 12248 10192 12257
rect 14372 12316 14424 12368
rect 14832 12316 14884 12368
rect 8484 12180 8536 12232
rect 14280 12180 14332 12232
rect 14924 12180 14976 12232
rect 17868 12223 17920 12232
rect 17868 12189 17877 12223
rect 17877 12189 17911 12223
rect 17911 12189 17920 12223
rect 17868 12180 17920 12189
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 4528 12112 4580 12164
rect 10140 12112 10192 12164
rect 11796 12112 11848 12164
rect 18236 12248 18288 12300
rect 19524 12248 19576 12300
rect 20536 12316 20588 12368
rect 20444 12248 20496 12300
rect 20628 12223 20680 12232
rect 3424 12044 3476 12096
rect 4620 12044 4672 12096
rect 4988 12044 5040 12096
rect 5816 12044 5868 12096
rect 6920 12044 6972 12096
rect 7288 12044 7340 12096
rect 8760 12044 8812 12096
rect 8944 12044 8996 12096
rect 9772 12044 9824 12096
rect 12164 12044 12216 12096
rect 18420 12112 18472 12164
rect 20628 12189 20637 12223
rect 20637 12189 20671 12223
rect 20671 12189 20680 12223
rect 20628 12180 20680 12189
rect 14188 12044 14240 12096
rect 14464 12044 14516 12096
rect 14740 12044 14792 12096
rect 17224 12044 17276 12096
rect 17408 12044 17460 12096
rect 20536 12112 20588 12164
rect 19984 12044 20036 12096
rect 21272 12087 21324 12096
rect 21272 12053 21281 12087
rect 21281 12053 21315 12087
rect 21315 12053 21324 12087
rect 21272 12044 21324 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 3056 11883 3108 11892
rect 3056 11849 3065 11883
rect 3065 11849 3099 11883
rect 3099 11849 3108 11883
rect 3056 11840 3108 11849
rect 4252 11840 4304 11892
rect 5172 11840 5224 11892
rect 5632 11883 5684 11892
rect 5632 11849 5641 11883
rect 5641 11849 5675 11883
rect 5675 11849 5684 11883
rect 5632 11840 5684 11849
rect 6644 11840 6696 11892
rect 6736 11840 6788 11892
rect 7932 11840 7984 11892
rect 8116 11840 8168 11892
rect 8668 11840 8720 11892
rect 9680 11840 9732 11892
rect 1584 11704 1636 11756
rect 2688 11747 2740 11756
rect 2688 11713 2697 11747
rect 2697 11713 2731 11747
rect 2731 11713 2740 11747
rect 2688 11704 2740 11713
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 4344 11704 4396 11756
rect 4988 11704 5040 11756
rect 7012 11704 7064 11756
rect 2044 11636 2096 11688
rect 2504 11636 2556 11688
rect 5816 11636 5868 11688
rect 6920 11679 6972 11688
rect 6920 11645 6929 11679
rect 6929 11645 6963 11679
rect 6963 11645 6972 11679
rect 6920 11636 6972 11645
rect 7104 11636 7156 11688
rect 7840 11636 7892 11688
rect 8116 11568 8168 11620
rect 8760 11772 8812 11824
rect 11980 11840 12032 11892
rect 14464 11883 14516 11892
rect 9772 11704 9824 11756
rect 8576 11636 8628 11688
rect 9036 11636 9088 11688
rect 11796 11772 11848 11824
rect 14464 11849 14473 11883
rect 14473 11849 14507 11883
rect 14507 11849 14516 11883
rect 14464 11840 14516 11849
rect 17316 11883 17368 11892
rect 17316 11849 17325 11883
rect 17325 11849 17359 11883
rect 17359 11849 17368 11883
rect 17316 11840 17368 11849
rect 17408 11883 17460 11892
rect 17408 11849 17417 11883
rect 17417 11849 17451 11883
rect 17451 11849 17460 11883
rect 17408 11840 17460 11849
rect 17592 11840 17644 11892
rect 19984 11840 20036 11892
rect 20904 11840 20956 11892
rect 21180 11840 21232 11892
rect 14188 11772 14240 11824
rect 10416 11747 10468 11756
rect 10416 11713 10425 11747
rect 10425 11713 10459 11747
rect 10459 11713 10468 11747
rect 10416 11704 10468 11713
rect 10508 11636 10560 11688
rect 12164 11679 12216 11688
rect 12164 11645 12173 11679
rect 12173 11645 12207 11679
rect 12207 11645 12216 11679
rect 12164 11636 12216 11645
rect 12532 11636 12584 11688
rect 13084 11679 13136 11688
rect 13084 11645 13093 11679
rect 13093 11645 13127 11679
rect 13127 11645 13136 11679
rect 13084 11636 13136 11645
rect 9864 11568 9916 11620
rect 14372 11636 14424 11688
rect 14740 11679 14792 11688
rect 14740 11645 14749 11679
rect 14749 11645 14783 11679
rect 14783 11645 14792 11679
rect 14740 11636 14792 11645
rect 20260 11815 20312 11824
rect 20260 11781 20269 11815
rect 20269 11781 20303 11815
rect 20303 11781 20312 11815
rect 20260 11772 20312 11781
rect 18604 11747 18656 11756
rect 18604 11713 18613 11747
rect 18613 11713 18647 11747
rect 18647 11713 18656 11747
rect 18604 11704 18656 11713
rect 19064 11747 19116 11756
rect 19064 11713 19073 11747
rect 19073 11713 19107 11747
rect 19107 11713 19116 11747
rect 19064 11704 19116 11713
rect 17224 11636 17276 11688
rect 17776 11636 17828 11688
rect 20628 11636 20680 11688
rect 20076 11568 20128 11620
rect 5908 11500 5960 11552
rect 7932 11500 7984 11552
rect 8024 11500 8076 11552
rect 11244 11500 11296 11552
rect 13636 11500 13688 11552
rect 16396 11500 16448 11552
rect 18052 11500 18104 11552
rect 18328 11500 18380 11552
rect 19524 11500 19576 11552
rect 20260 11500 20312 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 1676 11339 1728 11348
rect 1676 11305 1685 11339
rect 1685 11305 1719 11339
rect 1719 11305 1728 11339
rect 1676 11296 1728 11305
rect 2504 11339 2556 11348
rect 2504 11305 2513 11339
rect 2513 11305 2547 11339
rect 2547 11305 2556 11339
rect 2504 11296 2556 11305
rect 9496 11296 9548 11348
rect 9772 11339 9824 11348
rect 9772 11305 9781 11339
rect 9781 11305 9815 11339
rect 9815 11305 9824 11339
rect 9772 11296 9824 11305
rect 10140 11296 10192 11348
rect 11060 11339 11112 11348
rect 11060 11305 11069 11339
rect 11069 11305 11103 11339
rect 11103 11305 11112 11339
rect 11060 11296 11112 11305
rect 12992 11296 13044 11348
rect 13636 11296 13688 11348
rect 20628 11339 20680 11348
rect 3884 11228 3936 11280
rect 1492 11135 1544 11144
rect 1492 11101 1501 11135
rect 1501 11101 1535 11135
rect 1535 11101 1544 11135
rect 1492 11092 1544 11101
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 2964 11160 3016 11212
rect 3424 11160 3476 11212
rect 3792 11092 3844 11144
rect 4988 11092 5040 11144
rect 6000 11160 6052 11212
rect 11796 11228 11848 11280
rect 14740 11228 14792 11280
rect 17132 11228 17184 11280
rect 17776 11228 17828 11280
rect 8484 11203 8536 11212
rect 8484 11169 8493 11203
rect 8493 11169 8527 11203
rect 8527 11169 8536 11203
rect 8484 11160 8536 11169
rect 9220 11203 9272 11212
rect 9220 11169 9229 11203
rect 9229 11169 9263 11203
rect 9263 11169 9272 11203
rect 9220 11160 9272 11169
rect 9864 11160 9916 11212
rect 10048 11160 10100 11212
rect 17868 11160 17920 11212
rect 18236 11203 18288 11212
rect 18236 11169 18245 11203
rect 18245 11169 18279 11203
rect 18279 11169 18288 11203
rect 18236 11160 18288 11169
rect 2136 11024 2188 11076
rect 5264 10999 5316 11008
rect 5264 10965 5273 10999
rect 5273 10965 5307 10999
rect 5307 10965 5316 10999
rect 5264 10956 5316 10965
rect 5540 10956 5592 11008
rect 5908 10956 5960 11008
rect 6736 11024 6788 11076
rect 6644 10956 6696 11008
rect 7104 11092 7156 11144
rect 9404 11135 9456 11144
rect 7288 11024 7340 11076
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 15752 11092 15804 11144
rect 17040 11092 17092 11144
rect 19524 11135 19576 11144
rect 19524 11101 19558 11135
rect 19558 11101 19576 11135
rect 9864 11024 9916 11076
rect 11152 10956 11204 11008
rect 11980 11024 12032 11076
rect 13544 11067 13596 11076
rect 13544 11033 13553 11067
rect 13553 11033 13587 11067
rect 13587 11033 13596 11067
rect 13544 11024 13596 11033
rect 14372 11024 14424 11076
rect 15108 11024 15160 11076
rect 15936 11024 15988 11076
rect 19524 11092 19576 11101
rect 20628 11305 20637 11339
rect 20637 11305 20671 11339
rect 20671 11305 20680 11339
rect 20628 11296 20680 11305
rect 21180 11339 21232 11348
rect 21180 11305 21189 11339
rect 21189 11305 21223 11339
rect 21223 11305 21232 11339
rect 21180 11296 21232 11305
rect 21364 11092 21416 11144
rect 11704 10956 11756 11008
rect 12900 10956 12952 11008
rect 13820 10956 13872 11008
rect 16396 10956 16448 11008
rect 16948 10999 17000 11008
rect 16948 10965 16957 10999
rect 16957 10965 16991 10999
rect 16991 10965 17000 10999
rect 16948 10956 17000 10965
rect 17684 10999 17736 11008
rect 17684 10965 17693 10999
rect 17693 10965 17727 10999
rect 17727 10965 17736 10999
rect 17684 10956 17736 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 1584 10752 1636 10804
rect 2688 10752 2740 10804
rect 3056 10752 3108 10804
rect 3608 10752 3660 10804
rect 3792 10795 3844 10804
rect 3792 10761 3801 10795
rect 3801 10761 3835 10795
rect 3835 10761 3844 10795
rect 3792 10752 3844 10761
rect 4712 10752 4764 10804
rect 5908 10752 5960 10804
rect 6736 10795 6788 10804
rect 6736 10761 6745 10795
rect 6745 10761 6779 10795
rect 6779 10761 6788 10795
rect 6736 10752 6788 10761
rect 6920 10752 6972 10804
rect 7472 10752 7524 10804
rect 7656 10752 7708 10804
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 4436 10684 4488 10736
rect 8576 10752 8628 10804
rect 11704 10752 11756 10804
rect 11980 10752 12032 10804
rect 17684 10752 17736 10804
rect 18788 10752 18840 10804
rect 18972 10752 19024 10804
rect 10140 10684 10192 10736
rect 1676 10616 1728 10625
rect 3332 10616 3384 10668
rect 5080 10616 5132 10668
rect 6000 10616 6052 10668
rect 9772 10616 9824 10668
rect 3424 10548 3476 10600
rect 5172 10591 5224 10600
rect 5172 10557 5181 10591
rect 5181 10557 5215 10591
rect 5215 10557 5224 10591
rect 5172 10548 5224 10557
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 7380 10548 7432 10600
rect 9404 10548 9456 10600
rect 10324 10548 10376 10600
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 2504 10480 2556 10532
rect 2228 10412 2280 10464
rect 7472 10480 7524 10532
rect 8484 10480 8536 10532
rect 11152 10548 11204 10600
rect 12072 10684 12124 10736
rect 12716 10684 12768 10736
rect 18236 10684 18288 10736
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 15292 10616 15344 10668
rect 12808 10523 12860 10532
rect 12808 10489 12817 10523
rect 12817 10489 12851 10523
rect 12851 10489 12860 10523
rect 12808 10480 12860 10489
rect 14280 10480 14332 10532
rect 16304 10616 16356 10668
rect 19524 10684 19576 10736
rect 21272 10684 21324 10736
rect 15660 10591 15712 10600
rect 15660 10557 15669 10591
rect 15669 10557 15703 10591
rect 15703 10557 15712 10591
rect 15660 10548 15712 10557
rect 17132 10591 17184 10600
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17040 10480 17092 10532
rect 17684 10591 17736 10600
rect 5908 10455 5960 10464
rect 5908 10421 5917 10455
rect 5917 10421 5951 10455
rect 5951 10421 5960 10455
rect 5908 10412 5960 10421
rect 9220 10412 9272 10464
rect 11060 10412 11112 10464
rect 13820 10412 13872 10464
rect 14372 10455 14424 10464
rect 14372 10421 14381 10455
rect 14381 10421 14415 10455
rect 14415 10421 14424 10455
rect 14372 10412 14424 10421
rect 15844 10412 15896 10464
rect 16948 10412 17000 10464
rect 17684 10557 17693 10591
rect 17693 10557 17727 10591
rect 17727 10557 17736 10591
rect 17684 10548 17736 10557
rect 20352 10548 20404 10600
rect 21364 10591 21416 10600
rect 21364 10557 21373 10591
rect 21373 10557 21407 10591
rect 21407 10557 21416 10591
rect 21364 10548 21416 10557
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 19892 10412 19944 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1492 10208 1544 10260
rect 1952 10140 2004 10192
rect 4712 10208 4764 10260
rect 5080 10208 5132 10260
rect 5264 10208 5316 10260
rect 6644 10208 6696 10260
rect 4344 10140 4396 10192
rect 8668 10208 8720 10260
rect 9220 10208 9272 10260
rect 9772 10251 9824 10260
rect 8116 10140 8168 10192
rect 9772 10217 9781 10251
rect 9781 10217 9815 10251
rect 9815 10217 9824 10251
rect 9772 10208 9824 10217
rect 11428 10251 11480 10260
rect 11428 10217 11437 10251
rect 11437 10217 11471 10251
rect 11471 10217 11480 10251
rect 11428 10208 11480 10217
rect 14280 10208 14332 10260
rect 1860 10115 1912 10124
rect 1860 10081 1869 10115
rect 1869 10081 1903 10115
rect 1903 10081 1912 10115
rect 1860 10072 1912 10081
rect 3884 10072 3936 10124
rect 5264 10072 5316 10124
rect 6000 10115 6052 10124
rect 6000 10081 6009 10115
rect 6009 10081 6043 10115
rect 6043 10081 6052 10115
rect 6000 10072 6052 10081
rect 6644 10072 6696 10124
rect 7288 10072 7340 10124
rect 12072 10140 12124 10192
rect 17132 10208 17184 10260
rect 17960 10208 18012 10260
rect 19064 10208 19116 10260
rect 19524 10251 19576 10260
rect 19524 10217 19533 10251
rect 19533 10217 19567 10251
rect 19567 10217 19576 10251
rect 19524 10208 19576 10217
rect 1676 9979 1728 9988
rect 1676 9945 1685 9979
rect 1685 9945 1719 9979
rect 1719 9945 1728 9979
rect 1676 9936 1728 9945
rect 2780 9936 2832 9988
rect 3424 10004 3476 10056
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 5540 10004 5592 10056
rect 3516 9936 3568 9988
rect 5356 9936 5408 9988
rect 4068 9868 4120 9920
rect 4436 9911 4488 9920
rect 4436 9877 4445 9911
rect 4445 9877 4479 9911
rect 4479 9877 4488 9911
rect 4436 9868 4488 9877
rect 6736 9868 6788 9920
rect 6828 9911 6880 9920
rect 6828 9877 6837 9911
rect 6837 9877 6871 9911
rect 6871 9877 6880 9911
rect 8024 9936 8076 9988
rect 8944 9936 8996 9988
rect 9588 10072 9640 10124
rect 9772 10072 9824 10124
rect 18604 10140 18656 10192
rect 19432 10140 19484 10192
rect 19892 10140 19944 10192
rect 16304 10115 16356 10124
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 10140 10004 10192 10056
rect 11704 10004 11756 10056
rect 9588 9936 9640 9988
rect 11152 9936 11204 9988
rect 13636 10004 13688 10056
rect 13728 10004 13780 10056
rect 16304 10081 16313 10115
rect 16313 10081 16347 10115
rect 16347 10081 16356 10115
rect 16304 10072 16356 10081
rect 16396 10072 16448 10124
rect 18236 10072 18288 10124
rect 20536 10115 20588 10124
rect 20536 10081 20545 10115
rect 20545 10081 20579 10115
rect 20579 10081 20588 10115
rect 20536 10072 20588 10081
rect 20996 10072 21048 10124
rect 17684 10004 17736 10056
rect 18972 10004 19024 10056
rect 20352 10047 20404 10056
rect 20352 10013 20361 10047
rect 20361 10013 20395 10047
rect 20395 10013 20404 10047
rect 20352 10004 20404 10013
rect 20720 10004 20772 10056
rect 6828 9868 6880 9877
rect 7840 9911 7892 9920
rect 7840 9877 7849 9911
rect 7849 9877 7883 9911
rect 7883 9877 7892 9911
rect 7840 9868 7892 9877
rect 7932 9911 7984 9920
rect 7932 9877 7941 9911
rect 7941 9877 7975 9911
rect 7975 9877 7984 9911
rect 7932 9868 7984 9877
rect 8392 9868 8444 9920
rect 14096 9911 14148 9920
rect 14096 9877 14105 9911
rect 14105 9877 14139 9911
rect 14139 9877 14148 9911
rect 14096 9868 14148 9877
rect 14280 9936 14332 9988
rect 15844 9936 15896 9988
rect 16856 9936 16908 9988
rect 17592 9936 17644 9988
rect 18144 9979 18196 9988
rect 18144 9945 18153 9979
rect 18153 9945 18187 9979
rect 18187 9945 18196 9979
rect 18144 9936 18196 9945
rect 19156 9936 19208 9988
rect 15384 9868 15436 9920
rect 16120 9911 16172 9920
rect 16120 9877 16129 9911
rect 16129 9877 16163 9911
rect 16163 9877 16172 9911
rect 16120 9868 16172 9877
rect 17776 9868 17828 9920
rect 19708 9868 19760 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 1584 9571 1636 9580
rect 1584 9537 1593 9571
rect 1593 9537 1627 9571
rect 1627 9537 1636 9571
rect 2872 9664 2924 9716
rect 2228 9596 2280 9648
rect 3056 9664 3108 9716
rect 3332 9664 3384 9716
rect 6828 9664 6880 9716
rect 8944 9707 8996 9716
rect 1584 9528 1636 9537
rect 4436 9596 4488 9648
rect 6920 9596 6972 9648
rect 8944 9673 8953 9707
rect 8953 9673 8987 9707
rect 8987 9673 8996 9707
rect 8944 9664 8996 9673
rect 10600 9664 10652 9716
rect 10876 9664 10928 9716
rect 14280 9664 14332 9716
rect 14372 9664 14424 9716
rect 15660 9664 15712 9716
rect 15844 9707 15896 9716
rect 15844 9673 15853 9707
rect 15853 9673 15887 9707
rect 15887 9673 15896 9707
rect 15844 9664 15896 9673
rect 2596 9528 2648 9580
rect 2688 9528 2740 9580
rect 4620 9528 4672 9580
rect 5080 9528 5132 9580
rect 5908 9528 5960 9580
rect 7012 9528 7064 9580
rect 7564 9528 7616 9580
rect 10232 9528 10284 9580
rect 10600 9528 10652 9580
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 11980 9571 12032 9580
rect 11980 9537 12014 9571
rect 12014 9537 12032 9571
rect 11980 9528 12032 9537
rect 13728 9528 13780 9580
rect 15384 9596 15436 9648
rect 17684 9596 17736 9648
rect 18236 9664 18288 9716
rect 18788 9664 18840 9716
rect 19156 9664 19208 9716
rect 20260 9596 20312 9648
rect 16120 9528 16172 9580
rect 16764 9571 16816 9580
rect 16764 9537 16773 9571
rect 16773 9537 16807 9571
rect 16807 9537 16816 9571
rect 16764 9528 16816 9537
rect 18512 9528 18564 9580
rect 18604 9571 18656 9580
rect 18604 9537 18613 9571
rect 18613 9537 18647 9571
rect 18647 9537 18656 9571
rect 18604 9528 18656 9537
rect 4988 9460 5040 9512
rect 7380 9503 7432 9512
rect 7380 9469 7389 9503
rect 7389 9469 7423 9503
rect 7423 9469 7432 9503
rect 7380 9460 7432 9469
rect 10324 9503 10376 9512
rect 6552 9435 6604 9444
rect 6552 9401 6561 9435
rect 6561 9401 6595 9435
rect 6595 9401 6604 9435
rect 6552 9392 6604 9401
rect 6736 9392 6788 9444
rect 3240 9324 3292 9376
rect 3424 9367 3476 9376
rect 3424 9333 3433 9367
rect 3433 9333 3467 9367
rect 3467 9333 3476 9367
rect 3424 9324 3476 9333
rect 5356 9367 5408 9376
rect 5356 9333 5365 9367
rect 5365 9333 5399 9367
rect 5399 9333 5408 9367
rect 5356 9324 5408 9333
rect 6644 9324 6696 9376
rect 10324 9469 10333 9503
rect 10333 9469 10367 9503
rect 10367 9469 10376 9503
rect 10324 9460 10376 9469
rect 11152 9460 11204 9512
rect 14096 9460 14148 9512
rect 14280 9460 14332 9512
rect 16396 9460 16448 9512
rect 17776 9460 17828 9512
rect 19524 9528 19576 9580
rect 19800 9528 19852 9580
rect 20536 9528 20588 9580
rect 21364 9503 21416 9512
rect 13360 9392 13412 9444
rect 14648 9392 14700 9444
rect 15292 9392 15344 9444
rect 18052 9392 18104 9444
rect 19432 9392 19484 9444
rect 13084 9367 13136 9376
rect 13084 9333 13093 9367
rect 13093 9333 13127 9367
rect 13127 9333 13136 9367
rect 13084 9324 13136 9333
rect 13728 9324 13780 9376
rect 15476 9324 15528 9376
rect 15936 9324 15988 9376
rect 17960 9324 18012 9376
rect 19800 9324 19852 9376
rect 19984 9367 20036 9376
rect 19984 9333 19993 9367
rect 19993 9333 20027 9367
rect 20027 9333 20036 9367
rect 19984 9324 20036 9333
rect 21364 9469 21373 9503
rect 21373 9469 21407 9503
rect 21407 9469 21416 9503
rect 21364 9460 21416 9469
rect 20444 9324 20496 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 4712 9120 4764 9172
rect 6644 9163 6696 9172
rect 6644 9129 6653 9163
rect 6653 9129 6687 9163
rect 6687 9129 6696 9163
rect 6644 9120 6696 9129
rect 7840 9120 7892 9172
rect 10692 9120 10744 9172
rect 11152 9163 11204 9172
rect 11152 9129 11161 9163
rect 11161 9129 11195 9163
rect 11195 9129 11204 9163
rect 11152 9120 11204 9129
rect 11980 9120 12032 9172
rect 15936 9120 15988 9172
rect 2044 9052 2096 9104
rect 4988 9052 5040 9104
rect 6552 9052 6604 9104
rect 10600 9052 10652 9104
rect 12900 9052 12952 9104
rect 3424 8984 3476 9036
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 4712 9027 4764 9036
rect 4712 8993 4721 9027
rect 4721 8993 4755 9027
rect 4755 8993 4764 9027
rect 4712 8984 4764 8993
rect 3148 8916 3200 8968
rect 4620 8916 4672 8968
rect 5172 8916 5224 8968
rect 5356 8916 5408 8968
rect 9588 8984 9640 9036
rect 7104 8916 7156 8968
rect 7564 8916 7616 8968
rect 1676 8891 1728 8900
rect 1676 8857 1685 8891
rect 1685 8857 1719 8891
rect 1719 8857 1728 8891
rect 1676 8848 1728 8857
rect 1860 8891 1912 8900
rect 1860 8857 1869 8891
rect 1869 8857 1903 8891
rect 1903 8857 1912 8891
rect 1860 8848 1912 8857
rect 2596 8891 2648 8900
rect 2596 8857 2605 8891
rect 2605 8857 2639 8891
rect 2639 8857 2648 8891
rect 2596 8848 2648 8857
rect 3240 8848 3292 8900
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 11244 8916 11296 8968
rect 12440 8984 12492 9036
rect 13636 8984 13688 9036
rect 12992 8916 13044 8968
rect 13452 8916 13504 8968
rect 14280 8916 14332 8968
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 16764 8916 16816 8968
rect 18512 9120 18564 9172
rect 18880 9052 18932 9104
rect 17500 8984 17552 9036
rect 19800 9027 19852 9036
rect 19800 8993 19809 9027
rect 19809 8993 19843 9027
rect 19843 8993 19852 9027
rect 19800 8984 19852 8993
rect 19984 9027 20036 9036
rect 19984 8993 19993 9027
rect 19993 8993 20027 9027
rect 20027 8993 20036 9027
rect 19984 8984 20036 8993
rect 20536 8984 20588 9036
rect 17592 8916 17644 8968
rect 19708 8959 19760 8968
rect 19708 8925 19717 8959
rect 19717 8925 19751 8959
rect 19751 8925 19760 8959
rect 19708 8916 19760 8925
rect 2688 8823 2740 8832
rect 2688 8789 2697 8823
rect 2697 8789 2731 8823
rect 2731 8789 2740 8823
rect 2688 8780 2740 8789
rect 2780 8780 2832 8832
rect 2964 8780 3016 8832
rect 3148 8780 3200 8832
rect 3792 8780 3844 8832
rect 3976 8780 4028 8832
rect 5724 8780 5776 8832
rect 6828 8780 6880 8832
rect 6920 8780 6972 8832
rect 8116 8780 8168 8832
rect 8576 8780 8628 8832
rect 9404 8823 9456 8832
rect 9404 8789 9413 8823
rect 9413 8789 9447 8823
rect 9447 8789 9456 8823
rect 16396 8848 16448 8900
rect 17776 8848 17828 8900
rect 18788 8891 18840 8900
rect 18788 8857 18797 8891
rect 18797 8857 18831 8891
rect 18831 8857 18840 8891
rect 18788 8848 18840 8857
rect 18880 8848 18932 8900
rect 9404 8780 9456 8789
rect 12164 8780 12216 8832
rect 12716 8823 12768 8832
rect 12716 8789 12725 8823
rect 12725 8789 12759 8823
rect 12759 8789 12768 8823
rect 12716 8780 12768 8789
rect 13452 8780 13504 8832
rect 13636 8823 13688 8832
rect 13636 8789 13645 8823
rect 13645 8789 13679 8823
rect 13679 8789 13688 8823
rect 13636 8780 13688 8789
rect 14832 8823 14884 8832
rect 14832 8789 14841 8823
rect 14841 8789 14875 8823
rect 14875 8789 14884 8823
rect 14832 8780 14884 8789
rect 15292 8823 15344 8832
rect 15292 8789 15301 8823
rect 15301 8789 15335 8823
rect 15335 8789 15344 8823
rect 15292 8780 15344 8789
rect 17592 8780 17644 8832
rect 20904 8780 20956 8832
rect 21456 8780 21508 8832
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 2504 8576 2556 8628
rect 2596 8576 2648 8628
rect 3976 8619 4028 8628
rect 3976 8585 3985 8619
rect 3985 8585 4019 8619
rect 4019 8585 4028 8619
rect 3976 8576 4028 8585
rect 4068 8576 4120 8628
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 1952 8440 2004 8492
rect 3240 8440 3292 8492
rect 3792 8508 3844 8560
rect 4896 8576 4948 8628
rect 7104 8576 7156 8628
rect 7932 8576 7984 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 10048 8576 10100 8628
rect 6920 8508 6972 8560
rect 9680 8508 9732 8560
rect 3424 8372 3476 8424
rect 4068 8415 4120 8424
rect 3056 8236 3108 8288
rect 3332 8236 3384 8288
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4436 8372 4488 8424
rect 4896 8440 4948 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 6644 8440 6696 8492
rect 7472 8440 7524 8492
rect 4252 8304 4304 8356
rect 4896 8304 4948 8356
rect 5356 8304 5408 8356
rect 8116 8440 8168 8492
rect 18512 8576 18564 8628
rect 10048 8440 10100 8492
rect 9588 8415 9640 8424
rect 8668 8304 8720 8356
rect 9588 8381 9597 8415
rect 9597 8381 9631 8415
rect 9631 8381 9640 8415
rect 9588 8372 9640 8381
rect 10876 8372 10928 8424
rect 14832 8508 14884 8560
rect 17132 8508 17184 8560
rect 17684 8508 17736 8560
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 13544 8483 13596 8492
rect 12532 8440 12584 8449
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 13636 8483 13688 8492
rect 13636 8449 13645 8483
rect 13645 8449 13679 8483
rect 13679 8449 13688 8483
rect 14372 8483 14424 8492
rect 13636 8440 13688 8449
rect 11888 8415 11940 8424
rect 11888 8381 11897 8415
rect 11897 8381 11931 8415
rect 11931 8381 11940 8415
rect 11888 8372 11940 8381
rect 12256 8415 12308 8424
rect 12256 8381 12265 8415
rect 12265 8381 12299 8415
rect 12299 8381 12308 8415
rect 12256 8372 12308 8381
rect 12440 8415 12492 8424
rect 12440 8381 12449 8415
rect 12449 8381 12483 8415
rect 12483 8381 12492 8415
rect 12440 8372 12492 8381
rect 13728 8415 13780 8424
rect 13728 8381 13737 8415
rect 13737 8381 13771 8415
rect 13771 8381 13780 8415
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 16120 8483 16172 8492
rect 16120 8449 16129 8483
rect 16129 8449 16163 8483
rect 16163 8449 16172 8483
rect 16120 8440 16172 8449
rect 16396 8440 16448 8492
rect 17224 8440 17276 8492
rect 18696 8440 18748 8492
rect 20812 8508 20864 8560
rect 21364 8508 21416 8560
rect 20536 8483 20588 8492
rect 13728 8372 13780 8381
rect 12808 8304 12860 8356
rect 4620 8236 4672 8288
rect 8392 8236 8444 8288
rect 10876 8236 10928 8288
rect 13544 8304 13596 8356
rect 15844 8304 15896 8356
rect 16028 8304 16080 8356
rect 13176 8279 13228 8288
rect 13176 8245 13185 8279
rect 13185 8245 13219 8279
rect 13219 8245 13228 8279
rect 13176 8236 13228 8245
rect 17776 8304 17828 8356
rect 17960 8372 18012 8424
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 17132 8236 17184 8288
rect 17868 8236 17920 8288
rect 17960 8236 18012 8288
rect 20260 8279 20312 8288
rect 20260 8245 20269 8279
rect 20269 8245 20303 8279
rect 20303 8245 20312 8279
rect 20260 8236 20312 8245
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 2688 8032 2740 8084
rect 2504 7896 2556 7948
rect 3424 7896 3476 7948
rect 1952 7871 2004 7880
rect 1952 7837 1961 7871
rect 1961 7837 1995 7871
rect 1995 7837 2004 7871
rect 1952 7828 2004 7837
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 2412 7828 2464 7880
rect 2504 7692 2556 7744
rect 3332 7828 3384 7880
rect 4160 7964 4212 8016
rect 4528 7964 4580 8016
rect 4712 7896 4764 7948
rect 5632 7896 5684 7948
rect 7656 8032 7708 8084
rect 8116 8032 8168 8084
rect 12256 8032 12308 8084
rect 12440 8032 12492 8084
rect 7932 7964 7984 8016
rect 8484 7964 8536 8016
rect 12716 7964 12768 8016
rect 4436 7828 4488 7880
rect 13176 7896 13228 7948
rect 13452 7939 13504 7948
rect 13452 7905 13461 7939
rect 13461 7905 13495 7939
rect 13495 7905 13504 7939
rect 13452 7896 13504 7905
rect 7748 7871 7800 7880
rect 7748 7837 7757 7871
rect 7757 7837 7791 7871
rect 7791 7837 7800 7871
rect 7748 7828 7800 7837
rect 8392 7828 8444 7880
rect 9496 7828 9548 7880
rect 10324 7828 10376 7880
rect 14372 7828 14424 7880
rect 4620 7760 4672 7812
rect 5908 7760 5960 7812
rect 8300 7760 8352 7812
rect 8484 7760 8536 7812
rect 11244 7760 11296 7812
rect 11704 7760 11756 7812
rect 13452 7760 13504 7812
rect 20628 8032 20680 8084
rect 17684 7896 17736 7948
rect 17776 7896 17828 7948
rect 18880 7964 18932 8016
rect 18696 7939 18748 7948
rect 18696 7905 18705 7939
rect 18705 7905 18739 7939
rect 18739 7905 18748 7939
rect 18696 7896 18748 7905
rect 20260 7939 20312 7948
rect 20260 7905 20269 7939
rect 20269 7905 20303 7939
rect 20303 7905 20312 7939
rect 20260 7896 20312 7905
rect 15476 7828 15528 7880
rect 15568 7828 15620 7880
rect 17868 7828 17920 7880
rect 18788 7828 18840 7880
rect 19064 7828 19116 7880
rect 4436 7692 4488 7744
rect 4804 7735 4856 7744
rect 4804 7701 4813 7735
rect 4813 7701 4847 7735
rect 4847 7701 4856 7735
rect 4804 7692 4856 7701
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 10968 7735 11020 7744
rect 10968 7701 10977 7735
rect 10977 7701 11011 7735
rect 11011 7701 11020 7735
rect 10968 7692 11020 7701
rect 13268 7735 13320 7744
rect 13268 7701 13277 7735
rect 13277 7701 13311 7735
rect 13311 7701 13320 7735
rect 13268 7692 13320 7701
rect 14556 7692 14608 7744
rect 17776 7760 17828 7812
rect 20076 7828 20128 7880
rect 19064 7692 19116 7744
rect 19708 7735 19760 7744
rect 19708 7701 19717 7735
rect 19717 7701 19751 7735
rect 19751 7701 19760 7735
rect 19708 7692 19760 7701
rect 19800 7692 19852 7744
rect 21364 7735 21416 7744
rect 21364 7701 21373 7735
rect 21373 7701 21407 7735
rect 21407 7701 21416 7735
rect 21364 7692 21416 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 2504 7531 2556 7540
rect 2504 7497 2513 7531
rect 2513 7497 2547 7531
rect 2547 7497 2556 7531
rect 2504 7488 2556 7497
rect 2872 7531 2924 7540
rect 2872 7497 2881 7531
rect 2881 7497 2915 7531
rect 2915 7497 2924 7531
rect 2872 7488 2924 7497
rect 4344 7488 4396 7540
rect 4804 7488 4856 7540
rect 7196 7488 7248 7540
rect 9680 7488 9732 7540
rect 10232 7488 10284 7540
rect 11888 7531 11940 7540
rect 11888 7497 11897 7531
rect 11897 7497 11931 7531
rect 11931 7497 11940 7531
rect 11888 7488 11940 7497
rect 12532 7488 12584 7540
rect 1860 7463 1912 7472
rect 1860 7429 1869 7463
rect 1869 7429 1903 7463
rect 1903 7429 1912 7463
rect 1860 7420 1912 7429
rect 2780 7420 2832 7472
rect 1400 7352 1452 7404
rect 1676 7395 1728 7404
rect 1676 7361 1685 7395
rect 1685 7361 1719 7395
rect 1719 7361 1728 7395
rect 1676 7352 1728 7361
rect 7472 7420 7524 7472
rect 8392 7420 8444 7472
rect 3424 7352 3476 7404
rect 3884 7352 3936 7404
rect 9772 7420 9824 7472
rect 12072 7420 12124 7472
rect 13268 7488 13320 7540
rect 13820 7420 13872 7472
rect 3240 7284 3292 7336
rect 4160 7284 4212 7336
rect 5172 7284 5224 7336
rect 5540 7327 5592 7336
rect 2412 7148 2464 7200
rect 2596 7148 2648 7200
rect 5540 7293 5549 7327
rect 5549 7293 5583 7327
rect 5583 7293 5592 7327
rect 5540 7284 5592 7293
rect 14372 7352 14424 7404
rect 16948 7488 17000 7540
rect 17960 7488 18012 7540
rect 18696 7488 18748 7540
rect 19524 7488 19576 7540
rect 21180 7531 21232 7540
rect 21180 7497 21189 7531
rect 21189 7497 21223 7531
rect 21223 7497 21232 7531
rect 21180 7488 21232 7497
rect 16580 7352 16632 7404
rect 17684 7420 17736 7472
rect 18604 7420 18656 7472
rect 16948 7395 17000 7404
rect 16948 7361 16982 7395
rect 16982 7361 17000 7395
rect 16948 7352 17000 7361
rect 19524 7352 19576 7404
rect 21364 7420 21416 7472
rect 5908 7284 5960 7336
rect 5908 7148 5960 7200
rect 7012 7148 7064 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 9128 7284 9180 7336
rect 8300 7148 8352 7200
rect 9772 7148 9824 7200
rect 13452 7216 13504 7268
rect 15016 7284 15068 7336
rect 16120 7284 16172 7336
rect 16396 7284 16448 7336
rect 14648 7148 14700 7200
rect 15200 7191 15252 7200
rect 15200 7157 15209 7191
rect 15209 7157 15243 7191
rect 15243 7157 15252 7191
rect 15200 7148 15252 7157
rect 15936 7148 15988 7200
rect 19800 7284 19852 7336
rect 20812 7327 20864 7336
rect 20812 7293 20821 7327
rect 20821 7293 20855 7327
rect 20855 7293 20864 7327
rect 20812 7284 20864 7293
rect 21180 7284 21232 7336
rect 19524 7148 19576 7200
rect 20812 7148 20864 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 2320 6851 2372 6860
rect 2320 6817 2329 6851
rect 2329 6817 2363 6851
rect 2363 6817 2372 6851
rect 2320 6808 2372 6817
rect 2412 6808 2464 6860
rect 3792 6808 3844 6860
rect 5356 6944 5408 6996
rect 10692 6944 10744 6996
rect 13084 6944 13136 6996
rect 5632 6876 5684 6928
rect 5724 6808 5776 6860
rect 7012 6851 7064 6860
rect 940 6740 992 6792
rect 3240 6783 3292 6792
rect 3240 6749 3249 6783
rect 3249 6749 3283 6783
rect 3283 6749 3292 6783
rect 3240 6740 3292 6749
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 4620 6783 4672 6792
rect 4620 6749 4629 6783
rect 4629 6749 4663 6783
rect 4663 6749 4672 6783
rect 4620 6740 4672 6749
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 15660 6944 15712 6996
rect 16948 6987 17000 6996
rect 16948 6953 16957 6987
rect 16957 6953 16991 6987
rect 16991 6953 17000 6987
rect 16948 6944 17000 6953
rect 17776 6944 17828 6996
rect 17868 6944 17920 6996
rect 11244 6808 11296 6860
rect 1860 6715 1912 6724
rect 1860 6681 1869 6715
rect 1869 6681 1903 6715
rect 1903 6681 1912 6715
rect 1860 6672 1912 6681
rect 2228 6672 2280 6724
rect 5172 6672 5224 6724
rect 5632 6672 5684 6724
rect 5816 6672 5868 6724
rect 7196 6783 7248 6792
rect 7196 6749 7205 6783
rect 7205 6749 7239 6783
rect 7239 6749 7248 6783
rect 7196 6740 7248 6749
rect 9680 6740 9732 6792
rect 10324 6783 10376 6792
rect 10324 6749 10333 6783
rect 10333 6749 10367 6783
rect 10367 6749 10376 6783
rect 10324 6740 10376 6749
rect 12256 6740 12308 6792
rect 12348 6740 12400 6792
rect 15016 6808 15068 6860
rect 15476 6876 15528 6928
rect 17960 6876 18012 6928
rect 18052 6919 18104 6928
rect 18052 6885 18061 6919
rect 18061 6885 18095 6919
rect 18095 6885 18104 6919
rect 18052 6876 18104 6885
rect 14372 6740 14424 6792
rect 15660 6740 15712 6792
rect 16304 6783 16356 6792
rect 16304 6749 16313 6783
rect 16313 6749 16347 6783
rect 16347 6749 16356 6783
rect 16304 6740 16356 6749
rect 16580 6740 16632 6792
rect 17040 6740 17092 6792
rect 17316 6740 17368 6792
rect 17868 6740 17920 6792
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18328 6740 18380 6792
rect 18972 6740 19024 6792
rect 17960 6672 18012 6724
rect 18604 6715 18656 6724
rect 18604 6681 18613 6715
rect 18613 6681 18647 6715
rect 18647 6681 18656 6715
rect 18604 6672 18656 6681
rect 19432 6715 19484 6724
rect 19432 6681 19441 6715
rect 19441 6681 19475 6715
rect 19475 6681 19484 6715
rect 19432 6672 19484 6681
rect 2412 6647 2464 6656
rect 2412 6613 2421 6647
rect 2421 6613 2455 6647
rect 2455 6613 2464 6647
rect 2412 6604 2464 6613
rect 3056 6604 3108 6656
rect 3976 6604 4028 6656
rect 4712 6604 4764 6656
rect 5356 6604 5408 6656
rect 5908 6604 5960 6656
rect 6736 6604 6788 6656
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 7380 6604 7432 6656
rect 7748 6604 7800 6656
rect 8208 6647 8260 6656
rect 8208 6613 8217 6647
rect 8217 6613 8251 6647
rect 8251 6613 8260 6647
rect 8208 6604 8260 6613
rect 8852 6604 8904 6656
rect 9312 6604 9364 6656
rect 10876 6604 10928 6656
rect 12992 6604 13044 6656
rect 13176 6604 13228 6656
rect 13728 6647 13780 6656
rect 13728 6613 13737 6647
rect 13737 6613 13771 6647
rect 13771 6613 13780 6647
rect 13728 6604 13780 6613
rect 14740 6647 14792 6656
rect 14740 6613 14749 6647
rect 14749 6613 14783 6647
rect 14783 6613 14792 6647
rect 14740 6604 14792 6613
rect 15752 6604 15804 6656
rect 17316 6604 17368 6656
rect 17500 6604 17552 6656
rect 17776 6604 17828 6656
rect 20076 6672 20128 6724
rect 20260 6740 20312 6792
rect 20536 6740 20588 6792
rect 20812 6740 20864 6792
rect 21272 6740 21324 6792
rect 21824 6672 21876 6724
rect 19984 6647 20036 6656
rect 19984 6613 19993 6647
rect 19993 6613 20027 6647
rect 20027 6613 20036 6647
rect 19984 6604 20036 6613
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 2044 6400 2096 6452
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 2412 6400 2464 6452
rect 2688 6400 2740 6452
rect 2596 6332 2648 6384
rect 2964 6375 3016 6384
rect 2964 6341 2973 6375
rect 2973 6341 3007 6375
rect 3007 6341 3016 6375
rect 2964 6332 3016 6341
rect 3424 6264 3476 6316
rect 4712 6400 4764 6452
rect 5080 6400 5132 6452
rect 5540 6400 5592 6452
rect 6920 6400 6972 6452
rect 7840 6400 7892 6452
rect 8852 6443 8904 6452
rect 8852 6409 8861 6443
rect 8861 6409 8895 6443
rect 8895 6409 8904 6443
rect 8852 6400 8904 6409
rect 9128 6400 9180 6452
rect 9312 6443 9364 6452
rect 9312 6409 9321 6443
rect 9321 6409 9355 6443
rect 9355 6409 9364 6443
rect 9312 6400 9364 6409
rect 10416 6400 10468 6452
rect 10692 6443 10744 6452
rect 10692 6409 10701 6443
rect 10701 6409 10735 6443
rect 10735 6409 10744 6443
rect 10692 6400 10744 6409
rect 14648 6443 14700 6452
rect 14648 6409 14657 6443
rect 14657 6409 14691 6443
rect 14691 6409 14700 6443
rect 14648 6400 14700 6409
rect 4068 6332 4120 6384
rect 4896 6264 4948 6316
rect 5080 6264 5132 6316
rect 5540 6307 5592 6316
rect 5540 6273 5549 6307
rect 5549 6273 5583 6307
rect 5583 6273 5592 6307
rect 5540 6264 5592 6273
rect 6184 6332 6236 6384
rect 7748 6332 7800 6384
rect 2596 6128 2648 6180
rect 5264 6196 5316 6248
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 4988 6103 5040 6112
rect 4988 6069 4997 6103
rect 4997 6069 5031 6103
rect 5031 6069 5040 6103
rect 4988 6060 5040 6069
rect 5172 6128 5224 6180
rect 6092 6196 6144 6248
rect 6276 6196 6328 6248
rect 6644 6196 6696 6248
rect 7196 6264 7248 6316
rect 8024 6264 8076 6316
rect 8576 6332 8628 6384
rect 9680 6332 9732 6384
rect 9772 6264 9824 6316
rect 10692 6264 10744 6316
rect 11888 6307 11940 6316
rect 11888 6273 11897 6307
rect 11897 6273 11931 6307
rect 11931 6273 11940 6307
rect 11888 6264 11940 6273
rect 12164 6264 12216 6316
rect 6828 6128 6880 6180
rect 10968 6196 11020 6248
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 12716 6264 12768 6316
rect 15476 6332 15528 6384
rect 13268 6239 13320 6248
rect 5540 6060 5592 6112
rect 6276 6060 6328 6112
rect 6644 6060 6696 6112
rect 6736 6060 6788 6112
rect 10508 6128 10560 6180
rect 13268 6205 13277 6239
rect 13277 6205 13311 6239
rect 13311 6205 13320 6239
rect 13268 6196 13320 6205
rect 17960 6400 18012 6452
rect 19708 6400 19760 6452
rect 20628 6400 20680 6452
rect 16396 6332 16448 6384
rect 19984 6332 20036 6384
rect 20076 6332 20128 6384
rect 20720 6332 20772 6384
rect 14464 6196 14516 6248
rect 16948 6196 17000 6248
rect 17132 6239 17184 6248
rect 17132 6205 17141 6239
rect 17141 6205 17175 6239
rect 17175 6205 17184 6239
rect 17132 6196 17184 6205
rect 18512 6264 18564 6316
rect 18972 6264 19024 6316
rect 19800 6307 19852 6316
rect 19800 6273 19809 6307
rect 19809 6273 19843 6307
rect 19843 6273 19852 6307
rect 19800 6264 19852 6273
rect 12164 6128 12216 6180
rect 16304 6171 16356 6180
rect 10600 6060 10652 6112
rect 11152 6103 11204 6112
rect 11152 6069 11161 6103
rect 11161 6069 11195 6103
rect 11195 6069 11204 6103
rect 11152 6060 11204 6069
rect 11244 6060 11296 6112
rect 13636 6060 13688 6112
rect 13820 6103 13872 6112
rect 13820 6069 13829 6103
rect 13829 6069 13863 6103
rect 13863 6069 13872 6103
rect 13820 6060 13872 6069
rect 16304 6137 16313 6171
rect 16313 6137 16347 6171
rect 16347 6137 16356 6171
rect 16304 6128 16356 6137
rect 16396 6060 16448 6112
rect 16672 6103 16724 6112
rect 16672 6069 16681 6103
rect 16681 6069 16715 6103
rect 16715 6069 16724 6103
rect 16672 6060 16724 6069
rect 16948 6060 17000 6112
rect 18144 6060 18196 6112
rect 18696 6196 18748 6248
rect 19524 6196 19576 6248
rect 20904 6239 20956 6248
rect 20904 6205 20913 6239
rect 20913 6205 20947 6239
rect 20947 6205 20956 6239
rect 20904 6196 20956 6205
rect 18880 6128 18932 6180
rect 20628 6060 20680 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 2688 5856 2740 5908
rect 3976 5856 4028 5908
rect 5172 5899 5224 5908
rect 5172 5865 5181 5899
rect 5181 5865 5215 5899
rect 5215 5865 5224 5899
rect 5172 5856 5224 5865
rect 6736 5856 6788 5908
rect 7104 5899 7156 5908
rect 7104 5865 7113 5899
rect 7113 5865 7147 5899
rect 7147 5865 7156 5899
rect 7104 5856 7156 5865
rect 8208 5856 8260 5908
rect 9496 5856 9548 5908
rect 12164 5856 12216 5908
rect 13268 5856 13320 5908
rect 5724 5788 5776 5840
rect 6000 5788 6052 5840
rect 6920 5788 6972 5840
rect 7472 5788 7524 5840
rect 9680 5788 9732 5840
rect 11980 5831 12032 5840
rect 11980 5797 11989 5831
rect 11989 5797 12023 5831
rect 12023 5797 12032 5831
rect 11980 5788 12032 5797
rect 14372 5788 14424 5840
rect 5264 5720 5316 5772
rect 1584 5695 1636 5704
rect 1584 5661 1593 5695
rect 1593 5661 1627 5695
rect 1627 5661 1636 5695
rect 1584 5652 1636 5661
rect 4620 5652 4672 5704
rect 5448 5695 5500 5704
rect 5448 5661 5457 5695
rect 5457 5661 5491 5695
rect 5491 5661 5500 5695
rect 5448 5652 5500 5661
rect 5908 5695 5960 5704
rect 5908 5661 5917 5695
rect 5917 5661 5951 5695
rect 5951 5661 5960 5695
rect 5908 5652 5960 5661
rect 1860 5584 1912 5636
rect 2320 5627 2372 5636
rect 2320 5593 2332 5627
rect 2332 5593 2372 5627
rect 2320 5584 2372 5593
rect 2964 5584 3016 5636
rect 4160 5584 4212 5636
rect 5356 5584 5408 5636
rect 6644 5763 6696 5772
rect 6644 5729 6653 5763
rect 6653 5729 6687 5763
rect 6687 5729 6696 5763
rect 6644 5720 6696 5729
rect 7288 5720 7340 5772
rect 9496 5763 9548 5772
rect 7564 5695 7616 5704
rect 7564 5661 7573 5695
rect 7573 5661 7607 5695
rect 7607 5661 7616 5695
rect 7564 5652 7616 5661
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 11704 5720 11756 5772
rect 12348 5763 12400 5772
rect 12348 5729 12357 5763
rect 12357 5729 12391 5763
rect 12391 5729 12400 5763
rect 12348 5720 12400 5729
rect 13820 5720 13872 5772
rect 15844 5856 15896 5908
rect 18880 5899 18932 5908
rect 8116 5652 8168 5704
rect 8392 5652 8444 5704
rect 9680 5652 9732 5704
rect 10324 5695 10376 5704
rect 10324 5661 10333 5695
rect 10333 5661 10367 5695
rect 10367 5661 10376 5695
rect 10324 5652 10376 5661
rect 10968 5652 11020 5704
rect 11980 5652 12032 5704
rect 12440 5652 12492 5704
rect 12992 5652 13044 5704
rect 6184 5584 6236 5636
rect 2872 5516 2924 5568
rect 3424 5559 3476 5568
rect 3424 5525 3433 5559
rect 3433 5525 3467 5559
rect 3467 5525 3476 5559
rect 3424 5516 3476 5525
rect 4620 5516 4672 5568
rect 6736 5559 6788 5568
rect 6736 5525 6745 5559
rect 6745 5525 6779 5559
rect 6779 5525 6788 5559
rect 6736 5516 6788 5525
rect 6920 5516 6972 5568
rect 12072 5584 12124 5636
rect 12900 5584 12952 5636
rect 13268 5584 13320 5636
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 9404 5559 9456 5568
rect 9404 5525 9413 5559
rect 9413 5525 9447 5559
rect 9447 5525 9456 5559
rect 9404 5516 9456 5525
rect 11704 5559 11756 5568
rect 11704 5525 11713 5559
rect 11713 5525 11747 5559
rect 11747 5525 11756 5559
rect 11704 5516 11756 5525
rect 14280 5516 14332 5568
rect 16396 5763 16448 5772
rect 16396 5729 16405 5763
rect 16405 5729 16439 5763
rect 16439 5729 16448 5763
rect 16396 5720 16448 5729
rect 18880 5865 18889 5899
rect 18889 5865 18923 5899
rect 18923 5865 18932 5899
rect 18880 5856 18932 5865
rect 20168 5856 20220 5908
rect 20444 5856 20496 5908
rect 19248 5788 19300 5840
rect 15476 5695 15528 5704
rect 15476 5661 15485 5695
rect 15485 5661 15519 5695
rect 15519 5661 15528 5695
rect 15476 5652 15528 5661
rect 17500 5695 17552 5704
rect 17500 5661 17509 5695
rect 17509 5661 17543 5695
rect 17543 5661 17552 5695
rect 17500 5652 17552 5661
rect 17776 5695 17828 5704
rect 17776 5661 17810 5695
rect 17810 5661 17828 5695
rect 17776 5652 17828 5661
rect 19524 5652 19576 5704
rect 20720 5788 20772 5840
rect 20536 5720 20588 5772
rect 20628 5695 20680 5704
rect 20628 5661 20637 5695
rect 20637 5661 20671 5695
rect 20671 5661 20680 5695
rect 20628 5652 20680 5661
rect 15292 5584 15344 5636
rect 17592 5584 17644 5636
rect 17960 5584 18012 5636
rect 18696 5584 18748 5636
rect 17040 5516 17092 5568
rect 17868 5516 17920 5568
rect 18972 5516 19024 5568
rect 19524 5516 19576 5568
rect 20260 5516 20312 5568
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 3056 5355 3108 5364
rect 3056 5321 3065 5355
rect 3065 5321 3099 5355
rect 3099 5321 3108 5355
rect 3056 5312 3108 5321
rect 5908 5312 5960 5364
rect 6736 5312 6788 5364
rect 3332 5176 3384 5228
rect 5816 5244 5868 5296
rect 7840 5312 7892 5364
rect 11152 5312 11204 5364
rect 13544 5312 13596 5364
rect 8484 5244 8536 5296
rect 11244 5244 11296 5296
rect 12348 5244 12400 5296
rect 12992 5287 13044 5296
rect 12992 5253 13001 5287
rect 13001 5253 13035 5287
rect 13035 5253 13044 5287
rect 12992 5244 13044 5253
rect 15568 5244 15620 5296
rect 16120 5312 16172 5364
rect 16396 5312 16448 5364
rect 3976 5176 4028 5228
rect 1492 5108 1544 5160
rect 1860 5108 1912 5160
rect 2504 5108 2556 5160
rect 2872 5151 2924 5160
rect 2872 5117 2881 5151
rect 2881 5117 2915 5151
rect 2915 5117 2924 5151
rect 2872 5108 2924 5117
rect 4436 5176 4488 5228
rect 6000 5176 6052 5228
rect 6460 5176 6512 5228
rect 9496 5176 9548 5228
rect 11704 5219 11756 5228
rect 11704 5185 11713 5219
rect 11713 5185 11747 5219
rect 11747 5185 11756 5219
rect 11704 5176 11756 5185
rect 15844 5244 15896 5296
rect 2596 5040 2648 5092
rect 3332 4972 3384 5024
rect 5724 5040 5776 5092
rect 6828 5040 6880 5092
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 9220 5040 9272 5092
rect 9404 5040 9456 5092
rect 15292 5108 15344 5160
rect 13084 5040 13136 5092
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16948 5312 17000 5364
rect 17132 5312 17184 5364
rect 17592 5312 17644 5364
rect 18696 5355 18748 5364
rect 18696 5321 18705 5355
rect 18705 5321 18739 5355
rect 18739 5321 18748 5355
rect 18696 5312 18748 5321
rect 20536 5312 20588 5364
rect 17040 5287 17092 5296
rect 17040 5253 17049 5287
rect 17049 5253 17083 5287
rect 17083 5253 17092 5287
rect 17040 5244 17092 5253
rect 17500 5244 17552 5296
rect 17776 5176 17828 5228
rect 17960 5176 18012 5228
rect 18880 5176 18932 5228
rect 21180 5244 21232 5296
rect 19248 5219 19300 5228
rect 16948 5151 17000 5160
rect 16948 5117 16957 5151
rect 16957 5117 16991 5151
rect 16991 5117 17000 5151
rect 16948 5108 17000 5117
rect 19248 5185 19282 5219
rect 19282 5185 19300 5219
rect 19248 5176 19300 5185
rect 20536 5176 20588 5228
rect 17960 5040 18012 5092
rect 8300 5015 8352 5024
rect 8300 4981 8309 5015
rect 8309 4981 8343 5015
rect 8343 4981 8352 5015
rect 8300 4972 8352 4981
rect 9588 4972 9640 5024
rect 11244 4972 11296 5024
rect 11796 4972 11848 5024
rect 12440 4972 12492 5024
rect 13544 4972 13596 5024
rect 16120 5015 16172 5024
rect 16120 4981 16129 5015
rect 16129 4981 16163 5015
rect 16163 4981 16172 5015
rect 16120 4972 16172 4981
rect 21272 5015 21324 5024
rect 21272 4981 21281 5015
rect 21281 4981 21315 5015
rect 21315 4981 21324 5015
rect 21272 4972 21324 4981
rect 204 4836 256 4888
rect 940 4836 992 4888
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 2504 4811 2556 4820
rect 2504 4777 2513 4811
rect 2513 4777 2547 4811
rect 2547 4777 2556 4811
rect 2504 4768 2556 4777
rect 3884 4768 3936 4820
rect 4436 4768 4488 4820
rect 6828 4768 6880 4820
rect 8392 4768 8444 4820
rect 12256 4768 12308 4820
rect 12900 4811 12952 4820
rect 12900 4777 12909 4811
rect 12909 4777 12943 4811
rect 12943 4777 12952 4811
rect 12900 4768 12952 4777
rect 1952 4700 2004 4752
rect 2228 4675 2280 4684
rect 2228 4641 2237 4675
rect 2237 4641 2271 4675
rect 2271 4641 2280 4675
rect 2228 4632 2280 4641
rect 2596 4632 2648 4684
rect 2136 4564 2188 4616
rect 3976 4564 4028 4616
rect 4804 4632 4856 4684
rect 5908 4700 5960 4752
rect 10968 4700 11020 4752
rect 15292 4768 15344 4820
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 17776 4700 17828 4752
rect 18052 4743 18104 4752
rect 18052 4709 18061 4743
rect 18061 4709 18095 4743
rect 18095 4709 18104 4743
rect 18052 4700 18104 4709
rect 19984 4700 20036 4752
rect 6552 4632 6604 4684
rect 6736 4632 6788 4684
rect 9220 4632 9272 4684
rect 9588 4675 9640 4684
rect 9588 4641 9597 4675
rect 9597 4641 9631 4675
rect 9631 4641 9640 4675
rect 9588 4632 9640 4641
rect 12992 4632 13044 4684
rect 14096 4675 14148 4684
rect 14096 4641 14105 4675
rect 14105 4641 14139 4675
rect 14139 4641 14148 4675
rect 14096 4632 14148 4641
rect 16120 4632 16172 4684
rect 21180 4675 21232 4684
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7564 4564 7616 4616
rect 9128 4564 9180 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 11152 4564 11204 4616
rect 13820 4564 13872 4616
rect 14740 4564 14792 4616
rect 15752 4607 15804 4616
rect 15752 4573 15761 4607
rect 15761 4573 15795 4607
rect 15795 4573 15804 4607
rect 15752 4564 15804 4573
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 17408 4607 17460 4616
rect 17408 4573 17417 4607
rect 17417 4573 17451 4607
rect 17451 4573 17460 4607
rect 17408 4564 17460 4573
rect 3332 4496 3384 4548
rect 11796 4539 11848 4548
rect 11796 4505 11830 4539
rect 11830 4505 11848 4539
rect 11796 4496 11848 4505
rect 12072 4496 12124 4548
rect 19064 4564 19116 4616
rect 21180 4641 21189 4675
rect 21189 4641 21223 4675
rect 21223 4641 21232 4675
rect 21180 4632 21232 4641
rect 21272 4564 21324 4616
rect 3240 4428 3292 4480
rect 4068 4428 4120 4480
rect 4528 4471 4580 4480
rect 4528 4437 4537 4471
rect 4537 4437 4571 4471
rect 4571 4437 4580 4471
rect 4896 4471 4948 4480
rect 4528 4428 4580 4437
rect 4896 4437 4905 4471
rect 4905 4437 4939 4471
rect 4939 4437 4948 4471
rect 4896 4428 4948 4437
rect 5172 4471 5224 4480
rect 5172 4437 5181 4471
rect 5181 4437 5215 4471
rect 5215 4437 5224 4471
rect 5172 4428 5224 4437
rect 7104 4428 7156 4480
rect 8392 4428 8444 4480
rect 10784 4471 10836 4480
rect 10784 4437 10793 4471
rect 10793 4437 10827 4471
rect 10827 4437 10836 4471
rect 10784 4428 10836 4437
rect 11888 4428 11940 4480
rect 13820 4428 13872 4480
rect 14372 4428 14424 4480
rect 15200 4428 15252 4480
rect 15936 4471 15988 4480
rect 15936 4437 15945 4471
rect 15945 4437 15979 4471
rect 15979 4437 15988 4471
rect 15936 4428 15988 4437
rect 16948 4471 17000 4480
rect 16948 4437 16957 4471
rect 16957 4437 16991 4471
rect 16991 4437 17000 4471
rect 16948 4428 17000 4437
rect 18512 4428 18564 4480
rect 18696 4471 18748 4480
rect 18696 4437 18705 4471
rect 18705 4437 18739 4471
rect 18739 4437 18748 4471
rect 18696 4428 18748 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 1492 4267 1544 4276
rect 1492 4233 1501 4267
rect 1501 4233 1535 4267
rect 1535 4233 1544 4267
rect 1492 4224 1544 4233
rect 3332 4267 3384 4276
rect 3332 4233 3341 4267
rect 3341 4233 3375 4267
rect 3375 4233 3384 4267
rect 3332 4224 3384 4233
rect 1952 4156 2004 4208
rect 4620 4224 4672 4276
rect 8668 4224 8720 4276
rect 10508 4224 10560 4276
rect 10876 4224 10928 4276
rect 11152 4224 11204 4276
rect 14096 4224 14148 4276
rect 3884 4156 3936 4208
rect 4436 4156 4488 4208
rect 4804 4156 4856 4208
rect 5172 4156 5224 4208
rect 6644 4199 6696 4208
rect 6644 4165 6653 4199
rect 6653 4165 6687 4199
rect 6687 4165 6696 4199
rect 6644 4156 6696 4165
rect 1584 4088 1636 4140
rect 2596 4131 2648 4140
rect 2596 4097 2614 4131
rect 2614 4097 2648 4131
rect 2596 4088 2648 4097
rect 2964 4020 3016 4072
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 5724 4088 5776 4140
rect 6092 4088 6144 4140
rect 4896 4020 4948 4072
rect 5172 4063 5224 4072
rect 5172 4029 5181 4063
rect 5181 4029 5215 4063
rect 5215 4029 5224 4063
rect 7748 4088 7800 4140
rect 6552 4063 6604 4072
rect 5172 4020 5224 4029
rect 6552 4029 6561 4063
rect 6561 4029 6595 4063
rect 6595 4029 6604 4063
rect 6552 4020 6604 4029
rect 8484 4063 8536 4072
rect 8484 4029 8493 4063
rect 8493 4029 8527 4063
rect 8527 4029 8536 4063
rect 8484 4020 8536 4029
rect 9588 4156 9640 4208
rect 9404 4131 9456 4140
rect 9404 4097 9413 4131
rect 9413 4097 9447 4131
rect 9447 4097 9456 4131
rect 9404 4088 9456 4097
rect 10048 4088 10100 4140
rect 12072 4156 12124 4208
rect 9128 4063 9180 4072
rect 9128 4029 9137 4063
rect 9137 4029 9171 4063
rect 9171 4029 9180 4063
rect 9128 4020 9180 4029
rect 9680 4020 9732 4072
rect 10876 4063 10928 4072
rect 10876 4029 10885 4063
rect 10885 4029 10919 4063
rect 10919 4029 10928 4063
rect 10876 4020 10928 4029
rect 9588 3952 9640 4004
rect 12348 4088 12400 4140
rect 13084 4131 13136 4140
rect 13084 4097 13093 4131
rect 13093 4097 13127 4131
rect 13127 4097 13136 4131
rect 13084 4088 13136 4097
rect 13544 4131 13596 4140
rect 13544 4097 13553 4131
rect 13553 4097 13587 4131
rect 13587 4097 13596 4131
rect 13544 4088 13596 4097
rect 14556 4156 14608 4208
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 14740 4020 14792 4072
rect 15200 4131 15252 4140
rect 15200 4097 15234 4131
rect 15234 4097 15252 4131
rect 15200 4088 15252 4097
rect 17500 4156 17552 4208
rect 16948 4131 17000 4140
rect 16948 4097 16982 4131
rect 16982 4097 17000 4131
rect 16948 4088 17000 4097
rect 18144 4224 18196 4276
rect 18236 4156 18288 4208
rect 20168 4199 20220 4208
rect 20168 4165 20177 4199
rect 20177 4165 20211 4199
rect 20211 4165 20220 4199
rect 20168 4156 20220 4165
rect 12624 3995 12676 4004
rect 12624 3961 12633 3995
rect 12633 3961 12667 3995
rect 12667 3961 12676 3995
rect 12624 3952 12676 3961
rect 5448 3884 5500 3936
rect 6184 3884 6236 3936
rect 6920 3884 6972 3936
rect 7012 3884 7064 3936
rect 7288 3884 7340 3936
rect 8116 3884 8168 3936
rect 8208 3884 8260 3936
rect 10048 3884 10100 3936
rect 10140 3884 10192 3936
rect 11704 3927 11756 3936
rect 11704 3893 11713 3927
rect 11713 3893 11747 3927
rect 11747 3893 11756 3927
rect 11704 3884 11756 3893
rect 13728 3927 13780 3936
rect 13728 3893 13737 3927
rect 13737 3893 13771 3927
rect 13771 3893 13780 3927
rect 13728 3884 13780 3893
rect 14556 3884 14608 3936
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 19616 4020 19668 4072
rect 20536 4063 20588 4072
rect 20536 4029 20545 4063
rect 20545 4029 20579 4063
rect 20579 4029 20588 4063
rect 20536 4020 20588 4029
rect 20444 3952 20496 4004
rect 16304 3884 16356 3893
rect 19064 3884 19116 3936
rect 20076 3927 20128 3936
rect 20076 3893 20085 3927
rect 20085 3893 20119 3927
rect 20119 3893 20128 3927
rect 20076 3884 20128 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 1032 3680 1084 3732
rect 3056 3680 3108 3732
rect 3884 3680 3936 3732
rect 7104 3680 7156 3732
rect 8024 3680 8076 3732
rect 9404 3680 9456 3732
rect 9588 3680 9640 3732
rect 12900 3680 12952 3732
rect 14556 3680 14608 3732
rect 3792 3612 3844 3664
rect 6184 3612 6236 3664
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 572 3476 624 3528
rect 2320 3544 2372 3596
rect 2780 3544 2832 3596
rect 4344 3587 4396 3596
rect 4344 3553 4353 3587
rect 4353 3553 4387 3587
rect 4387 3553 4396 3587
rect 4344 3544 4396 3553
rect 4620 3587 4672 3596
rect 4620 3553 4629 3587
rect 4629 3553 4663 3587
rect 4663 3553 4672 3587
rect 4620 3544 4672 3553
rect 5724 3587 5776 3596
rect 5724 3553 5733 3587
rect 5733 3553 5767 3587
rect 5767 3553 5776 3587
rect 5724 3544 5776 3553
rect 6092 3544 6144 3596
rect 3240 3476 3292 3528
rect 5816 3519 5868 3528
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 6000 3476 6052 3528
rect 6920 3612 6972 3664
rect 7012 3587 7064 3596
rect 7012 3553 7021 3587
rect 7021 3553 7055 3587
rect 7055 3553 7064 3587
rect 7012 3544 7064 3553
rect 7288 3612 7340 3664
rect 7748 3612 7800 3664
rect 8944 3612 8996 3664
rect 10324 3612 10376 3664
rect 11612 3612 11664 3664
rect 13636 3655 13688 3664
rect 13636 3621 13645 3655
rect 13645 3621 13679 3655
rect 13679 3621 13688 3655
rect 13636 3612 13688 3621
rect 13728 3612 13780 3664
rect 8116 3587 8168 3596
rect 8116 3553 8125 3587
rect 8125 3553 8159 3587
rect 8159 3553 8168 3587
rect 8116 3544 8168 3553
rect 4252 3408 4304 3460
rect 4620 3408 4672 3460
rect 4988 3451 5040 3460
rect 4988 3417 4997 3451
rect 4997 3417 5031 3451
rect 5031 3417 5040 3451
rect 4988 3408 5040 3417
rect 6552 3476 6604 3528
rect 7656 3476 7708 3528
rect 8300 3476 8352 3528
rect 8392 3408 8444 3460
rect 8668 3408 8720 3460
rect 9772 3408 9824 3460
rect 10876 3544 10928 3596
rect 10600 3476 10652 3528
rect 3332 3340 3384 3392
rect 7932 3340 7984 3392
rect 8116 3340 8168 3392
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 10600 3383 10652 3392
rect 10600 3349 10609 3383
rect 10609 3349 10643 3383
rect 10643 3349 10652 3383
rect 10600 3340 10652 3349
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11244 3476 11296 3528
rect 12164 3519 12216 3528
rect 12164 3485 12173 3519
rect 12173 3485 12207 3519
rect 12207 3485 12216 3519
rect 12164 3476 12216 3485
rect 12808 3519 12860 3528
rect 12808 3485 12817 3519
rect 12817 3485 12851 3519
rect 12851 3485 12860 3519
rect 12808 3476 12860 3485
rect 14188 3519 14240 3528
rect 14188 3485 14197 3519
rect 14197 3485 14231 3519
rect 14231 3485 14240 3519
rect 14188 3476 14240 3485
rect 15200 3544 15252 3596
rect 16028 3476 16080 3528
rect 18696 3680 18748 3732
rect 22284 3680 22336 3732
rect 19524 3612 19576 3664
rect 19800 3544 19852 3596
rect 21640 3544 21692 3596
rect 11796 3383 11848 3392
rect 11796 3349 11805 3383
rect 11805 3349 11839 3383
rect 11839 3349 11848 3383
rect 11796 3340 11848 3349
rect 12624 3383 12676 3392
rect 12624 3349 12633 3383
rect 12633 3349 12667 3383
rect 12667 3349 12676 3383
rect 12624 3340 12676 3349
rect 14648 3408 14700 3460
rect 15844 3408 15896 3460
rect 15936 3408 15988 3460
rect 20352 3476 20404 3528
rect 18972 3408 19024 3460
rect 20628 3408 20680 3460
rect 15108 3340 15160 3392
rect 15384 3383 15436 3392
rect 15384 3349 15393 3383
rect 15393 3349 15427 3383
rect 15427 3349 15436 3383
rect 15384 3340 15436 3349
rect 15476 3340 15528 3392
rect 16028 3383 16080 3392
rect 16028 3349 16037 3383
rect 16037 3349 16071 3383
rect 16071 3349 16080 3383
rect 16028 3340 16080 3349
rect 16396 3340 16448 3392
rect 17132 3383 17184 3392
rect 17132 3349 17141 3383
rect 17141 3349 17175 3383
rect 17175 3349 17184 3383
rect 17132 3340 17184 3349
rect 17684 3383 17736 3392
rect 17684 3349 17693 3383
rect 17693 3349 17727 3383
rect 17727 3349 17736 3383
rect 17684 3340 17736 3349
rect 18604 3340 18656 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 1768 3000 1820 3052
rect 2780 3136 2832 3188
rect 3976 3179 4028 3188
rect 3976 3145 3985 3179
rect 3985 3145 4019 3179
rect 4019 3145 4028 3179
rect 3976 3136 4028 3145
rect 5172 3068 5224 3120
rect 6920 3136 6972 3188
rect 7472 3179 7524 3188
rect 7472 3145 7481 3179
rect 7481 3145 7515 3179
rect 7515 3145 7524 3179
rect 7472 3136 7524 3145
rect 5724 3000 5776 3052
rect 6920 3043 6972 3052
rect 6920 3009 6929 3043
rect 6929 3009 6963 3043
rect 6963 3009 6972 3043
rect 6920 3000 6972 3009
rect 7104 3000 7156 3052
rect 2964 2796 3016 2848
rect 6000 2932 6052 2984
rect 4068 2796 4120 2848
rect 7840 3000 7892 3052
rect 7748 2932 7800 2984
rect 8300 3068 8352 3120
rect 9128 3136 9180 3188
rect 9680 3179 9732 3188
rect 9680 3145 9689 3179
rect 9689 3145 9723 3179
rect 9723 3145 9732 3179
rect 9680 3136 9732 3145
rect 10600 3136 10652 3188
rect 10140 3111 10192 3120
rect 10140 3077 10149 3111
rect 10149 3077 10183 3111
rect 10183 3077 10192 3111
rect 10140 3068 10192 3077
rect 10876 3000 10928 3052
rect 12624 3136 12676 3188
rect 12716 3136 12768 3188
rect 14188 3136 14240 3188
rect 15292 3136 15344 3188
rect 15476 3179 15528 3188
rect 15476 3145 15485 3179
rect 15485 3145 15519 3179
rect 15519 3145 15528 3179
rect 15476 3136 15528 3145
rect 16028 3136 16080 3188
rect 17684 3136 17736 3188
rect 20904 3136 20956 3188
rect 11796 3068 11848 3120
rect 11060 3000 11112 3052
rect 11704 3000 11756 3052
rect 12532 3000 12584 3052
rect 12900 3043 12952 3052
rect 12900 3009 12909 3043
rect 12909 3009 12943 3043
rect 12943 3009 12952 3043
rect 12900 3000 12952 3009
rect 15384 3068 15436 3120
rect 17132 3068 17184 3120
rect 21364 3068 21416 3120
rect 14280 3043 14332 3052
rect 14280 3009 14289 3043
rect 14289 3009 14323 3043
rect 14323 3009 14332 3043
rect 14280 3000 14332 3009
rect 8944 2932 8996 2984
rect 7380 2864 7432 2916
rect 9680 2864 9732 2916
rect 10324 2864 10376 2916
rect 12164 2932 12216 2984
rect 15660 3000 15712 3052
rect 16304 2932 16356 2984
rect 17040 3000 17092 3052
rect 17316 3000 17368 3052
rect 18052 3043 18104 3052
rect 18052 3009 18061 3043
rect 18061 3009 18095 3043
rect 18095 3009 18104 3043
rect 18052 3000 18104 3009
rect 18328 3043 18380 3052
rect 18328 3009 18337 3043
rect 18337 3009 18371 3043
rect 18371 3009 18380 3043
rect 18328 3000 18380 3009
rect 19892 3000 19944 3052
rect 20076 3000 20128 3052
rect 21088 3043 21140 3052
rect 21088 3009 21097 3043
rect 21097 3009 21131 3043
rect 21131 3009 21140 3043
rect 21088 3000 21140 3009
rect 22744 3000 22796 3052
rect 17960 2932 18012 2984
rect 20720 2975 20772 2984
rect 20720 2941 20729 2975
rect 20729 2941 20763 2975
rect 20763 2941 20772 2975
rect 20720 2932 20772 2941
rect 13820 2864 13872 2916
rect 11152 2839 11204 2848
rect 11152 2805 11161 2839
rect 11161 2805 11195 2839
rect 11195 2805 11204 2839
rect 11152 2796 11204 2805
rect 12532 2796 12584 2848
rect 12992 2796 13044 2848
rect 16672 2864 16724 2916
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 14832 2796 14884 2848
rect 15936 2796 15988 2848
rect 17316 2796 17368 2848
rect 18236 2796 18288 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 1584 2635 1636 2644
rect 1584 2601 1593 2635
rect 1593 2601 1627 2635
rect 1627 2601 1636 2635
rect 1584 2592 1636 2601
rect 1308 2524 1360 2576
rect 3240 2592 3292 2644
rect 3884 2592 3936 2644
rect 2964 2499 3016 2508
rect 2964 2465 2973 2499
rect 2973 2465 3007 2499
rect 3007 2465 3016 2499
rect 2964 2456 3016 2465
rect 5356 2456 5408 2508
rect 5448 2499 5500 2508
rect 5448 2465 5457 2499
rect 5457 2465 5491 2499
rect 5491 2465 5500 2499
rect 6644 2592 6696 2644
rect 8024 2592 8076 2644
rect 9404 2635 9456 2644
rect 9404 2601 9413 2635
rect 9413 2601 9447 2635
rect 9447 2601 9456 2635
rect 9404 2592 9456 2601
rect 5448 2456 5500 2465
rect 7748 2499 7800 2508
rect 7748 2465 7757 2499
rect 7757 2465 7791 2499
rect 7791 2465 7800 2499
rect 7748 2456 7800 2465
rect 7932 2456 7984 2508
rect 4436 2388 4488 2440
rect 4528 2388 4580 2440
rect 6736 2388 6788 2440
rect 9220 2524 9272 2576
rect 9680 2592 9732 2644
rect 10048 2635 10100 2644
rect 10048 2601 10057 2635
rect 10057 2601 10091 2635
rect 10091 2601 10100 2635
rect 10048 2592 10100 2601
rect 10416 2592 10468 2644
rect 13176 2592 13228 2644
rect 10692 2524 10744 2576
rect 10968 2524 11020 2576
rect 9772 2456 9824 2508
rect 10416 2456 10468 2508
rect 11980 2524 12032 2576
rect 14096 2524 14148 2576
rect 15016 2524 15068 2576
rect 16396 2524 16448 2576
rect 11152 2456 11204 2508
rect 10876 2388 10928 2440
rect 11244 2388 11296 2440
rect 12532 2388 12584 2440
rect 12992 2388 13044 2440
rect 13820 2388 13872 2440
rect 14648 2431 14700 2440
rect 14648 2397 14657 2431
rect 14657 2397 14691 2431
rect 14691 2397 14700 2431
rect 14648 2388 14700 2397
rect 14740 2388 14792 2440
rect 15844 2456 15896 2508
rect 16672 2431 16724 2440
rect 16672 2397 16681 2431
rect 16681 2397 16715 2431
rect 16715 2397 16724 2431
rect 16672 2388 16724 2397
rect 12624 2320 12676 2372
rect 17776 2524 17828 2576
rect 21456 2456 21508 2508
rect 18512 2388 18564 2440
rect 20260 2431 20312 2440
rect 20260 2397 20269 2431
rect 20269 2397 20303 2431
rect 20303 2397 20312 2431
rect 20260 2388 20312 2397
rect 21272 2388 21324 2440
rect 3424 2295 3476 2304
rect 3424 2261 3433 2295
rect 3433 2261 3467 2295
rect 3467 2261 3476 2295
rect 3424 2252 3476 2261
rect 4068 2252 4120 2304
rect 6828 2252 6880 2304
rect 9128 2295 9180 2304
rect 9128 2261 9137 2295
rect 9137 2261 9171 2295
rect 9171 2261 9180 2295
rect 9128 2252 9180 2261
rect 9312 2252 9364 2304
rect 10784 2252 10836 2304
rect 12808 2252 12860 2304
rect 13268 2252 13320 2304
rect 13728 2252 13780 2304
rect 14556 2252 14608 2304
rect 15476 2252 15528 2304
rect 17224 2252 17276 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 2412 2048 2464 2100
rect 5264 2048 5316 2100
rect 5632 2048 5684 2100
rect 9312 2048 9364 2100
rect 16212 2048 16264 2100
rect 20536 2048 20588 2100
rect 3056 1980 3108 2032
rect 7564 1980 7616 2032
rect 15108 1980 15160 2032
rect 19800 1980 19852 2032
rect 9128 1912 9180 1964
rect 17040 1912 17092 1964
rect 3424 1300 3476 1352
rect 7196 1300 7248 1352
rect 14372 1300 14424 1352
rect 18328 1300 18380 1352
<< metal2 >>
rect 4526 22672 4582 22681
rect 4526 22607 4582 22616
rect 2042 22264 2098 22273
rect 2042 22199 2098 22208
rect 1490 21720 1546 21729
rect 1490 21655 1546 21664
rect 1504 20602 1532 21655
rect 1950 20768 2006 20777
rect 1950 20703 2006 20712
rect 1492 20596 1544 20602
rect 1492 20538 1544 20544
rect 1492 19712 1544 19718
rect 1492 19654 1544 19660
rect 1504 19417 1532 19654
rect 1964 19514 1992 20703
rect 2056 20602 2084 22199
rect 2870 21312 2926 21321
rect 2870 21247 2926 21256
rect 2044 20596 2096 20602
rect 2044 20538 2096 20544
rect 2778 20360 2834 20369
rect 2778 20295 2780 20304
rect 2832 20295 2834 20304
rect 2780 20266 2832 20272
rect 2884 20058 2912 21247
rect 2964 20596 3016 20602
rect 2964 20538 3016 20544
rect 2976 20398 3004 20538
rect 4540 20466 4568 22607
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 18694 22672 18750 22681
rect 18694 22607 18750 22616
rect 5736 20466 5764 22200
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 17236 20602 17264 22200
rect 9956 20596 10008 20602
rect 9956 20538 10008 20544
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 3884 20460 3936 20466
rect 3884 20402 3936 20408
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 2964 20392 3016 20398
rect 2964 20334 3016 20340
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 2136 19848 2188 19854
rect 2042 19816 2098 19825
rect 2136 19790 2188 19796
rect 2504 19848 2556 19854
rect 2504 19790 2556 19796
rect 2780 19848 2832 19854
rect 2780 19790 2832 19796
rect 2042 19751 2098 19760
rect 2056 19718 2084 19751
rect 2044 19712 2096 19718
rect 2044 19654 2096 19660
rect 1952 19508 2004 19514
rect 1952 19450 2004 19456
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1504 18873 1532 19110
rect 1688 18970 1716 19314
rect 2148 18970 2176 19790
rect 2516 19514 2544 19790
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2686 19408 2742 19417
rect 2686 19343 2688 19352
rect 2740 19343 2742 19352
rect 2688 19314 2740 19320
rect 2792 18970 2820 19790
rect 3896 19718 3924 20402
rect 4344 19848 4396 19854
rect 4344 19790 4396 19796
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3332 19712 3384 19718
rect 3332 19654 3384 19660
rect 3884 19712 3936 19718
rect 3884 19654 3936 19660
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 3160 19378 3188 19654
rect 3148 19372 3200 19378
rect 3148 19314 3200 19320
rect 3344 19310 3372 19654
rect 3332 19304 3384 19310
rect 3332 19246 3384 19252
rect 1676 18964 1728 18970
rect 1676 18906 1728 18912
rect 2136 18964 2188 18970
rect 2136 18906 2188 18912
rect 2780 18964 2832 18970
rect 2780 18906 2832 18912
rect 1490 18864 1546 18873
rect 1490 18799 1546 18808
rect 1676 18760 1728 18766
rect 1676 18702 1728 18708
rect 2136 18760 2188 18766
rect 2136 18702 2188 18708
rect 1308 18692 1360 18698
rect 1308 18634 1360 18640
rect 938 16280 994 16289
rect 32 16238 938 16266
rect 32 2281 60 16238
rect 938 16215 994 16224
rect 202 15872 258 15881
rect 202 15807 258 15816
rect 216 4894 244 15807
rect 938 15328 994 15337
rect 938 15263 994 15272
rect 952 6798 980 15263
rect 1216 14544 1268 14550
rect 1216 14486 1268 14492
rect 940 6792 992 6798
rect 938 6760 940 6769
rect 992 6760 994 6769
rect 938 6695 994 6704
rect 952 6669 980 6695
rect 204 4888 256 4894
rect 940 4888 992 4894
rect 204 4830 256 4836
rect 938 4856 940 4865
rect 992 4856 994 4865
rect 938 4791 994 4800
rect 1228 4593 1256 14486
rect 1214 4584 1270 4593
rect 1214 4519 1270 4528
rect 1032 3732 1084 3738
rect 1032 3674 1084 3680
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 202 3224 258 3233
rect 202 3159 258 3168
rect 18 2272 74 2281
rect 18 2207 74 2216
rect 216 800 244 3159
rect 584 800 612 3470
rect 1044 800 1072 3674
rect 1320 2582 1348 18634
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1504 18465 1532 18566
rect 1490 18456 1546 18465
rect 1688 18426 1716 18702
rect 1490 18391 1546 18400
rect 1676 18420 1728 18426
rect 1676 18362 1728 18368
rect 2148 18193 2176 18702
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2700 18290 2728 18634
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18358 3280 18566
rect 3240 18352 3292 18358
rect 3240 18294 3292 18300
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 3344 18222 3372 19246
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 3884 18624 3936 18630
rect 3884 18566 3936 18572
rect 3896 18426 3924 18566
rect 3884 18420 3936 18426
rect 3884 18362 3936 18368
rect 3896 18306 3924 18362
rect 3896 18290 4016 18306
rect 3424 18284 3476 18290
rect 3896 18284 4028 18290
rect 3896 18278 3976 18284
rect 3424 18226 3476 18232
rect 3976 18226 4028 18232
rect 3332 18216 3384 18222
rect 2134 18184 2190 18193
rect 3332 18158 3384 18164
rect 2134 18119 2190 18128
rect 2320 18148 2372 18154
rect 2320 18090 2372 18096
rect 1492 18080 1544 18086
rect 1490 18048 1492 18057
rect 1544 18048 1546 18057
rect 1490 17983 1546 17992
rect 1492 17536 1544 17542
rect 1490 17504 1492 17513
rect 2044 17536 2096 17542
rect 1544 17504 1546 17513
rect 2044 17478 2096 17484
rect 1490 17439 1546 17448
rect 1490 17096 1546 17105
rect 1490 17031 1492 17040
rect 1544 17031 1546 17040
rect 1492 17002 1544 17008
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1964 16590 1992 16934
rect 1676 16584 1728 16590
rect 1676 16526 1728 16532
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16153 1532 16390
rect 1490 16144 1546 16153
rect 1490 16079 1546 16088
rect 1492 15904 1544 15910
rect 1492 15846 1544 15852
rect 1504 15609 1532 15846
rect 1688 15706 1716 16526
rect 1676 15700 1728 15706
rect 1676 15642 1728 15648
rect 1490 15600 1546 15609
rect 2056 15570 2084 17478
rect 2332 16574 2360 18090
rect 2780 18080 2832 18086
rect 2780 18022 2832 18028
rect 2792 17746 2820 18022
rect 3240 17808 3292 17814
rect 3240 17750 3292 17756
rect 2780 17740 2832 17746
rect 2780 17682 2832 17688
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2504 16720 2556 16726
rect 2504 16662 2556 16668
rect 2134 16552 2190 16561
rect 2134 16487 2190 16496
rect 2240 16546 2360 16574
rect 2148 16454 2176 16487
rect 2136 16448 2188 16454
rect 2136 16390 2188 16396
rect 1490 15535 1546 15544
rect 2044 15564 2096 15570
rect 2044 15506 2096 15512
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 2136 15360 2188 15366
rect 2136 15302 2188 15308
rect 1504 15201 1532 15302
rect 1490 15192 1546 15201
rect 1490 15127 1546 15136
rect 2148 15026 2176 15302
rect 1952 15020 2004 15026
rect 1952 14962 2004 14968
rect 2136 15020 2188 15026
rect 2136 14962 2188 14968
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1676 14816 1728 14822
rect 1676 14758 1728 14764
rect 1504 14657 1532 14758
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1688 14414 1716 14758
rect 1964 14618 1992 14962
rect 1952 14612 2004 14618
rect 1952 14554 2004 14560
rect 1676 14408 1728 14414
rect 1676 14350 1728 14356
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1676 13932 1728 13938
rect 1676 13874 1728 13880
rect 1490 13832 1546 13841
rect 1490 13767 1492 13776
rect 1544 13767 1546 13776
rect 1492 13738 1544 13744
rect 1398 13424 1454 13433
rect 1398 13359 1454 13368
rect 1412 7410 1440 13359
rect 1490 13288 1546 13297
rect 1490 13223 1546 13232
rect 1504 13190 1532 13223
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1584 12844 1636 12850
rect 1584 12786 1636 12792
rect 1596 12345 1624 12786
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 1584 12164 1636 12170
rect 1584 12106 1636 12112
rect 1596 11937 1624 12106
rect 1582 11928 1638 11937
rect 1582 11863 1638 11872
rect 1584 11756 1636 11762
rect 1584 11698 1636 11704
rect 1596 11393 1624 11698
rect 1582 11384 1638 11393
rect 1688 11354 1716 13874
rect 2136 13864 2188 13870
rect 2136 13806 2188 13812
rect 2044 13388 2096 13394
rect 2044 13330 2096 13336
rect 1860 13184 1912 13190
rect 1860 13126 1912 13132
rect 1872 12850 1900 13126
rect 1950 12880 2006 12889
rect 1860 12844 1912 12850
rect 1950 12815 2006 12824
rect 1860 12786 1912 12792
rect 1766 12200 1822 12209
rect 1766 12135 1768 12144
rect 1820 12135 1822 12144
rect 1768 12106 1820 12112
rect 1582 11319 1638 11328
rect 1676 11348 1728 11354
rect 1492 11144 1544 11150
rect 1492 11086 1544 11092
rect 1504 10266 1532 11086
rect 1596 10810 1624 11319
rect 1676 11290 1728 11296
rect 1584 10804 1636 10810
rect 1584 10746 1636 10752
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1688 10441 1716 10610
rect 1674 10432 1730 10441
rect 1674 10367 1730 10376
rect 1872 10282 1900 12786
rect 1964 12646 1992 12815
rect 1952 12640 2004 12646
rect 1952 12582 2004 12588
rect 1964 11150 1992 12582
rect 2056 12102 2084 13330
rect 2148 13326 2176 13806
rect 2240 13462 2268 16546
rect 2516 15586 2544 16662
rect 2608 16250 2636 17138
rect 2792 16794 2820 17682
rect 3148 17604 3200 17610
rect 3148 17546 3200 17552
rect 2964 17196 3016 17202
rect 2964 17138 3016 17144
rect 2872 17060 2924 17066
rect 2872 17002 2924 17008
rect 2780 16788 2832 16794
rect 2780 16730 2832 16736
rect 2884 16658 2912 17002
rect 2872 16652 2924 16658
rect 2872 16594 2924 16600
rect 2596 16244 2648 16250
rect 2596 16186 2648 16192
rect 2688 16176 2740 16182
rect 2688 16118 2740 16124
rect 2424 15558 2544 15586
rect 2424 13546 2452 15558
rect 2504 15496 2556 15502
rect 2504 15438 2556 15444
rect 2516 14618 2544 15438
rect 2596 15360 2648 15366
rect 2596 15302 2648 15308
rect 2608 14822 2636 15302
rect 2596 14816 2648 14822
rect 2596 14758 2648 14764
rect 2504 14612 2556 14618
rect 2504 14554 2556 14560
rect 2608 14414 2636 14758
rect 2596 14408 2648 14414
rect 2596 14350 2648 14356
rect 2608 13870 2636 14350
rect 2596 13864 2648 13870
rect 2596 13806 2648 13812
rect 2424 13518 2544 13546
rect 2228 13456 2280 13462
rect 2228 13398 2280 13404
rect 2412 13456 2464 13462
rect 2412 13398 2464 13404
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 2056 11694 2084 12038
rect 2044 11688 2096 11694
rect 2044 11630 2096 11636
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 2136 11076 2188 11082
rect 2136 11018 2188 11024
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1780 10254 1900 10282
rect 1674 10024 1730 10033
rect 1674 9959 1676 9968
rect 1728 9959 1730 9968
rect 1676 9930 1728 9936
rect 1584 9580 1636 9586
rect 1584 9522 1636 9528
rect 1596 9489 1624 9522
rect 1582 9480 1638 9489
rect 1582 9415 1638 9424
rect 1676 8900 1728 8906
rect 1676 8842 1728 8848
rect 1688 8673 1716 8842
rect 1674 8664 1730 8673
rect 1674 8599 1730 8608
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1504 8129 1532 8434
rect 1490 8120 1546 8129
rect 1490 8055 1546 8064
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1676 7404 1728 7410
rect 1676 7346 1728 7352
rect 1582 6896 1638 6905
rect 1582 6831 1638 6840
rect 1596 6225 1624 6831
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 1596 5710 1624 6151
rect 1688 5817 1716 7346
rect 1674 5808 1730 5817
rect 1674 5743 1730 5752
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1492 5160 1544 5166
rect 1492 5102 1544 5108
rect 1504 4282 1532 5102
rect 1492 4276 1544 4282
rect 1492 4218 1544 4224
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 1584 4140 1636 4146
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 1504 800 1532 4111
rect 1584 4082 1636 4088
rect 1596 2650 1624 4082
rect 1780 3058 1808 10254
rect 1952 10192 2004 10198
rect 1858 10160 1914 10169
rect 1952 10134 2004 10140
rect 1858 10095 1860 10104
rect 1912 10095 1914 10104
rect 1860 10066 1912 10072
rect 1860 8900 1912 8906
rect 1860 8842 1912 8848
rect 1872 8401 1900 8842
rect 1964 8498 1992 10134
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 1858 8392 1914 8401
rect 1858 8327 1914 8336
rect 1952 7880 2004 7886
rect 1952 7822 2004 7828
rect 1858 7576 1914 7585
rect 1858 7511 1914 7520
rect 1872 7478 1900 7511
rect 1860 7472 1912 7478
rect 1964 7449 1992 7822
rect 1860 7414 1912 7420
rect 1950 7440 2006 7449
rect 1872 6882 1900 7414
rect 1950 7375 2006 7384
rect 1872 6854 1992 6882
rect 1860 6724 1912 6730
rect 1860 6666 1912 6672
rect 1872 6497 1900 6666
rect 1858 6488 1914 6497
rect 1858 6423 1914 6432
rect 1860 5636 1912 5642
rect 1860 5578 1912 5584
rect 1872 5166 1900 5578
rect 1860 5160 1912 5166
rect 1860 5102 1912 5108
rect 1964 4758 1992 6854
rect 2056 6458 2084 9046
rect 2044 6452 2096 6458
rect 2044 6394 2096 6400
rect 1952 4752 2004 4758
rect 1952 4694 2004 4700
rect 2148 4622 2176 11018
rect 2240 10470 2268 13194
rect 2320 12776 2372 12782
rect 2320 12718 2372 12724
rect 2332 12170 2360 12718
rect 2320 12164 2372 12170
rect 2320 12106 2372 12112
rect 2424 12050 2452 13398
rect 2516 12986 2544 13518
rect 2596 13184 2648 13190
rect 2596 13126 2648 13132
rect 2608 12986 2636 13126
rect 2504 12980 2556 12986
rect 2504 12922 2556 12928
rect 2596 12980 2648 12986
rect 2596 12922 2648 12928
rect 2332 12022 2452 12050
rect 2228 10464 2280 10470
rect 2228 10406 2280 10412
rect 2228 9648 2280 9654
rect 2228 9590 2280 9596
rect 2240 8945 2268 9590
rect 2226 8936 2282 8945
rect 2226 8871 2282 8880
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 2240 7721 2268 7822
rect 2226 7712 2282 7721
rect 2226 7647 2282 7656
rect 2332 7528 2360 12022
rect 2516 11778 2544 12922
rect 2700 11937 2728 16118
rect 2872 16040 2924 16046
rect 2872 15982 2924 15988
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13530 2820 13874
rect 2780 13524 2832 13530
rect 2780 13466 2832 13472
rect 2778 13288 2834 13297
rect 2778 13223 2834 13232
rect 2686 11928 2742 11937
rect 2686 11863 2742 11872
rect 2424 11750 2544 11778
rect 2688 11756 2740 11762
rect 2424 7886 2452 11750
rect 2688 11698 2740 11704
rect 2504 11688 2556 11694
rect 2504 11630 2556 11636
rect 2516 11354 2544 11630
rect 2504 11348 2556 11354
rect 2504 11290 2556 11296
rect 2700 10810 2728 11698
rect 2688 10804 2740 10810
rect 2688 10746 2740 10752
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2516 9625 2544 10474
rect 2792 9994 2820 13223
rect 2780 9988 2832 9994
rect 2780 9930 2832 9936
rect 2884 9722 2912 15982
rect 2976 11218 3004 17138
rect 3160 16590 3188 17546
rect 3252 17134 3280 17750
rect 3344 17746 3372 18158
rect 3332 17740 3384 17746
rect 3332 17682 3384 17688
rect 3240 17128 3292 17134
rect 3240 17070 3292 17076
rect 3240 16652 3292 16658
rect 3240 16594 3292 16600
rect 3148 16584 3200 16590
rect 3148 16526 3200 16532
rect 3148 15360 3200 15366
rect 3148 15302 3200 15308
rect 3160 15094 3188 15302
rect 3148 15088 3200 15094
rect 3148 15030 3200 15036
rect 3160 14482 3188 15030
rect 3148 14476 3200 14482
rect 3148 14418 3200 14424
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3068 14074 3096 14214
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3068 11898 3096 13806
rect 3148 13728 3200 13734
rect 3148 13670 3200 13676
rect 3160 13394 3188 13670
rect 3148 13388 3200 13394
rect 3148 13330 3200 13336
rect 3160 12782 3188 13330
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3146 12608 3202 12617
rect 3146 12543 3202 12552
rect 3056 11892 3108 11898
rect 3056 11834 3108 11840
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2502 9616 2558 9625
rect 2502 9551 2558 9560
rect 2596 9580 2648 9586
rect 2596 9522 2648 9528
rect 2688 9580 2740 9586
rect 2740 9540 2912 9568
rect 2688 9522 2740 9528
rect 2608 9024 2636 9522
rect 2516 8996 2636 9024
rect 2516 8634 2544 8996
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2608 8634 2636 8842
rect 2688 8832 2740 8838
rect 2688 8774 2740 8780
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2504 8628 2556 8634
rect 2504 8570 2556 8576
rect 2596 8628 2648 8634
rect 2596 8570 2648 8576
rect 2516 7954 2544 8570
rect 2700 8090 2728 8774
rect 2688 8084 2740 8090
rect 2688 8026 2740 8032
rect 2504 7948 2556 7954
rect 2504 7890 2556 7896
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2504 7744 2556 7750
rect 2504 7686 2556 7692
rect 2516 7546 2544 7686
rect 2240 7500 2360 7528
rect 2504 7540 2556 7546
rect 2240 6905 2268 7500
rect 2504 7482 2556 7488
rect 2792 7478 2820 8774
rect 2884 8004 2912 9540
rect 2976 8838 3004 11154
rect 3056 10804 3108 10810
rect 3056 10746 3108 10752
rect 3068 9722 3096 10746
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3160 9602 3188 12543
rect 3068 9574 3188 9602
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 3068 8294 3096 9574
rect 3252 9466 3280 16594
rect 3436 16454 3464 18226
rect 3884 18216 3936 18222
rect 3884 18158 3936 18164
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3896 17338 3924 18158
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 4080 16833 4108 19654
rect 4356 19446 4384 19790
rect 4540 19514 4568 20402
rect 6552 20392 6604 20398
rect 6552 20334 6604 20340
rect 4988 20256 5040 20262
rect 4988 20198 5040 20204
rect 4804 19780 4856 19786
rect 4804 19722 4856 19728
rect 4528 19508 4580 19514
rect 4528 19450 4580 19456
rect 4344 19440 4396 19446
rect 4344 19382 4396 19388
rect 4356 18766 4384 19382
rect 4620 18896 4672 18902
rect 4620 18838 4672 18844
rect 4344 18760 4396 18766
rect 4344 18702 4396 18708
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 4264 17678 4292 18022
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4066 16824 4122 16833
rect 4066 16759 4122 16768
rect 4356 16658 4384 18702
rect 4632 18630 4660 18838
rect 4620 18624 4672 18630
rect 4620 18566 4672 18572
rect 4712 18216 4764 18222
rect 4712 18158 4764 18164
rect 4724 17882 4752 18158
rect 4712 17876 4764 17882
rect 4712 17818 4764 17824
rect 4816 16998 4844 19722
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 18222 4936 19110
rect 4896 18216 4948 18222
rect 4896 18158 4948 18164
rect 5000 18034 5028 20198
rect 5264 19848 5316 19854
rect 5264 19790 5316 19796
rect 5276 19174 5304 19790
rect 5724 19712 5776 19718
rect 5724 19654 5776 19660
rect 5264 19168 5316 19174
rect 5264 19110 5316 19116
rect 5736 18766 5764 19654
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 5814 19408 5870 19417
rect 5814 19343 5870 19352
rect 5828 19174 5856 19343
rect 5816 19168 5868 19174
rect 5816 19110 5868 19116
rect 5264 18760 5316 18766
rect 5724 18760 5776 18766
rect 5316 18708 5580 18714
rect 5264 18702 5580 18708
rect 5724 18702 5776 18708
rect 5276 18686 5580 18702
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 4908 18006 5028 18034
rect 5264 18080 5316 18086
rect 5264 18022 5316 18028
rect 4908 17270 4936 18006
rect 4988 17536 5040 17542
rect 4988 17478 5040 17484
rect 5000 17338 5028 17478
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3332 16244 3384 16250
rect 3332 16186 3384 16192
rect 3344 13410 3372 16186
rect 3976 16040 4028 16046
rect 3976 15982 4028 15988
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 3884 14340 3936 14346
rect 3884 14282 3936 14288
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 3436 13530 3464 13806
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 3896 13530 3924 14282
rect 3424 13524 3476 13530
rect 3424 13466 3476 13472
rect 3884 13524 3936 13530
rect 3884 13466 3936 13472
rect 3344 13382 3556 13410
rect 3424 13320 3476 13326
rect 3424 13262 3476 13268
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3344 12918 3372 13126
rect 3332 12912 3384 12918
rect 3332 12854 3384 12860
rect 3436 12102 3464 13262
rect 3528 12753 3556 13382
rect 3514 12744 3570 12753
rect 3514 12679 3570 12688
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 3344 10985 3372 11698
rect 3436 11218 3464 12038
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3330 10976 3386 10985
rect 3330 10911 3386 10920
rect 3332 10668 3384 10674
rect 3332 10610 3384 10616
rect 3344 9722 3372 10610
rect 3436 10606 3464 11154
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3804 10810 3832 11086
rect 3608 10804 3660 10810
rect 3608 10746 3660 10752
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3620 10713 3648 10746
rect 3606 10704 3662 10713
rect 3606 10639 3662 10648
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3896 10130 3924 11222
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3424 10056 3476 10062
rect 3424 9998 3476 10004
rect 3332 9716 3384 9722
rect 3332 9658 3384 9664
rect 3160 9438 3280 9466
rect 3160 8974 3188 9438
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3252 8906 3280 9318
rect 3240 8900 3292 8906
rect 3240 8842 3292 8848
rect 3148 8832 3200 8838
rect 3148 8774 3200 8780
rect 3056 8288 3108 8294
rect 3056 8230 3108 8236
rect 2875 7976 2912 8004
rect 2875 7936 2903 7976
rect 2875 7908 2912 7936
rect 2884 7546 2912 7908
rect 2872 7540 2924 7546
rect 2872 7482 2924 7488
rect 2780 7472 2832 7478
rect 2780 7414 2832 7420
rect 2778 7304 2834 7313
rect 2778 7239 2834 7248
rect 2412 7200 2464 7206
rect 2412 7142 2464 7148
rect 2596 7200 2648 7206
rect 2596 7142 2648 7148
rect 2226 6896 2282 6905
rect 2424 6866 2452 7142
rect 2226 6831 2282 6840
rect 2320 6860 2372 6866
rect 2320 6802 2372 6808
rect 2412 6860 2464 6866
rect 2412 6802 2464 6808
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6458 2268 6666
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2332 5642 2360 6802
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 2424 6458 2452 6598
rect 2412 6452 2464 6458
rect 2412 6394 2464 6400
rect 2608 6390 2636 7142
rect 2688 6452 2740 6458
rect 2688 6394 2740 6400
rect 2596 6384 2648 6390
rect 2596 6326 2648 6332
rect 2596 6180 2648 6186
rect 2596 6122 2648 6128
rect 2320 5636 2372 5642
rect 2320 5578 2372 5584
rect 2504 5160 2556 5166
rect 2504 5102 2556 5108
rect 2516 4826 2544 5102
rect 2608 5098 2636 6122
rect 2700 5914 2728 6394
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2596 5092 2648 5098
rect 2596 5034 2648 5040
rect 2504 4820 2556 4826
rect 2504 4762 2556 4768
rect 2226 4720 2282 4729
rect 2608 4690 2636 5034
rect 2226 4655 2228 4664
rect 2280 4655 2282 4664
rect 2596 4684 2648 4690
rect 2228 4626 2280 4632
rect 2596 4626 2648 4632
rect 2136 4616 2188 4622
rect 1858 4584 1914 4593
rect 2136 4558 2188 4564
rect 1858 4519 1914 4528
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1872 2774 1900 4519
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1964 3602 1992 4150
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 2240 2774 2268 4626
rect 2608 4146 2636 4626
rect 2596 4140 2648 4146
rect 2596 4082 2648 4088
rect 2318 3632 2374 3641
rect 2792 3602 2820 7239
rect 3056 6656 3108 6662
rect 2962 6624 3018 6633
rect 3056 6598 3108 6604
rect 2962 6559 3018 6568
rect 2976 6390 3004 6559
rect 2964 6384 3016 6390
rect 2964 6326 3016 6332
rect 2964 5636 3016 5642
rect 2964 5578 3016 5584
rect 2872 5568 2924 5574
rect 2872 5510 2924 5516
rect 2884 5166 2912 5510
rect 2872 5160 2924 5166
rect 2872 5102 2924 5108
rect 2976 4078 3004 5578
rect 3068 5370 3096 6598
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3054 5264 3110 5273
rect 3054 5199 3110 5208
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2870 3632 2926 3641
rect 2318 3567 2320 3576
rect 2372 3567 2374 3576
rect 2780 3596 2832 3602
rect 2320 3538 2372 3544
rect 2870 3567 2926 3576
rect 2780 3538 2832 3544
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2792 2961 2820 3130
rect 2778 2952 2834 2961
rect 2778 2887 2834 2896
rect 1872 2746 1992 2774
rect 1584 2644 1636 2650
rect 1584 2586 1636 2592
rect 1964 800 1992 2746
rect 2148 2746 2268 2774
rect 2148 1057 2176 2746
rect 2412 2100 2464 2106
rect 2412 2042 2464 2048
rect 2134 1048 2190 1057
rect 2134 983 2190 992
rect 2424 800 2452 2042
rect 2884 800 2912 3567
rect 2976 2854 3004 4014
rect 3068 3738 3096 5199
rect 3160 4457 3188 8774
rect 3344 8537 3372 9658
rect 3436 9382 3464 9998
rect 3516 9988 3568 9994
rect 3516 9930 3568 9936
rect 3528 9489 3556 9930
rect 3514 9480 3570 9489
rect 3514 9415 3570 9424
rect 3424 9376 3476 9382
rect 3424 9318 3476 9324
rect 3436 9042 3464 9318
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3424 9036 3476 9042
rect 3424 8978 3476 8984
rect 3422 8936 3478 8945
rect 3988 8922 4016 15982
rect 4160 15904 4212 15910
rect 4160 15846 4212 15852
rect 4066 15736 4122 15745
rect 4066 15671 4122 15680
rect 4080 15201 4108 15671
rect 4172 15337 4200 15846
rect 4356 15502 4384 16594
rect 4804 16108 4856 16114
rect 4804 16050 4856 16056
rect 4344 15496 4396 15502
rect 4344 15438 4396 15444
rect 4158 15328 4214 15337
rect 4158 15263 4214 15272
rect 4066 15192 4122 15201
rect 4066 15127 4122 15136
rect 4068 15020 4120 15026
rect 4068 14962 4120 14968
rect 4252 15020 4304 15026
rect 4252 14962 4304 14968
rect 4080 13734 4108 14962
rect 4264 14482 4292 14962
rect 4356 14958 4384 15438
rect 4816 14958 4844 16050
rect 4344 14952 4396 14958
rect 4344 14894 4396 14900
rect 4804 14952 4856 14958
rect 4804 14894 4856 14900
rect 4252 14476 4304 14482
rect 4252 14418 4304 14424
rect 4356 14464 4384 14894
rect 4528 14816 4580 14822
rect 4528 14758 4580 14764
rect 4436 14476 4488 14482
rect 4356 14436 4436 14464
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 4080 13530 4108 13670
rect 4068 13524 4120 13530
rect 4068 13466 4120 13472
rect 4068 12980 4120 12986
rect 4172 12968 4200 14214
rect 4252 13728 4304 13734
rect 4252 13670 4304 13676
rect 4264 13462 4292 13670
rect 4252 13456 4304 13462
rect 4252 13398 4304 13404
rect 4356 13258 4384 14436
rect 4436 14418 4488 14424
rect 4540 13297 4568 14758
rect 4712 14408 4764 14414
rect 4712 14350 4764 14356
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 4526 13288 4582 13297
rect 4344 13252 4396 13258
rect 4526 13223 4582 13232
rect 4344 13194 4396 13200
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4264 12986 4292 13126
rect 4120 12940 4200 12968
rect 4252 12980 4304 12986
rect 4068 12922 4120 12928
rect 4252 12922 4304 12928
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 4080 12374 4108 12786
rect 4068 12368 4120 12374
rect 4068 12310 4120 12316
rect 4356 12238 4384 13194
rect 4526 13016 4582 13025
rect 4436 12980 4488 12986
rect 4526 12951 4582 12960
rect 4436 12922 4488 12928
rect 4448 12889 4476 12922
rect 4540 12918 4568 12951
rect 4528 12912 4580 12918
rect 4434 12880 4490 12889
rect 4528 12854 4580 12860
rect 4434 12815 4490 12824
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4448 12442 4476 12718
rect 4436 12436 4488 12442
rect 4436 12378 4488 12384
rect 4434 12336 4490 12345
rect 4434 12271 4490 12280
rect 4344 12232 4396 12238
rect 4344 12174 4396 12180
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 4068 9920 4120 9926
rect 4068 9862 4120 9868
rect 4080 9602 4108 9862
rect 4080 9574 4200 9602
rect 3422 8871 3478 8880
rect 3896 8894 4016 8922
rect 3330 8528 3386 8537
rect 3240 8492 3292 8498
rect 3330 8463 3386 8472
rect 3240 8434 3292 8440
rect 3252 7342 3280 8434
rect 3436 8430 3464 8871
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8566 3832 8774
rect 3792 8560 3844 8566
rect 3792 8502 3844 8508
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3332 8288 3384 8294
rect 3332 8230 3384 8236
rect 3344 8072 3372 8230
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 3344 8044 3464 8072
rect 3436 7954 3464 8044
rect 3424 7948 3476 7954
rect 3424 7890 3476 7896
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 3240 7336 3292 7342
rect 3240 7278 3292 7284
rect 3238 7032 3294 7041
rect 3238 6967 3294 6976
rect 3252 6798 3280 6967
rect 3240 6792 3292 6798
rect 3240 6734 3292 6740
rect 3252 5386 3280 6734
rect 3344 5545 3372 7822
rect 3896 7410 3924 8894
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3988 8634 4016 8774
rect 3976 8628 4028 8634
rect 3976 8570 4028 8576
rect 4068 8628 4120 8634
rect 4068 8570 4120 8576
rect 4080 8514 4108 8570
rect 3988 8486 4108 8514
rect 3424 7404 3476 7410
rect 3424 7346 3476 7352
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3436 7177 3464 7346
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5574 3464 6258
rect 3804 6225 3832 6802
rect 3988 6662 4016 8486
rect 4068 8424 4120 8430
rect 4068 8366 4120 8372
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 4080 6390 4108 8366
rect 4172 8344 4200 9574
rect 4264 8945 4292 11834
rect 4356 11762 4384 12174
rect 4344 11756 4396 11762
rect 4344 11698 4396 11704
rect 4448 10742 4476 12271
rect 4540 12170 4568 12854
rect 4632 12186 4660 14282
rect 4724 13938 4752 14350
rect 4804 14272 4856 14278
rect 4804 14214 4856 14220
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4724 13841 4752 13874
rect 4710 13832 4766 13841
rect 4710 13767 4766 13776
rect 4712 13728 4764 13734
rect 4712 13670 4764 13676
rect 4724 12306 4752 13670
rect 4816 12345 4844 14214
rect 4908 14090 4936 17206
rect 5080 16040 5132 16046
rect 5080 15982 5132 15988
rect 4988 15904 5040 15910
rect 5092 15881 5120 15982
rect 4988 15846 5040 15852
rect 5078 15872 5134 15881
rect 5000 14249 5028 15846
rect 5078 15807 5134 15816
rect 5276 15706 5304 18022
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5172 15360 5224 15366
rect 5172 15302 5224 15308
rect 5184 15026 5212 15302
rect 5172 15020 5224 15026
rect 5172 14962 5224 14968
rect 5080 14272 5132 14278
rect 4986 14240 5042 14249
rect 5080 14214 5132 14220
rect 4986 14175 5042 14184
rect 4908 14062 5028 14090
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4802 12336 4858 12345
rect 4712 12300 4764 12306
rect 4802 12271 4858 12280
rect 4712 12242 4764 12248
rect 4528 12164 4580 12170
rect 4632 12158 4844 12186
rect 4528 12106 4580 12112
rect 4620 12096 4672 12102
rect 4620 12038 4672 12044
rect 4632 11234 4660 12038
rect 4540 11206 4660 11234
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4344 10192 4396 10198
rect 4344 10134 4396 10140
rect 4250 8936 4306 8945
rect 4250 8871 4306 8880
rect 4252 8356 4304 8362
rect 4172 8316 4252 8344
rect 4252 8298 4304 8304
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4172 7342 4200 7958
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3790 6216 3846 6225
rect 4172 6202 4200 6734
rect 3790 6151 3846 6160
rect 4080 6174 4200 6202
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3976 5908 4028 5914
rect 3976 5850 4028 5856
rect 3424 5568 3476 5574
rect 3330 5536 3386 5545
rect 3424 5510 3476 5516
rect 3330 5471 3386 5480
rect 3252 5358 3464 5386
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3344 5030 3372 5170
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3332 4548 3384 4554
rect 3332 4490 3384 4496
rect 3240 4480 3292 4486
rect 3146 4448 3202 4457
rect 3240 4422 3292 4428
rect 3146 4383 3202 4392
rect 3056 3732 3108 3738
rect 3056 3674 3108 3680
rect 3252 3618 3280 4422
rect 3344 4282 3372 4490
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 3252 3590 3372 3618
rect 3240 3528 3292 3534
rect 3240 3470 3292 3476
rect 2964 2848 3016 2854
rect 2964 2790 3016 2796
rect 2976 2514 3004 2790
rect 3252 2650 3280 3470
rect 3344 3398 3372 3590
rect 3332 3392 3384 3398
rect 3332 3334 3384 3340
rect 3330 2680 3386 2689
rect 3240 2644 3292 2650
rect 3330 2615 3386 2624
rect 3240 2586 3292 2592
rect 3054 2544 3110 2553
rect 2964 2508 3016 2514
rect 3054 2479 3110 2488
rect 2964 2450 3016 2456
rect 3068 2038 3096 2479
rect 3056 2032 3108 2038
rect 3056 1974 3108 1980
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1950 0 2006 800
rect 2410 0 2466 800
rect 2870 0 2926 800
rect 3252 241 3280 2586
rect 3344 800 3372 2615
rect 3436 2530 3464 5358
rect 3988 5234 4016 5850
rect 4080 5522 4108 6174
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4172 5642 4200 6054
rect 4160 5636 4212 5642
rect 4160 5578 4212 5584
rect 4080 5494 4200 5522
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3974 4856 4030 4865
rect 3884 4820 3936 4826
rect 3974 4791 4030 4800
rect 3884 4762 3936 4768
rect 3896 4214 3924 4762
rect 3988 4622 4016 4791
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4068 4480 4120 4486
rect 4068 4422 4120 4428
rect 3884 4208 3936 4214
rect 3936 4156 4016 4162
rect 3884 4150 4016 4156
rect 3896 4134 4016 4150
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3896 3738 3924 4014
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3792 3664 3844 3670
rect 3792 3606 3844 3612
rect 3804 3505 3832 3606
rect 3790 3496 3846 3505
rect 3790 3431 3846 3440
rect 3988 3194 4016 4134
rect 3976 3188 4028 3194
rect 3976 3130 4028 3136
rect 4080 2854 4108 4422
rect 4172 4049 4200 5494
rect 4158 4040 4214 4049
rect 4158 3975 4214 3984
rect 4264 3466 4292 8298
rect 4356 7546 4384 10134
rect 4436 9920 4488 9926
rect 4436 9862 4488 9868
rect 4448 9654 4476 9862
rect 4436 9648 4488 9654
rect 4436 9590 4488 9596
rect 4540 9042 4568 11206
rect 4712 10804 4764 10810
rect 4712 10746 4764 10752
rect 4724 10266 4752 10746
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4632 8974 4660 9522
rect 4724 9178 4752 9998
rect 4712 9172 4764 9178
rect 4712 9114 4764 9120
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4436 8424 4488 8430
rect 4436 8366 4488 8372
rect 4448 7886 4476 8366
rect 4632 8294 4660 8910
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4528 8016 4580 8022
rect 4528 7958 4580 7964
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4436 7744 4488 7750
rect 4436 7686 4488 7692
rect 4344 7540 4396 7546
rect 4344 7482 4396 7488
rect 4342 6624 4398 6633
rect 4342 6559 4398 6568
rect 4356 3913 4384 6559
rect 4448 5953 4476 7686
rect 4434 5944 4490 5953
rect 4434 5879 4490 5888
rect 4436 5228 4488 5234
rect 4436 5170 4488 5176
rect 4448 4826 4476 5170
rect 4436 4820 4488 4826
rect 4436 4762 4488 4768
rect 4540 4486 4568 7958
rect 4632 7818 4660 8230
rect 4724 7954 4752 8978
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4710 7848 4766 7857
rect 4620 7812 4672 7818
rect 4816 7834 4844 12158
rect 4908 8634 4936 13670
rect 5000 12102 5028 14062
rect 4988 12096 5040 12102
rect 4988 12038 5040 12044
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11150 5028 11698
rect 4988 11144 5040 11150
rect 4988 11086 5040 11092
rect 5092 10792 5120 14214
rect 5276 13530 5304 15642
rect 5356 14884 5408 14890
rect 5356 14826 5408 14832
rect 5264 13524 5316 13530
rect 5264 13466 5316 13472
rect 5276 12986 5304 13466
rect 5264 12980 5316 12986
rect 5264 12922 5316 12928
rect 5264 12776 5316 12782
rect 5264 12718 5316 12724
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5184 11898 5212 12378
rect 5276 12306 5304 12718
rect 5264 12300 5316 12306
rect 5264 12242 5316 12248
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5264 11008 5316 11014
rect 5264 10950 5316 10956
rect 5000 10764 5120 10792
rect 5000 9897 5028 10764
rect 5080 10668 5132 10674
rect 5080 10610 5132 10616
rect 5092 10266 5120 10610
rect 5172 10600 5224 10606
rect 5172 10542 5224 10548
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 4986 9888 5042 9897
rect 4986 9823 5042 9832
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4988 9512 5040 9518
rect 4988 9454 5040 9460
rect 5000 9110 5028 9454
rect 4988 9104 5040 9110
rect 4988 9046 5040 9052
rect 4986 8936 5042 8945
rect 4986 8871 5042 8880
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4908 8362 4936 8434
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4816 7806 4936 7834
rect 4710 7783 4766 7792
rect 4620 7754 4672 7760
rect 4632 6798 4660 7754
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4632 5710 4660 6734
rect 4724 6662 4752 7783
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4816 7546 4844 7686
rect 4804 7540 4856 7546
rect 4804 7482 4856 7488
rect 4712 6656 4764 6662
rect 4712 6598 4764 6604
rect 4802 6488 4858 6497
rect 4712 6452 4764 6458
rect 4802 6423 4858 6432
rect 4712 6394 4764 6400
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4528 4480 4580 4486
rect 4528 4422 4580 4428
rect 4632 4282 4660 5510
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4342 3904 4398 3913
rect 4342 3839 4398 3848
rect 4356 3602 4384 3839
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4252 3460 4304 3466
rect 4252 3402 4304 3408
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 3884 2644 3936 2650
rect 3884 2586 3936 2592
rect 3436 2502 3556 2530
rect 3422 2408 3478 2417
rect 3422 2343 3478 2352
rect 3436 2310 3464 2343
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3424 1352 3476 1358
rect 3424 1294 3476 1300
rect 3238 232 3294 241
rect 3238 167 3294 176
rect 3330 0 3386 800
rect 3436 649 3464 1294
rect 3528 762 3556 2502
rect 3896 2009 3924 2586
rect 4448 2446 4476 4150
rect 4618 3632 4674 3641
rect 4618 3567 4620 3576
rect 4672 3567 4674 3576
rect 4620 3538 4672 3544
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 4526 2544 4582 2553
rect 4526 2479 4582 2488
rect 4540 2446 4568 2479
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 3882 2000 3938 2009
rect 3882 1935 3938 1944
rect 4080 1601 4108 2246
rect 4066 1592 4122 1601
rect 4066 1527 4122 1536
rect 3712 870 3832 898
rect 3712 762 3740 870
rect 3804 800 3832 870
rect 4264 870 4384 898
rect 4264 800 4292 870
rect 3528 734 3740 762
rect 3422 640 3478 649
rect 3422 575 3478 584
rect 3790 0 3846 800
rect 4250 0 4306 800
rect 4356 762 4384 870
rect 4632 762 4660 3402
rect 4724 800 4752 6394
rect 4816 4690 4844 6423
rect 4908 6322 4936 7806
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 5000 6118 5028 8871
rect 5092 6458 5120 9522
rect 5184 8974 5212 10542
rect 5276 10266 5304 10950
rect 5264 10260 5316 10266
rect 5264 10202 5316 10208
rect 5264 10124 5316 10130
rect 5264 10066 5316 10072
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5172 7336 5224 7342
rect 5172 7278 5224 7284
rect 5184 6730 5212 7278
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4816 4214 4844 4626
rect 4896 4480 4948 4486
rect 4896 4422 4948 4428
rect 4804 4208 4856 4214
rect 4804 4150 4856 4156
rect 4908 4078 4936 4422
rect 4896 4072 4948 4078
rect 4896 4014 4948 4020
rect 4986 3496 5042 3505
rect 4986 3431 4988 3440
rect 5040 3431 5042 3440
rect 4988 3402 5040 3408
rect 5000 3233 5028 3402
rect 4986 3224 5042 3233
rect 4986 3159 5042 3168
rect 5092 800 5120 6258
rect 5184 6186 5212 6666
rect 5276 6254 5304 10066
rect 5368 9994 5396 14826
rect 5460 12481 5488 18566
rect 5552 17542 5580 18686
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 6000 17808 6052 17814
rect 6000 17750 6052 17756
rect 5540 17536 5592 17542
rect 5540 17478 5592 17484
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5552 17270 5580 17478
rect 5540 17264 5592 17270
rect 5540 17206 5592 17212
rect 5816 17128 5868 17134
rect 5816 17070 5868 17076
rect 5828 16794 5856 17070
rect 5920 17066 5948 17478
rect 6012 17338 6040 17750
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6564 17354 6592 20334
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9404 19780 9456 19786
rect 9404 19722 9456 19728
rect 7748 19712 7800 19718
rect 7748 19654 7800 19660
rect 8392 19712 8444 19718
rect 8392 19654 8444 19660
rect 7760 19514 7788 19654
rect 7748 19508 7800 19514
rect 7748 19450 7800 19456
rect 7840 19372 7892 19378
rect 7840 19314 7892 19320
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 6644 18692 6696 18698
rect 6644 18634 6696 18640
rect 6656 18358 6684 18634
rect 7012 18624 7064 18630
rect 7012 18566 7064 18572
rect 6644 18352 6696 18358
rect 6644 18294 6696 18300
rect 6736 17604 6788 17610
rect 6736 17546 6788 17552
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6000 17332 6052 17338
rect 6564 17326 6684 17354
rect 6748 17338 6776 17546
rect 6000 17274 6052 17280
rect 5908 17060 5960 17066
rect 5908 17002 5960 17008
rect 5816 16788 5868 16794
rect 5816 16730 5868 16736
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5538 16008 5594 16017
rect 5538 15943 5540 15952
rect 5592 15943 5594 15952
rect 5540 15914 5592 15920
rect 5644 14464 5672 16594
rect 5828 16590 5856 16730
rect 5816 16584 5868 16590
rect 5816 16526 5868 16532
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5736 15162 5764 16458
rect 6012 16402 6040 17274
rect 6092 17264 6144 17270
rect 6092 17206 6144 17212
rect 6104 16998 6132 17206
rect 6552 17196 6604 17202
rect 6552 17138 6604 17144
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 5828 16374 6040 16402
rect 5724 15156 5776 15162
rect 5724 15098 5776 15104
rect 5828 15042 5856 16374
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 5908 15360 5960 15366
rect 5908 15302 5960 15308
rect 5552 14436 5672 14464
rect 5736 15014 5856 15042
rect 5446 12472 5502 12481
rect 5446 12407 5502 12416
rect 5446 11928 5502 11937
rect 5446 11863 5502 11872
rect 5356 9988 5408 9994
rect 5356 9930 5408 9936
rect 5356 9376 5408 9382
rect 5356 9318 5408 9324
rect 5368 8974 5396 9318
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5368 8362 5396 8910
rect 5356 8356 5408 8362
rect 5356 8298 5408 8304
rect 5460 7018 5488 11863
rect 5552 11014 5580 14436
rect 5736 12345 5764 15014
rect 5920 13802 5948 15302
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6000 15020 6052 15026
rect 6000 14962 6052 14968
rect 6012 14074 6040 14962
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6000 13932 6052 13938
rect 6000 13874 6052 13880
rect 5908 13796 5960 13802
rect 5908 13738 5960 13744
rect 6012 12986 6040 13874
rect 6460 13864 6512 13870
rect 6458 13832 6460 13841
rect 6512 13832 6514 13841
rect 6458 13767 6514 13776
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 6000 12980 6052 12986
rect 6000 12922 6052 12928
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12374 5948 12582
rect 5908 12368 5960 12374
rect 5722 12336 5778 12345
rect 5632 12300 5684 12306
rect 5908 12310 5960 12316
rect 6012 12306 6040 12718
rect 5722 12271 5778 12280
rect 6000 12300 6052 12306
rect 5632 12242 5684 12248
rect 6000 12242 6052 12248
rect 5644 11898 5672 12242
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10062 5580 10950
rect 5630 10568 5686 10577
rect 5630 10503 5686 10512
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5644 8072 5672 10503
rect 5736 8838 5764 12174
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5828 11694 5856 12038
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 5828 11506 5856 11630
rect 5908 11552 5960 11558
rect 5828 11500 5908 11506
rect 5828 11494 5960 11500
rect 5828 11478 5948 11494
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5644 8044 5764 8072
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5540 7336 5592 7342
rect 5540 7278 5592 7284
rect 5368 7002 5488 7018
rect 5356 6996 5488 7002
rect 5408 6990 5488 6996
rect 5356 6938 5408 6944
rect 5356 6656 5408 6662
rect 5356 6598 5408 6604
rect 5264 6248 5316 6254
rect 5264 6190 5316 6196
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5184 5914 5212 6122
rect 5172 5908 5224 5914
rect 5172 5850 5224 5856
rect 5264 5772 5316 5778
rect 5264 5714 5316 5720
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5184 4214 5212 4422
rect 5172 4208 5224 4214
rect 5172 4150 5224 4156
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5184 3126 5212 4014
rect 5172 3120 5224 3126
rect 5172 3062 5224 3068
rect 5276 2106 5304 5714
rect 5368 5642 5396 6598
rect 5446 6488 5502 6497
rect 5552 6458 5580 7278
rect 5644 6934 5672 7890
rect 5632 6928 5684 6934
rect 5632 6870 5684 6876
rect 5736 6866 5764 8044
rect 5724 6860 5776 6866
rect 5724 6802 5776 6808
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5446 6423 5502 6432
rect 5540 6452 5592 6458
rect 5460 6304 5488 6423
rect 5540 6394 5592 6400
rect 5540 6316 5592 6322
rect 5460 6276 5540 6304
rect 5540 6258 5592 6264
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5448 5704 5500 5710
rect 5448 5646 5500 5652
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 5368 2514 5396 4966
rect 5460 3942 5488 5646
rect 5448 3936 5500 3942
rect 5448 3878 5500 3884
rect 5446 3360 5502 3369
rect 5446 3295 5502 3304
rect 5460 2514 5488 3295
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5448 2508 5500 2514
rect 5448 2450 5500 2456
rect 5264 2100 5316 2106
rect 5264 2042 5316 2048
rect 5552 800 5580 6054
rect 5644 2106 5672 6666
rect 5736 6440 5764 6802
rect 5828 6730 5856 11478
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5920 10810 5948 10950
rect 5908 10804 5960 10810
rect 5908 10746 5960 10752
rect 6012 10674 6040 11154
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6000 10668 6052 10674
rect 6000 10610 6052 10616
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 9586 5948 10406
rect 6012 10130 6040 10610
rect 6000 10124 6052 10130
rect 6000 10066 6052 10072
rect 5998 9888 6054 9897
rect 5998 9823 6054 9832
rect 5908 9580 5960 9586
rect 5908 9522 5960 9528
rect 5908 7812 5960 7818
rect 5908 7754 5960 7760
rect 5920 7342 5948 7754
rect 5908 7336 5960 7342
rect 5908 7278 5960 7284
rect 5908 7200 5960 7206
rect 5908 7142 5960 7148
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 5920 6662 5948 7142
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5736 6412 5856 6440
rect 5724 5840 5776 5846
rect 5722 5808 5724 5817
rect 5776 5808 5778 5817
rect 5722 5743 5778 5752
rect 5828 5624 5856 6412
rect 6012 5930 6040 9823
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6564 9450 6592 17138
rect 6656 14278 6684 17326
rect 6736 17332 6788 17338
rect 6736 17274 6788 17280
rect 6932 16590 6960 17546
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 6736 16040 6788 16046
rect 6736 15982 6788 15988
rect 6644 14272 6696 14278
rect 6644 14214 6696 14220
rect 6656 14074 6684 14214
rect 6644 14068 6696 14074
rect 6644 14010 6696 14016
rect 6644 13932 6696 13938
rect 6644 13874 6696 13880
rect 6656 12458 6684 13874
rect 6748 13870 6776 15982
rect 7024 15434 7052 18566
rect 7208 17678 7236 18702
rect 7746 18184 7802 18193
rect 7746 18119 7802 18128
rect 7760 17882 7788 18119
rect 7748 17876 7800 17882
rect 7748 17818 7800 17824
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 15910 7144 16390
rect 7104 15904 7156 15910
rect 7104 15846 7156 15852
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 7012 15428 7064 15434
rect 7012 15370 7064 15376
rect 6932 14618 6960 15370
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6828 14340 6880 14346
rect 6828 14282 6880 14288
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 6748 13705 6776 13806
rect 6840 13802 6868 14282
rect 7024 14090 7052 15370
rect 7116 15348 7144 15846
rect 7208 15502 7236 17614
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7288 17196 7340 17202
rect 7288 17138 7340 17144
rect 7300 16794 7328 17138
rect 7380 17128 7432 17134
rect 7380 17070 7432 17076
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7392 16130 7420 17070
rect 7484 16697 7512 17478
rect 7656 16720 7708 16726
rect 7470 16688 7526 16697
rect 7656 16662 7708 16668
rect 7470 16623 7526 16632
rect 7564 16176 7616 16182
rect 7392 16102 7512 16130
rect 7564 16118 7616 16124
rect 7380 15972 7432 15978
rect 7380 15914 7432 15920
rect 7286 15736 7342 15745
rect 7286 15671 7288 15680
rect 7340 15671 7342 15680
rect 7288 15642 7340 15648
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7116 15320 7236 15348
rect 7024 14062 7144 14090
rect 7116 13802 7144 14062
rect 6828 13796 6880 13802
rect 6828 13738 6880 13744
rect 7104 13796 7156 13802
rect 7104 13738 7156 13744
rect 6734 13696 6790 13705
rect 6734 13631 6790 13640
rect 6840 13462 6868 13738
rect 6828 13456 6880 13462
rect 6828 13398 6880 13404
rect 7116 12782 7144 13738
rect 7208 13258 7236 15320
rect 7288 15020 7340 15026
rect 7288 14962 7340 14968
rect 7300 13530 7328 14962
rect 7288 13524 7340 13530
rect 7288 13466 7340 13472
rect 7196 13252 7248 13258
rect 7196 13194 7248 13200
rect 7288 13184 7340 13190
rect 7288 13126 7340 13132
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6656 12430 6776 12458
rect 6644 12368 6696 12374
rect 6644 12310 6696 12316
rect 6656 11898 6684 12310
rect 6748 11898 6776 12430
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 6736 11076 6788 11082
rect 6736 11018 6788 11024
rect 6644 11008 6696 11014
rect 6644 10950 6696 10956
rect 6656 10266 6684 10950
rect 6748 10810 6776 11018
rect 6736 10804 6788 10810
rect 6736 10746 6788 10752
rect 6644 10260 6696 10266
rect 6644 10202 6696 10208
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6552 9444 6604 9450
rect 6552 9386 6604 9392
rect 6656 9382 6684 10066
rect 6840 9926 6868 12718
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6932 11778 6960 12038
rect 6932 11762 7052 11778
rect 6932 11756 7064 11762
rect 6932 11750 7012 11756
rect 7012 11698 7064 11704
rect 6920 11688 6972 11694
rect 6920 11630 6972 11636
rect 6932 10810 6960 11630
rect 6920 10804 6972 10810
rect 6920 10746 6972 10752
rect 6736 9920 6788 9926
rect 6736 9862 6788 9868
rect 6828 9920 6880 9926
rect 6828 9862 6880 9868
rect 6748 9450 6776 9862
rect 6840 9722 6868 9862
rect 6828 9716 6880 9722
rect 6828 9658 6880 9664
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6644 9376 6696 9382
rect 6644 9318 6696 9324
rect 6656 9178 6684 9318
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6552 9104 6604 9110
rect 6552 9046 6604 9052
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6368 8492 6420 8498
rect 6564 8480 6592 9046
rect 6932 8838 6960 9590
rect 7024 9586 7052 11698
rect 7116 11694 7144 12718
rect 7300 12594 7328 13126
rect 7392 12918 7420 15914
rect 7484 13705 7512 16102
rect 7576 14822 7604 16118
rect 7564 14816 7616 14822
rect 7564 14758 7616 14764
rect 7470 13696 7526 13705
rect 7470 13631 7526 13640
rect 7472 13252 7524 13258
rect 7472 13194 7524 13200
rect 7380 12912 7432 12918
rect 7380 12854 7432 12860
rect 7208 12566 7328 12594
rect 7208 12306 7236 12566
rect 7288 12436 7340 12442
rect 7288 12378 7340 12384
rect 7196 12300 7248 12306
rect 7196 12242 7248 12248
rect 7300 12102 7328 12378
rect 7288 12096 7340 12102
rect 7288 12038 7340 12044
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7104 11144 7156 11150
rect 7392 11121 7420 12854
rect 7104 11086 7156 11092
rect 7378 11112 7434 11121
rect 7116 10713 7144 11086
rect 7288 11076 7340 11082
rect 7378 11047 7434 11056
rect 7288 11018 7340 11024
rect 7102 10704 7158 10713
rect 7158 10662 7236 10690
rect 7102 10639 7158 10648
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6420 8452 6592 8480
rect 6644 8492 6696 8498
rect 6368 8434 6420 8440
rect 6644 8434 6696 8440
rect 6380 8265 6408 8434
rect 6656 8378 6684 8434
rect 6564 8350 6684 8378
rect 6366 8256 6422 8265
rect 6366 8191 6422 8200
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 6184 6384 6236 6390
rect 6090 6352 6146 6361
rect 6184 6326 6236 6332
rect 6090 6287 6146 6296
rect 6104 6254 6132 6287
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6196 6089 6224 6326
rect 6276 6248 6328 6254
rect 6276 6190 6328 6196
rect 6288 6118 6316 6190
rect 6276 6112 6328 6118
rect 6182 6080 6238 6089
rect 6276 6054 6328 6060
rect 6182 6015 6238 6024
rect 5920 5902 6040 5930
rect 5920 5710 5948 5902
rect 6000 5840 6052 5846
rect 6000 5782 6052 5788
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5736 5596 5856 5624
rect 5736 5273 5764 5596
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5816 5296 5868 5302
rect 5722 5264 5778 5273
rect 5816 5238 5868 5244
rect 5722 5199 5778 5208
rect 5724 5092 5776 5098
rect 5724 5034 5776 5040
rect 5736 4146 5764 5034
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5724 3596 5776 3602
rect 5724 3538 5776 3544
rect 5736 3058 5764 3538
rect 5828 3534 5856 5238
rect 5920 4758 5948 5306
rect 6012 5234 6040 5782
rect 6196 5642 6224 6015
rect 6564 5658 6592 8350
rect 6736 6656 6788 6662
rect 6736 6598 6788 6604
rect 6644 6248 6696 6254
rect 6642 6216 6644 6225
rect 6696 6216 6698 6225
rect 6642 6151 6698 6160
rect 6748 6118 6776 6598
rect 6840 6440 6868 8774
rect 6932 8566 6960 8774
rect 6920 8560 6972 8566
rect 6920 8502 6972 8508
rect 7024 7313 7052 9522
rect 7104 8968 7156 8974
rect 7104 8910 7156 8916
rect 7116 8634 7144 8910
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 7208 7698 7236 10662
rect 7300 10606 7328 11018
rect 7484 10810 7512 13194
rect 7472 10804 7524 10810
rect 7472 10746 7524 10752
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7300 10130 7328 10542
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7392 9674 7420 10542
rect 7484 10538 7512 10746
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7576 9738 7604 14758
rect 7668 13870 7696 16662
rect 7852 16454 7880 19314
rect 8404 18970 8432 19654
rect 9416 19514 9444 19722
rect 9404 19508 9456 19514
rect 9404 19450 9456 19456
rect 8668 19372 8720 19378
rect 8668 19314 8720 19320
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8680 18834 8708 19314
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 8668 18828 8720 18834
rect 8668 18770 8720 18776
rect 8668 18692 8720 18698
rect 8668 18634 8720 18640
rect 8680 18222 8708 18634
rect 9312 18624 9364 18630
rect 9312 18566 9364 18572
rect 9404 18624 9456 18630
rect 9404 18566 9456 18572
rect 8668 18216 8720 18222
rect 8668 18158 8720 18164
rect 8392 17672 8444 17678
rect 8392 17614 8444 17620
rect 8116 17604 8168 17610
rect 8116 17546 8168 17552
rect 8128 17134 8156 17546
rect 8116 17128 8168 17134
rect 8116 17070 8168 17076
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 8208 16040 8260 16046
rect 8208 15982 8260 15988
rect 7932 15496 7984 15502
rect 7932 15438 7984 15444
rect 7840 14952 7892 14958
rect 7944 14906 7972 15438
rect 7892 14900 7972 14906
rect 7840 14894 7972 14900
rect 7852 14878 7972 14894
rect 7944 14618 7972 14878
rect 7932 14612 7984 14618
rect 7932 14554 7984 14560
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7748 13728 7800 13734
rect 7748 13670 7800 13676
rect 7760 13394 7788 13670
rect 7748 13388 7800 13394
rect 7748 13330 7800 13336
rect 7748 13184 7800 13190
rect 7748 13126 7800 13132
rect 7760 12986 7788 13126
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7932 12844 7984 12850
rect 7932 12786 7984 12792
rect 7656 12776 7708 12782
rect 7656 12718 7708 12724
rect 7668 12238 7696 12718
rect 7944 12434 7972 12786
rect 7760 12406 7972 12434
rect 7760 12374 7788 12406
rect 7748 12368 7800 12374
rect 7748 12310 7800 12316
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7116 7670 7236 7698
rect 7300 9646 7420 9674
rect 7484 9710 7604 9738
rect 7010 7304 7066 7313
rect 7010 7239 7066 7248
rect 7012 7200 7064 7206
rect 7012 7142 7064 7148
rect 7024 6866 7052 7142
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7116 6746 7144 7670
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7208 6798 7236 7482
rect 7024 6718 7144 6746
rect 7196 6792 7248 6798
rect 7196 6734 7248 6740
rect 6920 6452 6972 6458
rect 6840 6412 6920 6440
rect 6920 6394 6972 6400
rect 6828 6180 6880 6186
rect 6828 6122 6880 6128
rect 6644 6112 6696 6118
rect 6644 6054 6696 6060
rect 6736 6112 6788 6118
rect 6736 6054 6788 6060
rect 6656 5778 6684 6054
rect 6748 5914 6776 6054
rect 6736 5908 6788 5914
rect 6736 5850 6788 5856
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 6184 5636 6236 5642
rect 6564 5630 6684 5658
rect 6184 5578 6236 5584
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 6458 5264 6514 5273
rect 6000 5228 6052 5234
rect 6458 5199 6460 5208
rect 6000 5170 6052 5176
rect 6512 5199 6514 5208
rect 6460 5170 6512 5176
rect 5908 4752 5960 4758
rect 5908 4694 5960 4700
rect 6012 3534 6040 5170
rect 6552 4684 6604 4690
rect 6552 4626 6604 4632
rect 6148 4380 6456 4400
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 6092 4140 6144 4146
rect 6092 4082 6144 4088
rect 6104 3602 6132 4082
rect 6564 4078 6592 4626
rect 6656 4214 6684 5630
rect 6736 5568 6788 5574
rect 6736 5510 6788 5516
rect 6748 5370 6776 5510
rect 6736 5364 6788 5370
rect 6736 5306 6788 5312
rect 6840 5098 6868 6122
rect 6918 5944 6974 5953
rect 6918 5879 6974 5888
rect 6932 5846 6960 5879
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6920 5568 6972 5574
rect 6920 5510 6972 5516
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 6828 4820 6880 4826
rect 6828 4762 6880 4768
rect 6736 4684 6788 4690
rect 6736 4626 6788 4632
rect 6644 4208 6696 4214
rect 6644 4150 6696 4156
rect 6552 4072 6604 4078
rect 6552 4014 6604 4020
rect 6184 3936 6236 3942
rect 6184 3878 6236 3884
rect 6196 3670 6224 3878
rect 6564 3754 6592 4014
rect 6564 3726 6684 3754
rect 6184 3664 6236 3670
rect 6184 3606 6236 3612
rect 6092 3596 6144 3602
rect 6092 3538 6144 3544
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 6000 2984 6052 2990
rect 6000 2926 6052 2932
rect 5632 2100 5684 2106
rect 5632 2042 5684 2048
rect 6012 800 6040 2926
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 6564 1986 6592 3470
rect 6656 2650 6684 3726
rect 6644 2644 6696 2650
rect 6644 2586 6696 2592
rect 6748 2446 6776 4626
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6840 2310 6868 4762
rect 6932 3942 6960 5510
rect 7024 4740 7052 6718
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7116 5914 7144 6598
rect 7196 6316 7248 6322
rect 7196 6258 7248 6264
rect 7104 5908 7156 5914
rect 7104 5850 7156 5856
rect 7024 4712 7144 4740
rect 7012 4616 7064 4622
rect 7010 4584 7012 4593
rect 7064 4584 7066 4593
rect 7010 4519 7066 4528
rect 7116 4486 7144 4712
rect 7104 4480 7156 4486
rect 7104 4422 7156 4428
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 7012 3936 7064 3942
rect 7012 3878 7064 3884
rect 6920 3664 6972 3670
rect 6920 3606 6972 3612
rect 6932 3194 6960 3606
rect 7024 3602 7052 3878
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6918 3088 6974 3097
rect 7116 3058 7144 3674
rect 6918 3023 6920 3032
rect 6972 3023 6974 3032
rect 7104 3052 7156 3058
rect 6920 2994 6972 3000
rect 7104 2994 7156 3000
rect 6918 2952 6974 2961
rect 6918 2887 6974 2896
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6472 1958 6592 1986
rect 6472 800 6500 1958
rect 6932 800 6960 2887
rect 7208 1358 7236 6258
rect 7300 5778 7328 9646
rect 7380 9512 7432 9518
rect 7378 9480 7380 9489
rect 7432 9480 7434 9489
rect 7378 9415 7434 9424
rect 7484 8498 7512 9710
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 8974 7604 9522
rect 7564 8968 7616 8974
rect 7564 8910 7616 8916
rect 7668 8514 7696 10746
rect 7760 9058 7788 12310
rect 7840 12232 7892 12238
rect 7840 12174 7892 12180
rect 7852 11694 7880 12174
rect 7932 11892 7984 11898
rect 7932 11834 7984 11840
rect 7840 11688 7892 11694
rect 7840 11630 7892 11636
rect 7944 11558 7972 11834
rect 8036 11744 8064 15982
rect 8116 14612 8168 14618
rect 8116 14554 8168 14560
rect 8128 14278 8156 14554
rect 8116 14272 8168 14278
rect 8116 14214 8168 14220
rect 8220 13977 8248 15982
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8312 14074 8340 14418
rect 8404 14074 8432 17614
rect 8576 17128 8628 17134
rect 8576 17070 8628 17076
rect 8588 16794 8616 17070
rect 8680 17066 8708 18158
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 9324 17338 9352 18566
rect 9416 18426 9444 18566
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 9508 17678 9536 19790
rect 9588 17876 9640 17882
rect 9588 17818 9640 17824
rect 9496 17672 9548 17678
rect 9496 17614 9548 17620
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 8668 17060 8720 17066
rect 8668 17002 8720 17008
rect 8680 16794 8708 17002
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 8576 16788 8628 16794
rect 8576 16730 8628 16736
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8680 16658 8708 16730
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 9508 16590 9536 17614
rect 9600 17134 9628 17818
rect 9588 17128 9640 17134
rect 9586 17096 9588 17105
rect 9640 17096 9642 17105
rect 9586 17031 9642 17040
rect 9496 16584 9548 16590
rect 9496 16526 9548 16532
rect 9126 16144 9182 16153
rect 9126 16079 9128 16088
rect 9180 16079 9182 16088
rect 9128 16050 9180 16056
rect 8484 15904 8536 15910
rect 8484 15846 8536 15852
rect 9496 15904 9548 15910
rect 9496 15846 9548 15852
rect 9864 15904 9916 15910
rect 9864 15846 9916 15852
rect 8300 14068 8352 14074
rect 8300 14010 8352 14016
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8206 13968 8262 13977
rect 8206 13903 8262 13912
rect 8312 13870 8340 14010
rect 8300 13864 8352 13870
rect 8300 13806 8352 13812
rect 8116 13796 8168 13802
rect 8116 13738 8168 13744
rect 8128 11898 8156 13738
rect 8496 13410 8524 15846
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 8668 15632 8720 15638
rect 9508 15609 9536 15846
rect 9680 15700 9732 15706
rect 9680 15642 9732 15648
rect 8668 15574 8720 15580
rect 9494 15600 9550 15609
rect 8680 15366 8708 15574
rect 9494 15535 9550 15544
rect 9588 15496 9640 15502
rect 9310 15464 9366 15473
rect 9692 15473 9720 15642
rect 9588 15438 9640 15444
rect 9678 15464 9734 15473
rect 9310 15399 9312 15408
rect 9364 15399 9366 15408
rect 9312 15370 9364 15376
rect 8576 15360 8628 15366
rect 8576 15302 8628 15308
rect 8668 15360 8720 15366
rect 8668 15302 8720 15308
rect 8588 15094 8616 15302
rect 8576 15088 8628 15094
rect 8576 15030 8628 15036
rect 8680 14906 8708 15302
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9220 15020 9272 15026
rect 9220 14962 9272 14968
rect 8220 13382 8524 13410
rect 8588 14878 8708 14906
rect 8220 11937 8248 13382
rect 8300 13320 8352 13326
rect 8300 13262 8352 13268
rect 8312 12918 8340 13262
rect 8300 12912 8352 12918
rect 8300 12854 8352 12860
rect 8206 11928 8262 11937
rect 8116 11892 8168 11898
rect 8206 11863 8262 11872
rect 8116 11834 8168 11840
rect 8036 11716 8248 11744
rect 8116 11620 8168 11626
rect 8116 11562 8168 11568
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 10577 8064 11494
rect 8022 10568 8078 10577
rect 8022 10503 8078 10512
rect 8128 10198 8156 11562
rect 8116 10192 8168 10198
rect 8116 10134 8168 10140
rect 8024 9988 8076 9994
rect 8024 9930 8076 9936
rect 7840 9920 7892 9926
rect 7840 9862 7892 9868
rect 7932 9920 7984 9926
rect 7932 9862 7984 9868
rect 7852 9178 7880 9862
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7760 9030 7880 9058
rect 7472 8492 7524 8498
rect 7472 8434 7524 8440
rect 7576 8486 7696 8514
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7380 6656 7432 6662
rect 7380 6598 7432 6604
rect 7288 5772 7340 5778
rect 7288 5714 7340 5720
rect 7286 5672 7342 5681
rect 7286 5607 7342 5616
rect 7300 3942 7328 5607
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 7288 3664 7340 3670
rect 7288 3606 7340 3612
rect 7300 2774 7328 3606
rect 7392 2922 7420 6598
rect 7484 5846 7512 7414
rect 7472 5840 7524 5846
rect 7472 5782 7524 5788
rect 7576 5710 7604 8486
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 7564 5704 7616 5710
rect 7470 5672 7526 5681
rect 7564 5646 7616 5652
rect 7470 5607 7526 5616
rect 7484 3194 7512 5607
rect 7562 4720 7618 4729
rect 7562 4655 7618 4664
rect 7576 4622 7604 4655
rect 7564 4616 7616 4622
rect 7564 4558 7616 4564
rect 7472 3188 7524 3194
rect 7472 3130 7524 3136
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 7300 2746 7420 2774
rect 7196 1352 7248 1358
rect 7196 1294 7248 1300
rect 7392 800 7420 2746
rect 7576 2038 7604 4558
rect 7668 3534 7696 8026
rect 7748 7880 7800 7886
rect 7748 7822 7800 7828
rect 7760 7206 7788 7822
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6390 7788 6598
rect 7852 6458 7880 9030
rect 7944 8634 7972 9862
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7852 5370 7880 5510
rect 7840 5364 7892 5370
rect 7840 5306 7892 5312
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7760 4049 7788 4082
rect 7746 4040 7802 4049
rect 7746 3975 7802 3984
rect 7760 3670 7788 3975
rect 7748 3664 7800 3670
rect 7748 3606 7800 3612
rect 7944 3618 7972 7958
rect 8036 6322 8064 9930
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 8498 8156 8774
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 8128 8090 8156 8434
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8220 6746 8248 11716
rect 8312 7818 8340 12854
rect 8392 12708 8444 12714
rect 8392 12650 8444 12656
rect 8404 9926 8432 12650
rect 8484 12640 8536 12646
rect 8484 12582 8536 12588
rect 8496 12238 8524 12582
rect 8484 12232 8536 12238
rect 8484 12174 8536 12180
rect 8496 11218 8524 12174
rect 8588 11778 8616 14878
rect 9128 14816 9180 14822
rect 9128 14758 9180 14764
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 9140 14414 9168 14758
rect 9128 14408 9180 14414
rect 9128 14350 9180 14356
rect 8944 13932 8996 13938
rect 8680 13892 8944 13920
rect 8680 11898 8708 13892
rect 8944 13874 8996 13880
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 9140 12646 9168 14350
rect 9232 14226 9260 14962
rect 9508 14346 9536 15098
rect 9600 14822 9628 15438
rect 9678 15399 9734 15408
rect 9876 15337 9904 15846
rect 9862 15328 9918 15337
rect 9862 15263 9918 15272
rect 9588 14816 9640 14822
rect 9588 14758 9640 14764
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 9232 14198 9352 14226
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 9232 13530 9260 13738
rect 9220 13524 9272 13530
rect 9220 13466 9272 13472
rect 9220 12776 9272 12782
rect 9220 12718 9272 12724
rect 9128 12640 9180 12646
rect 9128 12582 9180 12588
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 9126 12472 9182 12481
rect 9048 12416 9126 12424
rect 9048 12407 9182 12416
rect 9048 12396 9168 12407
rect 8852 12368 8904 12374
rect 8852 12310 8904 12316
rect 8760 12096 8812 12102
rect 8760 12038 8812 12044
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8772 11830 8800 12038
rect 8760 11824 8812 11830
rect 8588 11750 8708 11778
rect 8760 11766 8812 11772
rect 8576 11688 8628 11694
rect 8576 11630 8628 11636
rect 8484 11212 8536 11218
rect 8484 11154 8536 11160
rect 8588 10810 8616 11630
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8484 10532 8536 10538
rect 8484 10474 8536 10480
rect 8392 9920 8444 9926
rect 8392 9862 8444 9868
rect 8496 9489 8524 10474
rect 8680 10266 8708 11750
rect 8864 11665 8892 12310
rect 8944 12096 8996 12102
rect 8942 12064 8944 12073
rect 8996 12064 8998 12073
rect 8942 11999 8998 12008
rect 9048 11694 9076 12396
rect 9232 12374 9260 12718
rect 9220 12368 9272 12374
rect 9126 12336 9182 12345
rect 9220 12310 9272 12316
rect 9126 12271 9182 12280
rect 9036 11688 9088 11694
rect 8850 11656 8906 11665
rect 9036 11630 9088 11636
rect 8850 11591 8906 11600
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 8668 10260 8720 10266
rect 8668 10202 8720 10208
rect 8944 9988 8996 9994
rect 8944 9930 8996 9936
rect 8956 9722 8984 9930
rect 8944 9716 8996 9722
rect 8944 9658 8996 9664
rect 8482 9480 8538 9489
rect 8482 9415 8538 9424
rect 8392 8288 8444 8294
rect 8392 8230 8444 8236
rect 8404 7886 8432 8230
rect 8496 8022 8524 9415
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 8576 8832 8628 8838
rect 8576 8774 8628 8780
rect 8484 8016 8536 8022
rect 8484 7958 8536 7964
rect 8392 7880 8444 7886
rect 8392 7822 8444 7828
rect 8300 7812 8352 7818
rect 8300 7754 8352 7760
rect 8484 7812 8536 7818
rect 8484 7754 8536 7760
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8404 7478 8432 7686
rect 8392 7472 8444 7478
rect 8392 7414 8444 7420
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8128 6718 8248 6746
rect 8024 6316 8076 6322
rect 8024 6258 8076 6264
rect 8128 5930 8156 6718
rect 8208 6656 8260 6662
rect 8208 6598 8260 6604
rect 8036 5902 8156 5930
rect 8220 5914 8248 6598
rect 8208 5908 8260 5914
rect 8036 3738 8064 5902
rect 8208 5850 8260 5856
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 8128 4185 8156 5646
rect 8312 5030 8340 7142
rect 8392 5704 8444 5710
rect 8392 5646 8444 5652
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8114 4176 8170 4185
rect 8114 4111 8170 4120
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 8208 3936 8260 3942
rect 8208 3878 8260 3884
rect 8024 3732 8076 3738
rect 8024 3674 8076 3680
rect 7944 3590 8064 3618
rect 8128 3602 8156 3878
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7932 3392 7984 3398
rect 7838 3360 7894 3369
rect 7932 3334 7984 3340
rect 7838 3295 7894 3304
rect 7852 3058 7880 3295
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 2514 7788 2926
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7852 800 7880 2994
rect 7944 2514 7972 3334
rect 8036 2650 8064 3590
rect 8116 3596 8168 3602
rect 8116 3538 8168 3544
rect 8116 3392 8168 3398
rect 8220 3380 8248 3878
rect 8312 3534 8340 4966
rect 8404 4826 8432 5646
rect 8496 5302 8524 7754
rect 8588 6390 8616 8774
rect 8668 8356 8720 8362
rect 8668 8298 8720 8304
rect 8576 6384 8628 6390
rect 8576 6326 8628 6332
rect 8484 5296 8536 5302
rect 8484 5238 8536 5244
rect 8392 4820 8444 4826
rect 8392 4762 8444 4768
rect 8392 4480 8444 4486
rect 8392 4422 8444 4428
rect 8300 3528 8352 3534
rect 8300 3470 8352 3476
rect 8168 3352 8248 3380
rect 8116 3334 8168 3340
rect 8312 3126 8340 3470
rect 8404 3466 8432 4422
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8496 3913 8524 4014
rect 8482 3904 8538 3913
rect 8482 3839 8538 3848
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8496 2961 8524 3839
rect 8482 2952 8538 2961
rect 8482 2887 8538 2896
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8312 870 8432 898
rect 8312 800 8340 870
rect 4356 734 4660 762
rect 4710 0 4766 800
rect 5078 0 5134 800
rect 5538 0 5594 800
rect 5998 0 6054 800
rect 6458 0 6514 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 8404 762 8432 870
rect 8588 762 8616 6326
rect 8680 4282 8708 8298
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 9140 7342 9168 12271
rect 9232 11218 9260 12310
rect 9220 11212 9272 11218
rect 9220 11154 9272 11160
rect 9220 10464 9272 10470
rect 9220 10406 9272 10412
rect 9232 10266 9260 10406
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9128 7336 9180 7342
rect 9128 7278 9180 7284
rect 8747 7100 9055 7120
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 8852 6656 8904 6662
rect 8852 6598 8904 6604
rect 8864 6458 8892 6598
rect 9140 6458 9168 7278
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8747 6012 9055 6032
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 9232 5098 9260 10202
rect 9324 6662 9352 14198
rect 9508 13802 9536 14282
rect 9600 13870 9628 14758
rect 9968 14521 9996 20538
rect 18708 20466 18736 22607
rect 20626 22264 20682 22273
rect 20626 22199 20682 22208
rect 19614 21720 19670 21729
rect 19614 21655 19670 21664
rect 19628 20602 19656 21655
rect 20258 21312 20314 21321
rect 20258 21247 20314 21256
rect 20166 20768 20222 20777
rect 20166 20703 20222 20712
rect 20180 20602 20208 20703
rect 19616 20596 19668 20602
rect 19616 20538 19668 20544
rect 20168 20596 20220 20602
rect 20168 20538 20220 20544
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 18696 20460 18748 20466
rect 18696 20402 18748 20408
rect 18788 20460 18840 20466
rect 18788 20402 18840 20408
rect 19524 20460 19576 20466
rect 19524 20402 19576 20408
rect 10336 20058 10364 20402
rect 11244 20324 11296 20330
rect 11244 20266 11296 20272
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 11256 19854 11284 20266
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 11244 19848 11296 19854
rect 11244 19790 11296 19796
rect 12624 19712 12676 19718
rect 12624 19654 12676 19660
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 12636 19378 12664 19654
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 12624 19372 12676 19378
rect 12624 19314 12676 19320
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 14280 19372 14332 19378
rect 14280 19314 14332 19320
rect 14464 19372 14516 19378
rect 14464 19314 14516 19320
rect 17960 19372 18012 19378
rect 17960 19314 18012 19320
rect 12900 19168 12952 19174
rect 12952 19116 13032 19122
rect 12900 19110 13032 19116
rect 12912 19094 13032 19110
rect 11244 18692 11296 18698
rect 11244 18634 11296 18640
rect 10048 18080 10100 18086
rect 10048 18022 10100 18028
rect 9954 14512 10010 14521
rect 9954 14447 10010 14456
rect 9772 14272 9824 14278
rect 9772 14214 9824 14220
rect 9588 13864 9640 13870
rect 9588 13806 9640 13812
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 12782 9536 13738
rect 9588 13728 9640 13734
rect 9588 13670 9640 13676
rect 9600 13394 9628 13670
rect 9784 13394 9812 14214
rect 9968 13938 9996 14447
rect 10060 13938 10088 18022
rect 10416 17740 10468 17746
rect 10416 17682 10468 17688
rect 10428 17134 10456 17682
rect 10508 17196 10560 17202
rect 10508 17138 10560 17144
rect 10416 17128 10468 17134
rect 10416 17070 10468 17076
rect 10520 16794 10548 17138
rect 11060 17128 11112 17134
rect 11060 17070 11112 17076
rect 10508 16788 10560 16794
rect 10508 16730 10560 16736
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10324 16516 10376 16522
rect 10324 16458 10376 16464
rect 10336 15706 10364 16458
rect 10704 15910 10732 16662
rect 10968 16652 11020 16658
rect 10968 16594 11020 16600
rect 10692 15904 10744 15910
rect 10690 15872 10692 15881
rect 10744 15872 10746 15881
rect 10690 15807 10746 15816
rect 10324 15700 10376 15706
rect 10324 15642 10376 15648
rect 10980 15502 11008 16594
rect 11072 16250 11100 17070
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11164 16590 11192 16934
rect 11152 16584 11204 16590
rect 11152 16526 11204 16532
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11060 16108 11112 16114
rect 11060 16050 11112 16056
rect 11072 15910 11100 16050
rect 11060 15904 11112 15910
rect 11060 15846 11112 15852
rect 11072 15570 11100 15846
rect 11256 15586 11284 18634
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11992 17542 12020 18226
rect 12900 18216 12952 18222
rect 12900 18158 12952 18164
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11980 17536 12032 17542
rect 11980 17478 12032 17484
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11060 15564 11112 15570
rect 11060 15506 11112 15512
rect 11164 15558 11284 15586
rect 10968 15496 11020 15502
rect 10968 15438 11020 15444
rect 11058 15464 11114 15473
rect 10600 15360 10652 15366
rect 10600 15302 10652 15308
rect 10508 14408 10560 14414
rect 10612 14385 10640 15302
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10508 14350 10560 14356
rect 10598 14376 10654 14385
rect 10520 14090 10548 14350
rect 10598 14311 10654 14320
rect 10704 14278 10732 14962
rect 10980 14958 11008 15438
rect 11058 15399 11114 15408
rect 10968 14952 11020 14958
rect 10968 14894 11020 14900
rect 10692 14272 10744 14278
rect 10692 14214 10744 14220
rect 10520 14062 10640 14090
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9968 13530 9996 13874
rect 9956 13524 10008 13530
rect 9956 13466 10008 13472
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9772 13388 9824 13394
rect 9772 13330 9824 13336
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9404 12708 9456 12714
rect 9404 12650 9456 12656
rect 9416 12306 9444 12650
rect 9494 12472 9550 12481
rect 9784 12434 9812 13330
rect 9864 13252 9916 13258
rect 9864 13194 9916 13200
rect 9494 12407 9550 12416
rect 9404 12300 9456 12306
rect 9404 12242 9456 12248
rect 9508 12186 9536 12407
rect 9692 12406 9812 12434
rect 9508 12158 9628 12186
rect 9600 12152 9628 12158
rect 9692 12152 9720 12406
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9600 12124 9720 12152
rect 9784 12102 9812 12242
rect 9772 12096 9824 12102
rect 9586 12064 9642 12073
rect 9642 12022 9720 12050
rect 9772 12038 9824 12044
rect 9586 11999 9642 12008
rect 9586 11928 9642 11937
rect 9692 11898 9720 12022
rect 9586 11863 9642 11872
rect 9680 11892 9732 11898
rect 9402 11656 9458 11665
rect 9402 11591 9458 11600
rect 9416 11150 9444 11591
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9404 10600 9456 10606
rect 9404 10542 9456 10548
rect 9416 10062 9444 10542
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9404 8832 9456 8838
rect 9508 8809 9536 11290
rect 9600 10130 9628 11863
rect 9680 11834 9732 11840
rect 9772 11756 9824 11762
rect 9772 11698 9824 11704
rect 9784 11354 9812 11698
rect 9876 11626 9904 13194
rect 10048 13184 10100 13190
rect 10048 13126 10100 13132
rect 10060 12986 10088 13126
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10508 12980 10560 12986
rect 10508 12922 10560 12928
rect 10140 12708 10192 12714
rect 10140 12650 10192 12656
rect 10152 12434 10180 12650
rect 9968 12406 10180 12434
rect 9864 11620 9916 11626
rect 9864 11562 9916 11568
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9876 11218 9904 11562
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9864 11076 9916 11082
rect 9864 11018 9916 11024
rect 9772 10668 9824 10674
rect 9772 10610 9824 10616
rect 9784 10266 9812 10610
rect 9772 10260 9824 10266
rect 9772 10202 9824 10208
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9588 9988 9640 9994
rect 9588 9930 9640 9936
rect 9600 9042 9628 9930
rect 9784 9489 9812 10066
rect 9770 9480 9826 9489
rect 9770 9415 9826 9424
rect 9588 9036 9640 9042
rect 9588 8978 9640 8984
rect 9404 8774 9456 8780
rect 9494 8800 9550 8809
rect 9416 7449 9444 8774
rect 9494 8735 9550 8744
rect 9784 8634 9812 9415
rect 9772 8628 9824 8634
rect 9772 8570 9824 8576
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9588 8424 9640 8430
rect 9692 8401 9720 8502
rect 9588 8366 9640 8372
rect 9678 8392 9734 8401
rect 9600 8294 9628 8366
rect 9678 8327 9734 8336
rect 9508 8276 9628 8294
rect 9508 8248 9720 8276
rect 9586 8120 9642 8129
rect 9586 8055 9642 8064
rect 9496 7880 9548 7886
rect 9496 7822 9548 7828
rect 9402 7440 9458 7449
rect 9402 7375 9458 7384
rect 9312 6656 9364 6662
rect 9312 6598 9364 6604
rect 9324 6458 9352 6598
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9508 5914 9536 7822
rect 9600 7426 9628 8055
rect 9692 7546 9720 8248
rect 9680 7540 9732 7546
rect 9680 7482 9732 7488
rect 9772 7472 9824 7478
rect 9600 7420 9772 7426
rect 9600 7414 9824 7420
rect 9600 7398 9812 7414
rect 9772 7200 9824 7206
rect 9772 7142 9824 7148
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 6390 9720 6734
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9496 5908 9548 5914
rect 9496 5850 9548 5856
rect 9508 5778 9536 5850
rect 9692 5846 9720 6326
rect 9784 6322 9812 7142
rect 9772 6316 9824 6322
rect 9772 6258 9824 6264
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9680 5704 9732 5710
rect 9600 5664 9680 5692
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5098 9444 5510
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9220 5092 9272 5098
rect 9220 5034 9272 5040
rect 9404 5092 9456 5098
rect 9404 5034 9456 5040
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 9232 4690 9260 5034
rect 9220 4684 9272 4690
rect 9220 4626 9272 4632
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 8668 4276 8720 4282
rect 8668 4218 8720 4224
rect 9140 4078 9168 4558
rect 9404 4140 9456 4146
rect 9404 4082 9456 4088
rect 9128 4072 9180 4078
rect 9128 4014 9180 4020
rect 9218 4040 9274 4049
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 8944 3664 8996 3670
rect 8944 3606 8996 3612
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8680 2632 8708 3402
rect 8956 3398 8984 3606
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 2990 8984 3334
rect 9140 3194 9168 4014
rect 9218 3975 9274 3984
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8944 2984 8996 2990
rect 8944 2926 8996 2932
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 8680 2604 8800 2632
rect 8772 800 8800 2604
rect 9232 2582 9260 3975
rect 9416 3738 9444 4082
rect 9404 3732 9456 3738
rect 9404 3674 9456 3680
rect 9508 2774 9536 5170
rect 9600 5030 9628 5664
rect 9680 5646 9732 5652
rect 9588 5024 9640 5030
rect 9588 4966 9640 4972
rect 9588 4684 9640 4690
rect 9588 4626 9640 4632
rect 9600 4214 9628 4626
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9588 4004 9640 4010
rect 9588 3946 9640 3952
rect 9600 3738 9628 3946
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9692 3194 9720 4014
rect 9784 3466 9812 6258
rect 9772 3460 9824 3466
rect 9772 3402 9824 3408
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 9508 2746 9628 2774
rect 9402 2680 9458 2689
rect 9402 2615 9404 2624
rect 9456 2615 9458 2624
rect 9404 2586 9456 2592
rect 9220 2576 9272 2582
rect 9220 2518 9272 2524
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 1970 9168 2246
rect 9128 1964 9180 1970
rect 9128 1906 9180 1912
rect 9232 800 9260 2518
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9324 2106 9352 2246
rect 9312 2100 9364 2106
rect 9312 2042 9364 2048
rect 9600 800 9628 2746
rect 9692 2650 9720 2858
rect 9876 2774 9904 11018
rect 9784 2746 9904 2774
rect 9968 2774 9996 12406
rect 10152 12306 10180 12406
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10152 11354 10180 12106
rect 10428 11762 10456 12922
rect 10416 11756 10468 11762
rect 10416 11698 10468 11704
rect 10140 11348 10192 11354
rect 10140 11290 10192 11296
rect 10048 11212 10100 11218
rect 10048 11154 10100 11160
rect 10060 9738 10088 11154
rect 10152 10742 10180 11290
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10305 10364 10542
rect 10322 10296 10378 10305
rect 10322 10231 10378 10240
rect 10140 10056 10192 10062
rect 10140 9998 10192 10004
rect 10152 9874 10180 9998
rect 10152 9846 10364 9874
rect 10060 9710 10180 9738
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10060 8634 10088 8910
rect 10048 8628 10100 8634
rect 10048 8570 10100 8576
rect 10048 8492 10100 8498
rect 10048 8434 10100 8440
rect 10060 4146 10088 8434
rect 10152 7426 10180 9710
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 10244 7546 10272 9522
rect 10336 9518 10364 9846
rect 10324 9512 10376 9518
rect 10324 9454 10376 9460
rect 10336 7886 10364 9454
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 10232 7540 10284 7546
rect 10232 7482 10284 7488
rect 10152 7398 10272 7426
rect 10138 5672 10194 5681
rect 10138 5607 10194 5616
rect 10152 4622 10180 5607
rect 10244 5522 10272 7398
rect 10336 6798 10364 7822
rect 10324 6792 10376 6798
rect 10324 6734 10376 6740
rect 10336 5710 10364 6734
rect 10428 6458 10456 11698
rect 10520 11694 10548 12922
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 6452 10468 6458
rect 10416 6394 10468 6400
rect 10520 6186 10548 11630
rect 10612 9722 10640 14062
rect 10784 13184 10836 13190
rect 10784 13126 10836 13132
rect 10692 10600 10744 10606
rect 10692 10542 10744 10548
rect 10600 9716 10652 9722
rect 10600 9658 10652 9664
rect 10598 9616 10654 9625
rect 10598 9551 10600 9560
rect 10652 9551 10654 9560
rect 10600 9522 10652 9528
rect 10612 9110 10640 9522
rect 10704 9178 10732 10542
rect 10692 9172 10744 9178
rect 10692 9114 10744 9120
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10704 6458 10732 6938
rect 10692 6452 10744 6458
rect 10692 6394 10744 6400
rect 10692 6316 10744 6322
rect 10612 6276 10692 6304
rect 10508 6180 10560 6186
rect 10508 6122 10560 6128
rect 10612 6118 10640 6276
rect 10692 6258 10744 6264
rect 10600 6112 10652 6118
rect 10600 6054 10652 6060
rect 10324 5704 10376 5710
rect 10324 5646 10376 5652
rect 10244 5494 10456 5522
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4140 10100 4146
rect 10048 4082 10100 4088
rect 10060 3942 10088 4082
rect 10048 3936 10100 3942
rect 10048 3878 10100 3884
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3126 10180 3878
rect 10324 3664 10376 3670
rect 10324 3606 10376 3612
rect 10140 3120 10192 3126
rect 10140 3062 10192 3068
rect 10336 2922 10364 3606
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 9968 2746 10088 2774
rect 9680 2644 9732 2650
rect 9680 2586 9732 2592
rect 9784 2514 9812 2746
rect 10060 2650 10088 2746
rect 10048 2644 10100 2650
rect 10048 2586 10100 2592
rect 9772 2508 9824 2514
rect 9772 2450 9824 2456
rect 10060 870 10180 898
rect 10060 800 10088 870
rect 8404 734 8616 762
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10152 762 10180 870
rect 10336 762 10364 2858
rect 10428 2650 10456 5494
rect 10508 4276 10560 4282
rect 10508 4218 10560 4224
rect 10520 3777 10548 4218
rect 10506 3768 10562 3777
rect 10506 3703 10562 3712
rect 10612 3534 10640 6054
rect 10796 5080 10824 13126
rect 11072 12986 11100 15399
rect 11060 12980 11112 12986
rect 11060 12922 11112 12928
rect 11058 12336 11114 12345
rect 11058 12271 11114 12280
rect 11072 11354 11100 12271
rect 11060 11348 11112 11354
rect 11060 11290 11112 11296
rect 11164 11014 11192 15558
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11808 14414 11836 16934
rect 11992 16658 12020 17478
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 11888 16108 11940 16114
rect 11888 16050 11940 16056
rect 11900 16017 11928 16050
rect 11886 16008 11942 16017
rect 11886 15943 11942 15952
rect 12084 15502 12112 18022
rect 12162 17640 12218 17649
rect 12162 17575 12164 17584
rect 12216 17575 12218 17584
rect 12164 17546 12216 17552
rect 12176 17134 12204 17546
rect 12256 17536 12308 17542
rect 12256 17478 12308 17484
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12164 17128 12216 17134
rect 12164 17070 12216 17076
rect 12176 16046 12204 17070
rect 12268 16658 12296 17478
rect 12636 17270 12664 17478
rect 12912 17338 12940 18158
rect 12900 17332 12952 17338
rect 12900 17274 12952 17280
rect 12624 17264 12676 17270
rect 12624 17206 12676 17212
rect 12348 17196 12400 17202
rect 12348 17138 12400 17144
rect 12256 16652 12308 16658
rect 12256 16594 12308 16600
rect 12164 16040 12216 16046
rect 12164 15982 12216 15988
rect 12254 16008 12310 16017
rect 12254 15943 12310 15952
rect 12072 15496 12124 15502
rect 12072 15438 12124 15444
rect 12268 14464 12296 15943
rect 12176 14436 12296 14464
rect 11796 14408 11848 14414
rect 11796 14350 11848 14356
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11888 14340 11940 14346
rect 11888 14282 11940 14288
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11256 14006 11284 14214
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11900 14074 11928 14282
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11244 14000 11296 14006
rect 11244 13942 11296 13948
rect 11888 13320 11940 13326
rect 11888 13262 11940 13268
rect 11244 13184 11296 13190
rect 11244 13126 11296 13132
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11256 12434 11284 13126
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11716 12889 11744 13126
rect 11702 12880 11758 12889
rect 11702 12815 11758 12824
rect 11796 12776 11848 12782
rect 11796 12718 11848 12724
rect 11256 12406 11744 12434
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 11244 11552 11296 11558
rect 11244 11494 11296 11500
rect 11256 11257 11284 11494
rect 11242 11248 11298 11257
rect 11242 11183 11298 11192
rect 11152 11008 11204 11014
rect 11152 10950 11204 10956
rect 11152 10600 11204 10606
rect 11152 10542 11204 10548
rect 11060 10464 11112 10470
rect 11060 10406 11112 10412
rect 10876 9716 10928 9722
rect 10876 9658 10928 9664
rect 10888 8430 10916 9658
rect 10876 8424 10928 8430
rect 10876 8366 10928 8372
rect 10888 8294 10916 8366
rect 10876 8288 10928 8294
rect 10876 8230 10928 8236
rect 10888 6905 10916 8230
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10874 6896 10930 6905
rect 10874 6831 10930 6840
rect 10876 6656 10928 6662
rect 10876 6598 10928 6604
rect 10704 5052 10824 5080
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10600 3392 10652 3398
rect 10600 3334 10652 3340
rect 10612 3194 10640 3334
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10704 2582 10732 5052
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10692 2576 10744 2582
rect 10692 2518 10744 2524
rect 10416 2508 10468 2514
rect 10416 2450 10468 2456
rect 10428 2394 10456 2450
rect 10428 2366 10548 2394
rect 10520 800 10548 2366
rect 10796 2310 10824 4422
rect 10888 4282 10916 6598
rect 10980 6254 11008 7686
rect 10968 6248 11020 6254
rect 10968 6190 11020 6196
rect 10980 5710 11008 6190
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 10968 4752 11020 4758
rect 10968 4694 11020 4700
rect 10876 4276 10928 4282
rect 10876 4218 10928 4224
rect 10876 4072 10928 4078
rect 10876 4014 10928 4020
rect 10888 3602 10916 4014
rect 10876 3596 10928 3602
rect 10876 3538 10928 3544
rect 10980 3534 11008 4694
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11072 3058 11100 10406
rect 11164 9994 11192 10542
rect 11256 10169 11284 11183
rect 11716 11098 11744 12406
rect 11808 12170 11836 12718
rect 11796 12164 11848 12170
rect 11796 12106 11848 12112
rect 11808 11830 11836 12106
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11808 11286 11836 11766
rect 11796 11280 11848 11286
rect 11796 11222 11848 11228
rect 11716 11070 11836 11098
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11716 10810 11744 10950
rect 11704 10804 11756 10810
rect 11704 10746 11756 10752
rect 11426 10296 11482 10305
rect 11426 10231 11428 10240
rect 11480 10231 11482 10240
rect 11428 10202 11480 10208
rect 11242 10160 11298 10169
rect 11242 10095 11298 10104
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 11164 9518 11192 9930
rect 11440 9908 11468 10202
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11256 9880 11468 9908
rect 11152 9512 11204 9518
rect 11152 9454 11204 9460
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11164 9081 11192 9114
rect 11150 9072 11206 9081
rect 11150 9007 11206 9016
rect 11256 8974 11284 9880
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11716 9586 11744 9998
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11244 8968 11296 8974
rect 11244 8910 11296 8916
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11716 7818 11744 9522
rect 11244 7812 11296 7818
rect 11244 7754 11296 7760
rect 11704 7812 11756 7818
rect 11704 7754 11756 7760
rect 11256 6866 11284 7754
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 11244 6860 11296 6866
rect 11244 6802 11296 6808
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 11152 6112 11204 6118
rect 11152 6054 11204 6060
rect 11244 6112 11296 6118
rect 11244 6054 11296 6060
rect 11164 5370 11192 6054
rect 11152 5364 11204 5370
rect 11152 5306 11204 5312
rect 11256 5302 11284 6054
rect 11716 5778 11744 7754
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 11244 5296 11296 5302
rect 11244 5238 11296 5244
rect 11716 5234 11744 5510
rect 11704 5228 11756 5234
rect 11704 5170 11756 5176
rect 11808 5114 11836 11070
rect 11900 8514 11928 13262
rect 11980 12708 12032 12714
rect 11980 12650 12032 12656
rect 11992 11898 12020 12650
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 11980 11076 12032 11082
rect 11980 11018 12032 11024
rect 11992 10810 12020 11018
rect 12084 10826 12112 14350
rect 12176 12186 12204 14436
rect 12256 14340 12308 14346
rect 12256 14282 12308 14288
rect 12268 14074 12296 14282
rect 12256 14068 12308 14074
rect 12256 14010 12308 14016
rect 12360 13530 12388 17138
rect 12532 17060 12584 17066
rect 12532 17002 12584 17008
rect 12544 16946 12572 17002
rect 12544 16918 12756 16946
rect 12624 16788 12676 16794
rect 12624 16730 12676 16736
rect 12532 13864 12584 13870
rect 12530 13832 12532 13841
rect 12584 13832 12586 13841
rect 12440 13796 12492 13802
rect 12530 13767 12586 13776
rect 12440 13738 12492 13744
rect 12348 13524 12400 13530
rect 12348 13466 12400 13472
rect 12254 13424 12310 13433
rect 12254 13359 12256 13368
rect 12308 13359 12310 13368
rect 12256 13330 12308 13336
rect 12346 13016 12402 13025
rect 12346 12951 12402 12960
rect 12360 12850 12388 12951
rect 12348 12844 12400 12850
rect 12348 12786 12400 12792
rect 12348 12436 12400 12442
rect 12348 12378 12400 12384
rect 12176 12158 12296 12186
rect 12164 12096 12216 12102
rect 12164 12038 12216 12044
rect 12176 11694 12204 12038
rect 12164 11688 12216 11694
rect 12164 11630 12216 11636
rect 11980 10804 12032 10810
rect 12084 10798 12204 10826
rect 11980 10746 12032 10752
rect 11992 9738 12020 10746
rect 12072 10736 12124 10742
rect 12072 10678 12124 10684
rect 12084 10198 12112 10678
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 11992 9710 12112 9738
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11992 9178 12020 9522
rect 11980 9172 12032 9178
rect 11980 9114 12032 9120
rect 11900 8486 12020 8514
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11900 7546 11928 8366
rect 11992 7993 12020 8486
rect 11978 7984 12034 7993
rect 11978 7919 12034 7928
rect 11888 7540 11940 7546
rect 11888 7482 11940 7488
rect 12084 7478 12112 9710
rect 12176 8838 12204 10798
rect 12164 8832 12216 8838
rect 12164 8774 12216 8780
rect 12268 8514 12296 12158
rect 12176 8486 12296 8514
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12176 6497 12204 8486
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12268 8090 12296 8366
rect 12256 8084 12308 8090
rect 12256 8026 12308 8032
rect 12268 6798 12296 8026
rect 12360 6882 12388 12378
rect 12452 9042 12480 13738
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12544 11694 12572 12582
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12544 7546 12572 8434
rect 12532 7540 12584 7546
rect 12532 7482 12584 7488
rect 12360 6854 12480 6882
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12162 6488 12218 6497
rect 12162 6423 12218 6432
rect 11888 6316 11940 6322
rect 12164 6316 12216 6322
rect 11888 6258 11940 6264
rect 12084 6276 12164 6304
rect 11716 5086 11836 5114
rect 11244 5024 11296 5030
rect 11244 4966 11296 4972
rect 11152 4616 11204 4622
rect 11152 4558 11204 4564
rect 11164 4282 11192 4558
rect 11152 4276 11204 4282
rect 11152 4218 11204 4224
rect 11256 3534 11284 4966
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 11716 4026 11744 5086
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11808 4554 11836 4966
rect 11796 4548 11848 4554
rect 11796 4490 11848 4496
rect 11900 4486 11928 6258
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11992 6089 12020 6190
rect 11978 6080 12034 6089
rect 11978 6015 12034 6024
rect 11992 5846 12020 6015
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11888 4480 11940 4486
rect 11888 4422 11940 4428
rect 11624 3998 11744 4026
rect 11624 3670 11652 3998
rect 11704 3936 11756 3942
rect 11704 3878 11756 3884
rect 11612 3664 11664 3670
rect 11612 3606 11664 3612
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 11716 3058 11744 3878
rect 11796 3392 11848 3398
rect 11796 3334 11848 3340
rect 11808 3126 11836 3334
rect 11796 3120 11848 3126
rect 11796 3062 11848 3068
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 11060 3052 11112 3058
rect 11060 2994 11112 3000
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 10888 2446 10916 2994
rect 11152 2848 11204 2854
rect 11152 2790 11204 2796
rect 10968 2576 11020 2582
rect 10968 2518 11020 2524
rect 10876 2440 10928 2446
rect 10876 2382 10928 2388
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10980 800 11008 2518
rect 11164 2514 11192 2790
rect 11992 2582 12020 5646
rect 12084 5642 12112 6276
rect 12164 6258 12216 6264
rect 12164 6180 12216 6186
rect 12164 6122 12216 6128
rect 12176 5914 12204 6122
rect 12164 5908 12216 5914
rect 12360 5896 12388 6734
rect 12164 5850 12216 5856
rect 12268 5868 12388 5896
rect 12072 5636 12124 5642
rect 12072 5578 12124 5584
rect 12268 4826 12296 5868
rect 12348 5772 12400 5778
rect 12348 5714 12400 5720
rect 12360 5302 12388 5714
rect 12452 5710 12480 6854
rect 12530 5808 12586 5817
rect 12530 5743 12586 5752
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12348 5296 12400 5302
rect 12348 5238 12400 5244
rect 12440 5024 12492 5030
rect 12440 4966 12492 4972
rect 12256 4820 12308 4826
rect 12256 4762 12308 4768
rect 12072 4548 12124 4554
rect 12072 4490 12124 4496
rect 12084 4214 12112 4490
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 12348 4140 12400 4146
rect 12452 4128 12480 4966
rect 12400 4100 12480 4128
rect 12348 4082 12400 4088
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12176 2990 12204 3470
rect 12164 2984 12216 2990
rect 12164 2926 12216 2932
rect 11980 2576 12032 2582
rect 11980 2518 12032 2524
rect 11152 2508 11204 2514
rect 11152 2450 11204 2456
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 11256 1986 11284 2382
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 11256 1958 11468 1986
rect 11440 800 11468 1958
rect 11992 1034 12020 2518
rect 11900 1006 12020 1034
rect 11900 800 11928 1006
rect 12360 800 12388 4082
rect 12544 3058 12572 5743
rect 12636 4010 12664 16730
rect 12728 13734 12756 16918
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 12912 16454 12940 16594
rect 12900 16448 12952 16454
rect 12900 16390 12952 16396
rect 12808 15972 12860 15978
rect 12808 15914 12860 15920
rect 12820 15706 12848 15914
rect 12808 15700 12860 15706
rect 12808 15642 12860 15648
rect 12820 15026 12848 15642
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 12820 14482 12848 14962
rect 12808 14476 12860 14482
rect 12808 14418 12860 14424
rect 12820 13938 12848 14418
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12912 13818 12940 16390
rect 12820 13790 12940 13818
rect 12716 13728 12768 13734
rect 12716 13670 12768 13676
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12889 12756 13126
rect 12714 12880 12770 12889
rect 12714 12815 12770 12824
rect 12820 12434 12848 13790
rect 12900 13524 12952 13530
rect 12900 13466 12952 13472
rect 12728 12406 12848 12434
rect 12728 10742 12756 12406
rect 12912 11014 12940 13466
rect 13004 13326 13032 19094
rect 13452 18964 13504 18970
rect 13452 18906 13504 18912
rect 13176 18420 13228 18426
rect 13176 18362 13228 18368
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13084 13864 13136 13870
rect 13082 13832 13084 13841
rect 13136 13832 13138 13841
rect 13082 13767 13138 13776
rect 13084 13388 13136 13394
rect 13084 13330 13136 13336
rect 12992 13320 13044 13326
rect 12992 13262 13044 13268
rect 13096 12918 13124 13330
rect 13084 12912 13136 12918
rect 13084 12854 13136 12860
rect 13096 12730 13124 12854
rect 13004 12702 13124 12730
rect 13004 11354 13032 12702
rect 13084 12436 13136 12442
rect 13084 12378 13136 12384
rect 13096 11694 13124 12378
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 12992 11348 13044 11354
rect 12992 11290 13044 11296
rect 12900 11008 12952 11014
rect 12900 10950 12952 10956
rect 12716 10736 12768 10742
rect 12716 10678 12768 10684
rect 12806 10568 12862 10577
rect 12806 10503 12808 10512
rect 12860 10503 12862 10512
rect 12808 10474 12860 10480
rect 12912 9674 12940 10950
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12728 9646 12940 9674
rect 12728 8838 12756 9646
rect 13096 9382 13124 10610
rect 13188 9625 13216 18362
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13280 17202 13308 18090
rect 13268 17196 13320 17202
rect 13268 17138 13320 17144
rect 13372 17082 13400 18362
rect 13464 18290 13492 18906
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13464 18086 13492 18226
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13280 17054 13400 17082
rect 13280 13190 13308 17054
rect 13360 15360 13412 15366
rect 13360 15302 13412 15308
rect 13372 14618 13400 15302
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13372 13841 13400 14214
rect 13358 13832 13414 13841
rect 13358 13767 13414 13776
rect 13360 13320 13412 13326
rect 13360 13262 13412 13268
rect 13372 13190 13400 13262
rect 13268 13184 13320 13190
rect 13268 13126 13320 13132
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13280 12617 13308 13126
rect 13372 12753 13400 13126
rect 13358 12744 13414 12753
rect 13358 12679 13414 12688
rect 13266 12608 13322 12617
rect 13266 12543 13322 12552
rect 13372 12434 13400 12679
rect 13280 12406 13400 12434
rect 13174 9616 13230 9625
rect 13174 9551 13230 9560
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 12900 9104 12952 9110
rect 12900 9046 12952 9052
rect 12716 8832 12768 8838
rect 12716 8774 12768 8780
rect 12728 8537 12756 8774
rect 12714 8528 12770 8537
rect 12714 8463 12770 8472
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12716 8016 12768 8022
rect 12716 7958 12768 7964
rect 12728 6322 12756 7958
rect 12716 6316 12768 6322
rect 12716 6258 12768 6264
rect 12624 4004 12676 4010
rect 12624 3946 12676 3952
rect 12820 3534 12848 8298
rect 12912 7993 12940 9046
rect 12992 8968 13044 8974
rect 12992 8910 13044 8916
rect 12898 7984 12954 7993
rect 12898 7919 12954 7928
rect 13004 6662 13032 8910
rect 13188 8378 13216 9551
rect 13280 8401 13308 12406
rect 13360 9444 13412 9450
rect 13360 9386 13412 9392
rect 13096 8350 13216 8378
rect 13266 8392 13322 8401
rect 13096 7002 13124 8350
rect 13266 8327 13322 8336
rect 13176 8288 13228 8294
rect 13176 8230 13228 8236
rect 13188 7954 13216 8230
rect 13176 7948 13228 7954
rect 13176 7890 13228 7896
rect 13268 7744 13320 7750
rect 13268 7686 13320 7692
rect 13280 7546 13308 7686
rect 13268 7540 13320 7546
rect 13268 7482 13320 7488
rect 13372 7313 13400 9386
rect 13464 8974 13492 18022
rect 13648 17134 13676 19314
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 14292 18766 14320 19314
rect 14476 19258 14504 19314
rect 14384 19230 14504 19258
rect 14384 19174 14412 19230
rect 14372 19168 14424 19174
rect 15108 19168 15160 19174
rect 14372 19110 14424 19116
rect 15028 19116 15108 19122
rect 15028 19110 15160 19116
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 14280 18760 14332 18766
rect 14280 18702 14332 18708
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 13820 17808 13872 17814
rect 13820 17750 13872 17756
rect 13636 17128 13688 17134
rect 13636 17070 13688 17076
rect 13648 16726 13676 17070
rect 13832 16998 13860 17750
rect 13820 16992 13872 16998
rect 13820 16934 13872 16940
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 13636 16720 13688 16726
rect 13636 16662 13688 16668
rect 13820 16040 13872 16046
rect 13820 15982 13872 15988
rect 13832 15910 13860 15982
rect 13820 15904 13872 15910
rect 13740 15864 13820 15892
rect 13636 15020 13688 15026
rect 13636 14962 13688 14968
rect 13648 14822 13676 14962
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13544 13864 13596 13870
rect 13544 13806 13596 13812
rect 13556 11200 13584 13806
rect 13636 12640 13688 12646
rect 13636 12582 13688 12588
rect 13648 11665 13676 12582
rect 13740 12209 13768 15864
rect 13820 15846 13872 15852
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 14188 15564 14240 15570
rect 14188 15506 14240 15512
rect 14200 15094 14228 15506
rect 14188 15088 14240 15094
rect 14188 15030 14240 15036
rect 14292 14822 14320 18702
rect 14384 18222 14412 19110
rect 15028 19094 15148 19110
rect 14924 18624 14976 18630
rect 14924 18566 14976 18572
rect 14936 18442 14964 18566
rect 14844 18414 14964 18442
rect 14844 18222 14872 18414
rect 14372 18216 14424 18222
rect 14372 18158 14424 18164
rect 14832 18216 14884 18222
rect 14832 18158 14884 18164
rect 14924 18216 14976 18222
rect 14924 18158 14976 18164
rect 14384 17746 14412 18158
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14372 17740 14424 17746
rect 14372 17682 14424 17688
rect 14384 17626 14412 17682
rect 14384 17598 14504 17626
rect 14372 17536 14424 17542
rect 14372 17478 14424 17484
rect 14384 17338 14412 17478
rect 14372 17332 14424 17338
rect 14372 17274 14424 17280
rect 14476 16658 14504 17598
rect 14568 17542 14596 17818
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14936 17338 14964 18158
rect 14924 17332 14976 17338
rect 14924 17274 14976 17280
rect 15028 17218 15056 19094
rect 15580 18766 15608 19110
rect 15568 18760 15620 18766
rect 15568 18702 15620 18708
rect 15108 18284 15160 18290
rect 15108 18226 15160 18232
rect 15120 17882 15148 18226
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15108 17876 15160 17882
rect 15108 17818 15160 17824
rect 15396 17678 15424 18022
rect 15580 17746 15608 18702
rect 17040 18624 17092 18630
rect 17040 18566 17092 18572
rect 17868 18624 17920 18630
rect 17868 18566 17920 18572
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 15568 17740 15620 17746
rect 15568 17682 15620 17688
rect 15384 17672 15436 17678
rect 15580 17626 15608 17682
rect 15384 17614 15436 17620
rect 15488 17598 15608 17626
rect 16212 17604 16264 17610
rect 15108 17536 15160 17542
rect 15108 17478 15160 17484
rect 15120 17338 15148 17478
rect 15108 17332 15160 17338
rect 15108 17274 15160 17280
rect 14844 17190 15056 17218
rect 14648 17128 14700 17134
rect 14648 17070 14700 17076
rect 14738 17096 14794 17105
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14556 16108 14608 16114
rect 14556 16050 14608 16056
rect 14464 15904 14516 15910
rect 14464 15846 14516 15852
rect 14476 15502 14504 15846
rect 14568 15570 14596 16050
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 14464 15496 14516 15502
rect 14660 15450 14688 17070
rect 14738 17031 14794 17040
rect 14464 15438 14516 15444
rect 14568 15422 14688 15450
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14280 14816 14332 14822
rect 14280 14758 14332 14764
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13832 12442 13860 13262
rect 14292 12646 14320 14758
rect 14384 14482 14412 15030
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14372 14272 14424 14278
rect 14372 14214 14424 14220
rect 14384 14074 14412 14214
rect 14372 14068 14424 14074
rect 14372 14010 14424 14016
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 13820 12436 13872 12442
rect 13820 12378 13872 12384
rect 14292 12238 14320 12582
rect 14476 12481 14504 13874
rect 14462 12472 14518 12481
rect 14462 12407 14518 12416
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14280 12232 14332 12238
rect 13726 12200 13782 12209
rect 14280 12174 14332 12180
rect 13726 12135 13782 12144
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14200 11830 14228 12038
rect 14188 11824 14240 11830
rect 14188 11766 14240 11772
rect 14384 11694 14412 12310
rect 14464 12096 14516 12102
rect 14464 12038 14516 12044
rect 14476 11898 14504 12038
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 11688 14424 11694
rect 13634 11656 13690 11665
rect 14372 11630 14424 11636
rect 13634 11591 13690 11600
rect 13636 11552 13688 11558
rect 13636 11494 13688 11500
rect 13648 11354 13676 11494
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 14384 11257 14412 11630
rect 14370 11248 14426 11257
rect 13556 11172 13676 11200
rect 14370 11183 14426 11192
rect 13648 11121 13676 11172
rect 13634 11112 13690 11121
rect 13544 11076 13596 11082
rect 14384 11082 14412 11183
rect 13634 11047 13690 11056
rect 14372 11076 14424 11082
rect 13544 11018 13596 11024
rect 14372 11018 14424 11024
rect 13556 10713 13584 11018
rect 13820 11008 13872 11014
rect 13820 10950 13872 10956
rect 13542 10704 13598 10713
rect 13542 10639 13598 10648
rect 13832 10554 13860 10950
rect 13648 10526 13860 10554
rect 14280 10532 14332 10538
rect 13648 10062 13676 10526
rect 14280 10474 14332 10480
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13636 10056 13688 10062
rect 13636 9998 13688 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13740 9586 13768 9998
rect 13728 9580 13780 9586
rect 13728 9522 13780 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13452 8968 13504 8974
rect 13452 8910 13504 8916
rect 13542 8936 13598 8945
rect 13542 8871 13598 8880
rect 13452 8832 13504 8838
rect 13556 8786 13584 8871
rect 13648 8838 13676 8978
rect 13504 8780 13584 8786
rect 13452 8774 13584 8780
rect 13636 8832 13688 8838
rect 13636 8774 13688 8780
rect 13464 8758 13584 8774
rect 13556 8673 13584 8758
rect 13542 8664 13598 8673
rect 13542 8599 13598 8608
rect 13556 8498 13584 8599
rect 13648 8498 13676 8774
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 13636 8492 13688 8498
rect 13636 8434 13688 8440
rect 13740 8430 13768 9318
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13544 8356 13596 8362
rect 13544 8298 13596 8304
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13464 7818 13492 7890
rect 13452 7812 13504 7818
rect 13452 7754 13504 7760
rect 13358 7304 13414 7313
rect 13464 7274 13492 7754
rect 13358 7239 13414 7248
rect 13452 7268 13504 7274
rect 13452 7210 13504 7216
rect 13084 6996 13136 7002
rect 13084 6938 13136 6944
rect 12992 6656 13044 6662
rect 12992 6598 13044 6604
rect 13176 6656 13228 6662
rect 13176 6598 13228 6604
rect 13004 5710 13032 6598
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5636 12952 5642
rect 12900 5578 12952 5584
rect 12912 4826 12940 5578
rect 12992 5296 13044 5302
rect 12992 5238 13044 5244
rect 12900 4820 12952 4826
rect 12900 4762 12952 4768
rect 13004 4690 13032 5238
rect 13084 5092 13136 5098
rect 13084 5034 13136 5040
rect 12992 4684 13044 4690
rect 12992 4626 13044 4632
rect 13096 4146 13124 5034
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 12808 3528 12860 3534
rect 12808 3470 12860 3476
rect 12624 3392 12676 3398
rect 12624 3334 12676 3340
rect 12636 3194 12664 3334
rect 12624 3188 12676 3194
rect 12624 3130 12676 3136
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12544 2446 12572 2790
rect 12728 2774 12756 3130
rect 12912 3058 12940 3674
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 12636 2746 12756 2774
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12636 2378 12664 2746
rect 13004 2446 13032 2790
rect 13188 2650 13216 6598
rect 13268 6248 13320 6254
rect 13268 6190 13320 6196
rect 13280 5914 13308 6190
rect 13268 5908 13320 5914
rect 13268 5850 13320 5856
rect 13280 5642 13308 5850
rect 13268 5636 13320 5642
rect 13268 5578 13320 5584
rect 13556 5370 13584 8298
rect 13832 7478 13860 10406
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 14292 10266 14320 10474
rect 14372 10464 14424 10470
rect 14372 10406 14424 10412
rect 14280 10260 14332 10266
rect 14280 10202 14332 10208
rect 14280 9988 14332 9994
rect 14280 9930 14332 9936
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14108 9518 14136 9862
rect 14292 9722 14320 9930
rect 14384 9722 14412 10406
rect 14280 9716 14332 9722
rect 14280 9658 14332 9664
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14096 9512 14148 9518
rect 14096 9454 14148 9460
rect 14280 9512 14332 9518
rect 14280 9454 14332 9460
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 14292 8974 14320 9454
rect 14280 8968 14332 8974
rect 14280 8910 14332 8916
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 14384 7886 14412 8434
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14568 7834 14596 15422
rect 14752 15042 14780 17031
rect 14660 15014 14780 15042
rect 14660 9450 14688 15014
rect 14740 13864 14792 13870
rect 14740 13806 14792 13812
rect 14752 12186 14780 13806
rect 14844 12374 14872 17190
rect 15488 17134 15516 17598
rect 16212 17546 16264 17552
rect 16304 17604 16356 17610
rect 16304 17546 16356 17552
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15476 17128 15528 17134
rect 15476 17070 15528 17076
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15120 16658 15148 17002
rect 15580 16794 15608 17478
rect 16132 17338 16160 17478
rect 16120 17332 16172 17338
rect 16120 17274 16172 17280
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 16224 16726 16252 17546
rect 16316 16794 16344 17546
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16408 17338 16436 17478
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 16396 17332 16448 17338
rect 16396 17274 16448 17280
rect 16304 16788 16356 16794
rect 16304 16730 16356 16736
rect 16028 16720 16080 16726
rect 16026 16688 16028 16697
rect 16212 16720 16264 16726
rect 16080 16688 16082 16697
rect 15108 16652 15160 16658
rect 16212 16662 16264 16668
rect 16026 16623 16082 16632
rect 15108 16594 15160 16600
rect 15016 16448 15068 16454
rect 15016 16390 15068 16396
rect 15028 15978 15056 16390
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 15016 15972 15068 15978
rect 15016 15914 15068 15920
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14922 14376 14978 14385
rect 14922 14311 14978 14320
rect 14936 14006 14964 14311
rect 14924 14000 14976 14006
rect 14924 13942 14976 13948
rect 14924 13184 14976 13190
rect 14924 13126 14976 13132
rect 14832 12368 14884 12374
rect 14832 12310 14884 12316
rect 14936 12238 14964 13126
rect 14924 12232 14976 12238
rect 14752 12158 14872 12186
rect 14924 12174 14976 12180
rect 14740 12096 14792 12102
rect 14844 12084 14872 12158
rect 14844 12056 14964 12084
rect 14740 12038 14792 12044
rect 14752 11694 14780 12038
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14752 11286 14780 11630
rect 14740 11280 14792 11286
rect 14740 11222 14792 11228
rect 14648 9444 14700 9450
rect 14648 9386 14700 9392
rect 14832 8832 14884 8838
rect 14832 8774 14884 8780
rect 14844 8566 14872 8774
rect 14832 8560 14884 8566
rect 14832 8502 14884 8508
rect 13820 7472 13872 7478
rect 13820 7414 13872 7420
rect 14384 7410 14412 7822
rect 14568 7806 14872 7834
rect 14556 7744 14608 7750
rect 14556 7686 14608 7692
rect 14372 7404 14424 7410
rect 14424 7364 14504 7392
rect 14372 7346 14424 7352
rect 13945 7100 14253 7120
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 13636 6112 13688 6118
rect 13636 6054 13688 6060
rect 13648 5817 13676 6054
rect 13634 5808 13690 5817
rect 13634 5743 13690 5752
rect 13544 5364 13596 5370
rect 13544 5306 13596 5312
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4146 13584 4966
rect 13544 4140 13596 4146
rect 13544 4082 13596 4088
rect 13740 4049 13768 6598
rect 13820 6112 13872 6118
rect 13820 6054 13872 6060
rect 13832 5778 13860 6054
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 14384 5846 14412 6734
rect 14476 6254 14504 7364
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 14462 5944 14518 5953
rect 14462 5879 14518 5888
rect 14372 5840 14424 5846
rect 14372 5782 14424 5788
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 14280 5568 14332 5574
rect 14280 5510 14332 5516
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 14096 4684 14148 4690
rect 14096 4626 14148 4632
rect 13820 4616 13872 4622
rect 13820 4558 13872 4564
rect 13832 4486 13860 4558
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 14108 4282 14136 4626
rect 14096 4276 14148 4282
rect 14096 4218 14148 4224
rect 13726 4040 13782 4049
rect 13726 3975 13782 3984
rect 13728 3936 13780 3942
rect 13728 3878 13780 3884
rect 13740 3670 13768 3878
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 13636 3664 13688 3670
rect 13634 3632 13636 3641
rect 13728 3664 13780 3670
rect 13688 3632 13690 3641
rect 13728 3606 13780 3612
rect 13634 3567 13690 3576
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14200 3194 14228 3470
rect 14188 3188 14240 3194
rect 14188 3130 14240 3136
rect 14292 3058 14320 5510
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 13820 2916 13872 2922
rect 13820 2858 13872 2864
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13832 2446 13860 2858
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 14096 2576 14148 2582
rect 14096 2518 14148 2524
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 12820 800 12848 2246
rect 13280 800 13308 2246
rect 13740 800 13768 2246
rect 14108 800 14136 2518
rect 14384 1358 14412 4422
rect 14476 4146 14504 5879
rect 14568 4214 14596 7686
rect 14648 7200 14700 7206
rect 14648 7142 14700 7148
rect 14660 7041 14688 7142
rect 14646 7032 14702 7041
rect 14646 6967 14702 6976
rect 14660 6458 14688 6967
rect 14740 6656 14792 6662
rect 14740 6598 14792 6604
rect 14648 6452 14700 6458
rect 14648 6394 14700 6400
rect 14752 4622 14780 6598
rect 14740 4616 14792 4622
rect 14740 4558 14792 4564
rect 14556 4208 14608 4214
rect 14556 4150 14608 4156
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 14740 4072 14792 4078
rect 14740 4014 14792 4020
rect 14556 3936 14608 3942
rect 14556 3878 14608 3884
rect 14568 3738 14596 3878
rect 14556 3732 14608 3738
rect 14556 3674 14608 3680
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14660 2446 14688 3402
rect 14752 2938 14780 4014
rect 14844 3097 14872 7806
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 14752 2910 14872 2938
rect 14844 2854 14872 2910
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14832 2848 14884 2854
rect 14832 2790 14884 2796
rect 14752 2446 14780 2790
rect 14936 2774 14964 12056
rect 15028 8945 15056 15302
rect 15212 15162 15240 16050
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 16212 15904 16264 15910
rect 16212 15846 16264 15852
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15672 15162 15700 15370
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15212 14958 15240 15098
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15568 14952 15620 14958
rect 15568 14894 15620 14900
rect 15580 14618 15608 14894
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15488 13977 15516 14214
rect 15474 13968 15530 13977
rect 15384 13932 15436 13938
rect 15474 13903 15530 13912
rect 15384 13874 15436 13880
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12850 15240 13194
rect 15200 12844 15252 12850
rect 15200 12786 15252 12792
rect 15396 12782 15424 13874
rect 15672 13433 15700 14350
rect 15658 13424 15714 13433
rect 15658 13359 15714 13368
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15474 13016 15530 13025
rect 15474 12951 15530 12960
rect 15488 12918 15516 12951
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15384 12776 15436 12782
rect 15384 12718 15436 12724
rect 15108 11076 15160 11082
rect 15108 11018 15160 11024
rect 15014 8936 15070 8945
rect 15014 8871 15070 8880
rect 15120 8786 15148 11018
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15304 9450 15332 10610
rect 15384 9920 15436 9926
rect 15384 9862 15436 9868
rect 15396 9654 15424 9862
rect 15384 9648 15436 9654
rect 15384 9590 15436 9596
rect 15292 9444 15344 9450
rect 15292 9386 15344 9392
rect 15476 9376 15528 9382
rect 15476 9318 15528 9324
rect 15488 8974 15516 9318
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 15028 8758 15148 8786
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15028 7342 15056 8758
rect 15106 8392 15162 8401
rect 15106 8327 15162 8336
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15016 6860 15068 6866
rect 15016 6802 15068 6808
rect 15028 4865 15056 6802
rect 15014 4856 15070 4865
rect 15014 4791 15070 4800
rect 15120 3398 15148 8327
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 4570 15240 7142
rect 15304 5953 15332 8774
rect 15580 7886 15608 13194
rect 15764 11150 15792 15846
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15948 12986 15976 13194
rect 15936 12980 15988 12986
rect 15936 12922 15988 12928
rect 15752 11144 15804 11150
rect 15752 11086 15804 11092
rect 15936 11076 15988 11082
rect 15936 11018 15988 11024
rect 15660 10600 15712 10606
rect 15660 10542 15712 10548
rect 15672 9722 15700 10542
rect 15844 10464 15896 10470
rect 15844 10406 15896 10412
rect 15856 9994 15884 10406
rect 15844 9988 15896 9994
rect 15844 9930 15896 9936
rect 15856 9722 15884 9930
rect 15660 9716 15712 9722
rect 15660 9658 15712 9664
rect 15844 9716 15896 9722
rect 15844 9658 15896 9664
rect 15948 9382 15976 11018
rect 16120 9920 16172 9926
rect 16120 9862 16172 9868
rect 16132 9586 16160 9862
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15936 9172 15988 9178
rect 15856 9132 15936 9160
rect 15856 8362 15884 9132
rect 15936 9114 15988 9120
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15844 8356 15896 8362
rect 15844 8298 15896 8304
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 15476 7880 15528 7886
rect 15476 7822 15528 7828
rect 15568 7880 15620 7886
rect 15568 7822 15620 7828
rect 15488 6934 15516 7822
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15476 6384 15528 6390
rect 15476 6326 15528 6332
rect 15290 5944 15346 5953
rect 15290 5879 15346 5888
rect 15488 5710 15516 6326
rect 15476 5704 15528 5710
rect 15476 5646 15528 5652
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5166 15332 5578
rect 15580 5302 15608 7822
rect 15660 6996 15712 7002
rect 15660 6938 15712 6944
rect 15672 6798 15700 6938
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15568 5296 15620 5302
rect 15568 5238 15620 5244
rect 15292 5160 15344 5166
rect 15292 5102 15344 5108
rect 15290 4856 15346 4865
rect 15290 4791 15292 4800
rect 15344 4791 15346 4800
rect 15292 4762 15344 4768
rect 15212 4542 15332 4570
rect 15200 4480 15252 4486
rect 15200 4422 15252 4428
rect 15212 4146 15240 4422
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15212 3602 15240 4082
rect 15200 3596 15252 3602
rect 15200 3538 15252 3544
rect 15108 3392 15160 3398
rect 15108 3334 15160 3340
rect 15304 3194 15332 4542
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 15396 3126 15424 3334
rect 15488 3194 15516 3334
rect 15476 3188 15528 3194
rect 15476 3130 15528 3136
rect 15384 3120 15436 3126
rect 15384 3062 15436 3068
rect 15672 3058 15700 6734
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15764 4622 15792 6598
rect 15856 5914 15884 8298
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15844 5296 15896 5302
rect 15844 5238 15896 5244
rect 15752 4616 15804 4622
rect 15856 4593 15884 5238
rect 15948 5234 15976 7142
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15752 4558 15804 4564
rect 15842 4584 15898 4593
rect 15842 4519 15898 4528
rect 15936 4480 15988 4486
rect 15936 4422 15988 4428
rect 15948 3466 15976 4422
rect 16040 3534 16068 8298
rect 16132 7857 16160 8434
rect 16118 7848 16174 7857
rect 16118 7783 16174 7792
rect 16120 7336 16172 7342
rect 16120 7278 16172 7284
rect 16132 5370 16160 7278
rect 16120 5364 16172 5370
rect 16120 5306 16172 5312
rect 16120 5024 16172 5030
rect 16120 4966 16172 4972
rect 16132 4690 16160 4966
rect 16120 4684 16172 4690
rect 16120 4626 16172 4632
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15936 3460 15988 3466
rect 15936 3402 15988 3408
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 14936 2746 15148 2774
rect 15016 2576 15068 2582
rect 15016 2518 15068 2524
rect 14648 2440 14700 2446
rect 14648 2382 14700 2388
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 14556 2304 14608 2310
rect 14556 2246 14608 2252
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 14568 800 14596 2246
rect 15028 800 15056 2518
rect 15120 2038 15148 2746
rect 15856 2514 15884 3402
rect 16028 3392 16080 3398
rect 16028 3334 16080 3340
rect 16040 3194 16068 3334
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15936 2848 15988 2854
rect 15936 2790 15988 2796
rect 15844 2508 15896 2514
rect 15844 2450 15896 2456
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15108 2032 15160 2038
rect 15108 1974 15160 1980
rect 15488 800 15516 2246
rect 15948 800 15976 2790
rect 16224 2106 16252 15846
rect 17052 15434 17080 18566
rect 17880 18290 17908 18566
rect 17132 18284 17184 18290
rect 17132 18226 17184 18232
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17144 17134 17172 18226
rect 17684 18216 17736 18222
rect 17684 18158 17736 18164
rect 17408 18080 17460 18086
rect 17408 18022 17460 18028
rect 17420 17270 17448 18022
rect 17498 17640 17554 17649
rect 17498 17575 17554 17584
rect 17512 17542 17540 17575
rect 17500 17536 17552 17542
rect 17552 17496 17632 17524
rect 17500 17478 17552 17484
rect 17408 17264 17460 17270
rect 17408 17206 17460 17212
rect 17132 17128 17184 17134
rect 17132 17070 17184 17076
rect 17224 17128 17276 17134
rect 17224 17070 17276 17076
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17144 16998 17172 17070
rect 17132 16992 17184 16998
rect 17132 16934 17184 16940
rect 17040 15428 17092 15434
rect 17040 15370 17092 15376
rect 17144 15314 17172 16934
rect 17236 16658 17264 17070
rect 17224 16652 17276 16658
rect 17224 16594 17276 16600
rect 17512 16114 17540 17070
rect 17604 16726 17632 17496
rect 17592 16720 17644 16726
rect 17592 16662 17644 16668
rect 17696 16590 17724 18158
rect 17868 18080 17920 18086
rect 17868 18022 17920 18028
rect 17776 17196 17828 17202
rect 17776 17138 17828 17144
rect 17788 16794 17816 17138
rect 17776 16788 17828 16794
rect 17776 16730 17828 16736
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 17500 16108 17552 16114
rect 17500 16050 17552 16056
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17052 15286 17172 15314
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 16580 15020 16632 15026
rect 16580 14962 16632 14968
rect 16948 15020 17000 15026
rect 16948 14962 17000 14968
rect 16592 14414 16620 14962
rect 16960 14618 16988 14962
rect 17052 14822 17080 15286
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16948 14612 17000 14618
rect 16948 14554 17000 14560
rect 16580 14408 16632 14414
rect 16580 14350 16632 14356
rect 16948 14408 17000 14414
rect 16948 14350 17000 14356
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 16304 13932 16356 13938
rect 16304 13874 16356 13880
rect 16316 12442 16344 13874
rect 16960 13546 16988 14350
rect 17052 14074 17080 14758
rect 17224 14544 17276 14550
rect 17316 14544 17368 14550
rect 17224 14486 17276 14492
rect 17314 14512 17316 14521
rect 17368 14512 17370 14521
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17144 13802 17172 14282
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 16960 13530 17080 13546
rect 16948 13524 17080 13530
rect 17000 13518 17080 13524
rect 16948 13466 17000 13472
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16960 12986 16988 13330
rect 17052 12986 17080 13518
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 17040 12980 17092 12986
rect 17040 12922 17092 12928
rect 17144 12782 17172 13738
rect 17132 12776 17184 12782
rect 17132 12718 17184 12724
rect 16396 12708 16448 12714
rect 16396 12650 16448 12656
rect 16304 12436 16356 12442
rect 16304 12378 16356 12384
rect 16408 11558 16436 12650
rect 16948 12436 17000 12442
rect 17236 12434 17264 14486
rect 17314 14447 17370 14456
rect 17328 14278 17356 14447
rect 17316 14272 17368 14278
rect 17316 14214 17368 14220
rect 17316 13728 17368 13734
rect 17316 13670 17368 13676
rect 17328 12866 17356 13670
rect 17420 13326 17448 15846
rect 17512 15502 17540 16050
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 17512 15094 17540 15438
rect 17500 15088 17552 15094
rect 17500 15030 17552 15036
rect 17500 13864 17552 13870
rect 17500 13806 17552 13812
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17408 13184 17460 13190
rect 17408 13126 17460 13132
rect 17420 12986 17448 13126
rect 17512 12986 17540 13806
rect 17408 12980 17460 12986
rect 17408 12922 17460 12928
rect 17500 12980 17552 12986
rect 17500 12922 17552 12928
rect 17328 12838 17540 12866
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 16948 12378 17000 12384
rect 17144 12406 17264 12434
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 16396 11552 16448 11558
rect 16396 11494 16448 11500
rect 16960 11014 16988 12378
rect 17038 12200 17094 12209
rect 17038 12135 17094 12144
rect 17052 11150 17080 12135
rect 17144 11286 17172 12406
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 11694 17264 12038
rect 17328 11898 17356 12582
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17420 11898 17448 12038
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17408 11892 17460 11898
rect 17408 11834 17460 11840
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 17132 11280 17184 11286
rect 17132 11222 17184 11228
rect 17040 11144 17092 11150
rect 17040 11086 17092 11092
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16304 10668 16356 10674
rect 16304 10610 16356 10616
rect 16316 10130 16344 10610
rect 16408 10130 16436 10950
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16960 10554 16988 10950
rect 16868 10526 16988 10554
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 17040 10532 17092 10538
rect 16304 10124 16356 10130
rect 16304 10066 16356 10072
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9518 16436 10066
rect 16868 9994 16896 10526
rect 17040 10474 17092 10480
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16856 9988 16908 9994
rect 16856 9930 16908 9936
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 16764 9580 16816 9586
rect 16764 9522 16816 9528
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16776 8974 16804 9522
rect 16764 8968 16816 8974
rect 16764 8910 16816 8916
rect 16396 8900 16448 8906
rect 16396 8842 16448 8848
rect 16408 8498 16436 8842
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16396 8492 16448 8498
rect 16396 8434 16448 8440
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 16960 7546 16988 10406
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 16580 7404 16632 7410
rect 16580 7346 16632 7352
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16396 7336 16448 7342
rect 16396 7278 16448 7284
rect 16304 6792 16356 6798
rect 16304 6734 16356 6740
rect 16316 6186 16344 6734
rect 16408 6390 16436 7278
rect 16592 6798 16620 7346
rect 16960 7002 16988 7346
rect 17052 7177 17080 10474
rect 17144 10266 17172 10542
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17512 10169 17540 12838
rect 17604 11898 17632 16526
rect 17696 16454 17724 16526
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17684 15700 17736 15706
rect 17684 15642 17736 15648
rect 17696 14550 17724 15642
rect 17684 14544 17736 14550
rect 17684 14486 17736 14492
rect 17788 13274 17816 16730
rect 17880 16658 17908 18022
rect 17972 17338 18000 19314
rect 18064 18222 18092 20198
rect 18800 20058 18828 20402
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 19536 20058 19564 20402
rect 18788 20052 18840 20058
rect 18788 19994 18840 20000
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 20272 19990 20300 21247
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20444 20392 20496 20398
rect 20444 20334 20496 20340
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 18328 19848 18380 19854
rect 18328 19790 18380 19796
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20076 19848 20128 19854
rect 20076 19790 20128 19796
rect 18340 19718 18368 19790
rect 18328 19712 18380 19718
rect 18328 19654 18380 19660
rect 18052 18216 18104 18222
rect 18052 18158 18104 18164
rect 18144 18216 18196 18222
rect 18144 18158 18196 18164
rect 18156 17338 18184 18158
rect 17960 17332 18012 17338
rect 17960 17274 18012 17280
rect 18144 17332 18196 17338
rect 18144 17274 18196 17280
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17868 16652 17920 16658
rect 17868 16594 17920 16600
rect 17972 16454 18000 17002
rect 17960 16448 18012 16454
rect 17880 16408 17960 16436
rect 17880 14074 17908 16408
rect 17960 16390 18012 16396
rect 18340 16250 18368 19654
rect 18708 19446 18736 19790
rect 19536 19718 19564 19790
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 18696 19440 18748 19446
rect 18696 19382 18748 19388
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19536 18850 19564 19654
rect 19628 18970 19656 19722
rect 19996 19514 20024 19790
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 20088 19378 20116 19790
rect 20076 19372 20128 19378
rect 20076 19314 20128 19320
rect 20260 19372 20312 19378
rect 20260 19314 20312 19320
rect 19616 18964 19668 18970
rect 19616 18906 19668 18912
rect 19536 18822 19656 18850
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 18972 18624 19024 18630
rect 18972 18566 19024 18572
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18524 17610 18552 18022
rect 18880 17672 18932 17678
rect 18880 17614 18932 17620
rect 18512 17604 18564 17610
rect 18512 17546 18564 17552
rect 18892 17202 18920 17614
rect 18880 17196 18932 17202
rect 18880 17138 18932 17144
rect 18512 16584 18564 16590
rect 18512 16526 18564 16532
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18236 16108 18288 16114
rect 18236 16050 18288 16056
rect 17960 15496 18012 15502
rect 17958 15464 17960 15473
rect 18012 15464 18014 15473
rect 17958 15399 18014 15408
rect 18064 15162 18092 16050
rect 18144 15428 18196 15434
rect 18144 15370 18196 15376
rect 18052 15156 18104 15162
rect 18052 15098 18104 15104
rect 17960 14612 18012 14618
rect 17960 14554 18012 14560
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17880 13530 17908 14010
rect 17972 13802 18000 14554
rect 18064 14482 18092 15098
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 18064 13870 18092 14418
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 17960 13796 18012 13802
rect 17960 13738 18012 13744
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17972 13394 18000 13738
rect 17960 13388 18012 13394
rect 17960 13330 18012 13336
rect 17696 13246 17816 13274
rect 17696 12442 17724 13246
rect 17868 12844 17920 12850
rect 17868 12786 17920 12792
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 17788 12646 17816 12718
rect 17776 12640 17828 12646
rect 17776 12582 17828 12588
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17880 12238 17908 12786
rect 17958 12472 18014 12481
rect 17958 12407 18014 12416
rect 17868 12232 17920 12238
rect 17868 12174 17920 12180
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17498 10160 17554 10169
rect 17498 10095 17554 10104
rect 17512 9160 17540 10095
rect 17604 9994 17632 11834
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17788 11286 17816 11630
rect 17776 11280 17828 11286
rect 17776 11222 17828 11228
rect 17684 11008 17736 11014
rect 17684 10950 17736 10956
rect 17696 10810 17724 10950
rect 17684 10804 17736 10810
rect 17684 10746 17736 10752
rect 17684 10600 17736 10606
rect 17684 10542 17736 10548
rect 17696 10062 17724 10542
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17696 9654 17724 9998
rect 17788 9926 17816 11222
rect 17880 11218 17908 12174
rect 17868 11212 17920 11218
rect 17868 11154 17920 11160
rect 17972 10266 18000 12407
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17776 9920 17828 9926
rect 17776 9862 17828 9868
rect 17684 9648 17736 9654
rect 17590 9616 17646 9625
rect 17684 9590 17736 9596
rect 17590 9551 17646 9560
rect 17328 9132 17540 9160
rect 17130 8664 17186 8673
rect 17328 8650 17356 9132
rect 17500 9036 17552 9042
rect 17186 8622 17356 8650
rect 17420 8996 17500 9024
rect 17130 8599 17186 8608
rect 17144 8566 17172 8599
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17224 8492 17276 8498
rect 17224 8434 17276 8440
rect 17132 8288 17184 8294
rect 17132 8230 17184 8236
rect 17038 7168 17094 7177
rect 17038 7103 17094 7112
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16580 6792 16632 6798
rect 16580 6734 16632 6740
rect 17040 6792 17092 6798
rect 17144 6769 17172 8230
rect 17040 6734 17092 6740
rect 17130 6760 17186 6769
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16396 6384 16448 6390
rect 16396 6326 16448 6332
rect 16948 6248 17000 6254
rect 16948 6190 17000 6196
rect 16304 6180 16356 6186
rect 16304 6122 16356 6128
rect 16960 6118 16988 6190
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16948 6112 17000 6118
rect 16948 6054 17000 6060
rect 16408 5778 16436 6054
rect 16396 5772 16448 5778
rect 16396 5714 16448 5720
rect 16684 5681 16712 6054
rect 16670 5672 16726 5681
rect 16670 5607 16726 5616
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 16960 5370 16988 6054
rect 17052 5574 17080 6734
rect 17130 6695 17186 6704
rect 17236 6497 17264 8434
rect 17314 7304 17370 7313
rect 17314 7239 17370 7248
rect 17328 6798 17356 7239
rect 17316 6792 17368 6798
rect 17316 6734 17368 6740
rect 17316 6656 17368 6662
rect 17314 6624 17316 6633
rect 17368 6624 17370 6633
rect 17314 6559 17370 6568
rect 17222 6488 17278 6497
rect 17222 6423 17278 6432
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 17144 5370 17172 6190
rect 16396 5364 16448 5370
rect 16396 5306 16448 5312
rect 16948 5364 17000 5370
rect 16948 5306 17000 5312
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16316 3942 16344 4558
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16316 2990 16344 3878
rect 16408 3398 16436 5306
rect 17040 5296 17092 5302
rect 17038 5264 17040 5273
rect 17092 5264 17094 5273
rect 17038 5199 17094 5208
rect 16948 5160 17000 5166
rect 16946 5128 16948 5137
rect 17000 5128 17002 5137
rect 16946 5063 17002 5072
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 16960 4146 16988 4422
rect 16948 4140 17000 4146
rect 16948 4082 17000 4088
rect 16396 3392 16448 3398
rect 16396 3334 16448 3340
rect 17132 3392 17184 3398
rect 17132 3334 17184 3340
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 17144 3126 17172 3334
rect 17132 3120 17184 3126
rect 17132 3062 17184 3068
rect 17040 3052 17092 3058
rect 17040 2994 17092 3000
rect 16304 2984 16356 2990
rect 16304 2926 16356 2932
rect 16672 2916 16724 2922
rect 16672 2858 16724 2864
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 16212 2100 16264 2106
rect 16212 2042 16264 2048
rect 16408 800 16436 2518
rect 16684 2446 16712 2858
rect 16672 2440 16724 2446
rect 16672 2382 16724 2388
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 17052 1970 17080 2994
rect 17236 2961 17264 6423
rect 17314 5808 17370 5817
rect 17314 5743 17370 5752
rect 17328 3058 17356 5743
rect 17420 4622 17448 8996
rect 17500 8978 17552 8984
rect 17604 8974 17632 9551
rect 17592 8968 17644 8974
rect 17592 8910 17644 8916
rect 17592 8832 17644 8838
rect 17592 8774 17644 8780
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 17512 6497 17540 6598
rect 17498 6488 17554 6497
rect 17498 6423 17554 6432
rect 17604 5760 17632 8774
rect 17696 8566 17724 9590
rect 18064 9568 18092 11494
rect 18156 11336 18184 15370
rect 18248 15094 18276 16050
rect 18524 15910 18552 16526
rect 18604 16176 18656 16182
rect 18604 16118 18656 16124
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18512 15904 18564 15910
rect 18512 15846 18564 15852
rect 18432 15638 18460 15846
rect 18328 15632 18380 15638
rect 18328 15574 18380 15580
rect 18420 15632 18472 15638
rect 18420 15574 18472 15580
rect 18236 15088 18288 15094
rect 18236 15030 18288 15036
rect 18340 13954 18368 15574
rect 18432 15434 18460 15574
rect 18420 15428 18472 15434
rect 18420 15370 18472 15376
rect 18524 14958 18552 15846
rect 18512 14952 18564 14958
rect 18512 14894 18564 14900
rect 18420 14816 18472 14822
rect 18420 14758 18472 14764
rect 18432 14074 18460 14758
rect 18512 14612 18564 14618
rect 18512 14554 18564 14560
rect 18420 14068 18472 14074
rect 18420 14010 18472 14016
rect 18524 14006 18552 14554
rect 18248 13926 18368 13954
rect 18512 14000 18564 14006
rect 18512 13942 18564 13948
rect 18248 12782 18276 13926
rect 18328 13864 18380 13870
rect 18328 13806 18380 13812
rect 18340 13530 18368 13806
rect 18328 13524 18380 13530
rect 18328 13466 18380 13472
rect 18328 13320 18380 13326
rect 18328 13262 18380 13268
rect 18236 12776 18288 12782
rect 18236 12718 18288 12724
rect 18248 12306 18276 12718
rect 18236 12300 18288 12306
rect 18236 12242 18288 12248
rect 18340 11558 18368 13262
rect 18616 12434 18644 16118
rect 18788 15020 18840 15026
rect 18788 14962 18840 14968
rect 18696 14408 18748 14414
rect 18694 14376 18696 14385
rect 18748 14376 18750 14385
rect 18694 14311 18750 14320
rect 18800 14074 18828 14962
rect 18880 14952 18932 14958
rect 18880 14894 18932 14900
rect 18892 14618 18920 14894
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18880 14476 18932 14482
rect 18880 14418 18932 14424
rect 18788 14068 18840 14074
rect 18788 14010 18840 14016
rect 18696 13932 18748 13938
rect 18696 13874 18748 13880
rect 18708 13326 18736 13874
rect 18696 13320 18748 13326
rect 18696 13262 18748 13268
rect 18708 12889 18736 13262
rect 18892 13190 18920 14418
rect 18880 13184 18932 13190
rect 18880 13126 18932 13132
rect 18694 12880 18750 12889
rect 18694 12815 18750 12824
rect 18616 12406 18736 12434
rect 18420 12164 18472 12170
rect 18420 12106 18472 12112
rect 18328 11552 18380 11558
rect 18328 11494 18380 11500
rect 18156 11308 18368 11336
rect 18236 11212 18288 11218
rect 18236 11154 18288 11160
rect 18248 10742 18276 11154
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 18248 10130 18276 10678
rect 18236 10124 18288 10130
rect 18236 10066 18288 10072
rect 18142 10024 18198 10033
rect 18142 9959 18144 9968
rect 18196 9959 18198 9968
rect 18144 9930 18196 9936
rect 18248 9722 18276 10066
rect 18236 9716 18288 9722
rect 18236 9658 18288 9664
rect 18064 9540 18184 9568
rect 17776 9512 17828 9518
rect 17774 9480 17776 9489
rect 17828 9480 17830 9489
rect 17774 9415 17830 9424
rect 18052 9444 18104 9450
rect 18052 9386 18104 9392
rect 17960 9376 18012 9382
rect 17960 9318 18012 9324
rect 17972 9081 18000 9318
rect 17774 9072 17830 9081
rect 17774 9007 17830 9016
rect 17958 9072 18014 9081
rect 17958 9007 18014 9016
rect 17788 8906 17816 9007
rect 17776 8900 17828 8906
rect 17776 8842 17828 8848
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17958 8528 18014 8537
rect 17696 7954 17724 8502
rect 17958 8463 18014 8472
rect 17972 8430 18000 8463
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17776 8356 17828 8362
rect 17776 8298 17828 8304
rect 17788 7954 17816 8298
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17960 8288 18012 8294
rect 17960 8230 18012 8236
rect 17684 7948 17736 7954
rect 17684 7890 17736 7896
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 17696 7478 17724 7890
rect 17880 7886 17908 8230
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17776 7812 17828 7818
rect 17776 7754 17828 7760
rect 17684 7472 17736 7478
rect 17684 7414 17736 7420
rect 17788 7002 17816 7754
rect 17972 7546 18000 8230
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 17958 7304 18014 7313
rect 17958 7239 18014 7248
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17868 6996 17920 7002
rect 17868 6938 17920 6944
rect 17880 6798 17908 6938
rect 17972 6934 18000 7239
rect 18064 7041 18092 9386
rect 18050 7032 18106 7041
rect 18050 6967 18106 6976
rect 17960 6928 18012 6934
rect 18052 6928 18104 6934
rect 17960 6870 18012 6876
rect 18050 6896 18052 6905
rect 18104 6896 18106 6905
rect 18050 6831 18106 6840
rect 17868 6792 17920 6798
rect 17868 6734 17920 6740
rect 17960 6724 18012 6730
rect 17960 6666 18012 6672
rect 17776 6656 17828 6662
rect 17774 6624 17776 6633
rect 17828 6624 17830 6633
rect 17774 6559 17830 6568
rect 17972 6458 18000 6666
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 18156 6202 18184 9540
rect 18340 7993 18368 11308
rect 18326 7984 18382 7993
rect 18326 7919 18382 7928
rect 18234 7712 18290 7721
rect 18234 7647 18290 7656
rect 18248 6798 18276 7647
rect 18340 6798 18368 7919
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 18156 6174 18276 6202
rect 18144 6112 18196 6118
rect 18144 6054 18196 6060
rect 17604 5732 17724 5760
rect 17500 5704 17552 5710
rect 17696 5692 17724 5732
rect 17776 5704 17828 5710
rect 17696 5664 17776 5692
rect 17500 5646 17552 5652
rect 17776 5646 17828 5652
rect 17512 5302 17540 5646
rect 17592 5636 17644 5642
rect 17592 5578 17644 5584
rect 17960 5636 18012 5642
rect 17960 5578 18012 5584
rect 17604 5370 17632 5578
rect 17868 5568 17920 5574
rect 17682 5536 17738 5545
rect 17868 5510 17920 5516
rect 17682 5471 17738 5480
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17500 5296 17552 5302
rect 17500 5238 17552 5244
rect 17408 4616 17460 4622
rect 17408 4558 17460 4564
rect 17512 4214 17540 5238
rect 17696 4826 17724 5471
rect 17880 5273 17908 5510
rect 17866 5264 17922 5273
rect 17776 5228 17828 5234
rect 17972 5234 18000 5578
rect 17866 5199 17922 5208
rect 17960 5228 18012 5234
rect 17776 5170 17828 5176
rect 17960 5170 18012 5176
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 17788 4758 17816 5170
rect 17960 5092 18012 5098
rect 17960 5034 18012 5040
rect 17776 4752 17828 4758
rect 17776 4694 17828 4700
rect 17500 4208 17552 4214
rect 17500 4150 17552 4156
rect 17972 3482 18000 5034
rect 18052 4752 18104 4758
rect 18050 4720 18052 4729
rect 18104 4720 18106 4729
rect 18050 4655 18106 4664
rect 18156 4282 18184 6054
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18248 4214 18276 6174
rect 18236 4208 18288 4214
rect 18236 4150 18288 4156
rect 18326 3904 18382 3913
rect 18326 3839 18382 3848
rect 18050 3496 18106 3505
rect 17972 3454 18050 3482
rect 18050 3431 18106 3440
rect 17684 3392 17736 3398
rect 17684 3334 17736 3340
rect 17696 3194 17724 3334
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 18064 3058 18092 3431
rect 18340 3058 18368 3839
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 18052 3052 18104 3058
rect 18052 2994 18104 3000
rect 18328 3052 18380 3058
rect 18328 2994 18380 3000
rect 17960 2984 18012 2990
rect 17222 2952 17278 2961
rect 17222 2887 17278 2896
rect 17958 2952 17960 2961
rect 18012 2952 18014 2961
rect 17958 2887 18014 2896
rect 17316 2848 17368 2854
rect 17316 2790 17368 2796
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 17224 2304 17276 2310
rect 17224 2246 17276 2252
rect 17040 1964 17092 1970
rect 17040 1906 17092 1912
rect 16868 870 16988 898
rect 16868 800 16896 870
rect 10152 734 10364 762
rect 10506 0 10562 800
rect 10966 0 11022 800
rect 11426 0 11482 800
rect 11886 0 11942 800
rect 12346 0 12402 800
rect 12806 0 12862 800
rect 13266 0 13322 800
rect 13726 0 13782 800
rect 14094 0 14150 800
rect 14554 0 14610 800
rect 15014 0 15070 800
rect 15474 0 15530 800
rect 15934 0 15990 800
rect 16394 0 16450 800
rect 16854 0 16910 800
rect 16960 762 16988 870
rect 17236 762 17264 2246
rect 17328 800 17356 2790
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 17788 800 17816 2518
rect 18248 800 18276 2790
rect 18432 2774 18460 12106
rect 18604 11756 18656 11762
rect 18604 11698 18656 11704
rect 18616 10985 18644 11698
rect 18602 10976 18658 10985
rect 18602 10911 18658 10920
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18616 9586 18644 10134
rect 18708 10033 18736 12406
rect 18878 11656 18934 11665
rect 18878 11591 18934 11600
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18694 10024 18750 10033
rect 18694 9959 18750 9968
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18524 9178 18552 9522
rect 18616 9489 18644 9522
rect 18602 9480 18658 9489
rect 18602 9415 18658 9424
rect 18512 9172 18564 9178
rect 18512 9114 18564 9120
rect 18708 8650 18736 9959
rect 18800 9722 18828 10746
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18892 9194 18920 11591
rect 18984 10810 19012 18566
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 19536 17882 19564 18702
rect 19524 17876 19576 17882
rect 19524 17818 19576 17824
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 19628 16250 19656 18822
rect 19708 18080 19760 18086
rect 19708 18022 19760 18028
rect 19720 17746 19748 18022
rect 19708 17740 19760 17746
rect 19708 17682 19760 17688
rect 19616 16244 19668 16250
rect 19616 16186 19668 16192
rect 19064 16040 19116 16046
rect 19064 15982 19116 15988
rect 19076 15502 19104 15982
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 19156 15564 19208 15570
rect 19156 15506 19208 15512
rect 19064 15496 19116 15502
rect 19064 15438 19116 15444
rect 19168 14804 19196 15506
rect 19432 15360 19484 15366
rect 19432 15302 19484 15308
rect 19444 15162 19472 15302
rect 19628 15178 19656 16186
rect 19720 16017 19748 17682
rect 19892 17672 19944 17678
rect 19892 17614 19944 17620
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19812 16590 19840 17206
rect 19904 17105 19932 17614
rect 19890 17096 19946 17105
rect 19890 17031 19946 17040
rect 19800 16584 19852 16590
rect 19800 16526 19852 16532
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20180 16250 20208 16526
rect 20168 16244 20220 16250
rect 20168 16186 20220 16192
rect 19706 16008 19762 16017
rect 19706 15943 19762 15952
rect 20272 15892 20300 19314
rect 20352 19168 20404 19174
rect 20352 19110 20404 19116
rect 20364 18426 20392 19110
rect 20456 18902 20484 20334
rect 20548 20058 20576 20402
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 20640 19666 20668 22199
rect 20718 20360 20774 20369
rect 20718 20295 20720 20304
rect 20772 20295 20774 20304
rect 20720 20266 20772 20272
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 20718 19816 20774 19825
rect 20718 19751 20774 19760
rect 20732 19718 20760 19751
rect 20548 19638 20668 19666
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 20548 19514 20576 19638
rect 20536 19508 20588 19514
rect 20536 19450 20588 19456
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20536 19372 20588 19378
rect 20536 19314 20588 19320
rect 20548 18970 20576 19314
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20444 18896 20496 18902
rect 20444 18838 20496 18844
rect 20640 18465 20668 19450
rect 21284 18873 21312 19654
rect 21376 19417 21404 20198
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21270 18864 21326 18873
rect 21270 18799 21326 18808
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 20626 18456 20682 18465
rect 20352 18420 20404 18426
rect 20626 18391 20682 18400
rect 20352 18362 20404 18368
rect 20628 18284 20680 18290
rect 20628 18226 20680 18232
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20364 17882 20392 18158
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20352 17604 20404 17610
rect 20352 17546 20404 17552
rect 20364 16794 20392 17546
rect 20640 17338 20668 18226
rect 20996 18080 21048 18086
rect 21284 18057 21312 18566
rect 21364 18080 21416 18086
rect 20996 18022 21048 18028
rect 21270 18048 21326 18057
rect 20628 17332 20680 17338
rect 20628 17274 20680 17280
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20824 16794 20852 17138
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20812 16788 20864 16794
rect 20812 16730 20864 16736
rect 20352 16652 20404 16658
rect 20352 16594 20404 16600
rect 20180 15864 20300 15892
rect 19432 15156 19484 15162
rect 19628 15150 19840 15178
rect 19432 15098 19484 15104
rect 19708 15020 19760 15026
rect 19708 14962 19760 14968
rect 19524 14952 19576 14958
rect 19524 14894 19576 14900
rect 19076 14776 19196 14804
rect 19076 14550 19104 14776
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19536 14618 19564 14894
rect 19524 14612 19576 14618
rect 19524 14554 19576 14560
rect 19064 14544 19116 14550
rect 19064 14486 19116 14492
rect 19340 14408 19392 14414
rect 19340 14350 19392 14356
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 19352 14006 19380 14350
rect 19340 14000 19392 14006
rect 19340 13942 19392 13948
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19352 12850 19380 12922
rect 19340 12844 19392 12850
rect 19340 12786 19392 12792
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19536 12306 19564 13874
rect 19628 12714 19656 14350
rect 19720 13274 19748 14962
rect 19812 14346 19840 15150
rect 19892 14952 19944 14958
rect 19892 14894 19944 14900
rect 19800 14340 19852 14346
rect 19800 14282 19852 14288
rect 19904 14090 19932 14894
rect 20076 14340 20128 14346
rect 20076 14282 20128 14288
rect 19812 14062 19932 14090
rect 19812 13802 19840 14062
rect 19800 13796 19852 13802
rect 19800 13738 19852 13744
rect 19812 13394 19840 13738
rect 19800 13388 19852 13394
rect 19800 13330 19852 13336
rect 19720 13246 19932 13274
rect 19708 13184 19760 13190
rect 19708 13126 19760 13132
rect 19720 12986 19748 13126
rect 19708 12980 19760 12986
rect 19708 12922 19760 12928
rect 19904 12782 19932 13246
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19616 12708 19668 12714
rect 19616 12650 19668 12656
rect 19904 12434 19932 12718
rect 19628 12406 19932 12434
rect 19524 12300 19576 12306
rect 19524 12242 19576 12248
rect 19064 11756 19116 11762
rect 19064 11698 19116 11704
rect 18972 10804 19024 10810
rect 18972 10746 19024 10752
rect 18970 10568 19026 10577
rect 18970 10503 19026 10512
rect 18984 10062 19012 10503
rect 19076 10470 19104 11698
rect 19524 11552 19576 11558
rect 19524 11494 19576 11500
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19536 11150 19564 11494
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19536 10266 19564 10678
rect 19064 10260 19116 10266
rect 19064 10202 19116 10208
rect 19524 10260 19576 10266
rect 19524 10202 19576 10208
rect 18972 10056 19024 10062
rect 18972 9998 19024 10004
rect 18892 9166 19012 9194
rect 18880 9104 18932 9110
rect 18880 9046 18932 9052
rect 18892 8906 18920 9046
rect 18788 8900 18840 8906
rect 18788 8842 18840 8848
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18800 8673 18828 8842
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18616 8622 18736 8650
rect 18786 8664 18842 8673
rect 18524 6322 18552 8570
rect 18616 7478 18644 8622
rect 18786 8599 18842 8608
rect 18696 8492 18748 8498
rect 18696 8434 18748 8440
rect 18708 7954 18736 8434
rect 18892 8022 18920 8842
rect 18880 8016 18932 8022
rect 18880 7958 18932 7964
rect 18696 7948 18748 7954
rect 18696 7890 18748 7896
rect 18788 7880 18840 7886
rect 18694 7848 18750 7857
rect 18788 7822 18840 7828
rect 18694 7783 18750 7792
rect 18708 7546 18736 7783
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18604 7472 18656 7478
rect 18604 7414 18656 7420
rect 18602 6760 18658 6769
rect 18602 6695 18604 6704
rect 18656 6695 18658 6704
rect 18604 6666 18656 6672
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18708 6254 18736 7482
rect 18800 6633 18828 7822
rect 18984 6798 19012 9166
rect 19076 7886 19104 10202
rect 19432 10192 19484 10198
rect 19432 10134 19484 10140
rect 19156 9988 19208 9994
rect 19156 9930 19208 9936
rect 19168 9722 19196 9930
rect 19156 9716 19208 9722
rect 19156 9658 19208 9664
rect 19444 9450 19472 10134
rect 19524 9580 19576 9586
rect 19524 9522 19576 9528
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 18972 6792 19024 6798
rect 18970 6760 18972 6769
rect 19024 6760 19026 6769
rect 18970 6695 19026 6704
rect 18786 6624 18842 6633
rect 18786 6559 18842 6568
rect 18696 6248 18748 6254
rect 18696 6190 18748 6196
rect 18696 5636 18748 5642
rect 18696 5578 18748 5584
rect 18708 5370 18736 5578
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18800 4706 18828 6559
rect 18970 6488 19026 6497
rect 18970 6423 19026 6432
rect 18984 6322 19012 6423
rect 18972 6316 19024 6322
rect 18972 6258 19024 6264
rect 18880 6180 18932 6186
rect 18880 6122 18932 6128
rect 18892 5914 18920 6122
rect 18880 5908 18932 5914
rect 18880 5850 18932 5856
rect 18984 5817 19012 6258
rect 18970 5808 19026 5817
rect 18970 5743 19026 5752
rect 18972 5568 19024 5574
rect 18972 5510 19024 5516
rect 18984 5250 19012 5510
rect 18892 5234 19012 5250
rect 18880 5228 19012 5234
rect 18932 5222 19012 5228
rect 18880 5170 18932 5176
rect 18524 4678 18828 4706
rect 18524 4486 18552 4678
rect 19076 4622 19104 7686
rect 19536 7546 19564 9522
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19524 7404 19576 7410
rect 19524 7346 19576 7352
rect 19536 7206 19564 7346
rect 19524 7200 19576 7206
rect 19524 7142 19576 7148
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 19432 6724 19484 6730
rect 19432 6666 19484 6672
rect 19444 6361 19472 6666
rect 19430 6352 19486 6361
rect 19430 6287 19486 6296
rect 19536 6254 19564 7142
rect 19524 6248 19576 6254
rect 19524 6190 19576 6196
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 19248 5840 19300 5846
rect 19248 5782 19300 5788
rect 19260 5234 19288 5782
rect 19524 5704 19576 5710
rect 19524 5646 19576 5652
rect 19536 5574 19564 5646
rect 19524 5568 19576 5574
rect 19524 5510 19576 5516
rect 19248 5228 19300 5234
rect 19248 5170 19300 5176
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 19064 4616 19116 4622
rect 19064 4558 19116 4564
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18696 4480 18748 4486
rect 18696 4422 18748 4428
rect 18708 3738 18736 4422
rect 19628 4078 19656 12406
rect 20088 12186 20116 14282
rect 19812 12158 20116 12186
rect 19708 9920 19760 9926
rect 19708 9862 19760 9868
rect 19720 8974 19748 9862
rect 19812 9586 19840 12158
rect 19984 12096 20036 12102
rect 19984 12038 20036 12044
rect 19996 11898 20024 12038
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 19892 10464 19944 10470
rect 19892 10406 19944 10412
rect 19904 10198 19932 10406
rect 19892 10192 19944 10198
rect 19892 10134 19944 10140
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19996 9466 20024 11834
rect 20076 11620 20128 11626
rect 20076 11562 20128 11568
rect 19904 9438 20024 9466
rect 19800 9376 19852 9382
rect 19800 9318 19852 9324
rect 19812 9042 19840 9318
rect 19800 9036 19852 9042
rect 19800 8978 19852 8984
rect 19708 8968 19760 8974
rect 19708 8910 19760 8916
rect 19798 8936 19854 8945
rect 19798 8871 19854 8880
rect 19812 7750 19840 8871
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19720 6458 19748 7686
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19708 6452 19760 6458
rect 19708 6394 19760 6400
rect 19812 6322 19840 7278
rect 19800 6316 19852 6322
rect 19800 6258 19852 6264
rect 19616 4072 19668 4078
rect 19616 4014 19668 4020
rect 19064 3936 19116 3942
rect 19064 3878 19116 3884
rect 18970 3768 19026 3777
rect 18696 3732 18748 3738
rect 18970 3703 19026 3712
rect 18696 3674 18748 3680
rect 18984 3466 19012 3703
rect 18972 3460 19024 3466
rect 18972 3402 19024 3408
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18432 2746 18552 2774
rect 18524 2446 18552 2746
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18328 1352 18380 1358
rect 18328 1294 18380 1300
rect 18340 1057 18368 1294
rect 18326 1048 18382 1057
rect 18326 983 18382 992
rect 18616 800 18644 3334
rect 19076 800 19104 3878
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19524 3664 19576 3670
rect 19524 3606 19576 3612
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19536 800 19564 3606
rect 19800 3596 19852 3602
rect 19800 3538 19852 3544
rect 19812 2038 19840 3538
rect 19904 3058 19932 9438
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9042 20024 9318
rect 19984 9036 20036 9042
rect 19984 8978 20036 8984
rect 20088 7886 20116 11562
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20076 6724 20128 6730
rect 20076 6666 20128 6672
rect 19984 6656 20036 6662
rect 19984 6598 20036 6604
rect 19996 6390 20024 6598
rect 20088 6390 20116 6666
rect 19984 6384 20036 6390
rect 19984 6326 20036 6332
rect 20076 6384 20128 6390
rect 20076 6326 20128 6332
rect 20180 5914 20208 15864
rect 20364 14074 20392 16594
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 15706 20760 16526
rect 20720 15700 20772 15706
rect 20720 15642 20772 15648
rect 20628 15496 20680 15502
rect 20628 15438 20680 15444
rect 20640 15162 20668 15438
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20732 15026 20760 15302
rect 20720 15020 20772 15026
rect 20720 14962 20772 14968
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20444 14000 20496 14006
rect 20444 13942 20496 13948
rect 20548 13954 20576 14418
rect 20456 13546 20484 13942
rect 20548 13926 20668 13954
rect 20640 13870 20668 13926
rect 20628 13864 20680 13870
rect 20628 13806 20680 13812
rect 20456 13518 20576 13546
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20260 13252 20312 13258
rect 20260 13194 20312 13200
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20272 12986 20300 13194
rect 20260 12980 20312 12986
rect 20260 12922 20312 12928
rect 20260 12844 20312 12850
rect 20260 12786 20312 12792
rect 20272 12050 20300 12786
rect 20364 12782 20392 13194
rect 20456 12782 20484 13398
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20444 12776 20496 12782
rect 20444 12718 20496 12724
rect 20456 12306 20484 12718
rect 20548 12374 20576 13518
rect 20640 13462 20668 13806
rect 20628 13456 20680 13462
rect 20628 13398 20680 13404
rect 20904 13388 20956 13394
rect 20904 13330 20956 13336
rect 20812 12912 20864 12918
rect 20812 12854 20864 12860
rect 20536 12368 20588 12374
rect 20536 12310 20588 12316
rect 20718 12336 20774 12345
rect 20444 12300 20496 12306
rect 20718 12271 20774 12280
rect 20444 12242 20496 12248
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20536 12164 20588 12170
rect 20536 12106 20588 12112
rect 20272 12022 20484 12050
rect 20258 11928 20314 11937
rect 20258 11863 20314 11872
rect 20272 11830 20300 11863
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20260 11552 20312 11558
rect 20260 11494 20312 11500
rect 20272 9654 20300 11494
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20364 10062 20392 10542
rect 20352 10056 20404 10062
rect 20352 9998 20404 10004
rect 20456 9738 20484 12022
rect 20548 11234 20576 12106
rect 20640 11694 20668 12174
rect 20628 11688 20680 11694
rect 20628 11630 20680 11636
rect 20640 11354 20668 11630
rect 20732 11393 20760 12271
rect 20718 11384 20774 11393
rect 20628 11348 20680 11354
rect 20718 11319 20774 11328
rect 20628 11290 20680 11296
rect 20548 11206 20668 11234
rect 20536 10124 20588 10130
rect 20536 10066 20588 10072
rect 20364 9710 20484 9738
rect 20260 9648 20312 9654
rect 20260 9590 20312 9596
rect 20260 8288 20312 8294
rect 20260 8230 20312 8236
rect 20272 7954 20300 8230
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20260 6792 20312 6798
rect 20260 6734 20312 6740
rect 20168 5908 20220 5914
rect 20168 5850 20220 5856
rect 20272 5574 20300 6734
rect 20260 5568 20312 5574
rect 20260 5510 20312 5516
rect 20166 4856 20222 4865
rect 20166 4791 20222 4800
rect 19984 4752 20036 4758
rect 19984 4694 20036 4700
rect 19892 3052 19944 3058
rect 19892 2994 19944 3000
rect 19800 2032 19852 2038
rect 19798 2000 19800 2009
rect 19852 2000 19854 2009
rect 19798 1935 19854 1944
rect 19812 1909 19840 1935
rect 19996 800 20024 4694
rect 20180 4214 20208 4791
rect 20168 4208 20220 4214
rect 20168 4150 20220 4156
rect 20076 3936 20128 3942
rect 20076 3878 20128 3884
rect 20088 3641 20116 3878
rect 20074 3632 20130 3641
rect 20074 3567 20130 3576
rect 20364 3534 20392 9710
rect 20548 9586 20576 10066
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20444 9376 20496 9382
rect 20444 9318 20496 9324
rect 20456 5914 20484 9318
rect 20536 9036 20588 9042
rect 20536 8978 20588 8984
rect 20548 8498 20576 8978
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20640 8378 20668 11206
rect 20732 10062 20760 11319
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20824 9738 20852 12854
rect 20916 11898 20944 13330
rect 21008 13326 21036 18022
rect 21364 18022 21416 18028
rect 21270 17983 21326 17992
rect 21088 17536 21140 17542
rect 21088 17478 21140 17484
rect 21272 17536 21324 17542
rect 21376 17513 21404 18022
rect 21272 17478 21324 17484
rect 21362 17504 21418 17513
rect 21100 17202 21128 17478
rect 21088 17196 21140 17202
rect 21088 17138 21140 17144
rect 21284 17105 21312 17478
rect 21362 17439 21418 17448
rect 21270 17096 21326 17105
rect 21270 17031 21326 17040
rect 21088 16992 21140 16998
rect 21088 16934 21140 16940
rect 21272 16992 21324 16998
rect 21272 16934 21324 16940
rect 21100 15502 21128 16934
rect 21284 16561 21312 16934
rect 21270 16552 21326 16561
rect 21270 16487 21326 16496
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21284 16153 21312 16390
rect 21270 16144 21326 16153
rect 21270 16079 21326 16088
rect 21272 15904 21324 15910
rect 21272 15846 21324 15852
rect 21284 15609 21312 15846
rect 21270 15600 21326 15609
rect 21270 15535 21326 15544
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21272 15360 21324 15366
rect 21272 15302 21324 15308
rect 21100 14414 21128 15302
rect 21284 15201 21312 15302
rect 21270 15192 21326 15201
rect 21270 15127 21326 15136
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21284 14657 21312 14758
rect 21270 14648 21326 14657
rect 21270 14583 21326 14592
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21088 14272 21140 14278
rect 21088 14214 21140 14220
rect 21100 13938 21128 14214
rect 21088 13932 21140 13938
rect 21088 13874 21140 13880
rect 20996 13320 21048 13326
rect 20996 13262 21048 13268
rect 20996 12912 21048 12918
rect 20996 12854 21048 12860
rect 21008 12442 21036 12854
rect 21086 12744 21142 12753
rect 21086 12679 21142 12688
rect 20996 12436 21048 12442
rect 20996 12378 21048 12384
rect 20904 11892 20956 11898
rect 20904 11834 20956 11840
rect 21008 10282 21036 12378
rect 20548 8350 20668 8378
rect 20732 9710 20852 9738
rect 20916 10254 21036 10282
rect 20548 6798 20576 8350
rect 20628 8084 20680 8090
rect 20628 8026 20680 8032
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20640 6458 20668 8026
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20732 6390 20760 9710
rect 20916 8838 20944 10254
rect 20994 10160 21050 10169
rect 20994 10095 20996 10104
rect 21048 10095 21050 10104
rect 20996 10066 21048 10072
rect 21100 9874 21128 12679
rect 21192 11898 21220 14282
rect 21272 14272 21324 14278
rect 21270 14240 21272 14249
rect 21324 14240 21326 14249
rect 21270 14175 21326 14184
rect 21272 14068 21324 14074
rect 21272 14010 21324 14016
rect 21284 13841 21312 14010
rect 21270 13832 21326 13841
rect 21270 13767 21326 13776
rect 21640 13524 21692 13530
rect 21640 13466 21692 13472
rect 21270 13288 21326 13297
rect 21270 13223 21326 13232
rect 21284 13190 21312 13223
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21362 12336 21418 12345
rect 21362 12271 21418 12280
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21180 11892 21232 11898
rect 21180 11834 21232 11840
rect 21192 11354 21220 11834
rect 21180 11348 21232 11354
rect 21180 11290 21232 11296
rect 21284 10742 21312 12038
rect 21376 11150 21404 12271
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 10736 21324 10742
rect 21272 10678 21324 10684
rect 21364 10600 21416 10606
rect 21364 10542 21416 10548
rect 21100 9846 21220 9874
rect 20904 8832 20956 8838
rect 20904 8774 20956 8780
rect 20812 8560 20864 8566
rect 20812 8502 20864 8508
rect 20824 7342 20852 8502
rect 21086 8392 21142 8401
rect 21086 8327 21142 8336
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6798 20852 7142
rect 20812 6792 20864 6798
rect 20812 6734 20864 6740
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20628 6112 20680 6118
rect 20628 6054 20680 6060
rect 20444 5908 20496 5914
rect 20444 5850 20496 5856
rect 20536 5772 20588 5778
rect 20536 5714 20588 5720
rect 20548 5370 20576 5714
rect 20640 5710 20668 6054
rect 20732 5846 20760 6326
rect 20904 6248 20956 6254
rect 20902 6216 20904 6225
rect 20956 6216 20958 6225
rect 20902 6151 20958 6160
rect 20720 5840 20772 5846
rect 20720 5782 20772 5788
rect 20628 5704 20680 5710
rect 20628 5646 20680 5652
rect 20536 5364 20588 5370
rect 20536 5306 20588 5312
rect 20548 5234 20576 5306
rect 20536 5228 20588 5234
rect 20536 5170 20588 5176
rect 20536 4072 20588 4078
rect 20536 4014 20588 4020
rect 20718 4040 20774 4049
rect 20444 4004 20496 4010
rect 20444 3946 20496 3952
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20074 3360 20130 3369
rect 20074 3295 20130 3304
rect 20088 3058 20116 3295
rect 20076 3052 20128 3058
rect 20076 2994 20128 3000
rect 20088 921 20116 2994
rect 20260 2440 20312 2446
rect 20260 2382 20312 2388
rect 20272 1329 20300 2382
rect 20258 1320 20314 1329
rect 20258 1255 20314 1264
rect 20074 912 20130 921
rect 20074 847 20130 856
rect 16960 734 17264 762
rect 17314 0 17370 800
rect 17774 0 17830 800
rect 18234 0 18290 800
rect 18602 0 18658 800
rect 19062 0 19118 800
rect 19522 0 19578 800
rect 19982 0 20038 800
rect 20272 241 20300 1255
rect 20456 800 20484 3946
rect 20548 2106 20576 4014
rect 20718 3975 20774 3984
rect 20626 3496 20682 3505
rect 20626 3431 20628 3440
rect 20680 3431 20682 3440
rect 20628 3402 20680 3408
rect 20732 2990 20760 3975
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 20720 2984 20772 2990
rect 20720 2926 20772 2932
rect 20536 2100 20588 2106
rect 20536 2042 20588 2048
rect 20548 1601 20576 2042
rect 20534 1592 20590 1601
rect 20534 1527 20590 1536
rect 20916 800 20944 3130
rect 21100 3058 21128 8327
rect 21192 7546 21220 9846
rect 21376 9518 21404 10542
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21376 8566 21404 9454
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21376 7478 21404 7686
rect 21364 7472 21416 7478
rect 21364 7414 21416 7420
rect 21180 7336 21232 7342
rect 21180 7278 21232 7284
rect 21192 6780 21220 7278
rect 21272 6792 21324 6798
rect 21192 6752 21272 6780
rect 21192 5302 21220 6752
rect 21272 6734 21324 6740
rect 21180 5296 21232 5302
rect 21180 5238 21232 5244
rect 21192 4690 21220 5238
rect 21272 5024 21324 5030
rect 21272 4966 21324 4972
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21284 4622 21312 4966
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21364 3120 21416 3126
rect 21364 3062 21416 3068
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21270 2544 21326 2553
rect 21270 2479 21326 2488
rect 21284 2446 21312 2479
rect 21272 2440 21324 2446
rect 21272 2382 21324 2388
rect 21376 800 21404 3062
rect 21468 2514 21496 8774
rect 21652 3602 21680 13466
rect 21824 6724 21876 6730
rect 21824 6666 21876 6672
rect 21640 3596 21692 3602
rect 21640 3538 21692 3544
rect 21456 2508 21508 2514
rect 21456 2450 21508 2456
rect 21836 800 21864 6666
rect 22284 3732 22336 3738
rect 22284 3674 22336 3680
rect 22296 800 22324 3674
rect 22744 3052 22796 3058
rect 22744 2994 22796 3000
rect 22756 800 22784 2994
rect 20258 232 20314 241
rect 20258 167 20314 176
rect 20442 0 20498 800
rect 20902 0 20958 800
rect 21362 0 21418 800
rect 21822 0 21878 800
rect 22282 0 22338 800
rect 22742 0 22798 800
<< via2 >>
rect 4526 22616 4582 22672
rect 2042 22208 2098 22264
rect 1490 21664 1546 21720
rect 1950 20712 2006 20768
rect 2870 21256 2926 21312
rect 2778 20324 2834 20360
rect 2778 20304 2780 20324
rect 2780 20304 2832 20324
rect 2832 20304 2834 20324
rect 18694 22616 18750 22672
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 2042 19760 2098 19816
rect 1490 19352 1546 19408
rect 2686 19372 2742 19408
rect 2686 19352 2688 19372
rect 2688 19352 2740 19372
rect 2740 19352 2742 19372
rect 1490 18808 1546 18864
rect 938 16224 994 16280
rect 202 15816 258 15872
rect 938 15272 994 15328
rect 938 6740 940 6760
rect 940 6740 992 6760
rect 992 6740 994 6760
rect 938 6704 994 6740
rect 938 4836 940 4856
rect 940 4836 992 4856
rect 992 4836 994 4856
rect 938 4800 994 4836
rect 1214 4528 1270 4584
rect 202 3168 258 3224
rect 18 2216 74 2272
rect 1490 18400 1546 18456
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 2134 18128 2190 18184
rect 1490 18028 1492 18048
rect 1492 18028 1544 18048
rect 1544 18028 1546 18048
rect 1490 17992 1546 18028
rect 1490 17484 1492 17504
rect 1492 17484 1544 17504
rect 1544 17484 1546 17504
rect 1490 17448 1546 17484
rect 1490 17060 1546 17096
rect 1490 17040 1492 17060
rect 1492 17040 1544 17060
rect 1544 17040 1546 17060
rect 1490 16088 1546 16144
rect 1490 15544 1546 15600
rect 2134 16496 2190 16552
rect 1490 15136 1546 15192
rect 1490 14592 1546 14648
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1490 13796 1546 13832
rect 1490 13776 1492 13796
rect 1492 13776 1544 13796
rect 1544 13776 1546 13796
rect 1398 13368 1454 13424
rect 1490 13232 1546 13288
rect 1582 12280 1638 12336
rect 1582 11872 1638 11928
rect 1582 11328 1638 11384
rect 1950 12824 2006 12880
rect 1766 12164 1822 12200
rect 1766 12144 1768 12164
rect 1768 12144 1820 12164
rect 1820 12144 1822 12164
rect 1674 10376 1730 10432
rect 1674 9988 1730 10024
rect 1674 9968 1676 9988
rect 1676 9968 1728 9988
rect 1728 9968 1730 9988
rect 1582 9424 1638 9480
rect 1674 8608 1730 8664
rect 1490 8064 1546 8120
rect 1582 6840 1638 6896
rect 1582 6160 1638 6216
rect 1674 5752 1730 5808
rect 1490 4120 1546 4176
rect 1858 10124 1914 10160
rect 1858 10104 1860 10124
rect 1860 10104 1912 10124
rect 1912 10104 1914 10124
rect 1858 8336 1914 8392
rect 1858 7520 1914 7576
rect 1950 7384 2006 7440
rect 1858 6432 1914 6488
rect 2226 8880 2282 8936
rect 2226 7656 2282 7712
rect 2778 13232 2834 13288
rect 2686 11872 2742 11928
rect 3146 12552 3202 12608
rect 2502 9560 2558 9616
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 4066 16768 4122 16824
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 5814 19352 5870 19408
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3514 12688 3570 12744
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3330 10920 3386 10976
rect 3606 10648 3662 10704
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 2778 7248 2834 7304
rect 2226 6840 2282 6896
rect 2226 4684 2282 4720
rect 2226 4664 2228 4684
rect 2228 4664 2280 4684
rect 2280 4664 2282 4684
rect 1858 4528 1914 4584
rect 2318 3596 2374 3632
rect 2962 6568 3018 6624
rect 3054 5208 3110 5264
rect 2318 3576 2320 3596
rect 2320 3576 2372 3596
rect 2372 3576 2374 3596
rect 2870 3576 2926 3632
rect 2778 2896 2834 2952
rect 2134 992 2190 1048
rect 3514 9424 3570 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3422 8880 3478 8936
rect 4066 15680 4122 15736
rect 4158 15272 4214 15328
rect 4066 15136 4122 15192
rect 4526 13232 4582 13288
rect 4526 12960 4582 13016
rect 4434 12824 4490 12880
rect 4434 12280 4490 12336
rect 3330 8472 3386 8528
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3238 6976 3294 7032
rect 3422 7112 3478 7168
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 4710 13776 4766 13832
rect 5078 15816 5134 15872
rect 4986 14184 5042 14240
rect 4802 12280 4858 12336
rect 4250 8880 4306 8936
rect 3790 6160 3846 6216
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3330 5480 3386 5536
rect 3146 4392 3202 4448
rect 3330 2624 3386 2680
rect 3054 2488 3110 2544
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3974 4800 4030 4856
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3790 3440 3846 3496
rect 4158 3984 4214 4040
rect 4342 6568 4398 6624
rect 4434 5888 4490 5944
rect 4710 7792 4766 7848
rect 4986 9832 5042 9888
rect 4986 8880 5042 8936
rect 4802 6432 4858 6488
rect 4342 3848 4398 3904
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 3422 2352 3478 2408
rect 3238 176 3294 232
rect 4618 3596 4674 3632
rect 4618 3576 4620 3596
rect 4620 3576 4672 3596
rect 4672 3576 4674 3596
rect 4526 2488 4582 2544
rect 3882 1944 3938 2000
rect 4066 1536 4122 1592
rect 3422 584 3478 640
rect 4986 3460 5042 3496
rect 4986 3440 4988 3460
rect 4988 3440 5040 3460
rect 5040 3440 5042 3460
rect 4986 3168 5042 3224
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 5538 15972 5594 16008
rect 5538 15952 5540 15972
rect 5540 15952 5592 15972
rect 5592 15952 5594 15972
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 5446 12416 5502 12472
rect 5446 11872 5502 11928
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6458 13812 6460 13832
rect 6460 13812 6512 13832
rect 6512 13812 6514 13832
rect 6458 13776 6514 13812
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5722 12280 5778 12336
rect 5630 10512 5686 10568
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 5446 6432 5502 6488
rect 5446 3304 5502 3360
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5998 9832 6054 9888
rect 5722 5788 5724 5808
rect 5724 5788 5776 5808
rect 5776 5788 5778 5808
rect 5722 5752 5778 5788
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 7746 18128 7802 18184
rect 7470 16632 7526 16688
rect 7286 15700 7342 15736
rect 7286 15680 7288 15700
rect 7288 15680 7340 15700
rect 7340 15680 7342 15700
rect 6734 13640 6790 13696
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 7470 13640 7526 13696
rect 7378 11056 7434 11112
rect 7102 10648 7158 10704
rect 6366 8200 6422 8256
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6090 6296 6146 6352
rect 6182 6024 6238 6080
rect 5722 5208 5778 5264
rect 6642 6196 6644 6216
rect 6644 6196 6696 6216
rect 6696 6196 6698 6216
rect 6642 6160 6698 6196
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 7010 7248 7066 7304
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6458 5228 6514 5264
rect 6458 5208 6460 5228
rect 6460 5208 6512 5228
rect 6512 5208 6514 5228
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6918 5888 6974 5944
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 7010 4564 7012 4584
rect 7012 4564 7064 4584
rect 7064 4564 7066 4584
rect 7010 4528 7066 4564
rect 6918 3052 6974 3088
rect 6918 3032 6920 3052
rect 6920 3032 6972 3052
rect 6972 3032 6974 3052
rect 6918 2896 6974 2952
rect 7378 9460 7380 9480
rect 7380 9460 7432 9480
rect 7432 9460 7434 9480
rect 7378 9424 7434 9460
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9586 17076 9588 17096
rect 9588 17076 9640 17096
rect 9640 17076 9642 17096
rect 9586 17040 9642 17076
rect 9126 16108 9182 16144
rect 9126 16088 9128 16108
rect 9128 16088 9180 16108
rect 9180 16088 9182 16108
rect 8206 13912 8262 13968
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9494 15544 9550 15600
rect 9310 15428 9366 15464
rect 9310 15408 9312 15428
rect 9312 15408 9364 15428
rect 9364 15408 9366 15428
rect 8206 11872 8262 11928
rect 8022 10512 8078 10568
rect 7286 5616 7342 5672
rect 7470 5616 7526 5672
rect 7562 4664 7618 4720
rect 7746 3984 7802 4040
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9678 15408 9734 15464
rect 9862 15272 9918 15328
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 9126 12416 9182 12472
rect 8942 12044 8944 12064
rect 8944 12044 8996 12064
rect 8996 12044 8998 12064
rect 8942 12008 8998 12044
rect 9126 12280 9182 12336
rect 8850 11600 8906 11656
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8482 9424 8538 9480
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8114 4120 8170 4176
rect 7838 3304 7894 3360
rect 8482 3848 8538 3904
rect 8482 2896 8538 2952
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 20626 22208 20682 22264
rect 19614 21664 19670 21720
rect 20258 21256 20314 21312
rect 20166 20712 20222 20768
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 9954 14456 10010 14512
rect 10690 15852 10692 15872
rect 10692 15852 10744 15872
rect 10744 15852 10746 15872
rect 10690 15816 10746 15852
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 10598 14320 10654 14376
rect 11058 15408 11114 15464
rect 9494 12416 9550 12472
rect 9586 12008 9642 12064
rect 9586 11872 9642 11928
rect 9402 11600 9458 11656
rect 9770 9424 9826 9480
rect 9494 8744 9550 8800
rect 9678 8336 9734 8392
rect 9586 8064 9642 8120
rect 9402 7384 9458 7440
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9218 3984 9274 4040
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 9402 2644 9458 2680
rect 9402 2624 9404 2644
rect 9404 2624 9456 2644
rect 9456 2624 9458 2644
rect 10322 10240 10378 10296
rect 10138 5616 10194 5672
rect 10598 9580 10654 9616
rect 10598 9560 10600 9580
rect 10600 9560 10652 9580
rect 10652 9560 10654 9580
rect 10506 3712 10562 3768
rect 11058 12280 11114 12336
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11886 15952 11942 16008
rect 12162 17604 12218 17640
rect 12162 17584 12164 17604
rect 12164 17584 12216 17604
rect 12216 17584 12218 17604
rect 12254 15952 12310 16008
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11702 12824 11758 12880
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11242 11192 11298 11248
rect 10874 6840 10930 6896
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11426 10260 11482 10296
rect 11426 10240 11428 10260
rect 11428 10240 11480 10260
rect 11480 10240 11482 10260
rect 11242 10104 11298 10160
rect 11150 9016 11206 9072
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 12530 13812 12532 13832
rect 12532 13812 12584 13832
rect 12584 13812 12586 13832
rect 12530 13776 12586 13812
rect 12254 13388 12310 13424
rect 12254 13368 12256 13388
rect 12256 13368 12308 13388
rect 12308 13368 12310 13388
rect 12346 12960 12402 13016
rect 11978 7928 12034 7984
rect 12162 6432 12218 6488
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11978 6024 12034 6080
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12530 5752 12586 5808
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 12714 12824 12770 12880
rect 13082 13812 13084 13832
rect 13084 13812 13136 13832
rect 13136 13812 13138 13832
rect 13082 13776 13138 13812
rect 12806 10532 12862 10568
rect 12806 10512 12808 10532
rect 12808 10512 12860 10532
rect 12860 10512 12862 10532
rect 13358 13776 13414 13832
rect 13358 12688 13414 12744
rect 13266 12552 13322 12608
rect 13174 9560 13230 9616
rect 12714 8472 12770 8528
rect 12898 7928 12954 7984
rect 13266 8336 13322 8392
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 14738 17040 14794 17096
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 14462 12416 14518 12472
rect 13726 12144 13782 12200
rect 13634 11600 13690 11656
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14370 11192 14426 11248
rect 13634 11056 13690 11112
rect 13542 10648 13598 10704
rect 13542 8880 13598 8936
rect 13542 8608 13598 8664
rect 13358 7248 13414 7304
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16026 16668 16028 16688
rect 16028 16668 16080 16688
rect 16080 16668 16082 16688
rect 16026 16632 16082 16668
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 14922 14320 14978 14376
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13634 5752 13690 5808
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 14462 5888 14518 5944
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13726 3984 13782 4040
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 13634 3612 13636 3632
rect 13636 3612 13688 3632
rect 13688 3612 13690 3632
rect 13634 3576 13690 3612
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14646 6976 14702 7032
rect 14830 3032 14886 3088
rect 15474 13912 15530 13968
rect 15658 13368 15714 13424
rect 15474 12960 15530 13016
rect 15014 8880 15070 8936
rect 15106 8336 15162 8392
rect 15014 4800 15070 4856
rect 15290 5888 15346 5944
rect 15290 4820 15346 4856
rect 15290 4800 15292 4820
rect 15292 4800 15344 4820
rect 15344 4800 15346 4820
rect 15842 4528 15898 4584
rect 16118 7792 16174 7848
rect 17498 17584 17554 17640
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 17314 14492 17316 14512
rect 17316 14492 17368 14512
rect 17368 14492 17370 14512
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 17314 14456 17370 14492
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 17038 12144 17094 12200
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 17958 15444 17960 15464
rect 17960 15444 18012 15464
rect 18012 15444 18014 15464
rect 17958 15408 18014 15444
rect 17958 12416 18014 12472
rect 17498 10104 17554 10160
rect 17590 9560 17646 9616
rect 17130 8608 17186 8664
rect 17038 7112 17094 7168
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16670 5616 16726 5672
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 17130 6704 17186 6760
rect 17314 7248 17370 7304
rect 17314 6604 17316 6624
rect 17316 6604 17368 6624
rect 17368 6604 17370 6624
rect 17314 6568 17370 6604
rect 17222 6432 17278 6488
rect 17038 5244 17040 5264
rect 17040 5244 17092 5264
rect 17092 5244 17094 5264
rect 17038 5208 17094 5244
rect 16946 5108 16948 5128
rect 16948 5108 17000 5128
rect 17000 5108 17002 5128
rect 16946 5072 17002 5108
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17314 5752 17370 5808
rect 17498 6432 17554 6488
rect 18694 14356 18696 14376
rect 18696 14356 18748 14376
rect 18748 14356 18750 14376
rect 18694 14320 18750 14356
rect 18694 12824 18750 12880
rect 18142 9988 18198 10024
rect 18142 9968 18144 9988
rect 18144 9968 18196 9988
rect 18196 9968 18198 9988
rect 17774 9460 17776 9480
rect 17776 9460 17828 9480
rect 17828 9460 17830 9480
rect 17774 9424 17830 9460
rect 17774 9016 17830 9072
rect 17958 9016 18014 9072
rect 17958 8472 18014 8528
rect 17958 7248 18014 7304
rect 18050 6976 18106 7032
rect 18050 6876 18052 6896
rect 18052 6876 18104 6896
rect 18104 6876 18106 6896
rect 18050 6840 18106 6876
rect 17774 6604 17776 6624
rect 17776 6604 17828 6624
rect 17828 6604 17830 6624
rect 17774 6568 17830 6604
rect 18326 7928 18382 7984
rect 18234 7656 18290 7712
rect 17682 5480 17738 5536
rect 17866 5208 17922 5264
rect 18050 4700 18052 4720
rect 18052 4700 18104 4720
rect 18104 4700 18106 4720
rect 18050 4664 18106 4700
rect 18326 3848 18382 3904
rect 18050 3440 18106 3496
rect 17222 2896 17278 2952
rect 17958 2932 17960 2952
rect 17960 2932 18012 2952
rect 18012 2932 18014 2952
rect 17958 2896 18014 2932
rect 18602 10920 18658 10976
rect 18878 11600 18934 11656
rect 18694 9968 18750 10024
rect 18602 9424 18658 9480
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19890 17040 19946 17096
rect 19706 15952 19762 16008
rect 20718 20324 20774 20360
rect 20718 20304 20720 20324
rect 20720 20304 20772 20324
rect 20772 20304 20774 20324
rect 20718 19760 20774 19816
rect 21362 19352 21418 19408
rect 21270 18808 21326 18864
rect 20626 18400 20682 18456
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18970 10512 19026 10568
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 18786 8608 18842 8664
rect 18694 7792 18750 7848
rect 18602 6724 18658 6760
rect 18602 6704 18604 6724
rect 18604 6704 18656 6724
rect 18656 6704 18658 6724
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 18970 6740 18972 6760
rect 18972 6740 19024 6760
rect 19024 6740 19026 6760
rect 18970 6704 19026 6740
rect 18786 6568 18842 6624
rect 18970 6432 19026 6488
rect 18970 5752 19026 5808
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19430 6296 19486 6352
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 19798 8880 19854 8936
rect 18970 3712 19026 3768
rect 18326 992 18382 1048
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 20718 12280 20774 12336
rect 20258 11872 20314 11928
rect 20718 11328 20774 11384
rect 20166 4800 20222 4856
rect 19798 1980 19800 2000
rect 19800 1980 19852 2000
rect 19852 1980 19854 2000
rect 19798 1944 19854 1980
rect 20074 3576 20130 3632
rect 21270 17992 21326 18048
rect 21362 17448 21418 17504
rect 21270 17040 21326 17096
rect 21270 16496 21326 16552
rect 21270 16088 21326 16144
rect 21270 15544 21326 15600
rect 21270 15136 21326 15192
rect 21270 14592 21326 14648
rect 21086 12688 21142 12744
rect 20994 10124 21050 10160
rect 20994 10104 20996 10124
rect 20996 10104 21048 10124
rect 21048 10104 21050 10124
rect 21270 14220 21272 14240
rect 21272 14220 21324 14240
rect 21324 14220 21326 14240
rect 21270 14184 21326 14220
rect 21270 13776 21326 13832
rect 21270 13232 21326 13288
rect 21362 12280 21418 12336
rect 21086 8336 21142 8392
rect 20902 6196 20904 6216
rect 20904 6196 20956 6216
rect 20956 6196 20958 6216
rect 20902 6160 20958 6196
rect 20074 3304 20130 3360
rect 20258 1264 20314 1320
rect 20074 856 20130 912
rect 20718 3984 20774 4040
rect 20626 3460 20682 3496
rect 20626 3440 20628 3460
rect 20628 3440 20680 3460
rect 20680 3440 20682 3460
rect 20534 1536 20590 1592
rect 21270 2488 21326 2544
rect 20258 176 20314 232
<< metal3 >>
rect 0 22674 800 22704
rect 4521 22674 4587 22677
rect 0 22672 4587 22674
rect 0 22616 4526 22672
rect 4582 22616 4587 22672
rect 0 22614 4587 22616
rect 0 22584 800 22614
rect 4521 22611 4587 22614
rect 18689 22674 18755 22677
rect 22200 22674 23000 22704
rect 18689 22672 23000 22674
rect 18689 22616 18694 22672
rect 18750 22616 23000 22672
rect 18689 22614 23000 22616
rect 18689 22611 18755 22614
rect 22200 22584 23000 22614
rect 0 22266 800 22296
rect 2037 22266 2103 22269
rect 0 22264 2103 22266
rect 0 22208 2042 22264
rect 2098 22208 2103 22264
rect 0 22206 2103 22208
rect 0 22176 800 22206
rect 2037 22203 2103 22206
rect 20621 22266 20687 22269
rect 22200 22266 23000 22296
rect 20621 22264 23000 22266
rect 20621 22208 20626 22264
rect 20682 22208 23000 22264
rect 20621 22206 23000 22208
rect 20621 22203 20687 22206
rect 22200 22176 23000 22206
rect 0 21722 800 21752
rect 1485 21722 1551 21725
rect 0 21720 1551 21722
rect 0 21664 1490 21720
rect 1546 21664 1551 21720
rect 0 21662 1551 21664
rect 0 21632 800 21662
rect 1485 21659 1551 21662
rect 19609 21722 19675 21725
rect 22200 21722 23000 21752
rect 19609 21720 23000 21722
rect 19609 21664 19614 21720
rect 19670 21664 23000 21720
rect 19609 21662 23000 21664
rect 19609 21659 19675 21662
rect 22200 21632 23000 21662
rect 0 21314 800 21344
rect 2865 21314 2931 21317
rect 0 21312 2931 21314
rect 0 21256 2870 21312
rect 2926 21256 2931 21312
rect 0 21254 2931 21256
rect 0 21224 800 21254
rect 2865 21251 2931 21254
rect 20253 21314 20319 21317
rect 22200 21314 23000 21344
rect 20253 21312 23000 21314
rect 20253 21256 20258 21312
rect 20314 21256 23000 21312
rect 20253 21254 23000 21256
rect 20253 21251 20319 21254
rect 22200 21224 23000 21254
rect 0 20770 800 20800
rect 1945 20770 2011 20773
rect 0 20768 2011 20770
rect 0 20712 1950 20768
rect 2006 20712 2011 20768
rect 0 20710 2011 20712
rect 0 20680 800 20710
rect 1945 20707 2011 20710
rect 20161 20770 20227 20773
rect 22200 20770 23000 20800
rect 20161 20768 23000 20770
rect 20161 20712 20166 20768
rect 20222 20712 23000 20768
rect 20161 20710 23000 20712
rect 20161 20707 20227 20710
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 22200 20680 23000 20710
rect 16538 20639 16858 20640
rect 0 20362 800 20392
rect 2773 20362 2839 20365
rect 0 20360 2839 20362
rect 0 20304 2778 20360
rect 2834 20304 2839 20360
rect 0 20302 2839 20304
rect 0 20272 800 20302
rect 2773 20299 2839 20302
rect 20713 20362 20779 20365
rect 22200 20362 23000 20392
rect 20713 20360 23000 20362
rect 20713 20304 20718 20360
rect 20774 20304 23000 20360
rect 20713 20302 23000 20304
rect 20713 20299 20779 20302
rect 22200 20272 23000 20302
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 0 19818 800 19848
rect 2037 19818 2103 19821
rect 0 19816 2103 19818
rect 0 19760 2042 19816
rect 2098 19760 2103 19816
rect 0 19758 2103 19760
rect 0 19728 800 19758
rect 2037 19755 2103 19758
rect 20713 19818 20779 19821
rect 22200 19818 23000 19848
rect 20713 19816 23000 19818
rect 20713 19760 20718 19816
rect 20774 19760 23000 19816
rect 20713 19758 23000 19760
rect 20713 19755 20779 19758
rect 22200 19728 23000 19758
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 0 19410 800 19440
rect 1485 19410 1551 19413
rect 0 19408 1551 19410
rect 0 19352 1490 19408
rect 1546 19352 1551 19408
rect 0 19350 1551 19352
rect 0 19320 800 19350
rect 1485 19347 1551 19350
rect 2681 19410 2747 19413
rect 5809 19410 5875 19413
rect 2681 19408 5875 19410
rect 2681 19352 2686 19408
rect 2742 19352 5814 19408
rect 5870 19352 5875 19408
rect 2681 19350 5875 19352
rect 2681 19347 2747 19350
rect 5809 19347 5875 19350
rect 21357 19410 21423 19413
rect 22200 19410 23000 19440
rect 21357 19408 23000 19410
rect 21357 19352 21362 19408
rect 21418 19352 23000 19408
rect 21357 19350 23000 19352
rect 21357 19347 21423 19350
rect 22200 19320 23000 19350
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 0 18866 800 18896
rect 1485 18866 1551 18869
rect 0 18864 1551 18866
rect 0 18808 1490 18864
rect 1546 18808 1551 18864
rect 0 18806 1551 18808
rect 0 18776 800 18806
rect 1485 18803 1551 18806
rect 21265 18866 21331 18869
rect 22200 18866 23000 18896
rect 21265 18864 23000 18866
rect 21265 18808 21270 18864
rect 21326 18808 23000 18864
rect 21265 18806 23000 18808
rect 21265 18803 21331 18806
rect 22200 18776 23000 18806
rect 6142 18528 6462 18529
rect 0 18458 800 18488
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 18463 16858 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 20621 18458 20687 18461
rect 22200 18458 23000 18488
rect 20621 18456 23000 18458
rect 20621 18400 20626 18456
rect 20682 18400 23000 18456
rect 20621 18398 23000 18400
rect 20621 18395 20687 18398
rect 22200 18368 23000 18398
rect 2129 18186 2195 18189
rect 7741 18186 7807 18189
rect 2129 18184 7807 18186
rect 2129 18128 2134 18184
rect 2190 18128 7746 18184
rect 7802 18128 7807 18184
rect 2129 18126 7807 18128
rect 2129 18123 2195 18126
rect 7741 18123 7807 18126
rect 0 18050 800 18080
rect 1485 18050 1551 18053
rect 0 18048 1551 18050
rect 0 17992 1490 18048
rect 1546 17992 1551 18048
rect 0 17990 1551 17992
rect 0 17960 800 17990
rect 1485 17987 1551 17990
rect 21265 18050 21331 18053
rect 22200 18050 23000 18080
rect 21265 18048 23000 18050
rect 21265 17992 21270 18048
rect 21326 17992 23000 18048
rect 21265 17990 23000 17992
rect 21265 17987 21331 17990
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 22200 17960 23000 17990
rect 19137 17919 19457 17920
rect 12157 17642 12223 17645
rect 17493 17642 17559 17645
rect 12157 17640 17559 17642
rect 12157 17584 12162 17640
rect 12218 17584 17498 17640
rect 17554 17584 17559 17640
rect 12157 17582 17559 17584
rect 12157 17579 12223 17582
rect 17493 17579 17559 17582
rect 0 17506 800 17536
rect 1485 17506 1551 17509
rect 0 17504 1551 17506
rect 0 17448 1490 17504
rect 1546 17448 1551 17504
rect 0 17446 1551 17448
rect 0 17416 800 17446
rect 1485 17443 1551 17446
rect 21357 17506 21423 17509
rect 22200 17506 23000 17536
rect 21357 17504 23000 17506
rect 21357 17448 21362 17504
rect 21418 17448 23000 17504
rect 21357 17446 23000 17448
rect 21357 17443 21423 17446
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 22200 17416 23000 17446
rect 16538 17375 16858 17376
rect 0 17098 800 17128
rect 1485 17098 1551 17101
rect 0 17096 1551 17098
rect 0 17040 1490 17096
rect 1546 17040 1551 17096
rect 0 17038 1551 17040
rect 0 17008 800 17038
rect 1485 17035 1551 17038
rect 9438 17036 9444 17100
rect 9508 17098 9514 17100
rect 9581 17098 9647 17101
rect 9508 17096 9647 17098
rect 9508 17040 9586 17096
rect 9642 17040 9647 17096
rect 9508 17038 9647 17040
rect 9508 17036 9514 17038
rect 9581 17035 9647 17038
rect 14733 17098 14799 17101
rect 19885 17098 19951 17101
rect 14733 17096 19951 17098
rect 14733 17040 14738 17096
rect 14794 17040 19890 17096
rect 19946 17040 19951 17096
rect 14733 17038 19951 17040
rect 14733 17035 14799 17038
rect 19885 17035 19951 17038
rect 21265 17098 21331 17101
rect 22200 17098 23000 17128
rect 21265 17096 23000 17098
rect 21265 17040 21270 17096
rect 21326 17040 23000 17096
rect 21265 17038 23000 17040
rect 21265 17035 21331 17038
rect 22200 17008 23000 17038
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 4061 16826 4127 16829
rect 4286 16826 4292 16828
rect 4061 16824 4292 16826
rect 4061 16768 4066 16824
rect 4122 16768 4292 16824
rect 4061 16766 4292 16768
rect 4061 16763 4127 16766
rect 4286 16764 4292 16766
rect 4356 16764 4362 16828
rect 2262 16628 2268 16692
rect 2332 16690 2338 16692
rect 7465 16690 7531 16693
rect 2332 16688 7531 16690
rect 2332 16632 7470 16688
rect 7526 16632 7531 16688
rect 2332 16630 7531 16632
rect 2332 16628 2338 16630
rect 7465 16627 7531 16630
rect 16021 16692 16087 16693
rect 16021 16688 16068 16692
rect 16132 16690 16138 16692
rect 16021 16632 16026 16688
rect 16021 16628 16068 16632
rect 16132 16630 16178 16690
rect 16132 16628 16138 16630
rect 16021 16627 16087 16628
rect 0 16554 800 16584
rect 2129 16554 2195 16557
rect 0 16552 2195 16554
rect 0 16496 2134 16552
rect 2190 16496 2195 16552
rect 0 16494 2195 16496
rect 0 16464 800 16494
rect 2129 16491 2195 16494
rect 21265 16554 21331 16557
rect 22200 16554 23000 16584
rect 21265 16552 23000 16554
rect 21265 16496 21270 16552
rect 21326 16496 23000 16552
rect 21265 16494 23000 16496
rect 21265 16491 21331 16494
rect 22200 16464 23000 16494
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 933 16282 999 16285
rect 933 16280 1778 16282
rect 933 16224 938 16280
rect 994 16224 1778 16280
rect 933 16222 1778 16224
rect 933 16219 999 16222
rect 0 16146 800 16176
rect 1485 16146 1551 16149
rect 0 16144 1551 16146
rect 0 16088 1490 16144
rect 1546 16088 1551 16144
rect 0 16086 1551 16088
rect 1718 16146 1778 16222
rect 9121 16146 9187 16149
rect 1718 16144 9187 16146
rect 1718 16088 9126 16144
rect 9182 16088 9187 16144
rect 1718 16086 9187 16088
rect 0 16056 800 16086
rect 1485 16083 1551 16086
rect 9121 16083 9187 16086
rect 21265 16146 21331 16149
rect 22200 16146 23000 16176
rect 21265 16144 23000 16146
rect 21265 16088 21270 16144
rect 21326 16088 23000 16144
rect 21265 16086 23000 16088
rect 21265 16083 21331 16086
rect 22200 16056 23000 16086
rect 5533 16010 5599 16013
rect 936 16008 5599 16010
rect 936 15952 5538 16008
rect 5594 15952 5599 16008
rect 936 15950 5599 15952
rect 197 15874 263 15877
rect 936 15874 996 15950
rect 5533 15947 5599 15950
rect 11881 16010 11947 16013
rect 12249 16010 12315 16013
rect 19701 16010 19767 16013
rect 11881 16008 19767 16010
rect 11881 15952 11886 16008
rect 11942 15952 12254 16008
rect 12310 15952 19706 16008
rect 19762 15952 19767 16008
rect 11881 15950 19767 15952
rect 11881 15947 11947 15950
rect 12249 15947 12315 15950
rect 19701 15947 19767 15950
rect 5073 15876 5139 15877
rect 197 15872 996 15874
rect 197 15816 202 15872
rect 258 15816 996 15872
rect 197 15814 996 15816
rect 197 15811 263 15814
rect 5022 15812 5028 15876
rect 5092 15874 5139 15876
rect 10685 15876 10751 15877
rect 10685 15874 10732 15876
rect 5092 15872 5184 15874
rect 5134 15816 5184 15872
rect 5092 15814 5184 15816
rect 10640 15872 10732 15874
rect 10640 15816 10690 15872
rect 10640 15814 10732 15816
rect 5092 15812 5139 15814
rect 5073 15811 5139 15812
rect 10685 15812 10732 15814
rect 10796 15812 10802 15876
rect 10685 15811 10751 15812
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 4061 15738 4127 15741
rect 7281 15738 7347 15741
rect 4061 15736 7347 15738
rect 4061 15680 4066 15736
rect 4122 15680 7286 15736
rect 7342 15680 7347 15736
rect 4061 15678 7347 15680
rect 4061 15675 4127 15678
rect 7281 15675 7347 15678
rect 0 15602 800 15632
rect 1485 15602 1551 15605
rect 0 15600 1551 15602
rect 0 15544 1490 15600
rect 1546 15544 1551 15600
rect 0 15542 1551 15544
rect 0 15512 800 15542
rect 1485 15539 1551 15542
rect 2630 15540 2636 15604
rect 2700 15602 2706 15604
rect 9489 15602 9555 15605
rect 2700 15600 9555 15602
rect 2700 15544 9494 15600
rect 9550 15544 9555 15600
rect 2700 15542 9555 15544
rect 2700 15540 2706 15542
rect 9489 15539 9555 15542
rect 21265 15602 21331 15605
rect 22200 15602 23000 15632
rect 21265 15600 23000 15602
rect 21265 15544 21270 15600
rect 21326 15544 23000 15600
rect 21265 15542 23000 15544
rect 21265 15539 21331 15542
rect 22200 15512 23000 15542
rect 9305 15466 9371 15469
rect 2730 15464 9371 15466
rect 2730 15408 9310 15464
rect 9366 15408 9371 15464
rect 2730 15406 9371 15408
rect 933 15330 999 15333
rect 2730 15330 2790 15406
rect 9305 15403 9371 15406
rect 9673 15466 9739 15469
rect 11053 15466 11119 15469
rect 17953 15466 18019 15469
rect 9673 15464 18019 15466
rect 9673 15408 9678 15464
rect 9734 15408 11058 15464
rect 11114 15408 17958 15464
rect 18014 15408 18019 15464
rect 9673 15406 18019 15408
rect 9673 15403 9739 15406
rect 11053 15403 11119 15406
rect 17953 15403 18019 15406
rect 933 15328 2790 15330
rect 933 15272 938 15328
rect 994 15272 2790 15328
rect 933 15270 2790 15272
rect 933 15267 999 15270
rect 3366 15268 3372 15332
rect 3436 15330 3442 15332
rect 4153 15330 4219 15333
rect 3436 15328 4219 15330
rect 3436 15272 4158 15328
rect 4214 15272 4219 15328
rect 3436 15270 4219 15272
rect 3436 15268 3442 15270
rect 4153 15267 4219 15270
rect 9254 15268 9260 15332
rect 9324 15330 9330 15332
rect 9857 15330 9923 15333
rect 9324 15328 9923 15330
rect 9324 15272 9862 15328
rect 9918 15272 9923 15328
rect 9324 15270 9923 15272
rect 9324 15268 9330 15270
rect 9857 15267 9923 15270
rect 6142 15264 6462 15265
rect 0 15194 800 15224
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 15199 16858 15200
rect 1485 15194 1551 15197
rect 4061 15194 4127 15197
rect 0 15192 1551 15194
rect 0 15136 1490 15192
rect 1546 15136 1551 15192
rect 0 15134 1551 15136
rect 0 15104 800 15134
rect 1485 15131 1551 15134
rect 2730 15192 4127 15194
rect 2730 15136 4066 15192
rect 4122 15136 4127 15192
rect 2730 15134 4127 15136
rect 2078 14996 2084 15060
rect 2148 15058 2154 15060
rect 2730 15058 2790 15134
rect 4061 15131 4127 15134
rect 21265 15194 21331 15197
rect 22200 15194 23000 15224
rect 21265 15192 23000 15194
rect 21265 15136 21270 15192
rect 21326 15136 23000 15192
rect 21265 15134 23000 15136
rect 21265 15131 21331 15134
rect 22200 15104 23000 15134
rect 2148 14998 2790 15058
rect 2148 14996 2154 14998
rect 3543 14720 3863 14721
rect 0 14650 800 14680
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 800 14590
rect 1485 14587 1551 14590
rect 21265 14650 21331 14653
rect 22200 14650 23000 14680
rect 21265 14648 23000 14650
rect 21265 14592 21270 14648
rect 21326 14592 23000 14648
rect 21265 14590 23000 14592
rect 21265 14587 21331 14590
rect 22200 14560 23000 14590
rect 9949 14514 10015 14517
rect 17309 14514 17375 14517
rect 9949 14512 17375 14514
rect 9949 14456 9954 14512
rect 10010 14456 17314 14512
rect 17370 14456 17375 14512
rect 9949 14454 17375 14456
rect 9949 14451 10015 14454
rect 17309 14451 17375 14454
rect 2446 14316 2452 14380
rect 2516 14378 2522 14380
rect 10593 14378 10659 14381
rect 2516 14376 10659 14378
rect 2516 14320 10598 14376
rect 10654 14320 10659 14376
rect 2516 14318 10659 14320
rect 2516 14316 2522 14318
rect 10593 14315 10659 14318
rect 14917 14378 14983 14381
rect 18689 14378 18755 14381
rect 14917 14376 18755 14378
rect 14917 14320 14922 14376
rect 14978 14320 18694 14376
rect 18750 14320 18755 14376
rect 14917 14318 18755 14320
rect 14917 14315 14983 14318
rect 18689 14315 18755 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 4470 14180 4476 14244
rect 4540 14242 4546 14244
rect 4981 14242 5047 14245
rect 4540 14240 5047 14242
rect 4540 14184 4986 14240
rect 5042 14184 5047 14240
rect 4540 14182 5047 14184
rect 4540 14180 4546 14182
rect 4981 14179 5047 14182
rect 21265 14242 21331 14245
rect 22200 14242 23000 14272
rect 21265 14240 23000 14242
rect 21265 14184 21270 14240
rect 21326 14184 23000 14240
rect 21265 14182 23000 14184
rect 21265 14179 21331 14182
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 22200 14152 23000 14182
rect 16538 14111 16858 14112
rect 3182 13908 3188 13972
rect 3252 13970 3258 13972
rect 8201 13970 8267 13973
rect 3252 13968 8267 13970
rect 3252 13912 8206 13968
rect 8262 13912 8267 13968
rect 3252 13910 8267 13912
rect 3252 13908 3258 13910
rect 8201 13907 8267 13910
rect 15469 13970 15535 13973
rect 19006 13970 19012 13972
rect 15469 13968 19012 13970
rect 15469 13912 15474 13968
rect 15530 13912 19012 13968
rect 15469 13910 19012 13912
rect 15469 13907 15535 13910
rect 19006 13908 19012 13910
rect 19076 13908 19082 13972
rect 0 13834 800 13864
rect 1485 13834 1551 13837
rect 0 13832 1551 13834
rect 0 13776 1490 13832
rect 1546 13776 1551 13832
rect 0 13774 1551 13776
rect 0 13744 800 13774
rect 1485 13771 1551 13774
rect 4705 13834 4771 13837
rect 5942 13834 5948 13836
rect 4705 13832 5948 13834
rect 4705 13776 4710 13832
rect 4766 13776 5948 13832
rect 4705 13774 5948 13776
rect 4705 13771 4771 13774
rect 5942 13772 5948 13774
rect 6012 13772 6018 13836
rect 6453 13834 6519 13837
rect 12525 13836 12591 13837
rect 13077 13836 13143 13837
rect 7598 13834 7604 13836
rect 6453 13832 7604 13834
rect 6453 13776 6458 13832
rect 6514 13776 7604 13832
rect 6453 13774 7604 13776
rect 6453 13771 6519 13774
rect 7598 13772 7604 13774
rect 7668 13772 7674 13836
rect 12525 13832 12572 13836
rect 12636 13834 12642 13836
rect 12525 13776 12530 13832
rect 12525 13772 12572 13776
rect 12636 13774 12682 13834
rect 13077 13832 13124 13836
rect 13188 13834 13194 13836
rect 13353 13834 13419 13837
rect 18822 13834 18828 13836
rect 13077 13776 13082 13832
rect 12636 13772 12642 13774
rect 13077 13772 13124 13776
rect 13188 13774 13234 13834
rect 13353 13832 18828 13834
rect 13353 13776 13358 13832
rect 13414 13776 18828 13832
rect 13353 13774 18828 13776
rect 13188 13772 13194 13774
rect 12525 13771 12591 13772
rect 13077 13771 13143 13772
rect 13353 13771 13419 13774
rect 18822 13772 18828 13774
rect 18892 13772 18898 13836
rect 21265 13834 21331 13837
rect 22200 13834 23000 13864
rect 21265 13832 23000 13834
rect 21265 13776 21270 13832
rect 21326 13776 23000 13832
rect 21265 13774 23000 13776
rect 21265 13771 21331 13774
rect 22200 13744 23000 13774
rect 4838 13636 4844 13700
rect 4908 13698 4914 13700
rect 6729 13698 6795 13701
rect 7465 13700 7531 13701
rect 4908 13696 6795 13698
rect 4908 13640 6734 13696
rect 6790 13640 6795 13696
rect 4908 13638 6795 13640
rect 4908 13636 4914 13638
rect 6729 13635 6795 13638
rect 7414 13636 7420 13700
rect 7484 13698 7531 13700
rect 7484 13696 7576 13698
rect 7526 13640 7576 13696
rect 7484 13638 7576 13640
rect 7484 13636 7531 13638
rect 7465 13635 7531 13636
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 1393 13426 1459 13429
rect 12249 13426 12315 13429
rect 1393 13424 12315 13426
rect 1393 13368 1398 13424
rect 1454 13368 12254 13424
rect 12310 13368 12315 13424
rect 1393 13366 12315 13368
rect 1393 13363 1459 13366
rect 12249 13363 12315 13366
rect 15653 13426 15719 13429
rect 18638 13426 18644 13428
rect 15653 13424 18644 13426
rect 15653 13368 15658 13424
rect 15714 13368 18644 13424
rect 15653 13366 18644 13368
rect 15653 13363 15719 13366
rect 18638 13364 18644 13366
rect 18708 13364 18714 13428
rect 0 13290 800 13320
rect 1485 13290 1551 13293
rect 0 13288 1551 13290
rect 0 13232 1490 13288
rect 1546 13232 1551 13288
rect 0 13230 1551 13232
rect 0 13200 800 13230
rect 1485 13227 1551 13230
rect 2773 13290 2839 13293
rect 4521 13290 4587 13293
rect 2773 13288 4587 13290
rect 2773 13232 2778 13288
rect 2834 13232 4526 13288
rect 4582 13232 4587 13288
rect 2773 13230 4587 13232
rect 2773 13227 2839 13230
rect 4521 13227 4587 13230
rect 21265 13290 21331 13293
rect 22200 13290 23000 13320
rect 21265 13288 23000 13290
rect 21265 13232 21270 13288
rect 21326 13232 23000 13288
rect 21265 13230 23000 13232
rect 21265 13227 21331 13230
rect 22200 13200 23000 13230
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 4286 12956 4292 13020
rect 4356 13018 4362 13020
rect 4521 13018 4587 13021
rect 4356 13016 4587 13018
rect 4356 12960 4526 13016
rect 4582 12960 4587 13016
rect 4356 12958 4587 12960
rect 4356 12956 4362 12958
rect 4521 12955 4587 12958
rect 12341 13018 12407 13021
rect 15469 13018 15535 13021
rect 12341 13016 15535 13018
rect 12341 12960 12346 13016
rect 12402 12960 15474 13016
rect 15530 12960 15535 13016
rect 12341 12958 15535 12960
rect 12341 12955 12407 12958
rect 15469 12955 15535 12958
rect 0 12882 800 12912
rect 1945 12882 2011 12885
rect 0 12880 2011 12882
rect 0 12824 1950 12880
rect 2006 12824 2011 12880
rect 0 12822 2011 12824
rect 0 12792 800 12822
rect 1945 12819 2011 12822
rect 4102 12820 4108 12884
rect 4172 12882 4178 12884
rect 4429 12882 4495 12885
rect 4172 12880 4495 12882
rect 4172 12824 4434 12880
rect 4490 12824 4495 12880
rect 4172 12822 4495 12824
rect 4172 12820 4178 12822
rect 4429 12819 4495 12822
rect 11094 12820 11100 12884
rect 11164 12882 11170 12884
rect 11697 12882 11763 12885
rect 11164 12880 11763 12882
rect 11164 12824 11702 12880
rect 11758 12824 11763 12880
rect 11164 12822 11763 12824
rect 11164 12820 11170 12822
rect 11697 12819 11763 12822
rect 12709 12884 12775 12885
rect 12709 12880 12756 12884
rect 12820 12882 12826 12884
rect 18689 12882 18755 12885
rect 22200 12882 23000 12912
rect 12709 12824 12714 12880
rect 12709 12820 12756 12824
rect 12820 12822 12866 12882
rect 18689 12880 23000 12882
rect 18689 12824 18694 12880
rect 18750 12824 23000 12880
rect 18689 12822 23000 12824
rect 12820 12820 12826 12822
rect 12709 12819 12775 12820
rect 18689 12819 18755 12822
rect 22200 12792 23000 12822
rect 3509 12746 3575 12749
rect 3190 12744 3575 12746
rect 3190 12688 3514 12744
rect 3570 12688 3575 12744
rect 3190 12686 3575 12688
rect 3190 12613 3250 12686
rect 3509 12683 3575 12686
rect 13353 12746 13419 12749
rect 21081 12746 21147 12749
rect 13353 12744 21147 12746
rect 13353 12688 13358 12744
rect 13414 12688 21086 12744
rect 21142 12688 21147 12744
rect 13353 12686 21147 12688
rect 13353 12683 13419 12686
rect 21081 12683 21147 12686
rect 3141 12608 3250 12613
rect 3141 12552 3146 12608
rect 3202 12552 3250 12608
rect 3141 12550 3250 12552
rect 3141 12547 3207 12550
rect 12014 12548 12020 12612
rect 12084 12610 12090 12612
rect 13261 12610 13327 12613
rect 12084 12608 13327 12610
rect 12084 12552 13266 12608
rect 13322 12552 13327 12608
rect 12084 12550 13327 12552
rect 12084 12548 12090 12550
rect 13261 12547 13327 12550
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 12479 19457 12480
rect 5441 12474 5507 12477
rect 9121 12474 9187 12477
rect 9489 12474 9555 12477
rect 5441 12472 6010 12474
rect 5441 12416 5446 12472
rect 5502 12416 6010 12472
rect 5441 12414 6010 12416
rect 5441 12411 5507 12414
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 4429 12338 4495 12341
rect 4797 12338 4863 12341
rect 5717 12340 5783 12341
rect 5717 12338 5764 12340
rect 4429 12336 4863 12338
rect 4429 12280 4434 12336
rect 4490 12280 4802 12336
rect 4858 12280 4863 12336
rect 4429 12278 4863 12280
rect 5672 12336 5764 12338
rect 5672 12280 5722 12336
rect 5672 12278 5764 12280
rect 4429 12275 4495 12278
rect 4797 12275 4863 12278
rect 5717 12276 5764 12278
rect 5828 12276 5834 12340
rect 5950 12338 6010 12414
rect 9121 12472 9555 12474
rect 9121 12416 9126 12472
rect 9182 12416 9494 12472
rect 9550 12416 9555 12472
rect 9121 12414 9555 12416
rect 9121 12411 9187 12414
rect 9489 12411 9555 12414
rect 14457 12474 14523 12477
rect 17953 12474 18019 12477
rect 14457 12472 18019 12474
rect 14457 12416 14462 12472
rect 14518 12416 17958 12472
rect 18014 12416 18019 12472
rect 14457 12414 18019 12416
rect 14457 12411 14523 12414
rect 17953 12411 18019 12414
rect 9121 12338 9187 12341
rect 5950 12336 9187 12338
rect 5950 12280 9126 12336
rect 9182 12280 9187 12336
rect 5950 12278 9187 12280
rect 5717 12275 5783 12276
rect 9121 12275 9187 12278
rect 11053 12338 11119 12341
rect 20713 12338 20779 12341
rect 11053 12336 20779 12338
rect 11053 12280 11058 12336
rect 11114 12280 20718 12336
rect 20774 12280 20779 12336
rect 11053 12278 20779 12280
rect 11053 12275 11119 12278
rect 20713 12275 20779 12278
rect 21357 12338 21423 12341
rect 22200 12338 23000 12368
rect 21357 12336 23000 12338
rect 21357 12280 21362 12336
rect 21418 12280 23000 12336
rect 21357 12278 23000 12280
rect 21357 12275 21423 12278
rect 22200 12248 23000 12278
rect 1761 12202 1827 12205
rect 13721 12202 13787 12205
rect 17033 12202 17099 12205
rect 1761 12200 17099 12202
rect 1761 12144 1766 12200
rect 1822 12144 13726 12200
rect 13782 12144 17038 12200
rect 17094 12144 17099 12200
rect 1761 12142 17099 12144
rect 1761 12139 1827 12142
rect 13721 12139 13787 12142
rect 17033 12139 17099 12142
rect 8937 12066 9003 12069
rect 9581 12066 9647 12069
rect 8937 12064 9647 12066
rect 8937 12008 8942 12064
rect 8998 12008 9586 12064
rect 9642 12008 9647 12064
rect 8937 12006 9647 12008
rect 8937 12003 9003 12006
rect 9581 12003 9647 12006
rect 6142 12000 6462 12001
rect 0 11930 800 11960
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 11935 16858 11936
rect 1577 11930 1643 11933
rect 0 11928 1643 11930
rect 0 11872 1582 11928
rect 1638 11872 1643 11928
rect 0 11870 1643 11872
rect 0 11840 800 11870
rect 1577 11867 1643 11870
rect 2681 11930 2747 11933
rect 5441 11930 5507 11933
rect 2681 11928 5507 11930
rect 2681 11872 2686 11928
rect 2742 11872 5446 11928
rect 5502 11872 5507 11928
rect 2681 11870 5507 11872
rect 2681 11867 2747 11870
rect 5441 11867 5507 11870
rect 8201 11930 8267 11933
rect 9581 11930 9647 11933
rect 8201 11928 9647 11930
rect 8201 11872 8206 11928
rect 8262 11872 9586 11928
rect 9642 11872 9647 11928
rect 8201 11870 9647 11872
rect 8201 11867 8267 11870
rect 9581 11867 9647 11870
rect 20253 11930 20319 11933
rect 22200 11930 23000 11960
rect 20253 11928 23000 11930
rect 20253 11872 20258 11928
rect 20314 11872 23000 11928
rect 20253 11870 23000 11872
rect 20253 11867 20319 11870
rect 22200 11840 23000 11870
rect 8845 11658 8911 11661
rect 9397 11658 9463 11661
rect 8845 11656 9463 11658
rect 8845 11600 8850 11656
rect 8906 11600 9402 11656
rect 9458 11600 9463 11656
rect 8845 11598 9463 11600
rect 8845 11595 8911 11598
rect 9397 11595 9463 11598
rect 13629 11658 13695 11661
rect 18873 11658 18939 11661
rect 13629 11656 18939 11658
rect 13629 11600 13634 11656
rect 13690 11600 18878 11656
rect 18934 11600 18939 11656
rect 13629 11598 18939 11600
rect 13629 11595 13695 11598
rect 18873 11595 18939 11598
rect 3543 11456 3863 11457
rect 0 11386 800 11416
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 1577 11386 1643 11389
rect 0 11384 1643 11386
rect 0 11328 1582 11384
rect 1638 11328 1643 11384
rect 0 11326 1643 11328
rect 0 11296 800 11326
rect 1577 11323 1643 11326
rect 20713 11386 20779 11389
rect 22200 11386 23000 11416
rect 20713 11384 23000 11386
rect 20713 11328 20718 11384
rect 20774 11328 23000 11384
rect 20713 11326 23000 11328
rect 20713 11323 20779 11326
rect 22200 11296 23000 11326
rect 11237 11250 11303 11253
rect 14365 11250 14431 11253
rect 11237 11248 14431 11250
rect 11237 11192 11242 11248
rect 11298 11192 14370 11248
rect 14426 11192 14431 11248
rect 11237 11190 14431 11192
rect 11237 11187 11303 11190
rect 14365 11187 14431 11190
rect 6862 11052 6868 11116
rect 6932 11114 6938 11116
rect 7373 11114 7439 11117
rect 6932 11112 7439 11114
rect 6932 11056 7378 11112
rect 7434 11056 7439 11112
rect 6932 11054 7439 11056
rect 6932 11052 6938 11054
rect 7373 11051 7439 11054
rect 13629 11114 13695 11117
rect 19926 11114 19932 11116
rect 13629 11112 19932 11114
rect 13629 11056 13634 11112
rect 13690 11056 19932 11112
rect 13629 11054 19932 11056
rect 13629 11051 13695 11054
rect 19926 11052 19932 11054
rect 19996 11052 20002 11116
rect 0 10978 800 11008
rect 3325 10978 3391 10981
rect 0 10976 3391 10978
rect 0 10920 3330 10976
rect 3386 10920 3391 10976
rect 0 10918 3391 10920
rect 0 10888 800 10918
rect 3325 10915 3391 10918
rect 18597 10978 18663 10981
rect 22200 10978 23000 11008
rect 18597 10976 23000 10978
rect 18597 10920 18602 10976
rect 18658 10920 23000 10976
rect 18597 10918 23000 10920
rect 18597 10915 18663 10918
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 22200 10888 23000 10918
rect 16538 10847 16858 10848
rect 3601 10706 3667 10709
rect 7097 10706 7163 10709
rect 3601 10704 7163 10706
rect 3601 10648 3606 10704
rect 3662 10648 7102 10704
rect 7158 10648 7163 10704
rect 3601 10646 7163 10648
rect 3601 10643 3667 10646
rect 7097 10643 7163 10646
rect 13537 10706 13603 10709
rect 17902 10706 17908 10708
rect 13537 10704 17908 10706
rect 13537 10648 13542 10704
rect 13598 10648 17908 10704
rect 13537 10646 17908 10648
rect 13537 10643 13603 10646
rect 17902 10644 17908 10646
rect 17972 10644 17978 10708
rect 5625 10570 5691 10573
rect 8017 10570 8083 10573
rect 5625 10568 8083 10570
rect 5625 10512 5630 10568
rect 5686 10512 8022 10568
rect 8078 10512 8083 10568
rect 5625 10510 8083 10512
rect 5625 10507 5691 10510
rect 8017 10507 8083 10510
rect 12801 10570 12867 10573
rect 18965 10570 19031 10573
rect 12801 10568 19626 10570
rect 12801 10512 12806 10568
rect 12862 10512 18970 10568
rect 19026 10512 19626 10568
rect 12801 10510 19626 10512
rect 12801 10507 12867 10510
rect 18965 10507 19031 10510
rect 0 10434 800 10464
rect 1669 10434 1735 10437
rect 0 10432 1735 10434
rect 0 10376 1674 10432
rect 1730 10376 1735 10432
rect 0 10374 1735 10376
rect 19566 10434 19626 10510
rect 22200 10434 23000 10464
rect 19566 10374 23000 10434
rect 0 10344 800 10374
rect 1669 10371 1735 10374
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 22200 10344 23000 10374
rect 19137 10303 19457 10304
rect 10317 10298 10383 10301
rect 11421 10298 11487 10301
rect 10317 10296 11487 10298
rect 10317 10240 10322 10296
rect 10378 10240 11426 10296
rect 11482 10240 11487 10296
rect 10317 10238 11487 10240
rect 10317 10235 10383 10238
rect 11421 10235 11487 10238
rect 1853 10162 1919 10165
rect 11237 10162 11303 10165
rect 1853 10160 11303 10162
rect 1853 10104 1858 10160
rect 1914 10104 11242 10160
rect 11298 10104 11303 10160
rect 1853 10102 11303 10104
rect 1853 10099 1919 10102
rect 11237 10099 11303 10102
rect 17493 10162 17559 10165
rect 20989 10162 21055 10165
rect 17493 10160 21055 10162
rect 17493 10104 17498 10160
rect 17554 10104 20994 10160
rect 21050 10104 21055 10160
rect 17493 10102 21055 10104
rect 17493 10099 17559 10102
rect 20989 10099 21055 10102
rect 0 10026 800 10056
rect 1669 10026 1735 10029
rect 0 10024 1735 10026
rect 0 9968 1674 10024
rect 1730 9968 1735 10024
rect 0 9966 1735 9968
rect 0 9936 800 9966
rect 1669 9963 1735 9966
rect 5022 9964 5028 10028
rect 5092 10026 5098 10028
rect 18137 10026 18203 10029
rect 5092 10024 18203 10026
rect 5092 9968 18142 10024
rect 18198 9968 18203 10024
rect 5092 9966 18203 9968
rect 5092 9964 5098 9966
rect 18137 9963 18203 9966
rect 18689 10026 18755 10029
rect 22200 10026 23000 10056
rect 18689 10024 23000 10026
rect 18689 9968 18694 10024
rect 18750 9968 23000 10024
rect 18689 9966 23000 9968
rect 18689 9963 18755 9966
rect 22200 9936 23000 9966
rect 4981 9890 5047 9893
rect 5993 9890 6059 9893
rect 4981 9888 6059 9890
rect 4981 9832 4986 9888
rect 5042 9832 5998 9888
rect 6054 9832 6059 9888
rect 4981 9830 6059 9832
rect 4981 9827 5047 9830
rect 5993 9827 6059 9830
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 2497 9618 2563 9621
rect 10593 9618 10659 9621
rect 2497 9616 10659 9618
rect 2497 9560 2502 9616
rect 2558 9560 10598 9616
rect 10654 9560 10659 9616
rect 2497 9558 10659 9560
rect 2497 9555 2563 9558
rect 10593 9555 10659 9558
rect 13169 9618 13235 9621
rect 17585 9618 17651 9621
rect 13169 9616 17651 9618
rect 13169 9560 13174 9616
rect 13230 9560 17590 9616
rect 17646 9560 17651 9616
rect 13169 9558 17651 9560
rect 13169 9555 13235 9558
rect 17585 9555 17651 9558
rect 0 9482 800 9512
rect 1577 9482 1643 9485
rect 3509 9482 3575 9485
rect 0 9480 1643 9482
rect 0 9424 1582 9480
rect 1638 9424 1643 9480
rect 0 9422 1643 9424
rect 0 9392 800 9422
rect 1577 9419 1643 9422
rect 2730 9480 3575 9482
rect 2730 9424 3514 9480
rect 3570 9424 3575 9480
rect 2730 9422 3575 9424
rect 0 9074 800 9104
rect 2730 9074 2790 9422
rect 3509 9419 3575 9422
rect 7373 9482 7439 9485
rect 8477 9482 8543 9485
rect 7373 9480 8543 9482
rect 7373 9424 7378 9480
rect 7434 9424 8482 9480
rect 8538 9424 8543 9480
rect 7373 9422 8543 9424
rect 7373 9419 7439 9422
rect 8477 9419 8543 9422
rect 9765 9482 9831 9485
rect 17769 9482 17835 9485
rect 9765 9480 17835 9482
rect 9765 9424 9770 9480
rect 9826 9424 17774 9480
rect 17830 9424 17835 9480
rect 9765 9422 17835 9424
rect 9765 9419 9831 9422
rect 17769 9419 17835 9422
rect 18597 9482 18663 9485
rect 22200 9482 23000 9512
rect 18597 9480 23000 9482
rect 18597 9424 18602 9480
rect 18658 9424 23000 9480
rect 18597 9422 23000 9424
rect 18597 9419 18663 9422
rect 22200 9392 23000 9422
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 9215 19457 9216
rect 0 9014 2790 9074
rect 11145 9074 11211 9077
rect 17769 9074 17835 9077
rect 11145 9072 17835 9074
rect 11145 9016 11150 9072
rect 11206 9016 17774 9072
rect 17830 9016 17835 9072
rect 11145 9014 17835 9016
rect 0 8984 800 9014
rect 11145 9011 11211 9014
rect 17769 9011 17835 9014
rect 17953 9074 18019 9077
rect 22200 9074 23000 9104
rect 17953 9072 23000 9074
rect 17953 9016 17958 9072
rect 18014 9016 23000 9072
rect 17953 9014 23000 9016
rect 17953 9011 18019 9014
rect 22200 8984 23000 9014
rect 2221 8938 2287 8941
rect 3417 8938 3483 8941
rect 2221 8936 3483 8938
rect 2221 8880 2226 8936
rect 2282 8880 3422 8936
rect 3478 8880 3483 8936
rect 2221 8878 3483 8880
rect 2221 8875 2287 8878
rect 3417 8875 3483 8878
rect 4245 8938 4311 8941
rect 4981 8938 5047 8941
rect 4245 8936 5047 8938
rect 4245 8880 4250 8936
rect 4306 8880 4986 8936
rect 5042 8880 5047 8936
rect 4245 8878 5047 8880
rect 4245 8875 4311 8878
rect 4981 8875 5047 8878
rect 13537 8938 13603 8941
rect 15009 8938 15075 8941
rect 19793 8938 19859 8941
rect 13537 8936 19859 8938
rect 13537 8880 13542 8936
rect 13598 8880 15014 8936
rect 15070 8880 19798 8936
rect 19854 8880 19859 8936
rect 13537 8878 19859 8880
rect 13537 8875 13603 8878
rect 15009 8875 15075 8878
rect 19793 8875 19859 8878
rect 9489 8802 9555 8805
rect 9622 8802 9628 8804
rect 9489 8800 9628 8802
rect 9489 8744 9494 8800
rect 9550 8744 9628 8800
rect 9489 8742 9628 8744
rect 9489 8739 9555 8742
rect 9622 8740 9628 8742
rect 9692 8740 9698 8804
rect 6142 8736 6462 8737
rect 0 8666 800 8696
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 1669 8666 1735 8669
rect 13537 8666 13603 8669
rect 17125 8668 17191 8669
rect 17125 8666 17172 8668
rect 0 8664 1735 8666
rect 0 8608 1674 8664
rect 1730 8608 1735 8664
rect 0 8606 1735 8608
rect 0 8576 800 8606
rect 1669 8603 1735 8606
rect 12390 8664 13603 8666
rect 12390 8608 13542 8664
rect 13598 8608 13603 8664
rect 12390 8606 13603 8608
rect 17080 8664 17172 8666
rect 17080 8608 17130 8664
rect 17080 8606 17172 8608
rect 3325 8530 3391 8533
rect 3918 8530 3924 8532
rect 3325 8528 3924 8530
rect 3325 8472 3330 8528
rect 3386 8472 3924 8528
rect 3325 8470 3924 8472
rect 3325 8467 3391 8470
rect 3918 8468 3924 8470
rect 3988 8468 3994 8532
rect 6862 8468 6868 8532
rect 6932 8530 6938 8532
rect 12390 8530 12450 8606
rect 13537 8603 13603 8606
rect 17125 8604 17172 8606
rect 17236 8604 17242 8668
rect 18781 8666 18847 8669
rect 22200 8666 23000 8696
rect 18781 8664 23000 8666
rect 18781 8608 18786 8664
rect 18842 8608 23000 8664
rect 18781 8606 23000 8608
rect 17125 8603 17191 8604
rect 18781 8603 18847 8606
rect 22200 8576 23000 8606
rect 6932 8470 12450 8530
rect 12709 8530 12775 8533
rect 17953 8530 18019 8533
rect 12709 8528 18019 8530
rect 12709 8472 12714 8528
rect 12770 8472 17958 8528
rect 18014 8472 18019 8528
rect 12709 8470 18019 8472
rect 6932 8468 6938 8470
rect 12709 8467 12775 8470
rect 17953 8467 18019 8470
rect 1853 8394 1919 8397
rect 9673 8394 9739 8397
rect 13261 8394 13327 8397
rect 15101 8394 15167 8397
rect 1853 8392 6930 8394
rect 1853 8336 1858 8392
rect 1914 8336 6930 8392
rect 1853 8334 6930 8336
rect 1853 8331 1919 8334
rect 6361 8258 6427 8261
rect 6678 8258 6684 8260
rect 6361 8256 6684 8258
rect 6361 8200 6366 8256
rect 6422 8200 6684 8256
rect 6361 8198 6684 8200
rect 6361 8195 6427 8198
rect 6678 8196 6684 8198
rect 6748 8196 6754 8260
rect 6870 8258 6930 8334
rect 8526 8334 9322 8394
rect 8526 8258 8586 8334
rect 6870 8198 8586 8258
rect 9262 8258 9322 8334
rect 9673 8392 15167 8394
rect 9673 8336 9678 8392
rect 9734 8336 13266 8392
rect 13322 8336 15106 8392
rect 15162 8336 15167 8392
rect 9673 8334 15167 8336
rect 9673 8331 9739 8334
rect 13261 8331 13327 8334
rect 15101 8331 15167 8334
rect 18822 8332 18828 8396
rect 18892 8394 18898 8396
rect 21081 8394 21147 8397
rect 18892 8392 21147 8394
rect 18892 8336 21086 8392
rect 21142 8336 21147 8392
rect 18892 8334 21147 8336
rect 18892 8332 18898 8334
rect 21081 8331 21147 8334
rect 11830 8258 11836 8260
rect 9262 8198 11836 8258
rect 11830 8196 11836 8198
rect 11900 8196 11906 8260
rect 3543 8192 3863 8193
rect 0 8122 800 8152
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 1485 8122 1551 8125
rect 9581 8124 9647 8125
rect 9581 8122 9628 8124
rect 0 8120 2790 8122
rect 0 8064 1490 8120
rect 1546 8064 2790 8120
rect 0 8062 2790 8064
rect 9536 8120 9628 8122
rect 9536 8064 9586 8120
rect 9536 8062 9628 8064
rect 0 8032 800 8062
rect 1485 8059 1551 8062
rect 2730 7986 2790 8062
rect 9581 8060 9628 8062
rect 9692 8060 9698 8124
rect 22200 8122 23000 8152
rect 19750 8062 23000 8122
rect 9581 8059 9647 8060
rect 4470 7986 4476 7988
rect 2730 7926 4476 7986
rect 4470 7924 4476 7926
rect 4540 7924 4546 7988
rect 8334 7924 8340 7988
rect 8404 7986 8410 7988
rect 11973 7986 12039 7989
rect 8404 7984 12039 7986
rect 8404 7928 11978 7984
rect 12034 7928 12039 7984
rect 8404 7926 12039 7928
rect 8404 7924 8410 7926
rect 11973 7923 12039 7926
rect 12893 7986 12959 7989
rect 18321 7986 18387 7989
rect 19750 7986 19810 8062
rect 22200 8032 23000 8062
rect 12893 7984 16314 7986
rect 12893 7928 12898 7984
rect 12954 7928 16314 7984
rect 12893 7926 16314 7928
rect 12893 7923 12959 7926
rect 4705 7850 4771 7853
rect 16113 7850 16179 7853
rect 4705 7848 16179 7850
rect 4705 7792 4710 7848
rect 4766 7792 16118 7848
rect 16174 7792 16179 7848
rect 4705 7790 16179 7792
rect 16254 7850 16314 7926
rect 18321 7984 19810 7986
rect 18321 7928 18326 7984
rect 18382 7928 19810 7984
rect 18321 7926 19810 7928
rect 18321 7923 18387 7926
rect 18689 7850 18755 7853
rect 16254 7848 18755 7850
rect 16254 7792 18694 7848
rect 18750 7792 18755 7848
rect 16254 7790 18755 7792
rect 4705 7787 4771 7790
rect 16113 7787 16179 7790
rect 18689 7787 18755 7790
rect 0 7714 800 7744
rect 2221 7714 2287 7717
rect 0 7712 2287 7714
rect 0 7656 2226 7712
rect 2282 7656 2287 7712
rect 0 7654 2287 7656
rect 0 7624 800 7654
rect 2221 7651 2287 7654
rect 18229 7714 18295 7717
rect 22200 7714 23000 7744
rect 18229 7712 23000 7714
rect 18229 7656 18234 7712
rect 18290 7656 23000 7712
rect 18229 7654 23000 7656
rect 18229 7651 18295 7654
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 22200 7624 23000 7654
rect 16538 7583 16858 7584
rect 1853 7578 1919 7581
rect 2078 7578 2084 7580
rect 1853 7576 2084 7578
rect 1853 7520 1858 7576
rect 1914 7520 2084 7576
rect 1853 7518 2084 7520
rect 1853 7515 1919 7518
rect 2078 7516 2084 7518
rect 2148 7516 2154 7580
rect 1945 7442 2011 7445
rect 9397 7442 9463 7445
rect 1945 7440 9463 7442
rect 1945 7384 1950 7440
rect 2006 7384 9402 7440
rect 9458 7384 9463 7440
rect 1945 7382 9463 7384
rect 1945 7379 2011 7382
rect 9397 7379 9463 7382
rect 2773 7306 2839 7309
rect 7005 7306 7071 7309
rect 2773 7304 7071 7306
rect 2773 7248 2778 7304
rect 2834 7248 7010 7304
rect 7066 7248 7071 7304
rect 2773 7246 7071 7248
rect 2773 7243 2839 7246
rect 7005 7243 7071 7246
rect 7966 7244 7972 7308
rect 8036 7306 8042 7308
rect 11094 7306 11100 7308
rect 8036 7246 11100 7306
rect 8036 7244 8042 7246
rect 11094 7244 11100 7246
rect 11164 7244 11170 7308
rect 13353 7306 13419 7309
rect 17309 7306 17375 7309
rect 13353 7304 17375 7306
rect 13353 7248 13358 7304
rect 13414 7248 17314 7304
rect 17370 7248 17375 7304
rect 13353 7246 17375 7248
rect 13353 7243 13419 7246
rect 17309 7243 17375 7246
rect 17953 7306 18019 7309
rect 17953 7304 19626 7306
rect 17953 7248 17958 7304
rect 18014 7248 19626 7304
rect 17953 7246 19626 7248
rect 17953 7243 18019 7246
rect 0 7170 800 7200
rect 3417 7170 3483 7173
rect 17033 7172 17099 7173
rect 16982 7170 16988 7172
rect 0 7168 3483 7170
rect 0 7112 3422 7168
rect 3478 7112 3483 7168
rect 0 7110 3483 7112
rect 16942 7110 16988 7170
rect 17052 7168 17099 7172
rect 17094 7112 17099 7168
rect 0 7080 800 7110
rect 3417 7107 3483 7110
rect 16982 7108 16988 7110
rect 17052 7108 17099 7112
rect 19566 7170 19626 7246
rect 22200 7170 23000 7200
rect 19566 7110 23000 7170
rect 17033 7107 17099 7108
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 22200 7080 23000 7110
rect 19137 7039 19457 7040
rect 3233 7034 3299 7037
rect 3366 7034 3372 7036
rect 3233 7032 3372 7034
rect 3233 6976 3238 7032
rect 3294 6976 3372 7032
rect 3233 6974 3372 6976
rect 3233 6971 3299 6974
rect 3366 6972 3372 6974
rect 3436 6972 3442 7036
rect 14641 7034 14707 7037
rect 18045 7034 18111 7037
rect 14641 7032 18111 7034
rect 14641 6976 14646 7032
rect 14702 6976 18050 7032
rect 18106 6976 18111 7032
rect 14641 6974 18111 6976
rect 14641 6971 14707 6974
rect 18045 6971 18111 6974
rect 1577 6898 1643 6901
rect 2221 6898 2287 6901
rect 1577 6896 2287 6898
rect 1577 6840 1582 6896
rect 1638 6840 2226 6896
rect 2282 6840 2287 6896
rect 1577 6838 2287 6840
rect 1577 6835 1643 6838
rect 2221 6835 2287 6838
rect 10869 6898 10935 6901
rect 18045 6898 18111 6901
rect 10869 6896 18111 6898
rect 10869 6840 10874 6896
rect 10930 6840 18050 6896
rect 18106 6840 18111 6896
rect 10869 6838 18111 6840
rect 10869 6835 10935 6838
rect 18045 6835 18111 6838
rect 0 6762 800 6792
rect 933 6762 999 6765
rect 0 6760 999 6762
rect 0 6704 938 6760
rect 994 6704 999 6760
rect 0 6702 999 6704
rect 0 6672 800 6702
rect 933 6699 999 6702
rect 17125 6762 17191 6765
rect 18597 6762 18663 6765
rect 17125 6760 18663 6762
rect 17125 6704 17130 6760
rect 17186 6704 18602 6760
rect 18658 6704 18663 6760
rect 17125 6702 18663 6704
rect 17125 6699 17191 6702
rect 18597 6699 18663 6702
rect 18965 6762 19031 6765
rect 22200 6762 23000 6792
rect 18965 6760 23000 6762
rect 18965 6704 18970 6760
rect 19026 6704 23000 6760
rect 18965 6702 23000 6704
rect 18965 6699 19031 6702
rect 22200 6672 23000 6702
rect 2957 6626 3023 6629
rect 4337 6626 4403 6629
rect 4838 6626 4844 6628
rect 2957 6624 4844 6626
rect 2957 6568 2962 6624
rect 3018 6568 4342 6624
rect 4398 6568 4844 6624
rect 2957 6566 4844 6568
rect 2957 6563 3023 6566
rect 4337 6563 4403 6566
rect 4838 6564 4844 6566
rect 4908 6564 4914 6628
rect 17309 6626 17375 6629
rect 17769 6626 17835 6629
rect 17309 6624 17835 6626
rect 17309 6568 17314 6624
rect 17370 6568 17774 6624
rect 17830 6568 17835 6624
rect 17309 6566 17835 6568
rect 17309 6563 17375 6566
rect 17769 6563 17835 6566
rect 18781 6626 18847 6629
rect 18781 6624 21098 6626
rect 18781 6568 18786 6624
rect 18842 6568 21098 6624
rect 18781 6566 21098 6568
rect 18781 6563 18847 6566
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 6495 16858 6496
rect 1853 6490 1919 6493
rect 4797 6490 4863 6493
rect 5022 6490 5028 6492
rect 1853 6488 2790 6490
rect 1853 6432 1858 6488
rect 1914 6432 2790 6488
rect 1853 6430 2790 6432
rect 1853 6427 1919 6430
rect 2730 6354 2790 6430
rect 4797 6488 5028 6490
rect 4797 6432 4802 6488
rect 4858 6432 5028 6488
rect 4797 6430 5028 6432
rect 4797 6427 4863 6430
rect 5022 6428 5028 6430
rect 5092 6490 5098 6492
rect 5441 6490 5507 6493
rect 12157 6490 12223 6493
rect 5092 6488 5507 6490
rect 5092 6432 5446 6488
rect 5502 6432 5507 6488
rect 5092 6430 5507 6432
rect 5092 6428 5098 6430
rect 5441 6427 5507 6430
rect 11838 6488 12223 6490
rect 11838 6432 12162 6488
rect 12218 6432 12223 6488
rect 11838 6430 12223 6432
rect 6085 6354 6151 6357
rect 11838 6354 11898 6430
rect 12157 6427 12223 6430
rect 17217 6490 17283 6493
rect 17493 6490 17559 6493
rect 18965 6492 19031 6493
rect 18965 6490 19012 6492
rect 17217 6488 17559 6490
rect 17217 6432 17222 6488
rect 17278 6432 17498 6488
rect 17554 6432 17559 6488
rect 17217 6430 17559 6432
rect 18920 6488 19012 6490
rect 18920 6432 18970 6488
rect 18920 6430 19012 6432
rect 17217 6427 17283 6430
rect 17493 6427 17559 6430
rect 18965 6428 19012 6430
rect 19076 6428 19082 6492
rect 18965 6427 19031 6428
rect 19425 6354 19491 6357
rect 2730 6352 11898 6354
rect 2730 6296 6090 6352
rect 6146 6296 11898 6352
rect 2730 6294 11898 6296
rect 12022 6352 19491 6354
rect 12022 6296 19430 6352
rect 19486 6296 19491 6352
rect 12022 6294 19491 6296
rect 6085 6291 6151 6294
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 3785 6218 3851 6221
rect 5758 6218 5764 6220
rect 3785 6216 5764 6218
rect 3785 6160 3790 6216
rect 3846 6160 5764 6216
rect 3785 6158 5764 6160
rect 3785 6155 3851 6158
rect 5758 6156 5764 6158
rect 5828 6218 5834 6220
rect 6637 6218 6703 6221
rect 12022 6218 12082 6294
rect 19425 6291 19491 6294
rect 20897 6218 20963 6221
rect 5828 6216 12082 6218
rect 5828 6160 6642 6216
rect 6698 6160 12082 6216
rect 5828 6158 12082 6160
rect 12390 6216 20963 6218
rect 12390 6160 20902 6216
rect 20958 6160 20963 6216
rect 12390 6158 20963 6160
rect 21038 6218 21098 6566
rect 22200 6218 23000 6248
rect 21038 6158 23000 6218
rect 5828 6156 5834 6158
rect 6637 6155 6703 6158
rect 6177 6082 6243 6085
rect 6862 6082 6868 6084
rect 6177 6080 6868 6082
rect 6177 6024 6182 6080
rect 6238 6024 6868 6080
rect 6177 6022 6868 6024
rect 6177 6019 6243 6022
rect 6862 6020 6868 6022
rect 6932 6020 6938 6084
rect 11830 6020 11836 6084
rect 11900 6082 11906 6084
rect 11973 6082 12039 6085
rect 12390 6082 12450 6158
rect 20897 6155 20963 6158
rect 22200 6128 23000 6158
rect 11900 6080 12450 6082
rect 11900 6024 11978 6080
rect 12034 6024 12450 6080
rect 11900 6022 12450 6024
rect 11900 6020 11906 6022
rect 11973 6019 12039 6022
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 5951 19457 5952
rect 4429 5946 4495 5949
rect 6913 5946 6979 5949
rect 4429 5944 6979 5946
rect 4429 5888 4434 5944
rect 4490 5888 6918 5944
rect 6974 5888 6979 5944
rect 4429 5886 6979 5888
rect 4429 5883 4495 5886
rect 6913 5883 6979 5886
rect 14457 5946 14523 5949
rect 15285 5946 15351 5949
rect 14457 5944 15351 5946
rect 14457 5888 14462 5944
rect 14518 5888 15290 5944
rect 15346 5888 15351 5944
rect 14457 5886 15351 5888
rect 14457 5883 14523 5886
rect 15285 5883 15351 5886
rect 0 5810 800 5840
rect 1669 5810 1735 5813
rect 0 5808 1735 5810
rect 0 5752 1674 5808
rect 1730 5752 1735 5808
rect 0 5750 1735 5752
rect 0 5720 800 5750
rect 1669 5747 1735 5750
rect 5717 5810 5783 5813
rect 12525 5810 12591 5813
rect 5717 5808 12591 5810
rect 5717 5752 5722 5808
rect 5778 5752 12530 5808
rect 12586 5752 12591 5808
rect 5717 5750 12591 5752
rect 5717 5747 5783 5750
rect 12525 5747 12591 5750
rect 13629 5810 13695 5813
rect 17309 5810 17375 5813
rect 13629 5808 17375 5810
rect 13629 5752 13634 5808
rect 13690 5752 17314 5808
rect 17370 5752 17375 5808
rect 13629 5750 17375 5752
rect 13629 5747 13695 5750
rect 17309 5747 17375 5750
rect 18965 5810 19031 5813
rect 22200 5810 23000 5840
rect 18965 5808 23000 5810
rect 18965 5752 18970 5808
rect 19026 5752 23000 5808
rect 18965 5750 23000 5752
rect 18965 5747 19031 5750
rect 22200 5720 23000 5750
rect 5942 5612 5948 5676
rect 6012 5674 6018 5676
rect 7281 5674 7347 5677
rect 7465 5676 7531 5677
rect 6012 5672 7347 5674
rect 6012 5616 7286 5672
rect 7342 5616 7347 5672
rect 6012 5614 7347 5616
rect 6012 5612 6018 5614
rect 7281 5611 7347 5614
rect 7414 5612 7420 5676
rect 7484 5674 7531 5676
rect 10133 5674 10199 5677
rect 16665 5674 16731 5677
rect 7484 5672 7576 5674
rect 7526 5616 7576 5672
rect 7484 5614 7576 5616
rect 10133 5672 16731 5674
rect 10133 5616 10138 5672
rect 10194 5616 16670 5672
rect 16726 5616 16731 5672
rect 10133 5614 16731 5616
rect 7484 5612 7531 5614
rect 7465 5611 7531 5612
rect 10133 5611 10199 5614
rect 16665 5611 16731 5614
rect 3325 5538 3391 5541
rect 2730 5536 3391 5538
rect 2730 5480 3330 5536
rect 3386 5480 3391 5536
rect 2730 5478 3391 5480
rect 0 5266 800 5296
rect 2730 5266 2790 5478
rect 3325 5475 3391 5478
rect 17166 5476 17172 5540
rect 17236 5538 17242 5540
rect 17677 5538 17743 5541
rect 17236 5536 17743 5538
rect 17236 5480 17682 5536
rect 17738 5480 17743 5536
rect 17236 5478 17743 5480
rect 17236 5476 17242 5478
rect 17677 5475 17743 5478
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 0 5206 2790 5266
rect 3049 5266 3115 5269
rect 5717 5266 5783 5269
rect 3049 5264 5783 5266
rect 3049 5208 3054 5264
rect 3110 5208 5722 5264
rect 5778 5208 5783 5264
rect 3049 5206 5783 5208
rect 0 5176 800 5206
rect 3049 5203 3115 5206
rect 5717 5203 5783 5206
rect 6453 5266 6519 5269
rect 17033 5266 17099 5269
rect 6453 5264 17099 5266
rect 6453 5208 6458 5264
rect 6514 5208 17038 5264
rect 17094 5208 17099 5264
rect 6453 5206 17099 5208
rect 6453 5203 6519 5206
rect 17033 5203 17099 5206
rect 17861 5266 17927 5269
rect 22200 5266 23000 5296
rect 17861 5264 23000 5266
rect 17861 5208 17866 5264
rect 17922 5208 23000 5264
rect 17861 5206 23000 5208
rect 17861 5203 17927 5206
rect 22200 5176 23000 5206
rect 16941 5132 17007 5133
rect 16941 5130 16988 5132
rect 16896 5128 16988 5130
rect 16896 5072 16946 5128
rect 16896 5070 16988 5072
rect 16941 5068 16988 5070
rect 17052 5068 17058 5132
rect 16941 5067 17007 5068
rect 3543 4928 3863 4929
rect 0 4858 800 4888
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 933 4858 999 4861
rect 0 4856 999 4858
rect 0 4800 938 4856
rect 994 4800 999 4856
rect 0 4798 999 4800
rect 0 4768 800 4798
rect 933 4795 999 4798
rect 3969 4858 4035 4861
rect 4102 4858 4108 4860
rect 3969 4856 4108 4858
rect 3969 4800 3974 4856
rect 4030 4800 4108 4856
rect 3969 4798 4108 4800
rect 3969 4795 4035 4798
rect 4102 4796 4108 4798
rect 4172 4858 4178 4860
rect 15009 4858 15075 4861
rect 15285 4858 15351 4861
rect 4172 4798 7850 4858
rect 4172 4796 4178 4798
rect 2221 4724 2287 4725
rect 7557 4724 7623 4725
rect 2221 4722 2268 4724
rect 2176 4720 2268 4722
rect 2176 4664 2226 4720
rect 2176 4662 2268 4664
rect 2221 4660 2268 4662
rect 2332 4660 2338 4724
rect 7557 4722 7604 4724
rect 7512 4720 7604 4722
rect 7512 4664 7562 4720
rect 7512 4662 7604 4664
rect 7557 4660 7604 4662
rect 7668 4660 7674 4724
rect 7790 4722 7850 4798
rect 15009 4856 15351 4858
rect 15009 4800 15014 4856
rect 15070 4800 15290 4856
rect 15346 4800 15351 4856
rect 15009 4798 15351 4800
rect 15009 4795 15075 4798
rect 15285 4795 15351 4798
rect 20161 4858 20227 4861
rect 22200 4858 23000 4888
rect 20161 4856 23000 4858
rect 20161 4800 20166 4856
rect 20222 4800 23000 4856
rect 20161 4798 23000 4800
rect 20161 4795 20227 4798
rect 22200 4768 23000 4798
rect 18045 4722 18111 4725
rect 7790 4720 18111 4722
rect 7790 4664 18050 4720
rect 18106 4664 18111 4720
rect 7790 4662 18111 4664
rect 2221 4659 2287 4660
rect 7557 4659 7623 4660
rect 18045 4659 18111 4662
rect 1209 4586 1275 4589
rect 1853 4586 1919 4589
rect 7005 4586 7071 4589
rect 1209 4584 7071 4586
rect 1209 4528 1214 4584
rect 1270 4528 1858 4584
rect 1914 4528 7010 4584
rect 7066 4528 7071 4584
rect 1209 4526 7071 4528
rect 1209 4523 1275 4526
rect 1853 4523 1919 4526
rect 7005 4523 7071 4526
rect 15837 4586 15903 4589
rect 15837 4584 19350 4586
rect 15837 4528 15842 4584
rect 15898 4528 19350 4584
rect 15837 4526 19350 4528
rect 15837 4523 15903 4526
rect 0 4450 800 4480
rect 3141 4450 3207 4453
rect 0 4448 3207 4450
rect 0 4392 3146 4448
rect 3202 4392 3207 4448
rect 0 4390 3207 4392
rect 19290 4450 19350 4526
rect 22200 4450 23000 4480
rect 19290 4390 23000 4450
rect 0 4360 800 4390
rect 3141 4387 3207 4390
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 22200 4360 23000 4390
rect 16538 4319 16858 4320
rect 1485 4178 1551 4181
rect 8109 4178 8175 4181
rect 1485 4176 8175 4178
rect 1485 4120 1490 4176
rect 1546 4120 8114 4176
rect 8170 4120 8175 4176
rect 1485 4118 8175 4120
rect 1485 4115 1551 4118
rect 8109 4115 8175 4118
rect 4153 4042 4219 4045
rect 2730 4040 4219 4042
rect 2730 3984 4158 4040
rect 4214 3984 4219 4040
rect 2730 3982 4219 3984
rect 0 3906 800 3936
rect 2730 3906 2790 3982
rect 4153 3979 4219 3982
rect 7741 4042 7807 4045
rect 9213 4044 9279 4045
rect 8334 4042 8340 4044
rect 7741 4040 8340 4042
rect 7741 3984 7746 4040
rect 7802 3984 8340 4040
rect 7741 3982 8340 3984
rect 7741 3979 7807 3982
rect 8334 3980 8340 3982
rect 8404 3980 8410 4044
rect 9213 4042 9260 4044
rect 9168 4040 9260 4042
rect 9168 3984 9218 4040
rect 9168 3982 9260 3984
rect 9213 3980 9260 3982
rect 9324 3980 9330 4044
rect 13721 4042 13787 4045
rect 13721 4040 17786 4042
rect 13721 3984 13726 4040
rect 13782 3984 17786 4040
rect 13721 3982 17786 3984
rect 9213 3979 9279 3980
rect 13721 3979 13787 3982
rect 0 3846 2790 3906
rect 4337 3906 4403 3909
rect 8477 3906 8543 3909
rect 4337 3904 8543 3906
rect 4337 3848 4342 3904
rect 4398 3848 8482 3904
rect 8538 3848 8543 3904
rect 4337 3846 8543 3848
rect 17726 3906 17786 3982
rect 17902 3980 17908 4044
rect 17972 4042 17978 4044
rect 20713 4042 20779 4045
rect 17972 4040 20779 4042
rect 17972 3984 20718 4040
rect 20774 3984 20779 4040
rect 17972 3982 20779 3984
rect 17972 3980 17978 3982
rect 20713 3979 20779 3982
rect 18321 3906 18387 3909
rect 22200 3906 23000 3936
rect 17726 3904 18387 3906
rect 17726 3848 18326 3904
rect 18382 3848 18387 3904
rect 17726 3846 18387 3848
rect 0 3816 800 3846
rect 4337 3843 4403 3846
rect 8477 3843 8543 3846
rect 18321 3843 18387 3846
rect 20302 3846 23000 3906
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 10501 3770 10567 3773
rect 10501 3768 13692 3770
rect 10501 3712 10506 3768
rect 10562 3712 13692 3768
rect 10501 3710 13692 3712
rect 10501 3707 10567 3710
rect 13632 3637 13692 3710
rect 18638 3708 18644 3772
rect 18708 3770 18714 3772
rect 18965 3770 19031 3773
rect 18708 3768 19031 3770
rect 18708 3712 18970 3768
rect 19026 3712 19031 3768
rect 18708 3710 19031 3712
rect 18708 3708 18714 3710
rect 18965 3707 19031 3710
rect 2313 3634 2379 3637
rect 2446 3634 2452 3636
rect 2313 3632 2452 3634
rect 2313 3576 2318 3632
rect 2374 3576 2452 3632
rect 2313 3574 2452 3576
rect 2313 3571 2379 3574
rect 2446 3572 2452 3574
rect 2516 3572 2522 3636
rect 2865 3634 2931 3637
rect 4613 3634 4679 3637
rect 12566 3634 12572 3636
rect 2865 3632 12572 3634
rect 2865 3576 2870 3632
rect 2926 3576 4618 3632
rect 4674 3576 12572 3632
rect 2865 3574 12572 3576
rect 2865 3571 2931 3574
rect 4613 3571 4679 3574
rect 12566 3572 12572 3574
rect 12636 3572 12642 3636
rect 13629 3634 13695 3637
rect 20069 3634 20135 3637
rect 13629 3632 20135 3634
rect 13629 3576 13634 3632
rect 13690 3576 20074 3632
rect 20130 3576 20135 3632
rect 13629 3574 20135 3576
rect 13629 3571 13695 3574
rect 20069 3571 20135 3574
rect 0 3498 800 3528
rect 3785 3498 3851 3501
rect 0 3496 3851 3498
rect 0 3440 3790 3496
rect 3846 3440 3851 3496
rect 0 3438 3851 3440
rect 0 3408 800 3438
rect 3785 3435 3851 3438
rect 4981 3498 5047 3501
rect 12750 3498 12756 3500
rect 4981 3496 12756 3498
rect 4981 3440 4986 3496
rect 5042 3440 12756 3496
rect 4981 3438 12756 3440
rect 4981 3435 5047 3438
rect 12750 3436 12756 3438
rect 12820 3436 12826 3500
rect 18045 3498 18111 3501
rect 20302 3498 20362 3846
rect 22200 3816 23000 3846
rect 18045 3496 20362 3498
rect 18045 3440 18050 3496
rect 18106 3440 20362 3496
rect 18045 3438 20362 3440
rect 20621 3498 20687 3501
rect 22200 3498 23000 3528
rect 20621 3496 23000 3498
rect 20621 3440 20626 3496
rect 20682 3440 23000 3496
rect 20621 3438 23000 3440
rect 18045 3435 18111 3438
rect 20621 3435 20687 3438
rect 22200 3408 23000 3438
rect 3918 3300 3924 3364
rect 3988 3362 3994 3364
rect 5441 3362 5507 3365
rect 3988 3360 5507 3362
rect 3988 3304 5446 3360
rect 5502 3304 5507 3360
rect 3988 3302 5507 3304
rect 3988 3300 3994 3302
rect 5441 3299 5507 3302
rect 7833 3362 7899 3365
rect 7966 3362 7972 3364
rect 7833 3360 7972 3362
rect 7833 3304 7838 3360
rect 7894 3304 7972 3360
rect 7833 3302 7972 3304
rect 7833 3299 7899 3302
rect 7966 3300 7972 3302
rect 8036 3300 8042 3364
rect 19926 3300 19932 3364
rect 19996 3362 20002 3364
rect 20069 3362 20135 3365
rect 19996 3360 20135 3362
rect 19996 3304 20074 3360
rect 20130 3304 20135 3360
rect 19996 3302 20135 3304
rect 19996 3300 20002 3302
rect 20069 3299 20135 3302
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 3231 16858 3232
rect 197 3226 263 3229
rect 4981 3226 5047 3229
rect 197 3224 5047 3226
rect 197 3168 202 3224
rect 258 3168 4986 3224
rect 5042 3168 5047 3224
rect 197 3166 5047 3168
rect 197 3163 263 3166
rect 4981 3163 5047 3166
rect 6913 3090 6979 3093
rect 14825 3090 14891 3093
rect 6913 3088 14891 3090
rect 6913 3032 6918 3088
rect 6974 3032 14830 3088
rect 14886 3032 14891 3088
rect 6913 3030 14891 3032
rect 6913 3027 6979 3030
rect 14825 3027 14891 3030
rect 0 2954 800 2984
rect 2773 2954 2839 2957
rect 3182 2954 3188 2956
rect 0 2952 3188 2954
rect 0 2896 2778 2952
rect 2834 2896 3188 2952
rect 0 2894 3188 2896
rect 0 2864 800 2894
rect 2773 2891 2839 2894
rect 3182 2892 3188 2894
rect 3252 2892 3258 2956
rect 6678 2892 6684 2956
rect 6748 2954 6754 2956
rect 6913 2954 6979 2957
rect 6748 2952 6979 2954
rect 6748 2896 6918 2952
rect 6974 2896 6979 2952
rect 6748 2894 6979 2896
rect 6748 2892 6754 2894
rect 6913 2891 6979 2894
rect 8477 2954 8543 2957
rect 17217 2954 17283 2957
rect 8477 2952 17283 2954
rect 8477 2896 8482 2952
rect 8538 2896 17222 2952
rect 17278 2896 17283 2952
rect 8477 2894 17283 2896
rect 8477 2891 8543 2894
rect 17217 2891 17283 2894
rect 17953 2954 18019 2957
rect 22200 2954 23000 2984
rect 17953 2952 23000 2954
rect 17953 2896 17958 2952
rect 18014 2896 23000 2952
rect 17953 2894 23000 2896
rect 17953 2891 18019 2894
rect 22200 2864 23000 2894
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 2630 2620 2636 2684
rect 2700 2682 2706 2684
rect 3325 2682 3391 2685
rect 2700 2680 3391 2682
rect 2700 2624 3330 2680
rect 3386 2624 3391 2680
rect 2700 2622 3391 2624
rect 2700 2620 2706 2622
rect 3325 2619 3391 2622
rect 9397 2682 9463 2685
rect 10726 2682 10732 2684
rect 9397 2680 10732 2682
rect 9397 2624 9402 2680
rect 9458 2624 10732 2680
rect 9397 2622 10732 2624
rect 9397 2619 9463 2622
rect 10726 2620 10732 2622
rect 10796 2620 10802 2684
rect 0 2546 800 2576
rect 3049 2546 3115 2549
rect 0 2544 3115 2546
rect 0 2488 3054 2544
rect 3110 2488 3115 2544
rect 0 2486 3115 2488
rect 3328 2546 3388 2619
rect 4521 2546 4587 2549
rect 3328 2544 4587 2546
rect 3328 2488 4526 2544
rect 4582 2488 4587 2544
rect 3328 2486 4587 2488
rect 0 2456 800 2486
rect 3049 2483 3115 2486
rect 4521 2483 4587 2486
rect 16062 2484 16068 2548
rect 16132 2546 16138 2548
rect 21265 2546 21331 2549
rect 22200 2546 23000 2576
rect 16132 2544 23000 2546
rect 16132 2488 21270 2544
rect 21326 2488 23000 2544
rect 16132 2486 23000 2488
rect 16132 2484 16138 2486
rect 21265 2483 21331 2486
rect 22200 2456 23000 2486
rect 3417 2410 3483 2413
rect 9438 2410 9444 2412
rect 3417 2408 9444 2410
rect 3417 2352 3422 2408
rect 3478 2352 9444 2408
rect 3417 2350 9444 2352
rect 3417 2347 3483 2350
rect 9438 2348 9444 2350
rect 9508 2348 9514 2412
rect 13 2274 79 2277
rect 13 2272 1042 2274
rect 13 2216 18 2272
rect 74 2216 1042 2272
rect 13 2214 1042 2216
rect 13 2211 79 2214
rect 0 2002 800 2032
rect 982 2002 1042 2214
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 3877 2002 3943 2005
rect 0 2000 3943 2002
rect 0 1944 3882 2000
rect 3938 1944 3943 2000
rect 0 1942 3943 1944
rect 0 1912 800 1942
rect 3877 1939 3943 1942
rect 19793 2002 19859 2005
rect 22200 2002 23000 2032
rect 19793 2000 23000 2002
rect 19793 1944 19798 2000
rect 19854 1944 23000 2000
rect 19793 1942 23000 1944
rect 19793 1939 19859 1942
rect 22200 1912 23000 1942
rect 0 1594 800 1624
rect 4061 1594 4127 1597
rect 0 1592 4127 1594
rect 0 1536 4066 1592
rect 4122 1536 4127 1592
rect 0 1534 4127 1536
rect 0 1504 800 1534
rect 4061 1531 4127 1534
rect 20529 1594 20595 1597
rect 22200 1594 23000 1624
rect 20529 1592 23000 1594
rect 20529 1536 20534 1592
rect 20590 1536 23000 1592
rect 20529 1534 23000 1536
rect 20529 1531 20595 1534
rect 22200 1504 23000 1534
rect 13118 1260 13124 1324
rect 13188 1322 13194 1324
rect 20253 1322 20319 1325
rect 13188 1320 20319 1322
rect 13188 1264 20258 1320
rect 20314 1264 20319 1320
rect 13188 1262 20319 1264
rect 13188 1260 13194 1262
rect 20253 1259 20319 1262
rect 0 1050 800 1080
rect 2129 1050 2195 1053
rect 0 1048 2195 1050
rect 0 992 2134 1048
rect 2190 992 2195 1048
rect 0 990 2195 992
rect 0 960 800 990
rect 2129 987 2195 990
rect 18321 1050 18387 1053
rect 22200 1050 23000 1080
rect 18321 1048 23000 1050
rect 18321 992 18326 1048
rect 18382 992 23000 1048
rect 18321 990 23000 992
rect 18321 987 18387 990
rect 22200 960 23000 990
rect 20069 914 20135 917
rect 20069 912 21282 914
rect 20069 856 20074 912
rect 20130 856 21282 912
rect 20069 854 21282 856
rect 20069 851 20135 854
rect 0 642 800 672
rect 3417 642 3483 645
rect 0 640 3483 642
rect 0 584 3422 640
rect 3478 584 3483 640
rect 0 582 3483 584
rect 21222 642 21282 854
rect 22200 642 23000 672
rect 21222 582 23000 642
rect 0 552 800 582
rect 3417 579 3483 582
rect 22200 552 23000 582
rect 0 234 800 264
rect 3233 234 3299 237
rect 0 232 3299 234
rect 0 176 3238 232
rect 3294 176 3299 232
rect 0 174 3299 176
rect 0 144 800 174
rect 3233 171 3299 174
rect 20253 234 20319 237
rect 22200 234 23000 264
rect 20253 232 23000 234
rect 20253 176 20258 232
rect 20314 176 23000 232
rect 20253 174 23000 176
rect 20253 171 20319 174
rect 22200 144 23000 174
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 9444 17036 9508 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 4292 16764 4356 16828
rect 2268 16628 2332 16692
rect 16068 16688 16132 16692
rect 16068 16632 16082 16688
rect 16082 16632 16132 16688
rect 16068 16628 16132 16632
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 5028 15872 5092 15876
rect 5028 15816 5078 15872
rect 5078 15816 5092 15872
rect 5028 15812 5092 15816
rect 10732 15872 10796 15876
rect 10732 15816 10746 15872
rect 10746 15816 10796 15872
rect 10732 15812 10796 15816
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 2636 15540 2700 15604
rect 3372 15268 3436 15332
rect 9260 15268 9324 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 2084 14996 2148 15060
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 2452 14316 2516 14380
rect 4476 14180 4540 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 3188 13908 3252 13972
rect 19012 13908 19076 13972
rect 5948 13772 6012 13836
rect 7604 13772 7668 13836
rect 12572 13832 12636 13836
rect 12572 13776 12586 13832
rect 12586 13776 12636 13832
rect 12572 13772 12636 13776
rect 13124 13832 13188 13836
rect 13124 13776 13138 13832
rect 13138 13776 13188 13832
rect 13124 13772 13188 13776
rect 18828 13772 18892 13836
rect 4844 13636 4908 13700
rect 7420 13696 7484 13700
rect 7420 13640 7470 13696
rect 7470 13640 7484 13696
rect 7420 13636 7484 13640
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 18644 13364 18708 13428
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 4292 12956 4356 13020
rect 4108 12820 4172 12884
rect 11100 12820 11164 12884
rect 12756 12880 12820 12884
rect 12756 12824 12770 12880
rect 12770 12824 12820 12880
rect 12756 12820 12820 12824
rect 12020 12548 12084 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 5764 12336 5828 12340
rect 5764 12280 5778 12336
rect 5778 12280 5828 12336
rect 5764 12276 5828 12280
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6868 11052 6932 11116
rect 19932 11052 19996 11116
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 17908 10644 17972 10708
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5028 9964 5092 10028
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 9628 8740 9692 8804
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 17172 8664 17236 8668
rect 17172 8608 17186 8664
rect 17186 8608 17236 8664
rect 3924 8468 3988 8532
rect 6868 8468 6932 8532
rect 17172 8604 17236 8608
rect 6684 8196 6748 8260
rect 18828 8332 18892 8396
rect 11836 8196 11900 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 9628 8120 9692 8124
rect 9628 8064 9642 8120
rect 9642 8064 9692 8120
rect 9628 8060 9692 8064
rect 4476 7924 4540 7988
rect 8340 7924 8404 7988
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 2084 7516 2148 7580
rect 7972 7244 8036 7308
rect 11100 7244 11164 7308
rect 16988 7168 17052 7172
rect 16988 7112 17038 7168
rect 17038 7112 17052 7168
rect 16988 7108 17052 7112
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 3372 6972 3436 7036
rect 4844 6564 4908 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 5028 6428 5092 6492
rect 19012 6488 19076 6492
rect 19012 6432 19026 6488
rect 19026 6432 19076 6488
rect 19012 6428 19076 6432
rect 5764 6156 5828 6220
rect 6868 6020 6932 6084
rect 11836 6020 11900 6084
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 5948 5612 6012 5676
rect 7420 5672 7484 5676
rect 7420 5616 7470 5672
rect 7470 5616 7484 5672
rect 7420 5612 7484 5616
rect 17172 5476 17236 5540
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 16988 5128 17052 5132
rect 16988 5072 17002 5128
rect 17002 5072 17052 5128
rect 16988 5068 17052 5072
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 4108 4796 4172 4860
rect 2268 4720 2332 4724
rect 2268 4664 2282 4720
rect 2282 4664 2332 4720
rect 2268 4660 2332 4664
rect 7604 4720 7668 4724
rect 7604 4664 7618 4720
rect 7618 4664 7668 4720
rect 7604 4660 7668 4664
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 8340 3980 8404 4044
rect 9260 4040 9324 4044
rect 9260 3984 9274 4040
rect 9274 3984 9324 4040
rect 9260 3980 9324 3984
rect 17908 3980 17972 4044
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 18644 3708 18708 3772
rect 2452 3572 2516 3636
rect 12572 3572 12636 3636
rect 12756 3436 12820 3500
rect 3924 3300 3988 3364
rect 7972 3300 8036 3364
rect 19932 3300 19996 3364
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 3188 2892 3252 2956
rect 6684 2892 6748 2956
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 2636 2620 2700 2684
rect 10732 2620 10796 2684
rect 16068 2484 16132 2548
rect 9444 2348 9508 2412
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 13124 1260 13188 1324
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 2267 16692 2333 16693
rect 2267 16628 2268 16692
rect 2332 16628 2333 16692
rect 2267 16627 2333 16628
rect 2083 15060 2149 15061
rect 2083 14996 2084 15060
rect 2148 14996 2149 15060
rect 2083 14995 2149 14996
rect 2086 7581 2146 14995
rect 2083 7580 2149 7581
rect 2083 7516 2084 7580
rect 2148 7516 2149 7580
rect 2083 7515 2149 7516
rect 2270 4725 2330 16627
rect 3543 15808 3863 16832
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 4291 16828 4357 16829
rect 4291 16764 4292 16828
rect 4356 16764 4357 16828
rect 4291 16763 4357 16764
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 2635 15604 2701 15605
rect 2635 15540 2636 15604
rect 2700 15540 2701 15604
rect 2635 15539 2701 15540
rect 2451 14380 2517 14381
rect 2451 14316 2452 14380
rect 2516 14316 2517 14380
rect 2451 14315 2517 14316
rect 2267 4724 2333 4725
rect 2267 4660 2268 4724
rect 2332 4660 2333 4724
rect 2267 4659 2333 4660
rect 2454 3637 2514 14315
rect 2451 3636 2517 3637
rect 2451 3572 2452 3636
rect 2516 3572 2517 3636
rect 2451 3571 2517 3572
rect 2638 2685 2698 15539
rect 3371 15332 3437 15333
rect 3371 15268 3372 15332
rect 3436 15268 3437 15332
rect 3371 15267 3437 15268
rect 3187 13972 3253 13973
rect 3187 13908 3188 13972
rect 3252 13908 3253 13972
rect 3187 13907 3253 13908
rect 3190 2957 3250 13907
rect 3374 7037 3434 15267
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 4294 13021 4354 16763
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 5027 15876 5093 15877
rect 5027 15812 5028 15876
rect 5092 15812 5093 15876
rect 5027 15811 5093 15812
rect 4475 14244 4541 14245
rect 4475 14180 4476 14244
rect 4540 14180 4541 14244
rect 4475 14179 4541 14180
rect 4291 13020 4357 13021
rect 4291 12956 4292 13020
rect 4356 12956 4357 13020
rect 4291 12955 4357 12956
rect 4107 12884 4173 12885
rect 4107 12820 4108 12884
rect 4172 12820 4173 12884
rect 4107 12819 4173 12820
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3923 8532 3989 8533
rect 3923 8468 3924 8532
rect 3988 8468 3989 8532
rect 3923 8467 3989 8468
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3371 7036 3437 7037
rect 3371 6972 3372 7036
rect 3436 6972 3437 7036
rect 3371 6971 3437 6972
rect 3543 6016 3863 7040
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3187 2956 3253 2957
rect 3187 2892 3188 2956
rect 3252 2892 3253 2956
rect 3187 2891 3253 2892
rect 3543 2752 3863 3776
rect 3926 3365 3986 8467
rect 4110 4861 4170 12819
rect 4478 7989 4538 14179
rect 4843 13700 4909 13701
rect 4843 13636 4844 13700
rect 4908 13636 4909 13700
rect 4843 13635 4909 13636
rect 4475 7988 4541 7989
rect 4475 7924 4476 7988
rect 4540 7924 4541 7988
rect 4475 7923 4541 7924
rect 4846 6629 4906 13635
rect 5030 10029 5090 15811
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 5947 13836 6013 13837
rect 5947 13772 5948 13836
rect 6012 13772 6013 13836
rect 5947 13771 6013 13772
rect 5763 12340 5829 12341
rect 5763 12276 5764 12340
rect 5828 12276 5829 12340
rect 5763 12275 5829 12276
rect 5027 10028 5093 10029
rect 5027 9964 5028 10028
rect 5092 9964 5093 10028
rect 5027 9963 5093 9964
rect 4843 6628 4909 6629
rect 4843 6564 4844 6628
rect 4908 6564 4909 6628
rect 4843 6563 4909 6564
rect 5030 6493 5090 9963
rect 5027 6492 5093 6493
rect 5027 6428 5028 6492
rect 5092 6428 5093 6492
rect 5027 6427 5093 6428
rect 5766 6221 5826 12275
rect 5763 6220 5829 6221
rect 5763 6156 5764 6220
rect 5828 6156 5829 6220
rect 5763 6155 5829 6156
rect 5950 5677 6010 13771
rect 6142 13088 6462 14112
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 9443 17100 9509 17101
rect 9443 17036 9444 17100
rect 9508 17036 9509 17100
rect 9443 17035 9509 17036
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 9259 15332 9325 15333
rect 9259 15268 9260 15332
rect 9324 15268 9325 15332
rect 9259 15267 9325 15268
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 7603 13836 7669 13837
rect 7603 13772 7604 13836
rect 7668 13772 7669 13836
rect 7603 13771 7669 13772
rect 7419 13700 7485 13701
rect 7419 13636 7420 13700
rect 7484 13636 7485 13700
rect 7419 13635 7485 13636
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6867 11116 6933 11117
rect 6867 11052 6868 11116
rect 6932 11052 6933 11116
rect 6867 11051 6933 11052
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6870 8533 6930 11051
rect 6867 8532 6933 8533
rect 6867 8468 6868 8532
rect 6932 8468 6933 8532
rect 6867 8467 6933 8468
rect 6683 8260 6749 8261
rect 6683 8196 6684 8260
rect 6748 8196 6749 8260
rect 6683 8195 6749 8196
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 5947 5676 6013 5677
rect 5947 5612 5948 5676
rect 6012 5612 6013 5676
rect 5947 5611 6013 5612
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 4107 4860 4173 4861
rect 4107 4796 4108 4860
rect 4172 4796 4173 4860
rect 4107 4795 4173 4796
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 3923 3364 3989 3365
rect 3923 3300 3924 3364
rect 3988 3300 3989 3364
rect 3923 3299 3989 3300
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 2635 2684 2701 2685
rect 2635 2620 2636 2684
rect 2700 2620 2701 2684
rect 2635 2619 2701 2620
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6686 2957 6746 8195
rect 6870 6085 6930 8467
rect 6867 6084 6933 6085
rect 6867 6020 6868 6084
rect 6932 6020 6933 6084
rect 6867 6019 6933 6020
rect 7422 5677 7482 13635
rect 7419 5676 7485 5677
rect 7419 5612 7420 5676
rect 7484 5612 7485 5676
rect 7419 5611 7485 5612
rect 7606 4725 7666 13771
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8339 7988 8405 7989
rect 8339 7924 8340 7988
rect 8404 7924 8405 7988
rect 8339 7923 8405 7924
rect 7971 7308 8037 7309
rect 7971 7244 7972 7308
rect 8036 7244 8037 7308
rect 7971 7243 8037 7244
rect 7603 4724 7669 4725
rect 7603 4660 7604 4724
rect 7668 4660 7669 4724
rect 7603 4659 7669 4660
rect 7974 3365 8034 7243
rect 8342 4045 8402 7923
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8339 4044 8405 4045
rect 8339 3980 8340 4044
rect 8404 3980 8405 4044
rect 8339 3979 8405 3980
rect 8741 3840 9061 4864
rect 9262 4045 9322 15267
rect 9259 4044 9325 4045
rect 9259 3980 9260 4044
rect 9324 3980 9325 4044
rect 9259 3979 9325 3980
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 7971 3364 8037 3365
rect 7971 3300 7972 3364
rect 8036 3300 8037 3364
rect 7971 3299 8037 3300
rect 6683 2956 6749 2957
rect 6683 2892 6684 2956
rect 6748 2892 6749 2956
rect 6683 2891 6749 2892
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 9446 2413 9506 17035
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 10731 15876 10797 15877
rect 10731 15812 10732 15876
rect 10796 15812 10797 15876
rect 10731 15811 10797 15812
rect 9627 8804 9693 8805
rect 9627 8740 9628 8804
rect 9692 8740 9693 8804
rect 9627 8739 9693 8740
rect 9630 8125 9690 8739
rect 9627 8124 9693 8125
rect 9627 8060 9628 8124
rect 9692 8060 9693 8124
rect 9627 8059 9693 8060
rect 10734 2685 10794 15811
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16067 16692 16133 16693
rect 16067 16628 16068 16692
rect 16132 16628 16133 16692
rect 16067 16627 16133 16628
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 12571 13836 12637 13837
rect 12571 13772 12572 13836
rect 12636 13772 12637 13836
rect 12571 13771 12637 13772
rect 13123 13836 13189 13837
rect 13123 13772 13124 13836
rect 13188 13772 13189 13836
rect 13123 13771 13189 13772
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11099 12884 11165 12885
rect 11099 12820 11100 12884
rect 11164 12820 11165 12884
rect 11099 12819 11165 12820
rect 11102 7309 11162 12819
rect 11340 12000 11660 13024
rect 12019 12612 12085 12613
rect 12019 12548 12020 12612
rect 12084 12548 12085 12612
rect 12019 12547 12085 12548
rect 12022 12450 12082 12547
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11838 12390 12082 12450
rect 11838 8261 11898 12390
rect 11835 8260 11901 8261
rect 11835 8196 11836 8260
rect 11900 8196 11901 8260
rect 11835 8195 11901 8196
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11099 7308 11165 7309
rect 11099 7244 11100 7308
rect 11164 7244 11165 7308
rect 11099 7243 11165 7244
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11838 6085 11898 8195
rect 11835 6084 11901 6085
rect 11835 6020 11836 6084
rect 11900 6020 11901 6084
rect 11835 6019 11901 6020
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 12574 3637 12634 13771
rect 12755 12884 12821 12885
rect 12755 12820 12756 12884
rect 12820 12820 12821 12884
rect 12755 12819 12821 12820
rect 12571 3636 12637 3637
rect 12571 3572 12572 3636
rect 12636 3572 12637 3636
rect 12571 3571 12637 3572
rect 12758 3501 12818 12819
rect 12755 3500 12821 3501
rect 12755 3436 12756 3500
rect 12820 3436 12821 3500
rect 12755 3435 12821 3436
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 10731 2684 10797 2685
rect 10731 2620 10732 2684
rect 10796 2620 10797 2684
rect 10731 2619 10797 2620
rect 9443 2412 9509 2413
rect 9443 2348 9444 2412
rect 9508 2348 9509 2412
rect 9443 2347 9509 2348
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13126 1325 13186 13771
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16070 2549 16130 16627
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19011 13972 19077 13973
rect 19011 13908 19012 13972
rect 19076 13908 19077 13972
rect 19011 13907 19077 13908
rect 18827 13836 18893 13837
rect 18827 13772 18828 13836
rect 18892 13772 18893 13836
rect 18827 13771 18893 13772
rect 18643 13428 18709 13429
rect 18643 13364 18644 13428
rect 18708 13364 18709 13428
rect 18643 13363 18709 13364
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 17907 10708 17973 10709
rect 17907 10644 17908 10708
rect 17972 10644 17973 10708
rect 17907 10643 17973 10644
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 17171 8668 17237 8669
rect 17171 8604 17172 8668
rect 17236 8604 17237 8668
rect 17171 8603 17237 8604
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16987 7172 17053 7173
rect 16987 7108 16988 7172
rect 17052 7108 17053 7172
rect 16987 7107 17053 7108
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16990 5133 17050 7107
rect 17174 5541 17234 8603
rect 17171 5540 17237 5541
rect 17171 5476 17172 5540
rect 17236 5476 17237 5540
rect 17171 5475 17237 5476
rect 16987 5132 17053 5133
rect 16987 5068 16988 5132
rect 17052 5068 17053 5132
rect 16987 5067 17053 5068
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 17910 4045 17970 10643
rect 17907 4044 17973 4045
rect 17907 3980 17908 4044
rect 17972 3980 17973 4044
rect 17907 3979 17973 3980
rect 18646 3773 18706 13363
rect 18830 8397 18890 13771
rect 18827 8396 18893 8397
rect 18827 8332 18828 8396
rect 18892 8332 18893 8396
rect 18827 8331 18893 8332
rect 19014 6493 19074 13907
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19931 11116 19997 11117
rect 19931 11052 19932 11116
rect 19996 11052 19997 11116
rect 19931 11051 19997 11052
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19011 6492 19077 6493
rect 19011 6428 19012 6492
rect 19076 6428 19077 6492
rect 19011 6427 19077 6428
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 18643 3772 18709 3773
rect 18643 3708 18644 3772
rect 18708 3708 18709 3772
rect 18643 3707 18709 3708
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16067 2548 16133 2549
rect 16067 2484 16068 2548
rect 16132 2484 16133 2548
rect 16067 2483 16133 2484
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 2752 19457 3776
rect 19934 3365 19994 11051
rect 19931 3364 19997 3365
rect 19931 3300 19932 3364
rect 19996 3300 19997 3364
rect 19931 3299 19997 3300
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
rect 13123 1324 13189 1325
rect 13123 1260 13124 1324
rect 13188 1260 13189 1324
rect 13123 1259 13189 1260
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__A
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A
timestamp 1649977179
transform 1 0 3220 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__A
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__A
timestamp 1649977179
transform -1 0 3036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A
timestamp 1649977179
transform -1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__A
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__A
timestamp 1649977179
transform -1 0 4692 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A
timestamp 1649977179
transform 1 0 5704 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__A
timestamp 1649977179
transform 1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A
timestamp 1649977179
transform -1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__A
timestamp 1649977179
transform 1 0 6716 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A
timestamp 1649977179
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A
timestamp 1649977179
transform 1 0 18400 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A
timestamp 1649977179
transform 1 0 18032 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__A
timestamp 1649977179
transform -1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A
timestamp 1649977179
transform -1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A
timestamp 1649977179
transform -1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__A
timestamp 1649977179
transform -1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A
timestamp 1649977179
transform 1 0 19412 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A
timestamp 1649977179
transform -1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__A
timestamp 1649977179
transform 1 0 18400 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A
timestamp 1649977179
transform -1 0 17664 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A
timestamp 1649977179
transform -1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A
timestamp 1649977179
transform -1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 12788 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 8740 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 5888 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 12696 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 3956 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 4784 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 3956 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3956 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 5612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 5796 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 5980 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 16284 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 18400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 17296 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform 1 0 17112 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 17480 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 4508 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 9108 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 7636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 12788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 5336 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 8464 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 6532 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 10396 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 9660 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 5520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 6716 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 8740 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 6532 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 7360 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_3.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 7544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 7360 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 5428 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_7.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 5060 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 9384 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12972 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_11.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 12880 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_13.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 14720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_15.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 13616 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10212 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_19.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 10672 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_21.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 12604 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_23.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__A0
timestamp 1649977179
transform -1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 17664 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10948 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10580 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4324 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 5888 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 1932 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5428 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_9.mux_l2_in_1__A0
timestamp 1649977179
transform 1 0 8096 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6992 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8188 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10396 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_25.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10580 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8280 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 6900 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 18400 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 17664 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 13248 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 15088 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_1__A0
timestamp 1649977179
transform -1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A0
timestamp 1649977179
transform -1 0 13432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 13340 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_2.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_2__A1
timestamp 1649977179
transform -1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_3__A1
timestamp 1649977179
transform -1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A0
timestamp 1649977179
transform 1 0 16192 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_4__A1
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_5__A0
timestamp 1649977179
transform -1 0 15180 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A0
timestamp 1649977179
transform 1 0 19320 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_6__A1
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 18492 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_0__A0
timestamp 1649977179
transform 1 0 18768 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_2__A1
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l2_in_3__A1
timestamp 1649977179
transform 1 0 11592 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11040 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 11040 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_16.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_2__A0
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_3__A1
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_32.mux_l2_in_1__A1
timestamp 1649977179
transform 1 0 13248 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp 1649977179
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_93
timestamp 1649977179
transform 1 0 9660 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_98
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_123
timestamp 1649977179
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_127
timestamp 1649977179
transform 1 0 12788 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_151
timestamp 1649977179
transform 1 0 14996 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_163
timestamp 1649977179
transform 1 0 16100 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1649977179
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_179
timestamp 1649977179
transform 1 0 17572 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_191
timestamp 1649977179
transform 1 0 18676 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_13 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_32
timestamp 1649977179
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_67
timestamp 1649977179
transform 1 0 7268 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_72
timestamp 1649977179
transform 1 0 7728 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_90
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_106
timestamp 1649977179
transform 1 0 10856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_116
timestamp 1649977179
transform 1 0 11776 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_121
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_131
timestamp 1649977179
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_136
timestamp 1649977179
transform 1 0 13616 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_140
timestamp 1649977179
transform 1 0 13984 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_144
timestamp 1649977179
transform 1 0 14352 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 1649977179
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_173
timestamp 1649977179
transform 1 0 17020 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_185
timestamp 1649977179
transform 1 0 18124 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_191
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1649977179
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_45
timestamp 1649977179
transform 1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_57
timestamp 1649977179
transform 1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_68
timestamp 1649977179
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_72
timestamp 1649977179
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_101
timestamp 1649977179
transform 1 0 10396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_112
timestamp 1649977179
transform 1 0 11408 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_117
timestamp 1649977179
transform 1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_123
timestamp 1649977179
transform 1 0 12420 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_128
timestamp 1649977179
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_134
timestamp 1649977179
transform 1 0 13432 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_145
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_156
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_167
timestamp 1649977179
transform 1 0 16468 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_171
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_176
timestamp 1649977179
transform 1 0 17296 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 1649977179
transform 1 0 17848 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_188
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_20
timestamp 1649977179
transform 1 0 2944 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1649977179
transform 1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_36
timestamp 1649977179
transform 1 0 4416 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_47
timestamp 1649977179
transform 1 0 5428 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_66
timestamp 1649977179
transform 1 0 7176 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_71
timestamp 1649977179
transform 1 0 7636 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_84
timestamp 1649977179
transform 1 0 8832 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_95
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_108
timestamp 1649977179
transform 1 0 11040 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_116
timestamp 1649977179
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_121
timestamp 1649977179
transform 1 0 12236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_126
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_3_133
timestamp 1649977179
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_138
timestamp 1649977179
transform 1 0 13800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_143
timestamp 1649977179
transform 1 0 14260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_148
timestamp 1649977179
transform 1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_189
timestamp 1649977179
transform 1 0 18492 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_194
timestamp 1649977179
transform 1 0 18952 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_200
timestamp 1649977179
transform 1 0 19504 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_204
timestamp 1649977179
transform 1 0 19872 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_209
timestamp 1649977179
transform 1 0 20332 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_42
timestamp 1649977179
transform 1 0 4968 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_57
timestamp 1649977179
transform 1 0 6348 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_62
timestamp 1649977179
transform 1 0 6808 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_72
timestamp 1649977179
transform 1 0 7728 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_94
timestamp 1649977179
transform 1 0 9752 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_101
timestamp 1649977179
transform 1 0 10396 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 1649977179
transform 1 0 10856 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_111
timestamp 1649977179
transform 1 0 11316 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_129
timestamp 1649977179
transform 1 0 12972 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_134
timestamp 1649977179
transform 1 0 13432 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_157
timestamp 1649977179
transform 1 0 15548 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp 1649977179
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_173
timestamp 1649977179
transform 1 0 17020 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_178
timestamp 1649977179
transform 1 0 17480 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_182
timestamp 1649977179
transform 1 0 17848 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_188
timestamp 1649977179
transform 1 0 18400 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_201
timestamp 1649977179
transform 1 0 19596 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_219
timestamp 1649977179
transform 1 0 21252 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_37
timestamp 1649977179
transform 1 0 4508 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_47
timestamp 1649977179
transform 1 0 5428 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_53
timestamp 1649977179
transform 1 0 5980 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_67
timestamp 1649977179
transform 1 0 7268 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_71
timestamp 1649977179
transform 1 0 7636 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_98
timestamp 1649977179
transform 1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_123
timestamp 1649977179
transform 1 0 12420 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_127
timestamp 1649977179
transform 1 0 12788 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_154
timestamp 1649977179
transform 1 0 15272 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_159
timestamp 1649977179
transform 1 0 15732 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_164
timestamp 1649977179
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1649977179
transform 1 0 17848 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_192
timestamp 1649977179
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_210
timestamp 1649977179
transform 1 0 20424 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 1649977179
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_8
timestamp 1649977179
transform 1 0 1840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 1649977179
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_45
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_76
timestamp 1649977179
transform 1 0 8096 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_81
timestamp 1649977179
transform 1 0 8556 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 1649977179
transform 1 0 11776 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 1649977179
transform 1 0 12144 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_150
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_161
timestamp 1649977179
transform 1 0 15916 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_172
timestamp 1649977179
transform 1 0 16928 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_176
timestamp 1649977179
transform 1 0 17296 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_206
timestamp 1649977179
transform 1 0 20056 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_217
timestamp 1649977179
transform 1 0 21068 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_13
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_24
timestamp 1649977179
transform 1 0 3312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_38
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_43
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_67
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_72
timestamp 1649977179
transform 1 0 7728 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_77
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_82
timestamp 1649977179
transform 1 0 8648 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_98
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_144
timestamp 1649977179
transform 1 0 14352 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_148
timestamp 1649977179
transform 1 0 14720 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 1649977179
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_178
timestamp 1649977179
transform 1 0 17480 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_189
timestamp 1649977179
transform 1 0 18492 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_197
timestamp 1649977179
transform 1 0 19228 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_208
timestamp 1649977179
transform 1 0 20240 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_219
timestamp 1649977179
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_9
timestamp 1649977179
transform 1 0 1932 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_20
timestamp 1649977179
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_36
timestamp 1649977179
transform 1 0 4416 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_54
timestamp 1649977179
transform 1 0 6072 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_59
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_71
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 1649977179
transform 1 0 10396 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_105
timestamp 1649977179
transform 1 0 10764 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_119
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_124
timestamp 1649977179
transform 1 0 12512 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_128
timestamp 1649977179
transform 1 0 12880 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_149
timestamp 1649977179
transform 1 0 14812 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_158
timestamp 1649977179
transform 1 0 15640 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_163
timestamp 1649977179
transform 1 0 16100 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_173
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_178
timestamp 1649977179
transform 1 0 17480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_182
timestamp 1649977179
transform 1 0 17848 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_188
timestamp 1649977179
transform 1 0 18400 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_203
timestamp 1649977179
transform 1 0 19780 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_9
timestamp 1649977179
transform 1 0 1932 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1649977179
transform 1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_24
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_29
timestamp 1649977179
transform 1 0 3772 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_33
timestamp 1649977179
transform 1 0 4140 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_43
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_101
timestamp 1649977179
transform 1 0 10396 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_109
timestamp 1649977179
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_122
timestamp 1649977179
transform 1 0 12328 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_128
timestamp 1649977179
transform 1 0 12880 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_146
timestamp 1649977179
transform 1 0 14536 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_151
timestamp 1649977179
transform 1 0 14996 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 1649977179
transform 1 0 15456 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_166
timestamp 1649977179
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_185
timestamp 1649977179
transform 1 0 18124 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_197
timestamp 1649977179
transform 1 0 19228 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_215
timestamp 1649977179
transform 1 0 20884 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_221
timestamp 1649977179
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_24
timestamp 1649977179
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_38
timestamp 1649977179
transform 1 0 4600 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp 1649977179
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 1649977179
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_108
timestamp 1649977179
transform 1 0 11040 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 1649977179
transform 1 0 12696 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_146
timestamp 1649977179
transform 1 0 14536 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1649977179
transform 1 0 14996 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_156
timestamp 1649977179
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_178
timestamp 1649977179
transform 1 0 17480 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_25
timestamp 1649977179
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_36
timestamp 1649977179
transform 1 0 4416 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_41
timestamp 1649977179
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_46
timestamp 1649977179
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_60
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_71
timestamp 1649977179
transform 1 0 7636 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_76
timestamp 1649977179
transform 1 0 8096 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_84
timestamp 1649977179
transform 1 0 8832 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_88
timestamp 1649977179
transform 1 0 9200 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_103
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_107
timestamp 1649977179
transform 1 0 10948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1649977179
transform 1 0 11960 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_129
timestamp 1649977179
transform 1 0 12972 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_140
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_11_160
timestamp 1649977179
transform 1 0 15824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1649977179
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_178
timestamp 1649977179
transform 1 0 17480 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_189
timestamp 1649977179
transform 1 0 18492 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_209
timestamp 1649977179
transform 1 0 20332 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_9
timestamp 1649977179
transform 1 0 1932 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_22
timestamp 1649977179
transform 1 0 3128 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_61
timestamp 1649977179
transform 1 0 6716 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1649977179
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_87
timestamp 1649977179
transform 1 0 9108 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1649977179
transform 1 0 9568 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_103
timestamp 1649977179
transform 1 0 10580 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_107
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_110
timestamp 1649977179
transform 1 0 11224 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_120
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_127
timestamp 1649977179
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_131
timestamp 1649977179
transform 1 0 13156 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_135
timestamp 1649977179
transform 1 0 13524 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_150
timestamp 1649977179
transform 1 0 14904 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_185
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_207
timestamp 1649977179
transform 1 0 20148 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_217
timestamp 1649977179
transform 1 0 21068 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_8
timestamp 1649977179
transform 1 0 1840 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_26
timestamp 1649977179
transform 1 0 3496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_30
timestamp 1649977179
transform 1 0 3864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_47
timestamp 1649977179
transform 1 0 5428 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_60
timestamp 1649977179
transform 1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_72
timestamp 1649977179
transform 1 0 7728 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_83
timestamp 1649977179
transform 1 0 8740 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_101
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_106
timestamp 1649977179
transform 1 0 10856 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_131
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1649977179
transform 1 0 14168 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_153
timestamp 1649977179
transform 1 0 15180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_164
timestamp 1649977179
transform 1 0 16192 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_186
timestamp 1649977179
transform 1 0 18216 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 1649977179
transform 1 0 18768 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_203
timestamp 1649977179
transform 1 0 19780 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_9
timestamp 1649977179
transform 1 0 1932 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_14
timestamp 1649977179
transform 1 0 2392 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_18
timestamp 1649977179
transform 1 0 2760 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_22
timestamp 1649977179
transform 1 0 3128 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_37
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_42
timestamp 1649977179
transform 1 0 4968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 1649977179
transform 1 0 5336 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_56
timestamp 1649977179
transform 1 0 6256 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_67
timestamp 1649977179
transform 1 0 7268 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_78
timestamp 1649977179
transform 1 0 8280 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_95
timestamp 1649977179
transform 1 0 9844 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_113
timestamp 1649977179
transform 1 0 11500 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_120
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1649977179
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_157
timestamp 1649977179
transform 1 0 15548 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_168
timestamp 1649977179
transform 1 0 16560 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_179
timestamp 1649977179
transform 1 0 17572 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_190
timestamp 1649977179
transform 1 0 18584 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_203
timestamp 1649977179
transform 1 0 19780 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_214
timestamp 1649977179
transform 1 0 20792 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_9
timestamp 1649977179
transform 1 0 1932 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 1649977179
transform 1 0 2300 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_28
timestamp 1649977179
transform 1 0 3680 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_45
timestamp 1649977179
transform 1 0 5244 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_50
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_70
timestamp 1649977179
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_80
timestamp 1649977179
transform 1 0 8464 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_85
timestamp 1649977179
transform 1 0 8924 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_89
timestamp 1649977179
transform 1 0 9292 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_99
timestamp 1649977179
transform 1 0 10212 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_128
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_138
timestamp 1649977179
transform 1 0 13800 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_142
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_163
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_178
timestamp 1649977179
transform 1 0 17480 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_196
timestamp 1649977179
transform 1 0 19136 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_15_203
timestamp 1649977179
transform 1 0 19780 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_7
timestamp 1649977179
transform 1 0 1748 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_12
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_38
timestamp 1649977179
transform 1 0 4600 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_49
timestamp 1649977179
transform 1 0 5612 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1649977179
transform 1 0 6716 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 1649977179
transform 1 0 8556 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_95
timestamp 1649977179
transform 1 0 9844 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_101
timestamp 1649977179
transform 1 0 10396 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_105
timestamp 1649977179
transform 1 0 10764 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_136
timestamp 1649977179
transform 1 0 13616 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_143
timestamp 1649977179
transform 1 0 14260 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_161
timestamp 1649977179
transform 1 0 15916 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_178
timestamp 1649977179
transform 1 0 17480 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 1649977179
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_213
timestamp 1649977179
transform 1 0 20700 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_9
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_22
timestamp 1649977179
transform 1 0 3128 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_31
timestamp 1649977179
transform 1 0 3956 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_50
timestamp 1649977179
transform 1 0 5704 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1649977179
transform 1 0 6532 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_64
timestamp 1649977179
transform 1 0 6992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 1649977179
transform 1 0 8004 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_79
timestamp 1649977179
transform 1 0 8372 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_83
timestamp 1649977179
transform 1 0 8740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_95
timestamp 1649977179
transform 1 0 9844 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_106
timestamp 1649977179
transform 1 0 10856 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_116
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_138
timestamp 1649977179
transform 1 0 13800 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_150
timestamp 1649977179
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1649977179
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_185
timestamp 1649977179
transform 1 0 18124 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1649977179
transform 1 0 18400 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_203
timestamp 1649977179
transform 1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_210
timestamp 1649977179
transform 1 0 20424 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_8
timestamp 1649977179
transform 1 0 1840 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_31
timestamp 1649977179
transform 1 0 3956 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_37
timestamp 1649977179
transform 1 0 4508 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_48
timestamp 1649977179
transform 1 0 5520 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1649977179
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_63
timestamp 1649977179
transform 1 0 6900 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_66
timestamp 1649977179
transform 1 0 7176 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_82
timestamp 1649977179
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1649977179
transform 1 0 9200 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_92
timestamp 1649977179
transform 1 0 9568 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_102
timestamp 1649977179
transform 1 0 10488 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_120
timestamp 1649977179
transform 1 0 12144 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_148
timestamp 1649977179
transform 1 0 14720 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_183
timestamp 1649977179
transform 1 0 17940 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_208
timestamp 1649977179
transform 1 0 20240 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_220
timestamp 1649977179
transform 1 0 21344 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_9
timestamp 1649977179
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_20
timestamp 1649977179
transform 1 0 2944 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_42
timestamp 1649977179
transform 1 0 4968 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_66
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_70
timestamp 1649977179
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_106
timestamp 1649977179
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_123
timestamp 1649977179
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_162
timestamp 1649977179
transform 1 0 16008 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_178
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_197
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_208
timestamp 1649977179
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1649977179
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_7
timestamp 1649977179
transform 1 0 1748 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_22
timestamp 1649977179
transform 1 0 3128 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_38
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_43
timestamp 1649977179
transform 1 0 5060 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_76
timestamp 1649977179
transform 1 0 8096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_20_103
timestamp 1649977179
transform 1 0 10580 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_107
timestamp 1649977179
transform 1 0 10948 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_111
timestamp 1649977179
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_115
timestamp 1649977179
transform 1 0 11684 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 1649977179
transform 1 0 12052 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_123
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_127
timestamp 1649977179
transform 1 0 12788 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_131
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_134
timestamp 1649977179
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_149
timestamp 1649977179
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 1649977179
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_206
timestamp 1649977179
transform 1 0 20056 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_212
timestamp 1649977179
transform 1 0 20608 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_216
timestamp 1649977179
transform 1 0 20976 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_12
timestamp 1649977179
transform 1 0 2208 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_23
timestamp 1649977179
transform 1 0 3220 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_29
timestamp 1649977179
transform 1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_33
timestamp 1649977179
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_43
timestamp 1649977179
transform 1 0 5060 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1649977179
transform 1 0 6532 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_63
timestamp 1649977179
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_78
timestamp 1649977179
transform 1 0 8280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_90
timestamp 1649977179
transform 1 0 9384 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_126
timestamp 1649977179
transform 1 0 12696 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_131
timestamp 1649977179
transform 1 0 13156 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_135
timestamp 1649977179
transform 1 0 13524 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_139
timestamp 1649977179
transform 1 0 13892 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_143
timestamp 1649977179
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_154
timestamp 1649977179
transform 1 0 15272 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_172
timestamp 1649977179
transform 1 0 16928 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_176
timestamp 1649977179
transform 1 0 17296 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_180
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_204
timestamp 1649977179
transform 1 0 19872 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_215
timestamp 1649977179
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_12
timestamp 1649977179
transform 1 0 2208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_16
timestamp 1649977179
transform 1 0 2576 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_38
timestamp 1649977179
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_42
timestamp 1649977179
transform 1 0 4968 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_46
timestamp 1649977179
transform 1 0 5336 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_52
timestamp 1649977179
transform 1 0 5888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_57
timestamp 1649977179
transform 1 0 6348 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_75
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_79
timestamp 1649977179
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_103
timestamp 1649977179
transform 1 0 10580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_107
timestamp 1649977179
transform 1 0 10948 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_110
timestamp 1649977179
transform 1 0 11224 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_22_121 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_129
timestamp 1649977179
transform 1 0 12972 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_134
timestamp 1649977179
transform 1 0 13432 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_138
timestamp 1649977179
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_150
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_154
timestamp 1649977179
transform 1 0 15272 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_157
timestamp 1649977179
transform 1 0 15548 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_179
timestamp 1649977179
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_183
timestamp 1649977179
transform 1 0 17940 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_215
timestamp 1649977179
transform 1 0 20884 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1649977179
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_32
timestamp 1649977179
transform 1 0 4048 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_36
timestamp 1649977179
transform 1 0 4416 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_40
timestamp 1649977179
transform 1 0 4784 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1649977179
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1649977179
transform 1 0 7176 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_70
timestamp 1649977179
transform 1 0 7544 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 1649977179
transform 1 0 9384 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1649977179
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_117
timestamp 1649977179
transform 1 0 11868 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_134
timestamp 1649977179
transform 1 0 13432 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_152
timestamp 1649977179
transform 1 0 15088 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_163
timestamp 1649977179
transform 1 0 16100 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_196
timestamp 1649977179
transform 1 0 19136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_207
timestamp 1649977179
transform 1 0 20148 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_212
timestamp 1649977179
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_216
timestamp 1649977179
transform 1 0 20976 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_12
timestamp 1649977179
transform 1 0 2208 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_21
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_45
timestamp 1649977179
transform 1 0 5244 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_49
timestamp 1649977179
transform 1 0 5612 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_68
timestamp 1649977179
transform 1 0 7360 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_72
timestamp 1649977179
transform 1 0 7728 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_87
timestamp 1649977179
transform 1 0 9108 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_91
timestamp 1649977179
transform 1 0 9476 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_101
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_24_105 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_111
timestamp 1649977179
transform 1 0 11316 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_128 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12880 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_150
timestamp 1649977179
transform 1 0 14904 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_155
timestamp 1649977179
transform 1 0 15364 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_173
timestamp 1649977179
transform 1 0 17020 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_182
timestamp 1649977179
transform 1 0 17848 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1649977179
transform 1 0 18216 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_200
timestamp 1649977179
transform 1 0 19504 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1649977179
transform 1 0 20424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_17
timestamp 1649977179
transform 1 0 2668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_21
timestamp 1649977179
transform 1 0 3036 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_25
timestamp 1649977179
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_33
timestamp 1649977179
transform 1 0 4140 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_37
timestamp 1649977179
transform 1 0 4508 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_43
timestamp 1649977179
transform 1 0 5060 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_49
timestamp 1649977179
transform 1 0 5612 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1649977179
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_59
timestamp 1649977179
transform 1 0 6532 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_65
timestamp 1649977179
transform 1 0 7084 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_73
timestamp 1649977179
transform 1 0 7820 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_77
timestamp 1649977179
transform 1 0 8188 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_85
timestamp 1649977179
transform 1 0 8924 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_89
timestamp 1649977179
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1649977179
transform 1 0 10028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_101
timestamp 1649977179
transform 1 0 10396 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_106
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 1649977179
transform 1 0 11224 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_122
timestamp 1649977179
transform 1 0 12328 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_134
timestamp 1649977179
transform 1 0 13432 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_140
timestamp 1649977179
transform 1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1649977179
transform 1 0 16928 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_176
timestamp 1649977179
transform 1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_194
timestamp 1649977179
transform 1 0 18952 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_200
timestamp 1649977179
transform 1 0 19504 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1649977179
transform 1 0 19872 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1649977179
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1649977179
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_31
timestamp 1649977179
transform 1 0 3956 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_35
timestamp 1649977179
transform 1 0 4324 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1649977179
transform 1 0 5888 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_62
timestamp 1649977179
transform 1 0 6808 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_74
timestamp 1649977179
transform 1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_105
timestamp 1649977179
transform 1 0 10764 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_134
timestamp 1649977179
transform 1 0 13432 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_138
timestamp 1649977179
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_150
timestamp 1649977179
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_154
timestamp 1649977179
transform 1 0 15272 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_164
timestamp 1649977179
transform 1 0 16192 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_175
timestamp 1649977179
transform 1 0 17204 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_186
timestamp 1649977179
transform 1 0 18216 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 1649977179
transform 1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_17
timestamp 1649977179
transform 1 0 2668 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_21
timestamp 1649977179
transform 1 0 3036 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_31
timestamp 1649977179
transform 1 0 3956 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_43
timestamp 1649977179
transform 1 0 5060 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_59
timestamp 1649977179
transform 1 0 6532 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_96
timestamp 1649977179
transform 1 0 9936 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_100
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_110
timestamp 1649977179
transform 1 0 11224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1649977179
transform 1 0 11776 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_131
timestamp 1649977179
transform 1 0 13156 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_134
timestamp 1649977179
transform 1 0 13432 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_145
timestamp 1649977179
transform 1 0 14444 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_157
timestamp 1649977179
transform 1 0 15548 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 1649977179
transform 1 0 16284 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_178
timestamp 1649977179
transform 1 0 17480 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_182
timestamp 1649977179
transform 1 0 17848 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_201
timestamp 1649977179
transform 1 0 19596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_211
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_7
timestamp 1649977179
transform 1 0 1748 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_12
timestamp 1649977179
transform 1 0 2208 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_17
timestamp 1649977179
transform 1 0 2668 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_22
timestamp 1649977179
transform 1 0 3128 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_32
timestamp 1649977179
transform 1 0 4048 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_49
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_67
timestamp 1649977179
transform 1 0 7268 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1649977179
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_101
timestamp 1649977179
transform 1 0 10396 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_119
timestamp 1649977179
transform 1 0 12052 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_130
timestamp 1649977179
transform 1 0 13064 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_161
timestamp 1649977179
transform 1 0 15916 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_172
timestamp 1649977179
transform 1 0 16928 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_200
timestamp 1649977179
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1649977179
transform 1 0 20424 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_17
timestamp 1649977179
transform 1 0 2668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_21
timestamp 1649977179
transform 1 0 3036 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_32
timestamp 1649977179
transform 1 0 4048 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_43
timestamp 1649977179
transform 1 0 5060 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_47
timestamp 1649977179
transform 1 0 5428 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_59
timestamp 1649977179
transform 1 0 6532 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_71
timestamp 1649977179
transform 1 0 7636 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_77
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_80
timestamp 1649977179
transform 1 0 8464 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_91
timestamp 1649977179
transform 1 0 9476 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_95
timestamp 1649977179
transform 1 0 9844 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_107
timestamp 1649977179
transform 1 0 10948 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_117
timestamp 1649977179
transform 1 0 11868 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_126
timestamp 1649977179
transform 1 0 12696 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1649977179
transform 1 0 13156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_135
timestamp 1649977179
transform 1 0 13524 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1649977179
transform 1 0 14536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_157
timestamp 1649977179
transform 1 0 15548 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_162
timestamp 1649977179
transform 1 0 16008 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_177
timestamp 1649977179
transform 1 0 17388 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_187
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_197
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 1649977179
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1649977179
transform 1 0 20424 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_12
timestamp 1649977179
transform 1 0 2208 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_17
timestamp 1649977179
transform 1 0 2668 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_22
timestamp 1649977179
transform 1 0 3128 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_31
timestamp 1649977179
transform 1 0 3956 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_35
timestamp 1649977179
transform 1 0 4324 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_39
timestamp 1649977179
transform 1 0 4692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_43
timestamp 1649977179
transform 1 0 5060 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_60
timestamp 1649977179
transform 1 0 6624 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_94
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_106
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_118
timestamp 1649977179
transform 1 0 11960 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_130
timestamp 1649977179
transform 1 0 13064 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1649977179
transform 1 0 13800 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_145
timestamp 1649977179
transform 1 0 14444 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_162
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_30_172
timestamp 1649977179
transform 1 0 16928 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_178
timestamp 1649977179
transform 1 0 17480 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_181
timestamp 1649977179
transform 1 0 17756 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_185
timestamp 1649977179
transform 1 0 18124 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_194
timestamp 1649977179
transform 1 0 18952 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_200
timestamp 1649977179
transform 1 0 19504 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 1649977179
transform 1 0 2760 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_23
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_44
timestamp 1649977179
transform 1 0 5152 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_48
timestamp 1649977179
transform 1 0 5520 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_91
timestamp 1649977179
transform 1 0 9476 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_96
timestamp 1649977179
transform 1 0 9936 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1649977179
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_121
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_140
timestamp 1649977179
transform 1 0 13984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_158
timestamp 1649977179
transform 1 0 15640 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_166
timestamp 1649977179
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_187
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_190
timestamp 1649977179
transform 1 0 18584 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_194
timestamp 1649977179
transform 1 0 18952 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_199
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_204
timestamp 1649977179
transform 1 0 19872 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1649977179
transform 1 0 20332 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_7
timestamp 1649977179
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_19
timestamp 1649977179
transform 1 0 2852 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1649977179
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_45
timestamp 1649977179
transform 1 0 5244 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_55
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_59
timestamp 1649977179
transform 1 0 6532 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_67
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1649977179
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_101
timestamp 1649977179
transform 1 0 10396 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_125
timestamp 1649977179
transform 1 0 12604 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_137
timestamp 1649977179
transform 1 0 13708 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1649977179
transform 1 0 1748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_13
timestamp 1649977179
transform 1 0 2300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_19
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_24
timestamp 1649977179
transform 1 0 3312 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_32
timestamp 1649977179
transform 1 0 4048 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_37
timestamp 1649977179
transform 1 0 4508 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_42
timestamp 1649977179
transform 1 0 4968 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_46
timestamp 1649977179
transform 1 0 5336 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_50
timestamp 1649977179
transform 1 0 5704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_63
timestamp 1649977179
transform 1 0 6900 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_75
timestamp 1649977179
transform 1 0 8004 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp 1649977179
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_180
timestamp 1649977179
transform 1 0 17664 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_186
timestamp 1649977179
transform 1 0 18216 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_189
timestamp 1649977179
transform 1 0 18492 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _056_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1649977179
transform -1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1649977179
transform 1 0 1932 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1649977179
transform 1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1649977179
transform 1 0 2392 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1649977179
transform 1 0 2392 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1649977179
transform 1 0 2392 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1649977179
transform 1 0 1932 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1649977179
transform 1 0 1932 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1649977179
transform 1 0 2392 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 1932 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 2392 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 3036 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 2944 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 20884 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform -1 0 20884 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform -1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform -1 0 20424 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 20424 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform -1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform -1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform -1 0 20424 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform -1 0 19872 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform -1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform -1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform -1 0 18492 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform -1 0 12236 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 12696 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform -1 0 13156 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 13432 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 13616 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 10856 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 13340 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform -1 0 12880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 14444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1649977179
transform -1 0 13800 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1649977179
transform -1 0 14720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1649977179
transform -1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 13340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1649977179
transform -1 0 13800 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1649977179
transform -1 0 16376 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13616 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 9660 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 7820 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 14812 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20608 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 16192 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 11684 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform -1 0 12052 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 7912 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 3864 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 14168 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform 1 0 6072 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform -1 0 19228 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 20516 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 11960 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform 1 0 20608 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform 1 0 5428 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform 1 0 19044 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform 1 0 7728 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform 1 0 13064 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform -1 0 19228 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform 1 0 9660 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform 1 0 5152 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform 1 0 8740 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 17480 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 6532 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 6164 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform -1 0 4692 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 4416 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1649977179
transform 1 0 1564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 3128 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1649977179
transform 1 0 1472 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1649977179
transform 1 0 1564 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1649977179
transform 1 0 1564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 3588 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1649977179
transform 1 0 1564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1649977179
transform 1 0 1472 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1649977179
transform 1 0 1564 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform 1 0 7268 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1649977179
transform 1 0 1564 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input26
timestamp 1649977179
transform 1 0 1472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1649977179
transform 1 0 1564 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform -1 0 2300 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 14996 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1649977179
transform -1 0 18952 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 15272 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1649977179
transform -1 0 18768 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1649977179
transform -1 0 21436 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1649977179
transform -1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input38
timestamp 1649977179
transform -1 0 21436 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input39
timestamp 1649977179
transform -1 0 20424 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1649977179
transform -1 0 21436 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 18952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 15456 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 20332 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 15916 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1649977179
transform -1 0 19228 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1649977179
transform -1 0 18400 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input47
timestamp 1649977179
transform -1 0 19780 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 18400 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform -1 0 18952 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 3496 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 10120 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform 1 0 8372 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1649977179
transform 1 0 10304 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform 1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 12696 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 5336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform -1 0 6624 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform -1 0 5060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform -1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input66
timestamp 1649977179
transform -1 0 7268 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform -1 0 8096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 6624 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1649977179
transform -1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input71
timestamp 1649977179
transform -1 0 3404 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform -1 0 7728 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input73
timestamp 1649977179
transform -1 0 2300 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1649977179
transform 1 0 8280 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input75
timestamp 1649977179
transform -1 0 5796 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1649977179
transform -1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform -1 0 4968 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1649977179
transform -1 0 20056 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input82
timestamp 1649977179
transform -1 0 13432 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1649977179
transform 1 0 20516 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1649977179
transform -1 0 21436 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform -1 0 16100 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input87
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21252 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7912 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7820 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 3036 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 2944 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 2024 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 4600 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8004 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11684 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 14536 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_11.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 12696 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9568 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10304 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12328 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14904 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14904 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16744 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17664 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 21436 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20884 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 10396 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3404 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 2024 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 3956 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 5244 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8556 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 5244 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4232 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 3496 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 4048 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4416 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7268 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 5244 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 3680 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7360 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 6532 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7912 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9108 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 11040 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7176 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14168 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 14536 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 17940 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10672 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 12328 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 17480 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19596 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform 1 0 10580 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11408 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11960 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 13616 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15916 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 15548 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14352 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 18952 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10580 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 8004 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l1_in_3__172 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 6808 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8648 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 9844 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7176 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 6348 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_2_
timestamp 1649977179
transform -1 0 4968 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l1_in_3_
timestamp 1649977179
transform 1 0 5152 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_3.mux_l1_in_3__182
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4600 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_3.mux_l3_in_0_
timestamp 1649977179
transform -1 0 4416 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 5704 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l1_in_3__155
timestamp 1649977179
transform 1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_3_
timestamp 1649977179
transform -1 0 2300 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform -1 0 2484 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 2944 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l3_in_0_
timestamp 1649977179
transform -1 0 3496 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6440 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_1_
timestamp 1649977179
transform 1 0 6440 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_2_
timestamp 1649977179
transform -1 0 6072 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_7.mux_l1_in_3__156
timestamp 1649977179
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l1_in_3_
timestamp 1649977179
transform -1 0 5060 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7176 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6072 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_7.mux_l3_in_0_
timestamp 1649977179
transform -1 0 7636 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12420 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10580 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_1__157
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_1_
timestamp 1649977179
transform -1 0 9844 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l3_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13156 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_11.mux_l2_in_1__173
timestamp 1649977179
transform -1 0 11960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_11.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12972 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12604 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_13.mux_l1_in_1__174
timestamp 1649977179
transform -1 0 11316 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_13.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11868 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13892 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_15.mux_l1_in_1__175
timestamp 1649977179
transform -1 0 14352 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15456 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15640 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_17.mux_l1_in_1__176
timestamp 1649977179
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 11960 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_19.mux_l1_in_1__177
timestamp 1649977179
transform -1 0 16376 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_19.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10396 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_21.mux_l1_in_1__178
timestamp 1649977179
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 14720 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17756 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_23.mux_l1_in_1__179
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 15180 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20608 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform -1 0 19780 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_1__180
timestamp 1649977179
transform -1 0 19780 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19964 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 19320 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 17204 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_27.mux_l2_in_0__181
timestamp 1649977179
transform -1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19412 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15640 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9016 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7820 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_2_
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_3__158
timestamp 1649977179
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_3_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_1_
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l4_in_0_
timestamp 1649977179
transform -1 0 3128 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 4968 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7636 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7728 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7452 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_2_
timestamp 1649977179
transform 1 0 6440 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_3__161
timestamp 1649977179
transform -1 0 6992 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_3_
timestamp 1649977179
transform 1 0 6716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5428 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_1_
timestamp 1649977179
transform 1 0 5888 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4784 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2116 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4140 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 4232 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 4692 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_3_
timestamp 1649977179
transform 1 0 5704 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_4_
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_5_
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_6_
timestamp 1649977179
transform -1 0 2944 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform -1 0 3956 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3128 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_3__163
timestamp 1649977179
transform -1 0 2208 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3128 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_1_
timestamp 1649977179
transform -1 0 3220 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l4_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5060 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6900 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_2_
timestamp 1649977179
transform -1 0 3956 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l2_in_3__164
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_3_
timestamp 1649977179
transform -1 0 3496 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_0_
timestamp 1649977179
transform 1 0 4416 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l3_in_1_
timestamp 1649977179
transform -1 0 4048 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l4_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_1_
timestamp 1649977179
transform 1 0 7360 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_2_
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l1_in_3__159
timestamp 1649977179
transform 1 0 8280 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_3_
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6072 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2668 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 9568 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 10028 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_3__160
timestamp 1649977179
transform -1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_3_
timestamp 1649977179
transform -1 0 9844 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9200 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_1_
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l3_in_0_
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 7820 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9476 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9108 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_2_
timestamp 1649977179
transform -1 0 7912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_1__162
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_1_
timestamp 1649977179
transform 1 0 7728 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7544 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3036 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16376 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 14444 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16100 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_2_
timestamp 1649977179
transform -1 0 14904 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_3__165
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_3_
timestamp 1649977179
transform -1 0 14536 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 14720 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 15088 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l4_in_0_
timestamp 1649977179
transform -1 0 15548 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18124 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17664 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 10856 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_2_
timestamp 1649977179
transform -1 0 12420 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_3__167
timestamp 1649977179
transform -1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_3_
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 15088 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_1_
timestamp 1649977179
transform -1 0 12788 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l4_in_0_
timestamp 1649977179
transform -1 0 13800 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19228 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20056 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19412 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 19412 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_3_
timestamp 1649977179
transform 1 0 20424 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_4_
timestamp 1649977179
transform -1 0 17480 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_5_
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_6_
timestamp 1649977179
transform 1 0 19504 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19044 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_2_
timestamp 1649977179
transform -1 0 18492 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_3__170
timestamp 1649977179
transform -1 0 19504 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_3_
timestamp 1649977179
transform 1 0 19320 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18952 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_1_
timestamp 1649977179
transform -1 0 18860 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l4_in_0_
timestamp 1649977179
transform -1 0 19136 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17480 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_1_
timestamp 1649977179
transform -1 0 8740 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_2_
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l2_in_3__171
timestamp 1649977179
transform 1 0 12880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_3_
timestamp 1649977179
transform 1 0 11960 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_0_
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l3_in_1_
timestamp 1649977179
transform -1 0 11224 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l4_in_0_
timestamp 1649977179
transform -1 0 12144 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_1_
timestamp 1649977179
transform -1 0 12328 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12236 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_3_
timestamp 1649977179
transform 1 0 14168 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l1_in_3__166
timestamp 1649977179
transform 1 0 15088 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16100 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16744 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8740 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_2_
timestamp 1649977179
transform -1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_3__168
timestamp 1649977179
transform -1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_3_
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15180 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_1_
timestamp 1649977179
transform -1 0 16928 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18768 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_1__169
timestamp 1649977179
transform -1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_1_
timestamp 1649977179
transform 1 0 20424 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20240 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20056 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output89 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 1748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 2852 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 2852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform -1 0 2300 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform -1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform -1 0 1748 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 1932 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform -1 0 1748 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform -1 0 1748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 12880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 18308 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 19136 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 18584 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 17480 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 14628 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output150
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  repeater151
timestamp 1649977179
transform 1 0 20240 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater152
timestamp 1649977179
transform -1 0 16376 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  repeater153
timestamp 1649977179
transform -1 0 3772 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  repeater154
timestamp 1649977179
transform -1 0 6072 0 -1 13056
box -38 -48 958 592
<< labels >>
rlabel metal2 s 21822 0 21878 800 6 SC_IN_BOT
port 0 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 3 nsew power input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_42_
port 4 nsew signal input
rlabel metal2 s 570 0 626 800 6 bottom_left_grid_pin_43_
port 5 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 bottom_left_grid_pin_44_
port 6 nsew signal input
rlabel metal2 s 1490 0 1546 800 6 bottom_left_grid_pin_45_
port 7 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 bottom_left_grid_pin_46_
port 8 nsew signal input
rlabel metal2 s 2410 0 2466 800 6 bottom_left_grid_pin_47_
port 9 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 bottom_left_grid_pin_48_
port 10 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 bottom_left_grid_pin_49_
port 11 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 ccff_head
port 12 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_tail
port 13 nsew signal tristate
rlabel metal3 s 0 3816 800 3936 6 chanx_left_in[0]
port 14 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[10]
port 15 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[11]
port 16 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[12]
port 17 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[13]
port 18 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[14]
port 19 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[15]
port 20 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[16]
port 21 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[17]
port 22 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[18]
port 23 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[19]
port 24 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[1]
port 25 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[2]
port 26 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[3]
port 27 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[4]
port 28 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[5]
port 29 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[6]
port 30 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[7]
port 31 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[8]
port 32 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[9]
port 33 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_out[0]
port 34 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[10]
port 35 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[11]
port 36 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[12]
port 37 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[13]
port 38 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[14]
port 39 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[15]
port 40 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[16]
port 41 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[17]
port 42 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[18]
port 43 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[19]
port 44 nsew signal tristate
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[1]
port 45 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[2]
port 46 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[3]
port 47 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[4]
port 48 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[5]
port 49 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[6]
port 50 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[7]
port 51 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[8]
port 52 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[9]
port 53 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 54 nsew signal input
rlabel metal3 s 22200 8576 23000 8696 6 chanx_right_in[10]
port 55 nsew signal input
rlabel metal3 s 22200 8984 23000 9104 6 chanx_right_in[11]
port 56 nsew signal input
rlabel metal3 s 22200 9392 23000 9512 6 chanx_right_in[12]
port 57 nsew signal input
rlabel metal3 s 22200 9936 23000 10056 6 chanx_right_in[13]
port 58 nsew signal input
rlabel metal3 s 22200 10344 23000 10464 6 chanx_right_in[14]
port 59 nsew signal input
rlabel metal3 s 22200 10888 23000 11008 6 chanx_right_in[15]
port 60 nsew signal input
rlabel metal3 s 22200 11296 23000 11416 6 chanx_right_in[16]
port 61 nsew signal input
rlabel metal3 s 22200 11840 23000 11960 6 chanx_right_in[17]
port 62 nsew signal input
rlabel metal3 s 22200 12248 23000 12368 6 chanx_right_in[18]
port 63 nsew signal input
rlabel metal3 s 22200 12792 23000 12912 6 chanx_right_in[19]
port 64 nsew signal input
rlabel metal3 s 22200 4360 23000 4480 6 chanx_right_in[1]
port 65 nsew signal input
rlabel metal3 s 22200 4768 23000 4888 6 chanx_right_in[2]
port 66 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 67 nsew signal input
rlabel metal3 s 22200 5720 23000 5840 6 chanx_right_in[4]
port 68 nsew signal input
rlabel metal3 s 22200 6128 23000 6248 6 chanx_right_in[5]
port 69 nsew signal input
rlabel metal3 s 22200 6672 23000 6792 6 chanx_right_in[6]
port 70 nsew signal input
rlabel metal3 s 22200 7080 23000 7200 6 chanx_right_in[7]
port 71 nsew signal input
rlabel metal3 s 22200 7624 23000 7744 6 chanx_right_in[8]
port 72 nsew signal input
rlabel metal3 s 22200 8032 23000 8152 6 chanx_right_in[9]
port 73 nsew signal input
rlabel metal3 s 22200 13200 23000 13320 6 chanx_right_out[0]
port 74 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[10]
port 75 nsew signal tristate
rlabel metal3 s 22200 18368 23000 18488 6 chanx_right_out[11]
port 76 nsew signal tristate
rlabel metal3 s 22200 18776 23000 18896 6 chanx_right_out[12]
port 77 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[13]
port 78 nsew signal tristate
rlabel metal3 s 22200 19728 23000 19848 6 chanx_right_out[14]
port 79 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[15]
port 80 nsew signal tristate
rlabel metal3 s 22200 20680 23000 20800 6 chanx_right_out[16]
port 81 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[17]
port 82 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[18]
port 83 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 chanx_right_out[19]
port 84 nsew signal tristate
rlabel metal3 s 22200 13744 23000 13864 6 chanx_right_out[1]
port 85 nsew signal tristate
rlabel metal3 s 22200 14152 23000 14272 6 chanx_right_out[2]
port 86 nsew signal tristate
rlabel metal3 s 22200 14560 23000 14680 6 chanx_right_out[3]
port 87 nsew signal tristate
rlabel metal3 s 22200 15104 23000 15224 6 chanx_right_out[4]
port 88 nsew signal tristate
rlabel metal3 s 22200 15512 23000 15632 6 chanx_right_out[5]
port 89 nsew signal tristate
rlabel metal3 s 22200 16056 23000 16176 6 chanx_right_out[6]
port 90 nsew signal tristate
rlabel metal3 s 22200 16464 23000 16584 6 chanx_right_out[7]
port 91 nsew signal tristate
rlabel metal3 s 22200 17008 23000 17128 6 chanx_right_out[8]
port 92 nsew signal tristate
rlabel metal3 s 22200 17416 23000 17536 6 chanx_right_out[9]
port 93 nsew signal tristate
rlabel metal2 s 3790 0 3846 800 6 chany_bottom_in[0]
port 94 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_in[10]
port 95 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[11]
port 96 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[12]
port 97 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[13]
port 98 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[14]
port 99 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[15]
port 100 nsew signal input
rlabel metal2 s 10966 0 11022 800 6 chany_bottom_in[16]
port 101 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 chany_bottom_in[17]
port 102 nsew signal input
rlabel metal2 s 11886 0 11942 800 6 chany_bottom_in[18]
port 103 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 chany_bottom_in[19]
port 104 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 chany_bottom_in[1]
port 105 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 chany_bottom_in[2]
port 106 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[3]
port 107 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 chany_bottom_in[4]
port 108 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 chany_bottom_in[5]
port 109 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 chany_bottom_in[6]
port 110 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 chany_bottom_in[7]
port 111 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 chany_bottom_in[8]
port 112 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[9]
port 113 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 chany_bottom_out[0]
port 114 nsew signal tristate
rlabel metal2 s 17314 0 17370 800 6 chany_bottom_out[10]
port 115 nsew signal tristate
rlabel metal2 s 17774 0 17830 800 6 chany_bottom_out[11]
port 116 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 117 nsew signal tristate
rlabel metal2 s 18602 0 18658 800 6 chany_bottom_out[13]
port 118 nsew signal tristate
rlabel metal2 s 19062 0 19118 800 6 chany_bottom_out[14]
port 119 nsew signal tristate
rlabel metal2 s 19522 0 19578 800 6 chany_bottom_out[15]
port 120 nsew signal tristate
rlabel metal2 s 19982 0 20038 800 6 chany_bottom_out[16]
port 121 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[17]
port 122 nsew signal tristate
rlabel metal2 s 20902 0 20958 800 6 chany_bottom_out[18]
port 123 nsew signal tristate
rlabel metal2 s 21362 0 21418 800 6 chany_bottom_out[19]
port 124 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[1]
port 125 nsew signal tristate
rlabel metal2 s 13726 0 13782 800 6 chany_bottom_out[2]
port 126 nsew signal tristate
rlabel metal2 s 14094 0 14150 800 6 chany_bottom_out[3]
port 127 nsew signal tristate
rlabel metal2 s 14554 0 14610 800 6 chany_bottom_out[4]
port 128 nsew signal tristate
rlabel metal2 s 15014 0 15070 800 6 chany_bottom_out[5]
port 129 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[6]
port 130 nsew signal tristate
rlabel metal2 s 15934 0 15990 800 6 chany_bottom_out[7]
port 131 nsew signal tristate
rlabel metal2 s 16394 0 16450 800 6 chany_bottom_out[8]
port 132 nsew signal tristate
rlabel metal2 s 16854 0 16910 800 6 chany_bottom_out[9]
port 133 nsew signal tristate
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_34_
port 134 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_35_
port 135 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_36_
port 136 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_37_
port 137 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_38_
port 138 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_39_
port 139 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_40_
port 140 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_41_
port 141 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 left_top_grid_pin_1_
port 142 nsew signal input
rlabel metal2 s 22742 0 22798 800 6 prog_clk_0_S_in
port 143 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 144 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 145 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 146 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 147 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 148 nsew signal input
rlabel metal3 s 22200 2456 23000 2576 6 right_bottom_grid_pin_39_
port 149 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 150 nsew signal input
rlabel metal3 s 22200 3408 23000 3528 6 right_bottom_grid_pin_41_
port 151 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 152 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
