magic
tech sky130A
magscale 1 2
timestamp 1650634230
<< viali >>
rect 1593 17289 1627 17323
rect 1961 17289 1995 17323
rect 2329 17289 2363 17323
rect 2697 17289 2731 17323
rect 3065 17289 3099 17323
rect 3433 17289 3467 17323
rect 4169 17289 4203 17323
rect 4537 17289 4571 17323
rect 4905 17289 4939 17323
rect 5273 17289 5307 17323
rect 5641 17289 5675 17323
rect 6009 17289 6043 17323
rect 6653 17289 6687 17323
rect 7021 17289 7055 17323
rect 7481 17289 7515 17323
rect 7941 17289 7975 17323
rect 8309 17289 8343 17323
rect 9045 17289 9079 17323
rect 9413 17289 9447 17323
rect 10609 17289 10643 17323
rect 13277 17289 13311 17323
rect 14381 17289 14415 17323
rect 14565 17289 14599 17323
rect 15577 17289 15611 17323
rect 12265 17221 12299 17255
rect 13093 17221 13127 17255
rect 15209 17221 15243 17255
rect 1777 17153 1811 17187
rect 2145 17153 2179 17187
rect 2513 17153 2547 17187
rect 2881 17153 2915 17187
rect 3249 17153 3283 17187
rect 3617 17153 3651 17187
rect 4353 17153 4387 17187
rect 4721 17153 4755 17187
rect 5089 17153 5123 17187
rect 5457 17153 5491 17187
rect 5825 17153 5859 17187
rect 6193 17153 6227 17187
rect 6837 17153 6871 17187
rect 7205 17153 7239 17187
rect 7665 17153 7699 17187
rect 8125 17153 8159 17187
rect 8493 17153 8527 17187
rect 8769 17153 8803 17187
rect 9229 17153 9263 17187
rect 9689 17153 9723 17187
rect 9873 17153 9907 17187
rect 10149 17153 10183 17187
rect 10517 17153 10551 17187
rect 10977 17153 11011 17187
rect 11345 17153 11379 17187
rect 11805 17153 11839 17187
rect 12173 17153 12207 17187
rect 12633 17153 12667 17187
rect 13001 17153 13035 17187
rect 13461 17153 13495 17187
rect 13829 17153 13863 17187
rect 14289 17153 14323 17187
rect 14749 17153 14783 17187
rect 15117 17153 15151 17187
rect 15393 17153 15427 17187
rect 10333 17017 10367 17051
rect 14933 17017 14967 17051
rect 8585 16949 8619 16983
rect 9505 16949 9539 16983
rect 10057 16949 10091 16983
rect 10793 16949 10827 16983
rect 11161 16949 11195 16983
rect 11621 16949 11655 16983
rect 11989 16949 12023 16983
rect 12449 16949 12483 16983
rect 12817 16949 12851 16983
rect 13645 16949 13679 16983
rect 14105 16949 14139 16983
rect 8953 16745 8987 16779
rect 10701 16745 10735 16779
rect 11069 16745 11103 16779
rect 11897 16745 11931 16779
rect 12725 16745 12759 16779
rect 13185 16745 13219 16779
rect 13461 16745 13495 16779
rect 14381 16745 14415 16779
rect 2329 16677 2363 16711
rect 14565 16677 14599 16711
rect 2421 16609 2455 16643
rect 14749 16609 14783 16643
rect 1685 16541 1719 16575
rect 2053 16541 2087 16575
rect 2145 16541 2179 16575
rect 15025 16541 15059 16575
rect 15301 16541 15335 16575
rect 15577 16541 15611 16575
rect 1501 16405 1535 16439
rect 1869 16405 1903 16439
rect 14841 16405 14875 16439
rect 15117 16405 15151 16439
rect 15393 16405 15427 16439
rect 15117 16133 15151 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 15393 16065 15427 16099
rect 15669 16065 15703 16099
rect 14933 15997 14967 16031
rect 1593 15929 1627 15963
rect 15209 15861 15243 15895
rect 15485 15861 15519 15895
rect 15485 15657 15519 15691
rect 4629 13889 4663 13923
rect 4169 13821 4203 13855
rect 4537 13685 4571 13719
rect 4169 13277 4203 13311
rect 4425 13277 4459 13311
rect 5549 13141 5583 13175
rect 4077 12937 4111 12971
rect 5273 12937 5307 12971
rect 7205 12937 7239 12971
rect 9413 12937 9447 12971
rect 14381 12937 14415 12971
rect 4261 12801 4295 12835
rect 4813 12801 4847 12835
rect 5457 12801 5491 12835
rect 7389 12801 7423 12835
rect 9597 12801 9631 12835
rect 14197 12801 14231 12835
rect 15393 12801 15427 12835
rect 4629 12665 4663 12699
rect 14013 12597 14047 12631
rect 15577 12597 15611 12631
rect 7941 11849 7975 11883
rect 1409 11713 1443 11747
rect 1685 11713 1719 11747
rect 7481 11713 7515 11747
rect 8125 11713 8159 11747
rect 7573 11645 7607 11679
rect 7665 11645 7699 11679
rect 1593 11509 1627 11543
rect 7113 11509 7147 11543
rect 8953 11237 8987 11271
rect 9505 11169 9539 11203
rect 9321 11101 9355 11135
rect 9781 11101 9815 11135
rect 6285 11033 6319 11067
rect 8033 11033 8067 11067
rect 9413 10965 9447 10999
rect 3065 10761 3099 10795
rect 7021 10761 7055 10795
rect 9137 10761 9171 10795
rect 9505 10761 9539 10795
rect 9965 10761 9999 10795
rect 10425 10761 10459 10795
rect 4353 10693 4387 10727
rect 5641 10625 5675 10659
rect 5917 10625 5951 10659
rect 6193 10625 6227 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 7645 10625 7679 10659
rect 10333 10625 10367 10659
rect 7389 10557 7423 10591
rect 9597 10557 9631 10591
rect 9689 10557 9723 10591
rect 10517 10557 10551 10591
rect 6561 10489 6595 10523
rect 5457 10421 5491 10455
rect 5733 10421 5767 10455
rect 6009 10421 6043 10455
rect 8769 10421 8803 10455
rect 10333 10217 10367 10251
rect 10885 10217 10919 10251
rect 13093 10217 13127 10251
rect 13369 10217 13403 10251
rect 13645 10217 13679 10251
rect 3387 10149 3421 10183
rect 8953 10149 8987 10183
rect 10609 10149 10643 10183
rect 12265 10149 12299 10183
rect 12541 10149 12575 10183
rect 5549 10081 5583 10115
rect 5733 10081 5767 10115
rect 5917 10081 5951 10115
rect 6101 10081 6135 10115
rect 7573 10081 7607 10115
rect 8125 10081 8159 10115
rect 9781 10081 9815 10115
rect 3316 10013 3350 10047
rect 4721 10013 4755 10047
rect 4997 10013 5031 10047
rect 8401 10013 8435 10047
rect 9137 10013 9171 10047
rect 9689 10013 9723 10047
rect 10241 10013 10275 10047
rect 10517 10013 10551 10047
rect 10793 10013 10827 10047
rect 11069 10013 11103 10047
rect 11345 10013 11379 10047
rect 11621 10013 11655 10047
rect 11897 10013 11931 10047
rect 12173 10013 12207 10047
rect 12449 10013 12483 10047
rect 12725 10013 12759 10047
rect 13001 10013 13035 10047
rect 13277 10013 13311 10047
rect 13553 10013 13587 10047
rect 13829 10013 13863 10047
rect 5457 9945 5491 9979
rect 4537 9877 4571 9911
rect 4813 9877 4847 9911
rect 5089 9877 5123 9911
rect 8309 9877 8343 9911
rect 8769 9877 8803 9911
rect 9229 9877 9263 9911
rect 9597 9877 9631 9911
rect 10057 9877 10091 9911
rect 11161 9877 11195 9911
rect 11437 9877 11471 9911
rect 11713 9877 11747 9911
rect 11989 9877 12023 9911
rect 12817 9877 12851 9911
rect 9321 9673 9355 9707
rect 3065 9605 3099 9639
rect 8953 9605 8987 9639
rect 5825 9537 5859 9571
rect 6193 9537 6227 9571
rect 6745 9537 6779 9571
rect 7961 9537 7995 9571
rect 9597 9537 9631 9571
rect 9873 9537 9907 9571
rect 2789 9469 2823 9503
rect 3249 9469 3283 9503
rect 8217 9469 8251 9503
rect 8677 9469 8711 9503
rect 8861 9469 8895 9503
rect 6009 9401 6043 9435
rect 5641 9333 5675 9367
rect 6561 9333 6595 9367
rect 6837 9333 6871 9367
rect 9413 9333 9447 9367
rect 9689 9333 9723 9367
rect 6101 9129 6135 9163
rect 7021 9129 7055 9163
rect 8953 9129 8987 9163
rect 8493 9061 8527 9095
rect 9413 8993 9447 9027
rect 9505 8993 9539 9027
rect 6285 8925 6319 8959
rect 6377 8925 6411 8959
rect 7113 8925 7147 8959
rect 8769 8925 8803 8959
rect 7380 8857 7414 8891
rect 8585 8789 8619 8823
rect 9321 8789 9355 8823
rect 6745 8585 6779 8619
rect 7858 8517 7892 8551
rect 11805 8517 11839 8551
rect 1685 8449 1719 8483
rect 8125 8449 8159 8483
rect 12633 8449 12667 8483
rect 1501 8313 1535 8347
rect 12817 8313 12851 8347
rect 7205 8041 7239 8075
rect 7021 7905 7055 7939
rect 7849 7905 7883 7939
rect 5273 7837 5307 7871
rect 7665 7837 7699 7871
rect 7573 7769 7607 7803
rect 4169 7361 4203 7395
rect 4721 7361 4755 7395
rect 5273 7361 5307 7395
rect 7297 7361 7331 7395
rect 9413 7361 9447 7395
rect 5089 7225 5123 7259
rect 3985 7157 4019 7191
rect 4537 7157 4571 7191
rect 7113 7157 7147 7191
rect 9229 7157 9263 7191
rect 3157 6749 3191 6783
rect 2973 6613 3007 6647
rect 1685 5185 1719 5219
rect 1501 4981 1535 5015
rect 15485 3689 15519 3723
rect 1685 3485 1719 3519
rect 15117 3485 15151 3519
rect 15669 3485 15703 3519
rect 14933 3417 14967 3451
rect 1501 3349 1535 3383
rect 15301 3349 15335 3383
rect 2329 3145 2363 3179
rect 14933 3145 14967 3179
rect 15209 3145 15243 3179
rect 1685 3009 1719 3043
rect 2053 3009 2087 3043
rect 2145 3009 2179 3043
rect 2421 3009 2455 3043
rect 14565 3009 14599 3043
rect 15117 3009 15151 3043
rect 15393 3009 15427 3043
rect 15669 3009 15703 3043
rect 1869 2873 1903 2907
rect 1501 2805 1535 2839
rect 8769 2805 8803 2839
rect 9229 2805 9263 2839
rect 10885 2805 10919 2839
rect 11529 2805 11563 2839
rect 12173 2805 12207 2839
rect 13461 2805 13495 2839
rect 13921 2805 13955 2839
rect 14749 2805 14783 2839
rect 15485 2805 15519 2839
rect 8953 2601 8987 2635
rect 9873 2601 9907 2635
rect 12725 2601 12759 2635
rect 14841 2601 14875 2635
rect 10149 2533 10183 2567
rect 13185 2533 13219 2567
rect 13553 2533 13587 2567
rect 12633 2465 12667 2499
rect 1869 2397 1903 2431
rect 2237 2397 2271 2431
rect 2697 2397 2731 2431
rect 3157 2397 3191 2431
rect 3525 2397 3559 2431
rect 4077 2397 4111 2431
rect 4445 2397 4479 2431
rect 4813 2397 4847 2431
rect 5266 2397 5300 2431
rect 5733 2397 5767 2431
rect 6101 2397 6135 2431
rect 6653 2397 6687 2431
rect 7021 2397 7055 2431
rect 7389 2397 7423 2431
rect 7849 2397 7883 2431
rect 8309 2397 8343 2431
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 9505 2397 9539 2431
rect 9689 2397 9723 2431
rect 9965 2397 9999 2431
rect 10333 2397 10367 2431
rect 10793 2397 10827 2431
rect 11161 2397 11195 2431
rect 11713 2397 11747 2431
rect 12081 2397 12115 2431
rect 12449 2397 12483 2431
rect 12909 2397 12943 2431
rect 13369 2397 13403 2431
rect 13737 2397 13771 2431
rect 14289 2397 14323 2431
rect 14657 2397 14691 2431
rect 15025 2397 15059 2431
rect 15485 2397 15519 2431
rect 10425 2329 10459 2363
rect 11253 2329 11287 2363
rect 13001 2329 13035 2363
rect 13829 2329 13863 2363
rect 15117 2329 15151 2363
rect 1685 2261 1719 2295
rect 2053 2261 2087 2295
rect 2513 2261 2547 2295
rect 2973 2261 3007 2295
rect 3341 2261 3375 2295
rect 3893 2261 3927 2295
rect 4261 2261 4295 2295
rect 4629 2261 4663 2295
rect 5089 2261 5123 2295
rect 5549 2261 5583 2295
rect 5917 2261 5951 2295
rect 6469 2261 6503 2295
rect 6837 2261 6871 2295
rect 7205 2261 7239 2295
rect 7665 2261 7699 2295
rect 8125 2261 8159 2295
rect 8493 2261 8527 2295
rect 9321 2261 9355 2295
rect 10609 2261 10643 2295
rect 10977 2261 11011 2295
rect 11529 2261 11563 2295
rect 11897 2261 11931 2295
rect 12265 2261 12299 2295
rect 14105 2261 14139 2295
rect 14473 2261 14507 2295
rect 15301 2261 15335 2295
rect 15669 2261 15703 2295
<< metal1 >>
rect 6178 17620 6184 17672
rect 6236 17660 6242 17672
rect 10870 17660 10876 17672
rect 6236 17632 10876 17660
rect 6236 17620 6242 17632
rect 10870 17620 10876 17632
rect 10928 17620 10934 17672
rect 9306 17552 9312 17604
rect 9364 17592 9370 17604
rect 13078 17592 13084 17604
rect 9364 17564 13084 17592
rect 9364 17552 9370 17564
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 9214 17484 9220 17536
rect 9272 17524 9278 17536
rect 13630 17524 13636 17536
rect 9272 17496 13636 17524
rect 9272 17484 9278 17496
rect 13630 17484 13636 17496
rect 13688 17484 13694 17536
rect 1104 17434 16008 17456
rect 1104 17382 4698 17434
rect 4750 17382 4762 17434
rect 4814 17382 4826 17434
rect 4878 17382 4890 17434
rect 4942 17382 4954 17434
rect 5006 17382 8446 17434
rect 8498 17382 8510 17434
rect 8562 17382 8574 17434
rect 8626 17382 8638 17434
rect 8690 17382 8702 17434
rect 8754 17382 12194 17434
rect 12246 17382 12258 17434
rect 12310 17382 12322 17434
rect 12374 17382 12386 17434
rect 12438 17382 12450 17434
rect 12502 17382 16008 17434
rect 1104 17360 16008 17382
rect 1394 17280 1400 17332
rect 1452 17320 1458 17332
rect 1581 17323 1639 17329
rect 1581 17320 1593 17323
rect 1452 17292 1593 17320
rect 1452 17280 1458 17292
rect 1581 17289 1593 17292
rect 1627 17289 1639 17323
rect 1581 17283 1639 17289
rect 1854 17280 1860 17332
rect 1912 17320 1918 17332
rect 1949 17323 2007 17329
rect 1949 17320 1961 17323
rect 1912 17292 1961 17320
rect 1912 17280 1918 17292
rect 1949 17289 1961 17292
rect 1995 17289 2007 17323
rect 1949 17283 2007 17289
rect 2222 17280 2228 17332
rect 2280 17320 2286 17332
rect 2317 17323 2375 17329
rect 2317 17320 2329 17323
rect 2280 17292 2329 17320
rect 2280 17280 2286 17292
rect 2317 17289 2329 17292
rect 2363 17289 2375 17323
rect 2682 17320 2688 17332
rect 2643 17292 2688 17320
rect 2317 17283 2375 17289
rect 2682 17280 2688 17292
rect 2740 17280 2746 17332
rect 3050 17320 3056 17332
rect 3011 17292 3056 17320
rect 3050 17280 3056 17292
rect 3108 17280 3114 17332
rect 3421 17323 3479 17329
rect 3421 17289 3433 17323
rect 3467 17320 3479 17323
rect 3510 17320 3516 17332
rect 3467 17292 3516 17320
rect 3467 17289 3479 17292
rect 3421 17283 3479 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 4154 17320 4160 17332
rect 4115 17292 4160 17320
rect 4154 17280 4160 17292
rect 4212 17280 4218 17332
rect 4338 17280 4344 17332
rect 4396 17320 4402 17332
rect 4525 17323 4583 17329
rect 4525 17320 4537 17323
rect 4396 17292 4537 17320
rect 4396 17280 4402 17292
rect 4525 17289 4537 17292
rect 4571 17289 4583 17323
rect 4525 17283 4583 17289
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 4893 17323 4951 17329
rect 4893 17320 4905 17323
rect 4672 17292 4905 17320
rect 4672 17280 4678 17292
rect 4893 17289 4905 17292
rect 4939 17289 4951 17323
rect 4893 17283 4951 17289
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 5261 17323 5319 17329
rect 5261 17320 5273 17323
rect 5224 17292 5273 17320
rect 5224 17280 5230 17292
rect 5261 17289 5273 17292
rect 5307 17289 5319 17323
rect 5626 17320 5632 17332
rect 5587 17292 5632 17320
rect 5261 17283 5319 17289
rect 5626 17280 5632 17292
rect 5684 17280 5690 17332
rect 5994 17320 6000 17332
rect 5955 17292 6000 17320
rect 5994 17280 6000 17292
rect 6052 17280 6058 17332
rect 6454 17280 6460 17332
rect 6512 17320 6518 17332
rect 6641 17323 6699 17329
rect 6641 17320 6653 17323
rect 6512 17292 6653 17320
rect 6512 17280 6518 17292
rect 6641 17289 6653 17292
rect 6687 17289 6699 17323
rect 6641 17283 6699 17289
rect 6914 17280 6920 17332
rect 6972 17320 6978 17332
rect 7009 17323 7067 17329
rect 7009 17320 7021 17323
rect 6972 17292 7021 17320
rect 6972 17280 6978 17292
rect 7009 17289 7021 17292
rect 7055 17289 7067 17323
rect 7009 17283 7067 17289
rect 7282 17280 7288 17332
rect 7340 17320 7346 17332
rect 7469 17323 7527 17329
rect 7469 17320 7481 17323
rect 7340 17292 7481 17320
rect 7340 17280 7346 17292
rect 7469 17289 7481 17292
rect 7515 17289 7527 17323
rect 7469 17283 7527 17289
rect 7742 17280 7748 17332
rect 7800 17320 7806 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7800 17292 7941 17320
rect 7800 17280 7806 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 8294 17320 8300 17332
rect 8255 17292 8300 17320
rect 7929 17283 7987 17289
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 9033 17323 9091 17329
rect 9033 17320 9045 17323
rect 8904 17292 9045 17320
rect 8904 17280 8910 17292
rect 9033 17289 9045 17292
rect 9079 17289 9091 17323
rect 9398 17320 9404 17332
rect 9359 17292 9404 17320
rect 9033 17283 9091 17289
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 10597 17323 10655 17329
rect 10597 17320 10609 17323
rect 10284 17292 10609 17320
rect 10284 17280 10290 17292
rect 3878 17252 3884 17264
rect 1780 17224 3884 17252
rect 1780 17193 1808 17224
rect 3878 17212 3884 17224
rect 3936 17212 3942 17264
rect 9306 17252 9312 17264
rect 8496 17224 9312 17252
rect 1765 17187 1823 17193
rect 1765 17153 1777 17187
rect 1811 17153 1823 17187
rect 2130 17184 2136 17196
rect 2091 17156 2136 17184
rect 1765 17147 1823 17153
rect 2130 17144 2136 17156
rect 2188 17144 2194 17196
rect 2501 17187 2559 17193
rect 2501 17153 2513 17187
rect 2547 17184 2559 17187
rect 2869 17187 2927 17193
rect 2547 17156 2774 17184
rect 2547 17153 2559 17156
rect 2501 17147 2559 17153
rect 2746 17116 2774 17156
rect 2869 17153 2881 17187
rect 2915 17184 2927 17187
rect 3142 17184 3148 17196
rect 2915 17156 3148 17184
rect 2915 17153 2927 17156
rect 2869 17147 2927 17153
rect 3142 17144 3148 17156
rect 3200 17144 3206 17196
rect 3237 17187 3295 17193
rect 3237 17153 3249 17187
rect 3283 17184 3295 17187
rect 3418 17184 3424 17196
rect 3283 17156 3424 17184
rect 3283 17153 3295 17156
rect 3237 17147 3295 17153
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 3602 17184 3608 17196
rect 3563 17156 3608 17184
rect 3602 17144 3608 17156
rect 3660 17144 3666 17196
rect 4341 17187 4399 17193
rect 4341 17153 4353 17187
rect 4387 17184 4399 17187
rect 4522 17184 4528 17196
rect 4387 17156 4528 17184
rect 4387 17153 4399 17156
rect 4341 17147 4399 17153
rect 4522 17144 4528 17156
rect 4580 17144 4586 17196
rect 4709 17187 4767 17193
rect 4709 17153 4721 17187
rect 4755 17153 4767 17187
rect 4709 17147 4767 17153
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5077 17147 5135 17153
rect 5445 17187 5503 17193
rect 5445 17153 5457 17187
rect 5491 17184 5503 17187
rect 5534 17184 5540 17196
rect 5491 17156 5540 17184
rect 5491 17153 5503 17156
rect 5445 17147 5503 17153
rect 3786 17116 3792 17128
rect 2746 17088 3792 17116
rect 3786 17076 3792 17088
rect 3844 17076 3850 17128
rect 4430 17076 4436 17128
rect 4488 17116 4494 17128
rect 4724 17116 4752 17147
rect 4488 17088 4752 17116
rect 5092 17116 5120 17147
rect 5534 17144 5540 17156
rect 5592 17144 5598 17196
rect 5810 17184 5816 17196
rect 5771 17156 5816 17184
rect 5810 17144 5816 17156
rect 5868 17144 5874 17196
rect 6178 17184 6184 17196
rect 6139 17156 6184 17184
rect 6178 17144 6184 17156
rect 6236 17144 6242 17196
rect 6362 17144 6368 17196
rect 6420 17184 6426 17196
rect 6825 17187 6883 17193
rect 6825 17184 6837 17187
rect 6420 17156 6837 17184
rect 6420 17144 6426 17156
rect 6825 17153 6837 17156
rect 6871 17153 6883 17187
rect 6825 17147 6883 17153
rect 7193 17187 7251 17193
rect 7193 17153 7205 17187
rect 7239 17153 7251 17187
rect 7193 17147 7251 17153
rect 7653 17187 7711 17193
rect 7653 17153 7665 17187
rect 7699 17184 7711 17187
rect 8113 17187 8171 17193
rect 7699 17156 8064 17184
rect 7699 17153 7711 17156
rect 7653 17147 7711 17153
rect 7098 17116 7104 17128
rect 5092 17088 7104 17116
rect 4488 17076 4494 17088
rect 7098 17076 7104 17088
rect 7156 17076 7162 17128
rect 7208 17116 7236 17147
rect 7834 17116 7840 17128
rect 7208 17088 7840 17116
rect 7834 17076 7840 17088
rect 7892 17076 7898 17128
rect 8036 17116 8064 17156
rect 8113 17153 8125 17187
rect 8159 17184 8171 17187
rect 8202 17184 8208 17196
rect 8159 17156 8208 17184
rect 8159 17153 8171 17156
rect 8113 17147 8171 17153
rect 8202 17144 8208 17156
rect 8260 17144 8266 17196
rect 8496 17193 8524 17224
rect 9306 17212 9312 17224
rect 9364 17212 9370 17264
rect 8481 17187 8539 17193
rect 8481 17153 8493 17187
rect 8527 17153 8539 17187
rect 8481 17147 8539 17153
rect 8757 17187 8815 17193
rect 8757 17153 8769 17187
rect 8803 17184 8815 17187
rect 8938 17184 8944 17196
rect 8803 17156 8944 17184
rect 8803 17153 8815 17156
rect 8757 17147 8815 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 9214 17184 9220 17196
rect 9175 17156 9220 17184
rect 9214 17144 9220 17156
rect 9272 17144 9278 17196
rect 9416 17184 9444 17280
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 9416 17156 9689 17184
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 9766 17144 9772 17196
rect 9824 17184 9830 17196
rect 10520 17193 10548 17292
rect 10597 17289 10609 17292
rect 10643 17289 10655 17323
rect 13265 17323 13323 17329
rect 13265 17320 13277 17323
rect 10597 17283 10655 17289
rect 10704 17292 13277 17320
rect 10704 17252 10732 17292
rect 13265 17289 13277 17292
rect 13311 17289 13323 17323
rect 13265 17283 13323 17289
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 14369 17323 14427 17329
rect 14369 17320 14381 17323
rect 14056 17292 14381 17320
rect 14056 17280 14062 17292
rect 12253 17255 12311 17261
rect 12253 17252 12265 17255
rect 10612 17224 10732 17252
rect 11808 17224 12265 17252
rect 9861 17187 9919 17193
rect 9861 17184 9873 17187
rect 9824 17156 9873 17184
rect 9824 17144 9830 17156
rect 9861 17153 9873 17156
rect 9907 17184 9919 17187
rect 10137 17187 10195 17193
rect 10137 17184 10149 17187
rect 9907 17156 10149 17184
rect 9907 17153 9919 17156
rect 9861 17147 9919 17153
rect 10137 17153 10149 17156
rect 10183 17153 10195 17187
rect 10137 17147 10195 17153
rect 10505 17187 10563 17193
rect 10505 17153 10517 17187
rect 10551 17153 10563 17187
rect 10505 17147 10563 17153
rect 9398 17116 9404 17128
rect 8036 17088 9404 17116
rect 9398 17076 9404 17088
rect 9456 17076 9462 17128
rect 9490 17076 9496 17128
rect 9548 17116 9554 17128
rect 10612 17116 10640 17224
rect 10686 17144 10692 17196
rect 10744 17184 10750 17196
rect 10965 17187 11023 17193
rect 10965 17184 10977 17187
rect 10744 17156 10977 17184
rect 10744 17144 10750 17156
rect 10965 17153 10977 17156
rect 11011 17153 11023 17187
rect 10965 17147 11023 17153
rect 11054 17144 11060 17196
rect 11112 17184 11118 17196
rect 11333 17187 11391 17193
rect 11333 17184 11345 17187
rect 11112 17156 11345 17184
rect 11112 17144 11118 17156
rect 11333 17153 11345 17156
rect 11379 17153 11391 17187
rect 11333 17147 11391 17153
rect 11514 17144 11520 17196
rect 11572 17184 11578 17196
rect 11808 17193 11836 17224
rect 12253 17221 12265 17224
rect 12299 17221 12311 17255
rect 13081 17255 13139 17261
rect 13081 17252 13093 17255
rect 12253 17215 12311 17221
rect 12636 17224 13093 17252
rect 11793 17187 11851 17193
rect 11793 17184 11805 17187
rect 11572 17156 11805 17184
rect 11572 17144 11578 17156
rect 11793 17153 11805 17156
rect 11839 17153 11851 17187
rect 11793 17147 11851 17153
rect 11882 17144 11888 17196
rect 11940 17184 11946 17196
rect 12161 17187 12219 17193
rect 12161 17184 12173 17187
rect 11940 17156 12173 17184
rect 11940 17144 11946 17156
rect 12161 17153 12173 17156
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12526 17144 12532 17196
rect 12584 17184 12590 17196
rect 12636 17193 12664 17224
rect 13081 17221 13093 17224
rect 13127 17221 13139 17255
rect 13081 17215 13139 17221
rect 12621 17187 12679 17193
rect 12621 17184 12633 17187
rect 12584 17156 12633 17184
rect 12584 17144 12590 17156
rect 12621 17153 12633 17156
rect 12667 17153 12679 17187
rect 12621 17147 12679 17153
rect 12710 17144 12716 17196
rect 12768 17184 12774 17196
rect 12989 17187 13047 17193
rect 12989 17184 13001 17187
rect 12768 17156 13001 17184
rect 12768 17144 12774 17156
rect 12989 17153 13001 17156
rect 13035 17153 13047 17187
rect 12989 17147 13047 17153
rect 13170 17144 13176 17196
rect 13228 17184 13234 17196
rect 13449 17187 13507 17193
rect 13449 17184 13461 17187
rect 13228 17156 13461 17184
rect 13228 17144 13234 17156
rect 13449 17153 13461 17156
rect 13495 17153 13507 17187
rect 13449 17147 13507 17153
rect 13538 17144 13544 17196
rect 13596 17184 13602 17196
rect 14292 17193 14320 17292
rect 14369 17289 14381 17292
rect 14415 17289 14427 17323
rect 14369 17283 14427 17289
rect 14553 17323 14611 17329
rect 14553 17289 14565 17323
rect 14599 17289 14611 17323
rect 15562 17320 15568 17332
rect 15523 17292 15568 17320
rect 14553 17283 14611 17289
rect 14568 17252 14596 17283
rect 15562 17280 15568 17292
rect 15620 17280 15626 17332
rect 15197 17255 15255 17261
rect 15197 17252 15209 17255
rect 14384 17224 14596 17252
rect 14752 17224 15209 17252
rect 13817 17187 13875 17193
rect 13817 17184 13829 17187
rect 13596 17156 13829 17184
rect 13596 17144 13602 17156
rect 13817 17153 13829 17156
rect 13863 17153 13875 17187
rect 13817 17147 13875 17153
rect 14277 17187 14335 17193
rect 14277 17153 14289 17187
rect 14323 17153 14335 17187
rect 14277 17147 14335 17153
rect 9548 17088 10640 17116
rect 9548 17076 9554 17088
rect 11238 17076 11244 17128
rect 11296 17116 11302 17128
rect 14384 17116 14412 17224
rect 14458 17144 14464 17196
rect 14516 17184 14522 17196
rect 14752 17193 14780 17224
rect 15197 17221 15209 17224
rect 15243 17221 15255 17255
rect 15197 17215 15255 17221
rect 14737 17187 14795 17193
rect 14737 17184 14749 17187
rect 14516 17156 14749 17184
rect 14516 17144 14522 17156
rect 14737 17153 14749 17156
rect 14783 17153 14795 17187
rect 14737 17147 14795 17153
rect 14826 17144 14832 17196
rect 14884 17184 14890 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 14884 17156 15117 17184
rect 14884 17144 14890 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 11296 17088 14412 17116
rect 11296 17076 11302 17088
rect 14550 17076 14556 17128
rect 14608 17116 14614 17128
rect 15396 17116 15424 17147
rect 14608 17088 15424 17116
rect 14608 17076 14614 17088
rect 9030 17008 9036 17060
rect 9088 17048 9094 17060
rect 10321 17051 10379 17057
rect 10321 17048 10333 17051
rect 9088 17020 10333 17048
rect 9088 17008 9094 17020
rect 10321 17017 10333 17020
rect 10367 17017 10379 17051
rect 10321 17011 10379 17017
rect 11698 17008 11704 17060
rect 11756 17048 11762 17060
rect 14921 17051 14979 17057
rect 14921 17048 14933 17051
rect 11756 17020 14933 17048
rect 11756 17008 11762 17020
rect 14921 17017 14933 17020
rect 14967 17017 14979 17051
rect 14921 17011 14979 17017
rect 8573 16983 8631 16989
rect 8573 16949 8585 16983
rect 8619 16980 8631 16983
rect 8846 16980 8852 16992
rect 8619 16952 8852 16980
rect 8619 16949 8631 16952
rect 8573 16943 8631 16949
rect 8846 16940 8852 16952
rect 8904 16940 8910 16992
rect 9306 16940 9312 16992
rect 9364 16980 9370 16992
rect 9493 16983 9551 16989
rect 9493 16980 9505 16983
rect 9364 16952 9505 16980
rect 9364 16940 9370 16952
rect 9493 16949 9505 16952
rect 9539 16949 9551 16983
rect 10042 16980 10048 16992
rect 10003 16952 10048 16980
rect 9493 16943 9551 16949
rect 10042 16940 10048 16952
rect 10100 16940 10106 16992
rect 10778 16980 10784 16992
rect 10739 16952 10784 16980
rect 10778 16940 10784 16952
rect 10836 16940 10842 16992
rect 11146 16980 11152 16992
rect 11107 16952 11152 16980
rect 11146 16940 11152 16952
rect 11204 16940 11210 16992
rect 11606 16980 11612 16992
rect 11567 16952 11612 16980
rect 11606 16940 11612 16952
rect 11664 16940 11670 16992
rect 11974 16980 11980 16992
rect 11935 16952 11980 16980
rect 11974 16940 11980 16952
rect 12032 16940 12038 16992
rect 12437 16983 12495 16989
rect 12437 16949 12449 16983
rect 12483 16980 12495 16983
rect 12618 16980 12624 16992
rect 12483 16952 12624 16980
rect 12483 16949 12495 16952
rect 12437 16943 12495 16949
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 12802 16980 12808 16992
rect 12763 16952 12808 16980
rect 12802 16940 12808 16952
rect 12860 16940 12866 16992
rect 13538 16940 13544 16992
rect 13596 16980 13602 16992
rect 13633 16983 13691 16989
rect 13633 16980 13645 16983
rect 13596 16952 13645 16980
rect 13596 16940 13602 16952
rect 13633 16949 13645 16952
rect 13679 16949 13691 16983
rect 13633 16943 13691 16949
rect 13722 16940 13728 16992
rect 13780 16980 13786 16992
rect 14093 16983 14151 16989
rect 14093 16980 14105 16983
rect 13780 16952 14105 16980
rect 13780 16940 13786 16952
rect 14093 16949 14105 16952
rect 14139 16949 14151 16983
rect 14093 16943 14151 16949
rect 1104 16890 16008 16912
rect 1104 16838 2824 16890
rect 2876 16838 2888 16890
rect 2940 16838 2952 16890
rect 3004 16838 3016 16890
rect 3068 16838 3080 16890
rect 3132 16838 6572 16890
rect 6624 16838 6636 16890
rect 6688 16838 6700 16890
rect 6752 16838 6764 16890
rect 6816 16838 6828 16890
rect 6880 16838 10320 16890
rect 10372 16838 10384 16890
rect 10436 16838 10448 16890
rect 10500 16838 10512 16890
rect 10564 16838 10576 16890
rect 10628 16838 14068 16890
rect 14120 16838 14132 16890
rect 14184 16838 14196 16890
rect 14248 16838 14260 16890
rect 14312 16838 14324 16890
rect 14376 16838 16008 16890
rect 1104 16816 16008 16838
rect 8938 16776 8944 16788
rect 8899 16748 8944 16776
rect 8938 16736 8944 16748
rect 8996 16736 9002 16788
rect 10686 16776 10692 16788
rect 10647 16748 10692 16776
rect 10686 16736 10692 16748
rect 10744 16736 10750 16788
rect 11054 16776 11060 16788
rect 11015 16748 11060 16776
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11882 16776 11888 16788
rect 11843 16748 11888 16776
rect 11882 16736 11888 16748
rect 11940 16736 11946 16788
rect 12710 16776 12716 16788
rect 12671 16748 12716 16776
rect 12710 16736 12716 16748
rect 12768 16736 12774 16788
rect 13170 16776 13176 16788
rect 13131 16748 13176 16776
rect 13170 16736 13176 16748
rect 13228 16736 13234 16788
rect 13446 16776 13452 16788
rect 13407 16748 13452 16776
rect 13446 16736 13452 16748
rect 13504 16736 13510 16788
rect 14369 16779 14427 16785
rect 14369 16745 14381 16779
rect 14415 16776 14427 16779
rect 14826 16776 14832 16788
rect 14415 16748 14832 16776
rect 14415 16745 14427 16748
rect 14369 16739 14427 16745
rect 14826 16736 14832 16748
rect 14884 16736 14890 16788
rect 2317 16711 2375 16717
rect 2317 16677 2329 16711
rect 2363 16708 2375 16711
rect 2363 16680 2912 16708
rect 2363 16677 2375 16680
rect 2317 16671 2375 16677
rect 1946 16600 1952 16652
rect 2004 16640 2010 16652
rect 2409 16643 2467 16649
rect 2409 16640 2421 16643
rect 2004 16612 2421 16640
rect 2004 16600 2010 16612
rect 2148 16581 2176 16612
rect 2409 16609 2421 16612
rect 2455 16609 2467 16643
rect 2409 16603 2467 16609
rect 1673 16575 1731 16581
rect 1673 16541 1685 16575
rect 1719 16572 1731 16575
rect 2041 16575 2099 16581
rect 1719 16544 1992 16572
rect 1719 16541 1731 16544
rect 1673 16535 1731 16541
rect 1026 16464 1032 16516
rect 1084 16504 1090 16516
rect 1084 16476 1900 16504
rect 1084 16464 1090 16476
rect 566 16396 572 16448
rect 624 16436 630 16448
rect 1872 16445 1900 16476
rect 1489 16439 1547 16445
rect 1489 16436 1501 16439
rect 624 16408 1501 16436
rect 624 16396 630 16408
rect 1489 16405 1501 16408
rect 1535 16405 1547 16439
rect 1489 16399 1547 16405
rect 1857 16439 1915 16445
rect 1857 16405 1869 16439
rect 1903 16405 1915 16439
rect 1964 16436 1992 16544
rect 2041 16541 2053 16575
rect 2087 16541 2099 16575
rect 2041 16535 2099 16541
rect 2133 16575 2191 16581
rect 2133 16541 2145 16575
rect 2179 16541 2191 16575
rect 2884 16572 2912 16680
rect 5810 16668 5816 16720
rect 5868 16708 5874 16720
rect 9950 16708 9956 16720
rect 5868 16680 9956 16708
rect 5868 16668 5874 16680
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 14553 16711 14611 16717
rect 14553 16677 14565 16711
rect 14599 16708 14611 16711
rect 15102 16708 15108 16720
rect 14599 16680 15108 16708
rect 14599 16677 14611 16680
rect 14553 16671 14611 16677
rect 15102 16668 15108 16680
rect 15160 16668 15166 16720
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 11974 16640 11980 16652
rect 6236 16612 11980 16640
rect 6236 16600 6242 16612
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 14737 16643 14795 16649
rect 14737 16609 14749 16643
rect 14783 16640 14795 16643
rect 14783 16612 15700 16640
rect 14783 16609 14795 16612
rect 14737 16603 14795 16609
rect 4246 16572 4252 16584
rect 2133 16535 2191 16541
rect 2240 16568 2636 16572
rect 2240 16544 2774 16568
rect 2884 16544 4252 16572
rect 2056 16504 2084 16535
rect 2240 16504 2268 16544
rect 2608 16540 2774 16544
rect 2056 16476 2268 16504
rect 2746 16504 2774 16540
rect 4246 16532 4252 16544
rect 4304 16532 4310 16584
rect 15028 16581 15056 16612
rect 15013 16575 15071 16581
rect 15013 16541 15025 16575
rect 15059 16574 15071 16575
rect 15289 16575 15347 16581
rect 15059 16546 15093 16574
rect 15059 16541 15071 16546
rect 15013 16535 15071 16541
rect 15289 16541 15301 16575
rect 15335 16541 15347 16575
rect 15289 16535 15347 16541
rect 3970 16504 3976 16516
rect 2746 16476 3976 16504
rect 3970 16464 3976 16476
rect 4028 16464 4034 16516
rect 9214 16464 9220 16516
rect 9272 16504 9278 16516
rect 15304 16504 15332 16535
rect 15378 16532 15384 16584
rect 15436 16572 15442 16584
rect 15565 16575 15623 16581
rect 15565 16572 15577 16575
rect 15436 16544 15577 16572
rect 15436 16532 15442 16544
rect 15565 16541 15577 16544
rect 15611 16541 15623 16575
rect 15672 16572 15700 16612
rect 16114 16572 16120 16584
rect 15672 16544 16120 16572
rect 15565 16535 15623 16541
rect 16114 16532 16120 16544
rect 16172 16532 16178 16584
rect 15654 16504 15660 16516
rect 9272 16476 15148 16504
rect 15304 16476 15660 16504
rect 9272 16464 9278 16476
rect 4062 16436 4068 16448
rect 1964 16408 4068 16436
rect 1857 16399 1915 16405
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 12618 16396 12624 16448
rect 12676 16436 12682 16448
rect 15120 16445 15148 16476
rect 15488 16448 15516 16476
rect 15654 16464 15660 16476
rect 15712 16464 15718 16516
rect 14829 16439 14887 16445
rect 14829 16436 14841 16439
rect 12676 16408 14841 16436
rect 12676 16396 12682 16408
rect 14829 16405 14841 16408
rect 14875 16405 14887 16439
rect 14829 16399 14887 16405
rect 15105 16439 15163 16445
rect 15105 16405 15117 16439
rect 15151 16405 15163 16439
rect 15378 16436 15384 16448
rect 15339 16408 15384 16436
rect 15105 16399 15163 16405
rect 15378 16396 15384 16408
rect 15436 16396 15442 16448
rect 15470 16396 15476 16448
rect 15528 16396 15534 16448
rect 1104 16346 16008 16368
rect 1104 16294 4698 16346
rect 4750 16294 4762 16346
rect 4814 16294 4826 16346
rect 4878 16294 4890 16346
rect 4942 16294 4954 16346
rect 5006 16294 8446 16346
rect 8498 16294 8510 16346
rect 8562 16294 8574 16346
rect 8626 16294 8638 16346
rect 8690 16294 8702 16346
rect 8754 16294 12194 16346
rect 12246 16294 12258 16346
rect 12310 16294 12322 16346
rect 12374 16294 12386 16346
rect 12438 16294 12450 16346
rect 12502 16294 16008 16346
rect 1104 16272 16008 16294
rect 15105 16167 15163 16173
rect 15105 16133 15117 16167
rect 15151 16164 15163 16167
rect 16942 16164 16948 16176
rect 15151 16136 16948 16164
rect 15151 16133 15163 16136
rect 15105 16127 15163 16133
rect 198 16056 204 16108
rect 256 16096 262 16108
rect 15396 16105 15424 16136
rect 16942 16124 16948 16136
rect 17000 16124 17006 16176
rect 1397 16099 1455 16105
rect 1397 16096 1409 16099
rect 256 16068 1409 16096
rect 256 16056 262 16068
rect 1397 16065 1409 16068
rect 1443 16096 1455 16099
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1443 16068 1685 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 15381 16099 15439 16105
rect 15381 16065 15393 16099
rect 15427 16065 15439 16099
rect 15381 16059 15439 16065
rect 15657 16099 15715 16105
rect 15657 16065 15669 16099
rect 15703 16096 15715 16099
rect 16482 16096 16488 16108
rect 15703 16068 16488 16096
rect 15703 16065 15715 16068
rect 15657 16059 15715 16065
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 16028 14979 16031
rect 15672 16028 15700 16059
rect 16482 16056 16488 16068
rect 16540 16056 16546 16108
rect 14967 16000 15700 16028
rect 14967 15997 14979 16000
rect 14921 15991 14979 15997
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 4614 15960 4620 15972
rect 1627 15932 4620 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 4614 15920 4620 15932
rect 4672 15920 4678 15972
rect 15194 15892 15200 15904
rect 15155 15864 15200 15892
rect 15194 15852 15200 15864
rect 15252 15852 15258 15904
rect 15286 15852 15292 15904
rect 15344 15892 15350 15904
rect 15473 15895 15531 15901
rect 15473 15892 15485 15895
rect 15344 15864 15485 15892
rect 15344 15852 15350 15864
rect 15473 15861 15485 15864
rect 15519 15861 15531 15895
rect 15473 15855 15531 15861
rect 1104 15802 16008 15824
rect 1104 15750 2824 15802
rect 2876 15750 2888 15802
rect 2940 15750 2952 15802
rect 3004 15750 3016 15802
rect 3068 15750 3080 15802
rect 3132 15750 6572 15802
rect 6624 15750 6636 15802
rect 6688 15750 6700 15802
rect 6752 15750 6764 15802
rect 6816 15750 6828 15802
rect 6880 15750 10320 15802
rect 10372 15750 10384 15802
rect 10436 15750 10448 15802
rect 10500 15750 10512 15802
rect 10564 15750 10576 15802
rect 10628 15750 14068 15802
rect 14120 15750 14132 15802
rect 14184 15750 14196 15802
rect 14248 15750 14260 15802
rect 14312 15750 14324 15802
rect 14376 15750 16008 15802
rect 1104 15728 16008 15750
rect 15470 15688 15476 15700
rect 15431 15660 15476 15688
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 1104 15258 16008 15280
rect 1104 15206 4698 15258
rect 4750 15206 4762 15258
rect 4814 15206 4826 15258
rect 4878 15206 4890 15258
rect 4942 15206 4954 15258
rect 5006 15206 8446 15258
rect 8498 15206 8510 15258
rect 8562 15206 8574 15258
rect 8626 15206 8638 15258
rect 8690 15206 8702 15258
rect 8754 15206 12194 15258
rect 12246 15206 12258 15258
rect 12310 15206 12322 15258
rect 12374 15206 12386 15258
rect 12438 15206 12450 15258
rect 12502 15206 16008 15258
rect 1104 15184 16008 15206
rect 1104 14714 16008 14736
rect 1104 14662 2824 14714
rect 2876 14662 2888 14714
rect 2940 14662 2952 14714
rect 3004 14662 3016 14714
rect 3068 14662 3080 14714
rect 3132 14662 6572 14714
rect 6624 14662 6636 14714
rect 6688 14662 6700 14714
rect 6752 14662 6764 14714
rect 6816 14662 6828 14714
rect 6880 14662 10320 14714
rect 10372 14662 10384 14714
rect 10436 14662 10448 14714
rect 10500 14662 10512 14714
rect 10564 14662 10576 14714
rect 10628 14662 14068 14714
rect 14120 14662 14132 14714
rect 14184 14662 14196 14714
rect 14248 14662 14260 14714
rect 14312 14662 14324 14714
rect 14376 14662 16008 14714
rect 1104 14640 16008 14662
rect 1104 14170 16008 14192
rect 1104 14118 4698 14170
rect 4750 14118 4762 14170
rect 4814 14118 4826 14170
rect 4878 14118 4890 14170
rect 4942 14118 4954 14170
rect 5006 14118 8446 14170
rect 8498 14118 8510 14170
rect 8562 14118 8574 14170
rect 8626 14118 8638 14170
rect 8690 14118 8702 14170
rect 8754 14118 12194 14170
rect 12246 14118 12258 14170
rect 12310 14118 12322 14170
rect 12374 14118 12386 14170
rect 12438 14118 12450 14170
rect 12502 14118 16008 14170
rect 1104 14096 16008 14118
rect 4614 13920 4620 13932
rect 4575 13892 4620 13920
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 3326 13812 3332 13864
rect 3384 13852 3390 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 3384 13824 4169 13852
rect 3384 13812 3390 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4525 13719 4583 13725
rect 4525 13685 4537 13719
rect 4571 13716 4583 13719
rect 8846 13716 8852 13728
rect 4571 13688 8852 13716
rect 4571 13685 4583 13688
rect 4525 13679 4583 13685
rect 8846 13676 8852 13688
rect 8904 13676 8910 13728
rect 1104 13626 16008 13648
rect 1104 13574 2824 13626
rect 2876 13574 2888 13626
rect 2940 13574 2952 13626
rect 3004 13574 3016 13626
rect 3068 13574 3080 13626
rect 3132 13574 6572 13626
rect 6624 13574 6636 13626
rect 6688 13574 6700 13626
rect 6752 13574 6764 13626
rect 6816 13574 6828 13626
rect 6880 13574 10320 13626
rect 10372 13574 10384 13626
rect 10436 13574 10448 13626
rect 10500 13574 10512 13626
rect 10564 13574 10576 13626
rect 10628 13574 14068 13626
rect 14120 13574 14132 13626
rect 14184 13574 14196 13626
rect 14248 13574 14260 13626
rect 14312 13574 14324 13626
rect 14376 13574 16008 13626
rect 1104 13552 16008 13574
rect 4154 13308 4160 13320
rect 4115 13280 4160 13308
rect 4154 13268 4160 13280
rect 4212 13268 4218 13320
rect 4246 13268 4252 13320
rect 4304 13308 4310 13320
rect 4413 13311 4471 13317
rect 4413 13308 4425 13311
rect 4304 13280 4425 13308
rect 4304 13268 4310 13280
rect 4413 13277 4425 13280
rect 4459 13277 4471 13311
rect 4413 13271 4471 13277
rect 5537 13175 5595 13181
rect 5537 13141 5549 13175
rect 5583 13172 5595 13175
rect 8018 13172 8024 13184
rect 5583 13144 8024 13172
rect 5583 13141 5595 13144
rect 5537 13135 5595 13141
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 1104 13082 16008 13104
rect 1104 13030 4698 13082
rect 4750 13030 4762 13082
rect 4814 13030 4826 13082
rect 4878 13030 4890 13082
rect 4942 13030 4954 13082
rect 5006 13030 8446 13082
rect 8498 13030 8510 13082
rect 8562 13030 8574 13082
rect 8626 13030 8638 13082
rect 8690 13030 8702 13082
rect 8754 13030 12194 13082
rect 12246 13030 12258 13082
rect 12310 13030 12322 13082
rect 12374 13030 12386 13082
rect 12438 13030 12450 13082
rect 12502 13030 16008 13082
rect 1104 13008 16008 13030
rect 4062 12968 4068 12980
rect 4023 12940 4068 12968
rect 4062 12928 4068 12940
rect 4120 12928 4126 12980
rect 5261 12971 5319 12977
rect 5261 12968 5273 12971
rect 4172 12940 5273 12968
rect 3786 12860 3792 12912
rect 3844 12900 3850 12912
rect 4172 12900 4200 12940
rect 5261 12937 5273 12940
rect 5307 12937 5319 12971
rect 5261 12931 5319 12937
rect 7098 12928 7104 12980
rect 7156 12968 7162 12980
rect 7193 12971 7251 12977
rect 7193 12968 7205 12971
rect 7156 12940 7205 12968
rect 7156 12928 7162 12940
rect 7193 12937 7205 12940
rect 7239 12937 7251 12971
rect 9398 12968 9404 12980
rect 9359 12940 9404 12968
rect 7193 12931 7251 12937
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 14369 12971 14427 12977
rect 14369 12937 14381 12971
rect 14415 12968 14427 12971
rect 14550 12968 14556 12980
rect 14415 12940 14556 12968
rect 14415 12937 14427 12940
rect 14369 12931 14427 12937
rect 14550 12928 14556 12940
rect 14608 12928 14614 12980
rect 10226 12900 10232 12912
rect 3844 12872 4200 12900
rect 4816 12872 10232 12900
rect 3844 12860 3850 12872
rect 4816 12841 4844 12872
rect 10226 12860 10232 12872
rect 10284 12860 10290 12912
rect 12406 12872 15424 12900
rect 4249 12835 4307 12841
rect 4249 12801 4261 12835
rect 4295 12801 4307 12835
rect 4249 12795 4307 12801
rect 4801 12835 4859 12841
rect 4801 12801 4813 12835
rect 4847 12801 4859 12835
rect 4801 12795 4859 12801
rect 5445 12835 5503 12841
rect 5445 12801 5457 12835
rect 5491 12832 5503 12835
rect 7374 12832 7380 12844
rect 5491 12804 7236 12832
rect 7335 12804 7380 12832
rect 5491 12801 5503 12804
rect 5445 12795 5503 12801
rect 4264 12764 4292 12795
rect 6086 12764 6092 12776
rect 4264 12736 6092 12764
rect 6086 12724 6092 12736
rect 6144 12724 6150 12776
rect 7208 12764 7236 12804
rect 7374 12792 7380 12804
rect 7432 12792 7438 12844
rect 9582 12832 9588 12844
rect 9543 12804 9588 12832
rect 9582 12792 9588 12804
rect 9640 12792 9646 12844
rect 8294 12764 8300 12776
rect 7208 12736 8300 12764
rect 8294 12724 8300 12736
rect 8352 12724 8358 12776
rect 8846 12724 8852 12776
rect 8904 12764 8910 12776
rect 12406 12764 12434 12872
rect 15396 12841 15424 12872
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 8904 12736 12434 12764
rect 14016 12804 14197 12832
rect 8904 12724 8910 12736
rect 3878 12656 3884 12708
rect 3936 12696 3942 12708
rect 4617 12699 4675 12705
rect 4617 12696 4629 12699
rect 3936 12668 4629 12696
rect 3936 12656 3942 12668
rect 4617 12665 4629 12668
rect 4663 12665 4675 12699
rect 4617 12659 4675 12665
rect 7650 12588 7656 12640
rect 7708 12628 7714 12640
rect 14016 12637 14044 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 15381 12835 15439 12841
rect 15381 12801 15393 12835
rect 15427 12801 15439 12835
rect 15381 12795 15439 12801
rect 14001 12631 14059 12637
rect 14001 12628 14013 12631
rect 7708 12600 14013 12628
rect 7708 12588 7714 12600
rect 14001 12597 14013 12600
rect 14047 12597 14059 12631
rect 15562 12628 15568 12640
rect 15523 12600 15568 12628
rect 14001 12591 14059 12597
rect 15562 12588 15568 12600
rect 15620 12588 15626 12640
rect 1104 12538 16008 12560
rect 1104 12486 2824 12538
rect 2876 12486 2888 12538
rect 2940 12486 2952 12538
rect 3004 12486 3016 12538
rect 3068 12486 3080 12538
rect 3132 12486 6572 12538
rect 6624 12486 6636 12538
rect 6688 12486 6700 12538
rect 6752 12486 6764 12538
rect 6816 12486 6828 12538
rect 6880 12486 10320 12538
rect 10372 12486 10384 12538
rect 10436 12486 10448 12538
rect 10500 12486 10512 12538
rect 10564 12486 10576 12538
rect 10628 12486 14068 12538
rect 14120 12486 14132 12538
rect 14184 12486 14196 12538
rect 14248 12486 14260 12538
rect 14312 12486 14324 12538
rect 14376 12486 16008 12538
rect 1104 12464 16008 12486
rect 1104 11994 16008 12016
rect 1104 11942 4698 11994
rect 4750 11942 4762 11994
rect 4814 11942 4826 11994
rect 4878 11942 4890 11994
rect 4942 11942 4954 11994
rect 5006 11942 8446 11994
rect 8498 11942 8510 11994
rect 8562 11942 8574 11994
rect 8626 11942 8638 11994
rect 8690 11942 8702 11994
rect 8754 11942 12194 11994
rect 12246 11942 12258 11994
rect 12310 11942 12322 11994
rect 12374 11942 12386 11994
rect 12438 11942 12450 11994
rect 12502 11942 16008 11994
rect 1104 11920 16008 11942
rect 4522 11840 4528 11892
rect 4580 11880 4586 11892
rect 7929 11883 7987 11889
rect 7929 11880 7941 11883
rect 4580 11852 7941 11880
rect 4580 11840 4586 11852
rect 7929 11849 7941 11852
rect 7975 11849 7987 11883
rect 7929 11843 7987 11849
rect 1394 11744 1400 11756
rect 1355 11716 1400 11744
rect 1394 11704 1400 11716
rect 1452 11744 1458 11756
rect 1673 11747 1731 11753
rect 1673 11744 1685 11747
rect 1452 11716 1685 11744
rect 1452 11704 1458 11716
rect 1673 11713 1685 11716
rect 1719 11713 1731 11747
rect 7466 11744 7472 11756
rect 7427 11716 7472 11744
rect 1673 11707 1731 11713
rect 7466 11704 7472 11716
rect 7524 11704 7530 11756
rect 8110 11744 8116 11756
rect 8071 11716 8116 11744
rect 8110 11704 8116 11716
rect 8168 11704 8174 11756
rect 7558 11676 7564 11688
rect 7519 11648 7564 11676
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 7653 11679 7711 11685
rect 7653 11645 7665 11679
rect 7699 11645 7711 11679
rect 7653 11639 7711 11645
rect 5442 11568 5448 11620
rect 5500 11608 5506 11620
rect 5500 11580 6040 11608
rect 5500 11568 5506 11580
rect 1581 11543 1639 11549
rect 1581 11509 1593 11543
rect 1627 11540 1639 11543
rect 5902 11540 5908 11552
rect 1627 11512 5908 11540
rect 1627 11509 1639 11512
rect 1581 11503 1639 11509
rect 5902 11500 5908 11512
rect 5960 11500 5966 11552
rect 6012 11540 6040 11580
rect 6914 11568 6920 11620
rect 6972 11608 6978 11620
rect 7668 11608 7696 11639
rect 6972 11580 7696 11608
rect 6972 11568 6978 11580
rect 7101 11543 7159 11549
rect 7101 11540 7113 11543
rect 6012 11512 7113 11540
rect 7101 11509 7113 11512
rect 7147 11509 7159 11543
rect 7101 11503 7159 11509
rect 1104 11450 16008 11472
rect 1104 11398 2824 11450
rect 2876 11398 2888 11450
rect 2940 11398 2952 11450
rect 3004 11398 3016 11450
rect 3068 11398 3080 11450
rect 3132 11398 6572 11450
rect 6624 11398 6636 11450
rect 6688 11398 6700 11450
rect 6752 11398 6764 11450
rect 6816 11398 6828 11450
rect 6880 11398 10320 11450
rect 10372 11398 10384 11450
rect 10436 11398 10448 11450
rect 10500 11398 10512 11450
rect 10564 11398 10576 11450
rect 10628 11398 14068 11450
rect 14120 11398 14132 11450
rect 14184 11398 14196 11450
rect 14248 11398 14260 11450
rect 14312 11398 14324 11450
rect 14376 11398 16008 11450
rect 1104 11376 16008 11398
rect 6454 11296 6460 11348
rect 6512 11336 6518 11348
rect 6512 11308 6914 11336
rect 6512 11296 6518 11308
rect 4338 11024 4344 11076
rect 4396 11064 4402 11076
rect 5258 11064 5264 11076
rect 4396 11036 5264 11064
rect 4396 11024 4402 11036
rect 5258 11024 5264 11036
rect 5316 11064 5322 11076
rect 6273 11067 6331 11073
rect 6273 11064 6285 11067
rect 5316 11036 6285 11064
rect 5316 11024 5322 11036
rect 6273 11033 6285 11036
rect 6319 11033 6331 11067
rect 6886 11064 6914 11308
rect 9122 11296 9128 11348
rect 9180 11336 9186 11348
rect 9490 11336 9496 11348
rect 9180 11308 9496 11336
rect 9180 11296 9186 11308
rect 9490 11296 9496 11308
rect 9548 11296 9554 11348
rect 7926 11228 7932 11280
rect 7984 11268 7990 11280
rect 8941 11271 8999 11277
rect 8941 11268 8953 11271
rect 7984 11240 8953 11268
rect 7984 11228 7990 11240
rect 8941 11237 8953 11240
rect 8987 11237 8999 11271
rect 8941 11231 8999 11237
rect 9490 11200 9496 11212
rect 9451 11172 9496 11200
rect 9490 11160 9496 11172
rect 9548 11160 9554 11212
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11132 9367 11135
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9355 11104 9781 11132
rect 9355 11101 9367 11104
rect 9309 11095 9367 11101
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 8021 11067 8079 11073
rect 6886 11036 7236 11064
rect 6273 11027 6331 11033
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 7098 10996 7104 11008
rect 5684 10968 7104 10996
rect 5684 10956 5690 10968
rect 7098 10956 7104 10968
rect 7156 10956 7162 11008
rect 7208 10996 7236 11036
rect 8021 11033 8033 11067
rect 8067 11064 8079 11067
rect 9674 11064 9680 11076
rect 8067 11036 9680 11064
rect 8067 11033 8079 11036
rect 8021 11027 8079 11033
rect 9674 11024 9680 11036
rect 9732 11024 9738 11076
rect 9306 10996 9312 11008
rect 7208 10968 9312 10996
rect 9306 10956 9312 10968
rect 9364 10956 9370 11008
rect 9398 10956 9404 11008
rect 9456 10996 9462 11008
rect 9456 10968 9501 10996
rect 9456 10956 9462 10968
rect 12710 10956 12716 11008
rect 12768 10996 12774 11008
rect 13722 10996 13728 11008
rect 12768 10968 13728 10996
rect 12768 10956 12774 10968
rect 13722 10956 13728 10968
rect 13780 10956 13786 11008
rect 1104 10906 16008 10928
rect 1104 10854 4698 10906
rect 4750 10854 4762 10906
rect 4814 10854 4826 10906
rect 4878 10854 4890 10906
rect 4942 10854 4954 10906
rect 5006 10854 8446 10906
rect 8498 10854 8510 10906
rect 8562 10854 8574 10906
rect 8626 10854 8638 10906
rect 8690 10854 8702 10906
rect 8754 10854 12194 10906
rect 12246 10854 12258 10906
rect 12310 10854 12322 10906
rect 12374 10854 12386 10906
rect 12438 10854 12450 10906
rect 12502 10854 16008 10906
rect 1104 10832 16008 10854
rect 3053 10795 3111 10801
rect 3053 10761 3065 10795
rect 3099 10792 3111 10795
rect 4154 10792 4160 10804
rect 3099 10764 4160 10792
rect 3099 10761 3111 10764
rect 3053 10755 3111 10761
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 7009 10795 7067 10801
rect 7009 10792 7021 10795
rect 4448 10764 7021 10792
rect 4338 10724 4344 10736
rect 4299 10696 4344 10724
rect 4338 10684 4344 10696
rect 4396 10684 4402 10736
rect 3418 10616 3424 10668
rect 3476 10656 3482 10668
rect 4448 10656 4476 10764
rect 7009 10761 7021 10764
rect 7055 10761 7067 10795
rect 7009 10755 7067 10761
rect 7558 10752 7564 10804
rect 7616 10792 7622 10804
rect 9125 10795 9183 10801
rect 9125 10792 9137 10795
rect 7616 10764 9137 10792
rect 7616 10752 7622 10764
rect 9125 10761 9137 10764
rect 9171 10761 9183 10795
rect 9125 10755 9183 10761
rect 9493 10795 9551 10801
rect 9493 10761 9505 10795
rect 9539 10792 9551 10795
rect 9953 10795 10011 10801
rect 9953 10792 9965 10795
rect 9539 10764 9965 10792
rect 9539 10761 9551 10764
rect 9493 10755 9551 10761
rect 9953 10761 9965 10764
rect 9999 10761 10011 10795
rect 9953 10755 10011 10761
rect 10226 10752 10232 10804
rect 10284 10792 10290 10804
rect 10413 10795 10471 10801
rect 10413 10792 10425 10795
rect 10284 10764 10425 10792
rect 10284 10752 10290 10764
rect 10413 10761 10425 10764
rect 10459 10792 10471 10795
rect 10686 10792 10692 10804
rect 10459 10764 10692 10792
rect 10459 10761 10471 10764
rect 10413 10755 10471 10761
rect 10686 10752 10692 10764
rect 10744 10752 10750 10804
rect 7742 10724 7748 10736
rect 5920 10696 6914 10724
rect 5626 10656 5632 10668
rect 3476 10628 4476 10656
rect 5587 10628 5632 10656
rect 3476 10616 3482 10628
rect 5626 10616 5632 10628
rect 5684 10616 5690 10668
rect 5920 10665 5948 10696
rect 5905 10659 5963 10665
rect 5905 10625 5917 10659
rect 5951 10625 5963 10659
rect 6178 10656 6184 10668
rect 6139 10628 6184 10656
rect 5905 10619 5963 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6270 10616 6276 10668
rect 6328 10656 6334 10668
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 6328 10628 6745 10656
rect 6328 10616 6334 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 3234 10548 3240 10600
rect 3292 10588 3298 10600
rect 3292 10560 6592 10588
rect 3292 10548 3298 10560
rect 5534 10480 5540 10532
rect 5592 10520 5598 10532
rect 6178 10520 6184 10532
rect 5592 10492 6184 10520
rect 5592 10480 5598 10492
rect 6178 10480 6184 10492
rect 6236 10480 6242 10532
rect 6564 10529 6592 10560
rect 6549 10523 6607 10529
rect 6549 10489 6561 10523
rect 6595 10489 6607 10523
rect 6549 10483 6607 10489
rect 5074 10412 5080 10464
rect 5132 10452 5138 10464
rect 5445 10455 5503 10461
rect 5445 10452 5457 10455
rect 5132 10424 5457 10452
rect 5132 10412 5138 10424
rect 5445 10421 5457 10424
rect 5491 10421 5503 10455
rect 5718 10452 5724 10464
rect 5679 10424 5724 10452
rect 5445 10415 5503 10421
rect 5718 10412 5724 10424
rect 5776 10412 5782 10464
rect 5994 10452 6000 10464
rect 5955 10424 6000 10452
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6886 10452 6914 10696
rect 7208 10696 7748 10724
rect 7208 10665 7236 10696
rect 7742 10684 7748 10696
rect 7800 10684 7806 10736
rect 7834 10684 7840 10736
rect 7892 10724 7898 10736
rect 11790 10724 11796 10736
rect 7892 10696 11796 10724
rect 7892 10684 7898 10696
rect 11790 10684 11796 10696
rect 11848 10684 11854 10736
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 7282 10616 7288 10668
rect 7340 10656 7346 10668
rect 7633 10659 7691 10665
rect 7633 10656 7645 10659
rect 7340 10628 7645 10656
rect 7340 10616 7346 10628
rect 7633 10625 7645 10628
rect 7679 10625 7691 10659
rect 7633 10619 7691 10625
rect 9490 10616 9496 10668
rect 9548 10656 9554 10668
rect 9548 10628 9720 10656
rect 9548 10616 9554 10628
rect 7006 10548 7012 10600
rect 7064 10588 7070 10600
rect 7377 10591 7435 10597
rect 7377 10588 7389 10591
rect 7064 10560 7389 10588
rect 7064 10548 7070 10560
rect 7377 10557 7389 10560
rect 7423 10557 7435 10591
rect 7377 10551 7435 10557
rect 9306 10548 9312 10600
rect 9364 10588 9370 10600
rect 9692 10597 9720 10628
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 10321 10659 10379 10665
rect 10321 10656 10333 10659
rect 10192 10628 10333 10656
rect 10192 10616 10198 10628
rect 10321 10625 10333 10628
rect 10367 10625 10379 10659
rect 10321 10619 10379 10625
rect 9585 10591 9643 10597
rect 9585 10588 9597 10591
rect 9364 10560 9597 10588
rect 9364 10548 9370 10560
rect 9585 10557 9597 10560
rect 9631 10557 9643 10591
rect 9585 10551 9643 10557
rect 9677 10591 9735 10597
rect 9677 10557 9689 10591
rect 9723 10557 9735 10591
rect 9677 10551 9735 10557
rect 10226 10548 10232 10600
rect 10284 10588 10290 10600
rect 10505 10591 10563 10597
rect 10505 10588 10517 10591
rect 10284 10560 10517 10588
rect 10284 10548 10290 10560
rect 10505 10557 10517 10560
rect 10551 10557 10563 10591
rect 10505 10551 10563 10557
rect 11146 10520 11152 10532
rect 8312 10492 11152 10520
rect 8312 10452 8340 10492
rect 11146 10480 11152 10492
rect 11204 10480 11210 10532
rect 6886 10424 8340 10452
rect 8757 10455 8815 10461
rect 8757 10421 8769 10455
rect 8803 10452 8815 10455
rect 8846 10452 8852 10464
rect 8803 10424 8852 10452
rect 8803 10421 8815 10424
rect 8757 10415 8815 10421
rect 8846 10412 8852 10424
rect 8904 10412 8910 10464
rect 9858 10412 9864 10464
rect 9916 10452 9922 10464
rect 10778 10452 10784 10464
rect 9916 10424 10784 10452
rect 9916 10412 9922 10424
rect 10778 10412 10784 10424
rect 10836 10412 10842 10464
rect 12894 10412 12900 10464
rect 12952 10452 12958 10464
rect 15378 10452 15384 10464
rect 12952 10424 15384 10452
rect 12952 10412 12958 10424
rect 15378 10412 15384 10424
rect 15436 10412 15442 10464
rect 1104 10362 16008 10384
rect 1104 10310 2824 10362
rect 2876 10310 2888 10362
rect 2940 10310 2952 10362
rect 3004 10310 3016 10362
rect 3068 10310 3080 10362
rect 3132 10310 6572 10362
rect 6624 10310 6636 10362
rect 6688 10310 6700 10362
rect 6752 10310 6764 10362
rect 6816 10310 6828 10362
rect 6880 10310 10320 10362
rect 10372 10310 10384 10362
rect 10436 10310 10448 10362
rect 10500 10310 10512 10362
rect 10564 10310 10576 10362
rect 10628 10310 14068 10362
rect 14120 10310 14132 10362
rect 14184 10310 14196 10362
rect 14248 10310 14260 10362
rect 14312 10310 14324 10362
rect 14376 10310 16008 10362
rect 1104 10288 16008 10310
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 6454 10248 6460 10260
rect 4764 10220 6460 10248
rect 4764 10208 4770 10220
rect 6454 10208 6460 10220
rect 6512 10208 6518 10260
rect 7098 10208 7104 10260
rect 7156 10248 7162 10260
rect 9030 10248 9036 10260
rect 7156 10220 9036 10248
rect 7156 10208 7162 10220
rect 9030 10208 9036 10220
rect 9088 10208 9094 10260
rect 9950 10208 9956 10260
rect 10008 10248 10014 10260
rect 10321 10251 10379 10257
rect 10321 10248 10333 10251
rect 10008 10220 10333 10248
rect 10008 10208 10014 10220
rect 10321 10217 10333 10220
rect 10367 10217 10379 10251
rect 10870 10248 10876 10260
rect 10831 10220 10876 10248
rect 10321 10211 10379 10217
rect 10870 10208 10876 10220
rect 10928 10208 10934 10260
rect 12710 10248 12716 10260
rect 11808 10220 12716 10248
rect 3375 10183 3433 10189
rect 3375 10149 3387 10183
rect 3421 10180 3433 10183
rect 3421 10152 6132 10180
rect 3421 10149 3433 10152
rect 3375 10143 3433 10149
rect 5442 10072 5448 10124
rect 5500 10112 5506 10124
rect 5537 10115 5595 10121
rect 5537 10112 5549 10115
rect 5500 10084 5549 10112
rect 5500 10072 5506 10084
rect 5537 10081 5549 10084
rect 5583 10081 5595 10115
rect 5537 10075 5595 10081
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 5810 10112 5816 10124
rect 5767 10084 5816 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 5810 10072 5816 10084
rect 5868 10072 5874 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 6104 10121 6132 10152
rect 6178 10140 6184 10192
rect 6236 10180 6242 10192
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 6236 10152 8953 10180
rect 6236 10140 6242 10152
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 9858 10180 9864 10192
rect 8941 10143 8999 10149
rect 9048 10152 9864 10180
rect 6089 10115 6147 10121
rect 5960 10084 6005 10112
rect 5960 10072 5966 10084
rect 6089 10081 6101 10115
rect 6135 10081 6147 10115
rect 7558 10112 7564 10124
rect 7519 10084 7564 10112
rect 6089 10075 6147 10081
rect 7558 10072 7564 10084
rect 7616 10072 7622 10124
rect 8018 10072 8024 10124
rect 8076 10112 8082 10124
rect 8113 10115 8171 10121
rect 8113 10112 8125 10115
rect 8076 10084 8125 10112
rect 8076 10072 8082 10084
rect 8113 10081 8125 10084
rect 8159 10081 8171 10115
rect 9048 10112 9076 10152
rect 9858 10140 9864 10152
rect 9916 10140 9922 10192
rect 10042 10140 10048 10192
rect 10100 10180 10106 10192
rect 10597 10183 10655 10189
rect 10597 10180 10609 10183
rect 10100 10152 10609 10180
rect 10100 10140 10106 10152
rect 10597 10149 10609 10152
rect 10643 10149 10655 10183
rect 11808 10180 11836 10220
rect 12710 10208 12716 10220
rect 12768 10208 12774 10260
rect 13078 10248 13084 10260
rect 13039 10220 13084 10248
rect 13078 10208 13084 10220
rect 13136 10208 13142 10260
rect 13354 10248 13360 10260
rect 13315 10220 13360 10248
rect 13354 10208 13360 10220
rect 13412 10208 13418 10260
rect 13630 10248 13636 10260
rect 13591 10220 13636 10248
rect 13630 10208 13636 10220
rect 13688 10208 13694 10260
rect 10597 10143 10655 10149
rect 10704 10152 11836 10180
rect 8113 10075 8171 10081
rect 8404 10084 9076 10112
rect 3326 10053 3332 10056
rect 3304 10047 3332 10053
rect 3304 10013 3316 10047
rect 3304 10007 3332 10013
rect 3326 10004 3332 10007
rect 3384 10004 3390 10056
rect 4706 10004 4712 10056
rect 4764 10044 4770 10056
rect 4764 10016 4809 10044
rect 4764 10004 4770 10016
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 4985 10047 5043 10053
rect 4985 10044 4997 10047
rect 4948 10016 4997 10044
rect 4948 10004 4954 10016
rect 4985 10013 4997 10016
rect 5031 10013 5043 10047
rect 4985 10007 5043 10013
rect 8294 10004 8300 10056
rect 8352 10044 8358 10056
rect 8404 10053 8432 10084
rect 9490 10072 9496 10124
rect 9548 10112 9554 10124
rect 9769 10115 9827 10121
rect 9769 10112 9781 10115
rect 9548 10084 9781 10112
rect 9548 10072 9554 10084
rect 9769 10081 9781 10084
rect 9815 10081 9827 10115
rect 10704 10112 10732 10152
rect 11882 10140 11888 10192
rect 11940 10180 11946 10192
rect 12253 10183 12311 10189
rect 12253 10180 12265 10183
rect 11940 10152 12265 10180
rect 11940 10140 11946 10152
rect 12253 10149 12265 10152
rect 12299 10149 12311 10183
rect 12526 10180 12532 10192
rect 12487 10152 12532 10180
rect 12253 10143 12311 10149
rect 12526 10140 12532 10152
rect 12584 10140 12590 10192
rect 15286 10180 15292 10192
rect 13004 10152 15292 10180
rect 11238 10112 11244 10124
rect 9769 10075 9827 10081
rect 10244 10084 10732 10112
rect 10796 10084 11244 10112
rect 8389 10047 8447 10053
rect 8389 10044 8401 10047
rect 8352 10016 8401 10044
rect 8352 10004 8358 10016
rect 8389 10013 8401 10016
rect 8435 10013 8447 10047
rect 9122 10044 9128 10056
rect 9083 10016 9128 10044
rect 8389 10007 8447 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 9214 10004 9220 10056
rect 9272 10044 9278 10056
rect 10244 10053 10272 10084
rect 10796 10053 10824 10084
rect 11238 10072 11244 10084
rect 11296 10072 11302 10124
rect 11698 10112 11704 10124
rect 11348 10084 11704 10112
rect 9677 10047 9735 10053
rect 9677 10044 9689 10047
rect 9272 10016 9689 10044
rect 9272 10004 9278 10016
rect 9677 10013 9689 10016
rect 9723 10013 9735 10047
rect 9677 10007 9735 10013
rect 10229 10047 10287 10053
rect 10229 10013 10241 10047
rect 10275 10013 10287 10047
rect 10229 10007 10287 10013
rect 10505 10047 10563 10053
rect 10505 10013 10517 10047
rect 10551 10013 10563 10047
rect 10505 10007 10563 10013
rect 10781 10047 10839 10053
rect 10781 10013 10793 10047
rect 10827 10013 10839 10047
rect 11054 10044 11060 10056
rect 11015 10016 11060 10044
rect 10781 10007 10839 10013
rect 3970 9936 3976 9988
rect 4028 9976 4034 9988
rect 5445 9979 5503 9985
rect 4028 9948 4844 9976
rect 4028 9936 4034 9948
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 4816 9917 4844 9948
rect 5445 9945 5457 9979
rect 5491 9976 5503 9979
rect 5491 9948 6040 9976
rect 5491 9945 5503 9948
rect 5445 9939 5503 9945
rect 4525 9911 4583 9917
rect 4525 9908 4537 9911
rect 2096 9880 4537 9908
rect 2096 9868 2102 9880
rect 4525 9877 4537 9880
rect 4571 9877 4583 9911
rect 4525 9871 4583 9877
rect 4801 9911 4859 9917
rect 4801 9877 4813 9911
rect 4847 9877 4859 9911
rect 4801 9871 4859 9877
rect 5077 9911 5135 9917
rect 5077 9877 5089 9911
rect 5123 9908 5135 9911
rect 5166 9908 5172 9920
rect 5123 9880 5172 9908
rect 5123 9877 5135 9880
rect 5077 9871 5135 9877
rect 5166 9868 5172 9880
rect 5224 9868 5230 9920
rect 6012 9908 6040 9948
rect 9766 9936 9772 9988
rect 9824 9976 9830 9988
rect 10520 9976 10548 10007
rect 11054 10004 11060 10016
rect 11112 10004 11118 10056
rect 11348 10053 11376 10084
rect 11698 10072 11704 10084
rect 11756 10072 11762 10124
rect 12894 10112 12900 10124
rect 11900 10084 12900 10112
rect 11900 10053 11928 10084
rect 12894 10072 12900 10084
rect 12952 10072 12958 10124
rect 11333 10047 11391 10053
rect 11333 10013 11345 10047
rect 11379 10013 11391 10047
rect 11333 10007 11391 10013
rect 11609 10047 11667 10053
rect 11609 10013 11621 10047
rect 11655 10013 11667 10047
rect 11609 10007 11667 10013
rect 11885 10047 11943 10053
rect 11885 10013 11897 10047
rect 11931 10013 11943 10047
rect 11885 10007 11943 10013
rect 9824 9948 10548 9976
rect 11624 9976 11652 10007
rect 11974 10004 11980 10056
rect 12032 10044 12038 10056
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 12032 10016 12173 10044
rect 12032 10004 12038 10016
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12437 10047 12495 10053
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 12618 10044 12624 10056
rect 12483 10016 12624 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 13004 10053 13032 10152
rect 15286 10140 15292 10152
rect 15344 10140 15350 10192
rect 15194 10112 15200 10124
rect 13556 10084 15200 10112
rect 13556 10053 13584 10084
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 12713 10047 12771 10053
rect 12713 10013 12725 10047
rect 12759 10013 12771 10047
rect 12713 10007 12771 10013
rect 12989 10047 13047 10053
rect 12989 10013 13001 10047
rect 13035 10013 13047 10047
rect 12989 10007 13047 10013
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10013 13323 10047
rect 13265 10007 13323 10013
rect 13541 10047 13599 10053
rect 13541 10013 13553 10047
rect 13587 10013 13599 10047
rect 13814 10044 13820 10056
rect 13775 10016 13820 10044
rect 13541 10007 13599 10013
rect 12728 9976 12756 10007
rect 13280 9976 13308 10007
rect 13814 10004 13820 10016
rect 13872 10004 13878 10056
rect 14918 9976 14924 9988
rect 11624 9948 12664 9976
rect 12728 9948 13216 9976
rect 13280 9948 14924 9976
rect 9824 9936 9830 9948
rect 12636 9920 12664 9948
rect 7190 9908 7196 9920
rect 6012 9880 7196 9908
rect 7190 9868 7196 9880
rect 7248 9868 7254 9920
rect 8202 9868 8208 9920
rect 8260 9908 8266 9920
rect 8297 9911 8355 9917
rect 8297 9908 8309 9911
rect 8260 9880 8309 9908
rect 8260 9868 8266 9880
rect 8297 9877 8309 9880
rect 8343 9877 8355 9911
rect 8297 9871 8355 9877
rect 8757 9911 8815 9917
rect 8757 9877 8769 9911
rect 8803 9908 8815 9911
rect 9030 9908 9036 9920
rect 8803 9880 9036 9908
rect 8803 9877 8815 9880
rect 8757 9871 8815 9877
rect 9030 9868 9036 9880
rect 9088 9868 9094 9920
rect 9214 9908 9220 9920
rect 9175 9880 9220 9908
rect 9214 9868 9220 9880
rect 9272 9868 9278 9920
rect 9582 9908 9588 9920
rect 9543 9880 9588 9908
rect 9582 9868 9588 9880
rect 9640 9868 9646 9920
rect 9950 9868 9956 9920
rect 10008 9908 10014 9920
rect 10045 9911 10103 9917
rect 10045 9908 10057 9911
rect 10008 9880 10057 9908
rect 10008 9868 10014 9880
rect 10045 9877 10057 9880
rect 10091 9877 10103 9911
rect 10045 9871 10103 9877
rect 11149 9911 11207 9917
rect 11149 9877 11161 9911
rect 11195 9908 11207 9911
rect 11238 9908 11244 9920
rect 11195 9880 11244 9908
rect 11195 9877 11207 9880
rect 11149 9871 11207 9877
rect 11238 9868 11244 9880
rect 11296 9868 11302 9920
rect 11422 9908 11428 9920
rect 11383 9880 11428 9908
rect 11422 9868 11428 9880
rect 11480 9868 11486 9920
rect 11514 9868 11520 9920
rect 11572 9908 11578 9920
rect 11701 9911 11759 9917
rect 11701 9908 11713 9911
rect 11572 9880 11713 9908
rect 11572 9868 11578 9880
rect 11701 9877 11713 9880
rect 11747 9877 11759 9911
rect 11701 9871 11759 9877
rect 11790 9868 11796 9920
rect 11848 9908 11854 9920
rect 11977 9911 12035 9917
rect 11977 9908 11989 9911
rect 11848 9880 11989 9908
rect 11848 9868 11854 9880
rect 11977 9877 11989 9880
rect 12023 9877 12035 9911
rect 11977 9871 12035 9877
rect 12618 9868 12624 9920
rect 12676 9868 12682 9920
rect 12710 9868 12716 9920
rect 12768 9908 12774 9920
rect 12805 9911 12863 9917
rect 12805 9908 12817 9911
rect 12768 9880 12817 9908
rect 12768 9868 12774 9880
rect 12805 9877 12817 9880
rect 12851 9877 12863 9911
rect 13188 9908 13216 9948
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 14734 9908 14740 9920
rect 13188 9880 14740 9908
rect 12805 9871 12863 9877
rect 14734 9868 14740 9880
rect 14792 9868 14798 9920
rect 1104 9818 16008 9840
rect 1104 9766 4698 9818
rect 4750 9766 4762 9818
rect 4814 9766 4826 9818
rect 4878 9766 4890 9818
rect 4942 9766 4954 9818
rect 5006 9766 8446 9818
rect 8498 9766 8510 9818
rect 8562 9766 8574 9818
rect 8626 9766 8638 9818
rect 8690 9766 8702 9818
rect 8754 9766 12194 9818
rect 12246 9766 12258 9818
rect 12310 9766 12322 9818
rect 12374 9766 12386 9818
rect 12438 9766 12450 9818
rect 12502 9766 16008 9818
rect 1104 9744 16008 9766
rect 3418 9664 3424 9716
rect 3476 9704 3482 9716
rect 5166 9704 5172 9716
rect 3476 9676 5172 9704
rect 3476 9664 3482 9676
rect 5166 9664 5172 9676
rect 5224 9664 5230 9716
rect 5442 9664 5448 9716
rect 5500 9704 5506 9716
rect 5500 9676 5764 9704
rect 5500 9664 5506 9676
rect 3053 9639 3111 9645
rect 3053 9605 3065 9639
rect 3099 9636 3111 9639
rect 3326 9636 3332 9648
rect 3099 9608 3332 9636
rect 3099 9605 3111 9608
rect 3053 9599 3111 9605
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 5736 9636 5764 9676
rect 5810 9664 5816 9716
rect 5868 9704 5874 9716
rect 6362 9704 6368 9716
rect 5868 9676 6368 9704
rect 5868 9664 5874 9676
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 8294 9704 8300 9716
rect 6472 9676 8300 9704
rect 6472 9636 6500 9676
rect 8294 9664 8300 9676
rect 8352 9664 8358 9716
rect 9306 9704 9312 9716
rect 9267 9676 9312 9704
rect 9306 9664 9312 9676
rect 9364 9664 9370 9716
rect 10226 9704 10232 9716
rect 9508 9676 10232 9704
rect 5736 9608 6500 9636
rect 6656 9608 7328 9636
rect 5810 9568 5816 9580
rect 5771 9540 5816 9568
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 6181 9571 6239 9577
rect 6181 9537 6193 9571
rect 6227 9568 6239 9571
rect 6656 9568 6684 9608
rect 6227 9540 6684 9568
rect 6733 9571 6791 9577
rect 6227 9537 6239 9540
rect 6181 9531 6239 9537
rect 6733 9537 6745 9571
rect 6779 9552 6791 9571
rect 7098 9568 7104 9580
rect 6840 9552 7104 9568
rect 6779 9540 7104 9552
rect 6779 9537 6868 9540
rect 6733 9531 6868 9537
rect 6748 9524 6868 9531
rect 7098 9528 7104 9540
rect 7156 9528 7162 9580
rect 7300 9568 7328 9608
rect 7374 9596 7380 9648
rect 7432 9636 7438 9648
rect 8754 9636 8760 9648
rect 7432 9608 8760 9636
rect 7432 9596 7438 9608
rect 8754 9596 8760 9608
rect 8812 9596 8818 9648
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 8941 9639 8999 9645
rect 8941 9636 8953 9639
rect 8904 9608 8953 9636
rect 8904 9596 8910 9608
rect 8941 9605 8953 9608
rect 8987 9636 8999 9639
rect 9122 9636 9128 9648
rect 8987 9608 9128 9636
rect 8987 9605 8999 9608
rect 8941 9599 8999 9605
rect 9122 9596 9128 9608
rect 9180 9596 9186 9648
rect 7650 9568 7656 9580
rect 7300 9540 7656 9568
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7949 9571 8007 9577
rect 7949 9537 7961 9571
rect 7995 9568 8007 9571
rect 8478 9568 8484 9580
rect 7995 9540 8484 9568
rect 7995 9537 8007 9540
rect 7949 9531 8007 9537
rect 8478 9528 8484 9540
rect 8536 9528 8542 9580
rect 9508 9568 9536 9676
rect 10226 9664 10232 9676
rect 10284 9664 10290 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 13630 9704 13636 9716
rect 12676 9676 13636 9704
rect 12676 9664 12682 9676
rect 13630 9664 13636 9676
rect 13688 9664 13694 9716
rect 13538 9636 13544 9648
rect 9600 9608 13544 9636
rect 9600 9577 9628 9608
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 8680 9540 9536 9568
rect 9585 9571 9643 9577
rect 2777 9503 2835 9509
rect 2777 9469 2789 9503
rect 2823 9500 2835 9503
rect 3234 9500 3240 9512
rect 2823 9472 3004 9500
rect 3195 9472 3240 9500
rect 2823 9469 2835 9472
rect 2777 9463 2835 9469
rect 2976 9432 3004 9472
rect 3234 9460 3240 9472
rect 3292 9460 3298 9512
rect 4246 9460 4252 9512
rect 4304 9500 4310 9512
rect 8202 9500 8208 9512
rect 4304 9472 6132 9500
rect 8163 9472 8208 9500
rect 4304 9460 4310 9472
rect 3142 9432 3148 9444
rect 2976 9404 3148 9432
rect 3142 9392 3148 9404
rect 3200 9392 3206 9444
rect 4154 9392 4160 9444
rect 4212 9432 4218 9444
rect 5997 9435 6055 9441
rect 5997 9432 6009 9435
rect 4212 9404 6009 9432
rect 4212 9392 4218 9404
rect 5997 9401 6009 9404
rect 6043 9401 6055 9435
rect 5997 9395 6055 9401
rect 2130 9324 2136 9376
rect 2188 9364 2194 9376
rect 5629 9367 5687 9373
rect 5629 9364 5641 9367
rect 2188 9336 5641 9364
rect 2188 9324 2194 9336
rect 5629 9333 5641 9336
rect 5675 9333 5687 9367
rect 6104 9364 6132 9472
rect 8202 9460 8208 9472
rect 8260 9460 8266 9512
rect 8680 9509 8708 9540
rect 9585 9537 9597 9571
rect 9631 9537 9643 9571
rect 9585 9531 9643 9537
rect 9861 9571 9919 9577
rect 9861 9537 9873 9571
rect 9907 9568 9919 9571
rect 12802 9568 12808 9580
rect 9907 9540 12808 9568
rect 9907 9537 9919 9540
rect 9861 9531 9919 9537
rect 12802 9528 12808 9540
rect 12860 9528 12866 9580
rect 8665 9503 8723 9509
rect 8665 9469 8677 9503
rect 8711 9469 8723 9503
rect 8846 9500 8852 9512
rect 8807 9472 8852 9500
rect 8665 9463 8723 9469
rect 6638 9392 6644 9444
rect 6696 9392 6702 9444
rect 8680 9432 8708 9463
rect 8846 9460 8852 9472
rect 8904 9460 8910 9512
rect 9306 9460 9312 9512
rect 9364 9500 9370 9512
rect 11606 9500 11612 9512
rect 9364 9472 11612 9500
rect 9364 9460 9370 9472
rect 11606 9460 11612 9472
rect 11664 9460 11670 9512
rect 8220 9404 8708 9432
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 6104 9336 6561 9364
rect 5629 9327 5687 9333
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6656 9364 6684 9392
rect 6825 9367 6883 9373
rect 6825 9364 6837 9367
rect 6656 9336 6837 9364
rect 6549 9327 6607 9333
rect 6825 9333 6837 9336
rect 6871 9364 6883 9367
rect 7834 9364 7840 9376
rect 6871 9336 7840 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7834 9324 7840 9336
rect 7892 9324 7898 9376
rect 8018 9324 8024 9376
rect 8076 9364 8082 9376
rect 8220 9364 8248 9404
rect 8754 9392 8760 9444
rect 8812 9432 8818 9444
rect 9858 9432 9864 9444
rect 8812 9404 9864 9432
rect 8812 9392 8818 9404
rect 9858 9392 9864 9404
rect 9916 9392 9922 9444
rect 8076 9336 8248 9364
rect 8076 9324 8082 9336
rect 8294 9324 8300 9376
rect 8352 9364 8358 9376
rect 9401 9367 9459 9373
rect 9401 9364 9413 9367
rect 8352 9336 9413 9364
rect 8352 9324 8358 9336
rect 9401 9333 9413 9336
rect 9447 9333 9459 9367
rect 9401 9327 9459 9333
rect 9677 9367 9735 9373
rect 9677 9333 9689 9367
rect 9723 9364 9735 9367
rect 10226 9364 10232 9376
rect 9723 9336 10232 9364
rect 9723 9333 9735 9336
rect 9677 9327 9735 9333
rect 10226 9324 10232 9336
rect 10284 9324 10290 9376
rect 1104 9274 16008 9296
rect 1104 9222 2824 9274
rect 2876 9222 2888 9274
rect 2940 9222 2952 9274
rect 3004 9222 3016 9274
rect 3068 9222 3080 9274
rect 3132 9222 6572 9274
rect 6624 9222 6636 9274
rect 6688 9222 6700 9274
rect 6752 9222 6764 9274
rect 6816 9222 6828 9274
rect 6880 9222 10320 9274
rect 10372 9222 10384 9274
rect 10436 9222 10448 9274
rect 10500 9222 10512 9274
rect 10564 9222 10576 9274
rect 10628 9222 14068 9274
rect 14120 9222 14132 9274
rect 14184 9222 14196 9274
rect 14248 9222 14260 9274
rect 14312 9222 14324 9274
rect 14376 9222 16008 9274
rect 1104 9200 16008 9222
rect 3602 9120 3608 9172
rect 3660 9160 3666 9172
rect 6089 9163 6147 9169
rect 6089 9160 6101 9163
rect 3660 9132 6101 9160
rect 3660 9120 3666 9132
rect 6089 9129 6101 9132
rect 6135 9129 6147 9163
rect 6089 9123 6147 9129
rect 7009 9163 7067 9169
rect 7009 9129 7021 9163
rect 7055 9160 7067 9163
rect 7282 9160 7288 9172
rect 7055 9132 7288 9160
rect 7055 9129 7067 9132
rect 7009 9123 7067 9129
rect 7282 9120 7288 9132
rect 7340 9120 7346 9172
rect 7466 9120 7472 9172
rect 7524 9160 7530 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 7524 9132 8953 9160
rect 7524 9120 7530 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 8478 9092 8484 9104
rect 8391 9064 8484 9092
rect 8478 9052 8484 9064
rect 8536 9092 8542 9104
rect 8536 9064 9536 9092
rect 8536 9052 8542 9064
rect 9508 9036 9536 9064
rect 5810 8984 5816 9036
rect 5868 9024 5874 9036
rect 5868 8996 7236 9024
rect 5868 8984 5874 8996
rect 6273 8959 6331 8965
rect 6273 8925 6285 8959
rect 6319 8925 6331 8959
rect 6273 8919 6331 8925
rect 6288 8888 6316 8919
rect 6362 8916 6368 8968
rect 6420 8956 6426 8968
rect 6420 8928 6465 8956
rect 6420 8916 6426 8928
rect 7006 8916 7012 8968
rect 7064 8956 7070 8968
rect 7101 8959 7159 8965
rect 7101 8956 7113 8959
rect 7064 8928 7113 8956
rect 7064 8916 7070 8928
rect 7101 8925 7113 8928
rect 7147 8925 7159 8959
rect 7208 8956 7236 8996
rect 9030 8984 9036 9036
rect 9088 9024 9094 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 9088 8996 9413 9024
rect 9088 8984 9094 8996
rect 9401 8993 9413 8996
rect 9447 8993 9459 9027
rect 9401 8987 9459 8993
rect 9490 8984 9496 9036
rect 9548 9024 9554 9036
rect 9548 8996 9593 9024
rect 9548 8984 9554 8996
rect 8757 8959 8815 8965
rect 7208 8928 8708 8956
rect 7101 8919 7159 8925
rect 6914 8888 6920 8900
rect 6288 8860 6920 8888
rect 6914 8848 6920 8860
rect 6972 8848 6978 8900
rect 7368 8891 7426 8897
rect 7368 8857 7380 8891
rect 7414 8888 7426 8891
rect 8018 8888 8024 8900
rect 7414 8860 8024 8888
rect 7414 8857 7426 8860
rect 7368 8851 7426 8857
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 8680 8888 8708 8928
rect 8757 8925 8769 8959
rect 8803 8956 8815 8959
rect 12066 8956 12072 8968
rect 8803 8928 12072 8956
rect 8803 8925 8815 8928
rect 8757 8919 8815 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 9398 8888 9404 8900
rect 8680 8860 9404 8888
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 8573 8823 8631 8829
rect 8573 8820 8585 8823
rect 4580 8792 8585 8820
rect 4580 8780 4586 8792
rect 8573 8789 8585 8792
rect 8619 8789 8631 8823
rect 8573 8783 8631 8789
rect 9309 8823 9367 8829
rect 9309 8789 9321 8823
rect 9355 8820 9367 8823
rect 9858 8820 9864 8832
rect 9355 8792 9864 8820
rect 9355 8789 9367 8792
rect 9309 8783 9367 8789
rect 9858 8780 9864 8792
rect 9916 8820 9922 8832
rect 10778 8820 10784 8832
rect 9916 8792 10784 8820
rect 9916 8780 9922 8792
rect 10778 8780 10784 8792
rect 10836 8780 10842 8832
rect 1104 8730 16008 8752
rect 1104 8678 4698 8730
rect 4750 8678 4762 8730
rect 4814 8678 4826 8730
rect 4878 8678 4890 8730
rect 4942 8678 4954 8730
rect 5006 8678 8446 8730
rect 8498 8678 8510 8730
rect 8562 8678 8574 8730
rect 8626 8678 8638 8730
rect 8690 8678 8702 8730
rect 8754 8678 12194 8730
rect 12246 8678 12258 8730
rect 12310 8678 12322 8730
rect 12374 8678 12386 8730
rect 12438 8678 12450 8730
rect 12502 8678 16008 8730
rect 1104 8656 16008 8678
rect 6362 8576 6368 8628
rect 6420 8616 6426 8628
rect 6733 8619 6791 8625
rect 6733 8616 6745 8619
rect 6420 8588 6745 8616
rect 6420 8576 6426 8588
rect 6733 8585 6745 8588
rect 6779 8585 6791 8619
rect 8846 8616 8852 8628
rect 6733 8579 6791 8585
rect 6886 8588 8852 8616
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 3326 8480 3332 8492
rect 1719 8452 3332 8480
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3142 8372 3148 8424
rect 3200 8412 3206 8424
rect 3418 8412 3424 8424
rect 3200 8384 3424 8412
rect 3200 8372 3206 8384
rect 3418 8372 3424 8384
rect 3476 8372 3482 8424
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 6086 8304 6092 8356
rect 6144 8344 6150 8356
rect 6886 8344 6914 8588
rect 8846 8576 8852 8588
rect 8904 8576 8910 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10686 8616 10692 8628
rect 9916 8588 10692 8616
rect 9916 8576 9922 8588
rect 10686 8576 10692 8588
rect 10744 8576 10750 8628
rect 7834 8508 7840 8560
rect 7892 8557 7898 8560
rect 7892 8548 7904 8557
rect 7892 8520 7937 8548
rect 7892 8511 7904 8520
rect 7892 8508 7898 8511
rect 9674 8508 9680 8560
rect 9732 8548 9738 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 9732 8520 11805 8548
rect 9732 8508 9738 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 11793 8511 11851 8517
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 8113 8483 8171 8489
rect 7156 8452 8064 8480
rect 7156 8440 7162 8452
rect 8036 8412 8064 8452
rect 8113 8449 8125 8483
rect 8159 8480 8171 8483
rect 8202 8480 8208 8492
rect 8159 8452 8208 8480
rect 8159 8449 8171 8452
rect 8113 8443 8171 8449
rect 8202 8440 8208 8452
rect 8260 8440 8266 8492
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8480 12679 8483
rect 12667 8452 12848 8480
rect 12667 8449 12679 8452
rect 12621 8443 12679 8449
rect 12526 8412 12532 8424
rect 8036 8384 12532 8412
rect 12526 8372 12532 8384
rect 12584 8372 12590 8424
rect 12820 8356 12848 8452
rect 12802 8344 12808 8356
rect 6144 8316 6914 8344
rect 12763 8316 12808 8344
rect 6144 8304 6150 8316
rect 12802 8304 12808 8316
rect 12860 8304 12866 8356
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 8202 8276 8208 8288
rect 7064 8248 8208 8276
rect 7064 8236 7070 8248
rect 8202 8236 8208 8248
rect 8260 8236 8266 8288
rect 1104 8186 16008 8208
rect 1104 8134 2824 8186
rect 2876 8134 2888 8186
rect 2940 8134 2952 8186
rect 3004 8134 3016 8186
rect 3068 8134 3080 8186
rect 3132 8134 6572 8186
rect 6624 8134 6636 8186
rect 6688 8134 6700 8186
rect 6752 8134 6764 8186
rect 6816 8134 6828 8186
rect 6880 8134 10320 8186
rect 10372 8134 10384 8186
rect 10436 8134 10448 8186
rect 10500 8134 10512 8186
rect 10564 8134 10576 8186
rect 10628 8134 14068 8186
rect 14120 8134 14132 8186
rect 14184 8134 14196 8186
rect 14248 8134 14260 8186
rect 14312 8134 14324 8186
rect 14376 8134 16008 8186
rect 1104 8112 16008 8134
rect 7190 8072 7196 8084
rect 7151 8044 7196 8072
rect 7190 8032 7196 8044
rect 7248 8032 7254 8084
rect 7558 8032 7564 8084
rect 7616 8072 7622 8084
rect 8202 8072 8208 8084
rect 7616 8044 8208 8072
rect 7616 8032 7622 8044
rect 8202 8032 8208 8044
rect 8260 8032 8266 8084
rect 7006 7936 7012 7948
rect 6967 7908 7012 7936
rect 7006 7896 7012 7908
rect 7064 7896 7070 7948
rect 7834 7936 7840 7948
rect 7795 7908 7840 7936
rect 7834 7896 7840 7908
rect 7892 7896 7898 7948
rect 5258 7868 5264 7880
rect 5219 7840 5264 7868
rect 5258 7828 5264 7840
rect 5316 7828 5322 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 9214 7868 9220 7880
rect 7699 7840 9220 7868
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 9214 7828 9220 7840
rect 9272 7828 9278 7880
rect 7561 7803 7619 7809
rect 7561 7769 7573 7803
rect 7607 7800 7619 7803
rect 7926 7800 7932 7812
rect 7607 7772 7932 7800
rect 7607 7769 7619 7772
rect 7561 7763 7619 7769
rect 7926 7760 7932 7772
rect 7984 7760 7990 7812
rect 1104 7642 16008 7664
rect 1104 7590 4698 7642
rect 4750 7590 4762 7642
rect 4814 7590 4826 7642
rect 4878 7590 4890 7642
rect 4942 7590 4954 7642
rect 5006 7590 8446 7642
rect 8498 7590 8510 7642
rect 8562 7590 8574 7642
rect 8626 7590 8638 7642
rect 8690 7590 8702 7642
rect 8754 7590 12194 7642
rect 12246 7590 12258 7642
rect 12310 7590 12322 7642
rect 12374 7590 12386 7642
rect 12438 7590 12450 7642
rect 12502 7590 16008 7642
rect 1104 7568 16008 7590
rect 9122 7528 9128 7540
rect 4172 7500 9128 7528
rect 4172 7401 4200 7500
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 10134 7460 10140 7472
rect 4724 7432 10140 7460
rect 4724 7401 4752 7432
rect 10134 7420 10140 7432
rect 10192 7420 10198 7472
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4709 7395 4767 7401
rect 4709 7361 4721 7395
rect 4755 7361 4767 7395
rect 4709 7355 4767 7361
rect 5261 7395 5319 7401
rect 5261 7361 5273 7395
rect 5307 7392 5319 7395
rect 5442 7392 5448 7404
rect 5307 7364 5448 7392
rect 5307 7361 5319 7364
rect 5261 7355 5319 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 7285 7395 7343 7401
rect 7285 7361 7297 7395
rect 7331 7392 7343 7395
rect 8938 7392 8944 7404
rect 7331 7364 8944 7392
rect 7331 7361 7343 7364
rect 7285 7355 7343 7361
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9306 7352 9312 7404
rect 9364 7392 9370 7404
rect 9401 7395 9459 7401
rect 9401 7392 9413 7395
rect 9364 7364 9413 7392
rect 9364 7352 9370 7364
rect 9401 7361 9413 7364
rect 9447 7361 9459 7395
rect 9401 7355 9459 7361
rect 3602 7216 3608 7268
rect 3660 7256 3666 7268
rect 5077 7259 5135 7265
rect 5077 7256 5089 7259
rect 3660 7228 5089 7256
rect 3660 7216 3666 7228
rect 5077 7225 5089 7228
rect 5123 7225 5135 7259
rect 5077 7219 5135 7225
rect 3970 7188 3976 7200
rect 3931 7160 3976 7188
rect 3970 7148 3976 7160
rect 4028 7148 4034 7200
rect 4522 7188 4528 7200
rect 4483 7160 4528 7188
rect 4522 7148 4528 7160
rect 4580 7148 4586 7200
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 7101 7191 7159 7197
rect 7101 7188 7113 7191
rect 5684 7160 7113 7188
rect 5684 7148 5690 7160
rect 7101 7157 7113 7160
rect 7147 7157 7159 7191
rect 7101 7151 7159 7157
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9217 7191 9275 7197
rect 9217 7188 9229 7191
rect 9088 7160 9229 7188
rect 9088 7148 9094 7160
rect 9217 7157 9229 7160
rect 9263 7157 9275 7191
rect 9217 7151 9275 7157
rect 1104 7098 16008 7120
rect 1104 7046 2824 7098
rect 2876 7046 2888 7098
rect 2940 7046 2952 7098
rect 3004 7046 3016 7098
rect 3068 7046 3080 7098
rect 3132 7046 6572 7098
rect 6624 7046 6636 7098
rect 6688 7046 6700 7098
rect 6752 7046 6764 7098
rect 6816 7046 6828 7098
rect 6880 7046 10320 7098
rect 10372 7046 10384 7098
rect 10436 7046 10448 7098
rect 10500 7046 10512 7098
rect 10564 7046 10576 7098
rect 10628 7046 14068 7098
rect 14120 7046 14132 7098
rect 14184 7046 14196 7098
rect 14248 7046 14260 7098
rect 14312 7046 14324 7098
rect 14376 7046 16008 7098
rect 1104 7024 16008 7046
rect 3142 6780 3148 6792
rect 3103 6752 3148 6780
rect 3142 6740 3148 6752
rect 3200 6740 3206 6792
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3142 6644 3148 6656
rect 3007 6616 3148 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 3142 6604 3148 6616
rect 3200 6604 3206 6656
rect 1104 6554 16008 6576
rect 1104 6502 4698 6554
rect 4750 6502 4762 6554
rect 4814 6502 4826 6554
rect 4878 6502 4890 6554
rect 4942 6502 4954 6554
rect 5006 6502 8446 6554
rect 8498 6502 8510 6554
rect 8562 6502 8574 6554
rect 8626 6502 8638 6554
rect 8690 6502 8702 6554
rect 8754 6502 12194 6554
rect 12246 6502 12258 6554
rect 12310 6502 12322 6554
rect 12374 6502 12386 6554
rect 12438 6502 12450 6554
rect 12502 6502 16008 6554
rect 1104 6480 16008 6502
rect 1104 6010 16008 6032
rect 1104 5958 2824 6010
rect 2876 5958 2888 6010
rect 2940 5958 2952 6010
rect 3004 5958 3016 6010
rect 3068 5958 3080 6010
rect 3132 5958 6572 6010
rect 6624 5958 6636 6010
rect 6688 5958 6700 6010
rect 6752 5958 6764 6010
rect 6816 5958 6828 6010
rect 6880 5958 10320 6010
rect 10372 5958 10384 6010
rect 10436 5958 10448 6010
rect 10500 5958 10512 6010
rect 10564 5958 10576 6010
rect 10628 5958 14068 6010
rect 14120 5958 14132 6010
rect 14184 5958 14196 6010
rect 14248 5958 14260 6010
rect 14312 5958 14324 6010
rect 14376 5958 16008 6010
rect 1104 5936 16008 5958
rect 1104 5466 16008 5488
rect 1104 5414 4698 5466
rect 4750 5414 4762 5466
rect 4814 5414 4826 5466
rect 4878 5414 4890 5466
rect 4942 5414 4954 5466
rect 5006 5414 8446 5466
rect 8498 5414 8510 5466
rect 8562 5414 8574 5466
rect 8626 5414 8638 5466
rect 8690 5414 8702 5466
rect 8754 5414 12194 5466
rect 12246 5414 12258 5466
rect 12310 5414 12322 5466
rect 12374 5414 12386 5466
rect 12438 5414 12450 5466
rect 12502 5414 16008 5466
rect 1104 5392 16008 5414
rect 1673 5219 1731 5225
rect 1673 5185 1685 5219
rect 1719 5216 1731 5219
rect 3142 5216 3148 5228
rect 1719 5188 3148 5216
rect 1719 5185 1731 5188
rect 1673 5179 1731 5185
rect 3142 5176 3148 5188
rect 3200 5176 3206 5228
rect 1486 5012 1492 5024
rect 1447 4984 1492 5012
rect 1486 4972 1492 4984
rect 1544 4972 1550 5024
rect 1104 4922 16008 4944
rect 1104 4870 2824 4922
rect 2876 4870 2888 4922
rect 2940 4870 2952 4922
rect 3004 4870 3016 4922
rect 3068 4870 3080 4922
rect 3132 4870 6572 4922
rect 6624 4870 6636 4922
rect 6688 4870 6700 4922
rect 6752 4870 6764 4922
rect 6816 4870 6828 4922
rect 6880 4870 10320 4922
rect 10372 4870 10384 4922
rect 10436 4870 10448 4922
rect 10500 4870 10512 4922
rect 10564 4870 10576 4922
rect 10628 4870 14068 4922
rect 14120 4870 14132 4922
rect 14184 4870 14196 4922
rect 14248 4870 14260 4922
rect 14312 4870 14324 4922
rect 14376 4870 16008 4922
rect 1104 4848 16008 4870
rect 1104 4378 16008 4400
rect 1104 4326 4698 4378
rect 4750 4326 4762 4378
rect 4814 4326 4826 4378
rect 4878 4326 4890 4378
rect 4942 4326 4954 4378
rect 5006 4326 8446 4378
rect 8498 4326 8510 4378
rect 8562 4326 8574 4378
rect 8626 4326 8638 4378
rect 8690 4326 8702 4378
rect 8754 4326 12194 4378
rect 12246 4326 12258 4378
rect 12310 4326 12322 4378
rect 12374 4326 12386 4378
rect 12438 4326 12450 4378
rect 12502 4326 16008 4378
rect 1104 4304 16008 4326
rect 1104 3834 16008 3856
rect 1104 3782 2824 3834
rect 2876 3782 2888 3834
rect 2940 3782 2952 3834
rect 3004 3782 3016 3834
rect 3068 3782 3080 3834
rect 3132 3782 6572 3834
rect 6624 3782 6636 3834
rect 6688 3782 6700 3834
rect 6752 3782 6764 3834
rect 6816 3782 6828 3834
rect 6880 3782 10320 3834
rect 10372 3782 10384 3834
rect 10436 3782 10448 3834
rect 10500 3782 10512 3834
rect 10564 3782 10576 3834
rect 10628 3782 14068 3834
rect 14120 3782 14132 3834
rect 14184 3782 14196 3834
rect 14248 3782 14260 3834
rect 14312 3782 14324 3834
rect 14376 3782 16008 3834
rect 1104 3760 16008 3782
rect 13814 3680 13820 3732
rect 13872 3720 13878 3732
rect 15473 3723 15531 3729
rect 15473 3720 15485 3723
rect 13872 3692 15485 3720
rect 13872 3680 13878 3692
rect 15473 3689 15485 3692
rect 15519 3689 15531 3723
rect 15473 3683 15531 3689
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3516 1731 3519
rect 4522 3516 4528 3528
rect 1719 3488 4528 3516
rect 1719 3485 1731 3488
rect 1673 3479 1731 3485
rect 4522 3476 4528 3488
rect 4580 3476 4586 3528
rect 15105 3519 15163 3525
rect 15105 3485 15117 3519
rect 15151 3516 15163 3519
rect 15657 3519 15715 3525
rect 15657 3516 15669 3519
rect 15151 3488 15669 3516
rect 15151 3485 15163 3488
rect 15105 3479 15163 3485
rect 15657 3485 15669 3488
rect 15703 3516 15715 3519
rect 16942 3516 16948 3528
rect 15703 3488 16948 3516
rect 15703 3485 15715 3488
rect 15657 3479 15715 3485
rect 16942 3476 16948 3488
rect 17000 3476 17006 3528
rect 14921 3451 14979 3457
rect 14921 3417 14933 3451
rect 14967 3448 14979 3451
rect 14967 3420 15700 3448
rect 14967 3417 14979 3420
rect 14921 3411 14979 3417
rect 15672 3392 15700 3420
rect 1026 3340 1032 3392
rect 1084 3380 1090 3392
rect 1489 3383 1547 3389
rect 1489 3380 1501 3383
rect 1084 3352 1501 3380
rect 1084 3340 1090 3352
rect 1489 3349 1501 3352
rect 1535 3349 1547 3383
rect 15286 3380 15292 3392
rect 15247 3352 15292 3380
rect 1489 3343 1547 3349
rect 15286 3340 15292 3352
rect 15344 3340 15350 3392
rect 15654 3340 15660 3392
rect 15712 3340 15718 3392
rect 1104 3290 16008 3312
rect 1104 3238 4698 3290
rect 4750 3238 4762 3290
rect 4814 3238 4826 3290
rect 4878 3238 4890 3290
rect 4942 3238 4954 3290
rect 5006 3238 8446 3290
rect 8498 3238 8510 3290
rect 8562 3238 8574 3290
rect 8626 3238 8638 3290
rect 8690 3238 8702 3290
rect 8754 3238 12194 3290
rect 12246 3238 12258 3290
rect 12310 3238 12322 3290
rect 12374 3238 12386 3290
rect 12438 3238 12450 3290
rect 12502 3238 16008 3290
rect 1104 3216 16008 3238
rect 2317 3179 2375 3185
rect 2317 3145 2329 3179
rect 2363 3176 2375 3179
rect 3234 3176 3240 3188
rect 2363 3148 3240 3176
rect 2363 3145 2375 3148
rect 2317 3139 2375 3145
rect 3234 3136 3240 3148
rect 3292 3136 3298 3188
rect 14918 3176 14924 3188
rect 14879 3148 14924 3176
rect 14918 3136 14924 3148
rect 14976 3136 14982 3188
rect 15197 3179 15255 3185
rect 15197 3145 15209 3179
rect 15243 3145 15255 3179
rect 15197 3139 15255 3145
rect 3970 3108 3976 3120
rect 1688 3080 3976 3108
rect 1688 3049 1716 3080
rect 3970 3068 3976 3080
rect 4028 3068 4034 3120
rect 14734 3068 14740 3120
rect 14792 3108 14798 3120
rect 15212 3108 15240 3139
rect 14792 3080 15240 3108
rect 14792 3068 14798 3080
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 2038 3040 2044 3052
rect 1999 3012 2044 3040
rect 1673 3003 1731 3009
rect 2038 3000 2044 3012
rect 2096 3000 2102 3052
rect 2130 3000 2136 3052
rect 2188 3040 2194 3052
rect 2409 3043 2467 3049
rect 2409 3040 2421 3043
rect 2188 3012 2421 3040
rect 2188 3000 2194 3012
rect 2409 3009 2421 3012
rect 2455 3009 2467 3043
rect 2409 3003 2467 3009
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 15105 3043 15163 3049
rect 14599 3012 15056 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 9582 2932 9588 2984
rect 9640 2972 9646 2984
rect 9640 2944 14872 2972
rect 9640 2932 9646 2944
rect 566 2864 572 2916
rect 624 2904 630 2916
rect 1857 2907 1915 2913
rect 1857 2904 1869 2907
rect 624 2876 1869 2904
rect 624 2864 630 2876
rect 1857 2873 1869 2876
rect 1903 2873 1915 2907
rect 1857 2867 1915 2873
rect 198 2796 204 2848
rect 256 2836 262 2848
rect 1489 2839 1547 2845
rect 1489 2836 1501 2839
rect 256 2808 1501 2836
rect 256 2796 262 2808
rect 1489 2805 1501 2808
rect 1535 2805 1547 2839
rect 8754 2836 8760 2848
rect 8715 2808 8760 2836
rect 1489 2799 1547 2805
rect 8754 2796 8760 2808
rect 8812 2796 8818 2848
rect 9214 2836 9220 2848
rect 9175 2808 9220 2836
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 10870 2836 10876 2848
rect 10831 2808 10876 2836
rect 10870 2796 10876 2808
rect 10928 2796 10934 2848
rect 11330 2796 11336 2848
rect 11388 2836 11394 2848
rect 11517 2839 11575 2845
rect 11517 2836 11529 2839
rect 11388 2808 11529 2836
rect 11388 2796 11394 2808
rect 11517 2805 11529 2808
rect 11563 2805 11575 2839
rect 11517 2799 11575 2805
rect 12161 2839 12219 2845
rect 12161 2805 12173 2839
rect 12207 2836 12219 2839
rect 12526 2836 12532 2848
rect 12207 2808 12532 2836
rect 12207 2805 12219 2808
rect 12161 2799 12219 2805
rect 12526 2796 12532 2808
rect 12584 2796 12590 2848
rect 13446 2836 13452 2848
rect 13407 2808 13452 2836
rect 13446 2796 13452 2808
rect 13504 2796 13510 2848
rect 13906 2836 13912 2848
rect 13867 2808 13912 2836
rect 13906 2796 13912 2808
rect 13964 2796 13970 2848
rect 14734 2836 14740 2848
rect 14695 2808 14740 2836
rect 14734 2796 14740 2808
rect 14792 2796 14798 2848
rect 14844 2836 14872 2944
rect 15028 2904 15056 3012
rect 15105 3009 15117 3043
rect 15151 3009 15163 3043
rect 15378 3040 15384 3052
rect 15339 3012 15384 3040
rect 15105 3003 15163 3009
rect 15120 2972 15148 3003
rect 15378 3000 15384 3012
rect 15436 3000 15442 3052
rect 15654 3040 15660 3052
rect 15615 3012 15660 3040
rect 15654 3000 15660 3012
rect 15712 3000 15718 3052
rect 15286 2972 15292 2984
rect 15120 2944 15292 2972
rect 15286 2932 15292 2944
rect 15344 2972 15350 2984
rect 16482 2972 16488 2984
rect 15344 2944 16488 2972
rect 15344 2932 15350 2944
rect 16482 2932 16488 2944
rect 16540 2932 16546 2984
rect 15194 2904 15200 2916
rect 15028 2876 15200 2904
rect 15194 2864 15200 2876
rect 15252 2864 15258 2916
rect 15473 2839 15531 2845
rect 15473 2836 15485 2839
rect 14844 2808 15485 2836
rect 15473 2805 15485 2808
rect 15519 2805 15531 2839
rect 15473 2799 15531 2805
rect 1104 2746 16008 2768
rect 1104 2694 2824 2746
rect 2876 2694 2888 2746
rect 2940 2694 2952 2746
rect 3004 2694 3016 2746
rect 3068 2694 3080 2746
rect 3132 2694 6572 2746
rect 6624 2694 6636 2746
rect 6688 2694 6700 2746
rect 6752 2694 6764 2746
rect 6816 2694 6828 2746
rect 6880 2694 10320 2746
rect 10372 2694 10384 2746
rect 10436 2694 10448 2746
rect 10500 2694 10512 2746
rect 10564 2694 10576 2746
rect 10628 2694 14068 2746
rect 14120 2694 14132 2746
rect 14184 2694 14196 2746
rect 14248 2694 14260 2746
rect 14312 2694 14324 2746
rect 14376 2694 16008 2746
rect 1104 2672 16008 2694
rect 5074 2632 5080 2644
rect 1872 2604 5080 2632
rect 1872 2437 1900 2604
rect 5074 2592 5080 2604
rect 5132 2592 5138 2644
rect 5258 2592 5264 2644
rect 5316 2632 5322 2644
rect 8294 2632 8300 2644
rect 5316 2604 8300 2632
rect 5316 2592 5322 2604
rect 8294 2592 8300 2604
rect 8352 2592 8358 2644
rect 8846 2592 8852 2644
rect 8904 2632 8910 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8904 2604 8953 2632
rect 8904 2592 8910 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 9858 2632 9864 2644
rect 9819 2604 9864 2632
rect 8941 2595 8999 2601
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 12066 2592 12072 2644
rect 12124 2632 12130 2644
rect 12713 2635 12771 2641
rect 12713 2632 12725 2635
rect 12124 2604 12725 2632
rect 12124 2592 12130 2604
rect 12713 2601 12725 2604
rect 12759 2601 12771 2635
rect 12713 2595 12771 2601
rect 13630 2592 13636 2644
rect 13688 2632 13694 2644
rect 14829 2635 14887 2641
rect 14829 2632 14841 2635
rect 13688 2604 14841 2632
rect 13688 2592 13694 2604
rect 14829 2601 14841 2604
rect 14875 2601 14887 2635
rect 14829 2595 14887 2601
rect 3602 2564 3608 2576
rect 2240 2536 3608 2564
rect 2240 2437 2268 2536
rect 3602 2524 3608 2536
rect 3660 2524 3666 2576
rect 5626 2564 5632 2576
rect 4816 2536 5632 2564
rect 4154 2496 4160 2508
rect 3160 2468 4160 2496
rect 1857 2431 1915 2437
rect 1857 2397 1869 2431
rect 1903 2397 1915 2431
rect 1857 2391 1915 2397
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2682 2428 2688 2440
rect 2643 2400 2688 2428
rect 2225 2391 2283 2397
rect 2682 2388 2688 2400
rect 2740 2388 2746 2440
rect 3160 2437 3188 2468
rect 4154 2456 4160 2468
rect 4212 2456 4218 2508
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2397 3203 2431
rect 3145 2391 3203 2397
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 4065 2431 4123 2437
rect 4065 2397 4077 2431
rect 4111 2428 4123 2431
rect 4246 2428 4252 2440
rect 4111 2400 4252 2428
rect 4111 2397 4123 2400
rect 4065 2391 4123 2397
rect 3528 2360 3556 2391
rect 4246 2388 4252 2400
rect 4304 2388 4310 2440
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 4614 2428 4620 2440
rect 4479 2400 4620 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4816 2437 4844 2536
rect 5626 2524 5632 2536
rect 5684 2524 5690 2576
rect 6886 2536 9168 2564
rect 6886 2496 6914 2536
rect 9030 2496 9036 2508
rect 5736 2468 6914 2496
rect 7392 2468 9036 2496
rect 5258 2437 5264 2440
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5254 2391 5264 2437
rect 5316 2428 5322 2440
rect 5736 2437 5764 2468
rect 5721 2431 5779 2437
rect 5316 2400 5354 2428
rect 5258 2388 5264 2391
rect 5316 2388 5322 2400
rect 5721 2397 5733 2431
rect 5767 2397 5779 2431
rect 6086 2428 6092 2440
rect 6047 2400 6092 2428
rect 5721 2391 5779 2397
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 6638 2428 6644 2440
rect 6599 2400 6644 2428
rect 6638 2388 6644 2400
rect 6696 2388 6702 2440
rect 7009 2431 7067 2437
rect 7009 2397 7021 2431
rect 7055 2428 7067 2431
rect 7282 2428 7288 2440
rect 7055 2400 7288 2428
rect 7055 2397 7067 2400
rect 7009 2391 7067 2397
rect 7282 2388 7288 2400
rect 7340 2388 7346 2440
rect 7392 2437 7420 2468
rect 9030 2456 9036 2468
rect 9088 2456 9094 2508
rect 9140 2496 9168 2536
rect 9398 2524 9404 2576
rect 9456 2564 9462 2576
rect 10137 2567 10195 2573
rect 10137 2564 10149 2567
rect 9456 2536 10149 2564
rect 9456 2524 9462 2536
rect 10137 2533 10149 2536
rect 10183 2533 10195 2567
rect 10137 2527 10195 2533
rect 10778 2524 10784 2576
rect 10836 2564 10842 2576
rect 13173 2567 13231 2573
rect 13173 2564 13185 2567
rect 10836 2536 13185 2564
rect 10836 2524 10842 2536
rect 13173 2533 13185 2536
rect 13219 2533 13231 2567
rect 13173 2527 13231 2533
rect 13262 2524 13268 2576
rect 13320 2564 13326 2576
rect 13541 2567 13599 2573
rect 13541 2564 13553 2567
rect 13320 2536 13553 2564
rect 13320 2524 13326 2536
rect 13541 2533 13553 2536
rect 13587 2533 13599 2567
rect 13541 2527 13599 2533
rect 9858 2496 9864 2508
rect 9140 2468 9864 2496
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 12621 2499 12679 2505
rect 12621 2496 12633 2499
rect 12084 2468 12633 2496
rect 7377 2431 7435 2437
rect 7377 2397 7389 2431
rect 7423 2397 7435 2431
rect 7834 2428 7840 2440
rect 7795 2400 7840 2428
rect 7377 2391 7435 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 8297 2431 8355 2437
rect 8297 2397 8309 2431
rect 8343 2397 8355 2431
rect 8662 2428 8668 2440
rect 8623 2400 8668 2428
rect 8297 2391 8355 2397
rect 5994 2360 6000 2372
rect 3528 2332 6000 2360
rect 5994 2320 6000 2332
rect 6052 2320 6058 2372
rect 8312 2360 8340 2391
rect 8662 2388 8668 2400
rect 8720 2388 8726 2440
rect 8846 2388 8852 2440
rect 8904 2428 8910 2440
rect 9125 2431 9183 2437
rect 9125 2428 9137 2431
rect 8904 2400 9137 2428
rect 8904 2388 8910 2400
rect 9125 2397 9137 2400
rect 9171 2397 9183 2431
rect 9125 2391 9183 2397
rect 9214 2388 9220 2440
rect 9272 2428 9278 2440
rect 9493 2431 9551 2437
rect 9493 2428 9505 2431
rect 9272 2400 9505 2428
rect 9272 2388 9278 2400
rect 9493 2397 9505 2400
rect 9539 2397 9551 2431
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 9493 2391 9551 2397
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9732 2400 9965 2428
rect 9732 2388 9738 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 10321 2431 10379 2437
rect 10321 2397 10333 2431
rect 10367 2428 10379 2431
rect 10367 2400 10401 2428
rect 10367 2397 10379 2400
rect 10321 2391 10379 2397
rect 8312 2332 8892 2360
rect 1486 2252 1492 2304
rect 1544 2292 1550 2304
rect 1673 2295 1731 2301
rect 1673 2292 1685 2295
rect 1544 2264 1685 2292
rect 1544 2252 1550 2264
rect 1673 2261 1685 2264
rect 1719 2261 1731 2295
rect 1673 2255 1731 2261
rect 1854 2252 1860 2304
rect 1912 2292 1918 2304
rect 2041 2295 2099 2301
rect 2041 2292 2053 2295
rect 1912 2264 2053 2292
rect 1912 2252 1918 2264
rect 2041 2261 2053 2264
rect 2087 2261 2099 2295
rect 2041 2255 2099 2261
rect 2314 2252 2320 2304
rect 2372 2292 2378 2304
rect 2501 2295 2559 2301
rect 2501 2292 2513 2295
rect 2372 2264 2513 2292
rect 2372 2252 2378 2264
rect 2501 2261 2513 2264
rect 2547 2261 2559 2295
rect 2501 2255 2559 2261
rect 2774 2252 2780 2304
rect 2832 2292 2838 2304
rect 2961 2295 3019 2301
rect 2961 2292 2973 2295
rect 2832 2264 2973 2292
rect 2832 2252 2838 2264
rect 2961 2261 2973 2264
rect 3007 2261 3019 2295
rect 2961 2255 3019 2261
rect 3142 2252 3148 2304
rect 3200 2292 3206 2304
rect 3329 2295 3387 2301
rect 3329 2292 3341 2295
rect 3200 2264 3341 2292
rect 3200 2252 3206 2264
rect 3329 2261 3341 2264
rect 3375 2261 3387 2295
rect 3329 2255 3387 2261
rect 3602 2252 3608 2304
rect 3660 2292 3666 2304
rect 3881 2295 3939 2301
rect 3881 2292 3893 2295
rect 3660 2264 3893 2292
rect 3660 2252 3666 2264
rect 3881 2261 3893 2264
rect 3927 2261 3939 2295
rect 3881 2255 3939 2261
rect 4062 2252 4068 2304
rect 4120 2292 4126 2304
rect 4249 2295 4307 2301
rect 4249 2292 4261 2295
rect 4120 2264 4261 2292
rect 4120 2252 4126 2264
rect 4249 2261 4261 2264
rect 4295 2261 4307 2295
rect 4249 2255 4307 2261
rect 4430 2252 4436 2304
rect 4488 2292 4494 2304
rect 4617 2295 4675 2301
rect 4617 2292 4629 2295
rect 4488 2264 4629 2292
rect 4488 2252 4494 2264
rect 4617 2261 4629 2264
rect 4663 2261 4675 2295
rect 5074 2292 5080 2304
rect 5035 2264 5080 2292
rect 4617 2255 4675 2261
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 5350 2252 5356 2304
rect 5408 2292 5414 2304
rect 5537 2295 5595 2301
rect 5537 2292 5549 2295
rect 5408 2264 5549 2292
rect 5408 2252 5414 2264
rect 5537 2261 5549 2264
rect 5583 2261 5595 2295
rect 5537 2255 5595 2261
rect 5718 2252 5724 2304
rect 5776 2292 5782 2304
rect 5905 2295 5963 2301
rect 5905 2292 5917 2295
rect 5776 2264 5917 2292
rect 5776 2252 5782 2264
rect 5905 2261 5917 2264
rect 5951 2261 5963 2295
rect 5905 2255 5963 2261
rect 6178 2252 6184 2304
rect 6236 2292 6242 2304
rect 6457 2295 6515 2301
rect 6457 2292 6469 2295
rect 6236 2264 6469 2292
rect 6236 2252 6242 2264
rect 6457 2261 6469 2264
rect 6503 2261 6515 2295
rect 6457 2255 6515 2261
rect 6638 2252 6644 2304
rect 6696 2292 6702 2304
rect 6825 2295 6883 2301
rect 6825 2292 6837 2295
rect 6696 2264 6837 2292
rect 6696 2252 6702 2264
rect 6825 2261 6837 2264
rect 6871 2261 6883 2295
rect 6825 2255 6883 2261
rect 7006 2252 7012 2304
rect 7064 2292 7070 2304
rect 7193 2295 7251 2301
rect 7193 2292 7205 2295
rect 7064 2264 7205 2292
rect 7064 2252 7070 2264
rect 7193 2261 7205 2264
rect 7239 2261 7251 2295
rect 7193 2255 7251 2261
rect 7466 2252 7472 2304
rect 7524 2292 7530 2304
rect 7653 2295 7711 2301
rect 7653 2292 7665 2295
rect 7524 2264 7665 2292
rect 7524 2252 7530 2264
rect 7653 2261 7665 2264
rect 7699 2261 7711 2295
rect 7653 2255 7711 2261
rect 7926 2252 7932 2304
rect 7984 2292 7990 2304
rect 8113 2295 8171 2301
rect 8113 2292 8125 2295
rect 7984 2264 8125 2292
rect 7984 2252 7990 2264
rect 8113 2261 8125 2264
rect 8159 2261 8171 2295
rect 8113 2255 8171 2261
rect 8294 2252 8300 2304
rect 8352 2292 8358 2304
rect 8481 2295 8539 2301
rect 8481 2292 8493 2295
rect 8352 2264 8493 2292
rect 8352 2252 8358 2264
rect 8481 2261 8493 2264
rect 8527 2261 8539 2295
rect 8864 2292 8892 2332
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 8996 2332 9812 2360
rect 8996 2320 9002 2332
rect 9122 2292 9128 2304
rect 8864 2264 9128 2292
rect 8481 2255 8539 2261
rect 9122 2252 9128 2264
rect 9180 2252 9186 2304
rect 9306 2292 9312 2304
rect 9267 2264 9312 2292
rect 9306 2252 9312 2264
rect 9364 2252 9370 2304
rect 9784 2292 9812 2332
rect 10042 2320 10048 2372
rect 10100 2360 10106 2372
rect 10336 2360 10364 2391
rect 10502 2388 10508 2440
rect 10560 2428 10566 2440
rect 10781 2431 10839 2437
rect 10781 2428 10793 2431
rect 10560 2400 10793 2428
rect 10560 2388 10566 2400
rect 10781 2397 10793 2400
rect 10827 2397 10839 2431
rect 10781 2391 10839 2397
rect 10413 2363 10471 2369
rect 10413 2360 10425 2363
rect 10100 2332 10425 2360
rect 10100 2320 10106 2332
rect 10413 2329 10425 2332
rect 10459 2329 10471 2363
rect 10796 2360 10824 2391
rect 11054 2388 11060 2440
rect 11112 2428 11118 2440
rect 11149 2431 11207 2437
rect 11149 2428 11161 2431
rect 11112 2400 11161 2428
rect 11112 2388 11118 2400
rect 11149 2397 11161 2400
rect 11195 2397 11207 2431
rect 11149 2391 11207 2397
rect 11330 2388 11336 2440
rect 11388 2428 11394 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11388 2400 11713 2428
rect 11388 2388 11394 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 11701 2391 11759 2397
rect 11790 2388 11796 2440
rect 11848 2428 11854 2440
rect 12084 2437 12112 2468
rect 12621 2465 12633 2468
rect 12667 2465 12679 2499
rect 12621 2459 12679 2465
rect 12069 2431 12127 2437
rect 12069 2428 12081 2431
rect 11848 2400 12081 2428
rect 11848 2388 11854 2400
rect 12069 2397 12081 2400
rect 12115 2397 12127 2431
rect 12069 2391 12127 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12526 2428 12532 2440
rect 12483 2400 12532 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 12526 2388 12532 2400
rect 12584 2388 12590 2440
rect 12897 2431 12955 2437
rect 12897 2397 12909 2431
rect 12943 2428 12955 2431
rect 12943 2400 12977 2428
rect 12943 2397 12955 2400
rect 12897 2391 12955 2397
rect 11241 2363 11299 2369
rect 11241 2360 11253 2363
rect 10796 2332 11253 2360
rect 10413 2323 10471 2329
rect 11241 2329 11253 2332
rect 11287 2329 11299 2363
rect 11241 2323 11299 2329
rect 11440 2332 12572 2360
rect 10597 2295 10655 2301
rect 10597 2292 10609 2295
rect 9784 2264 10609 2292
rect 10597 2261 10609 2264
rect 10643 2261 10655 2295
rect 10962 2292 10968 2304
rect 10923 2264 10968 2292
rect 10597 2255 10655 2261
rect 10962 2252 10968 2264
rect 11020 2252 11026 2304
rect 11146 2252 11152 2304
rect 11204 2292 11210 2304
rect 11440 2292 11468 2332
rect 11204 2264 11468 2292
rect 11204 2252 11210 2264
rect 11514 2252 11520 2304
rect 11572 2292 11578 2304
rect 11882 2292 11888 2304
rect 11572 2264 11617 2292
rect 11843 2264 11888 2292
rect 11572 2252 11578 2264
rect 11882 2252 11888 2264
rect 11940 2252 11946 2304
rect 12066 2252 12072 2304
rect 12124 2292 12130 2304
rect 12253 2295 12311 2301
rect 12253 2292 12265 2295
rect 12124 2264 12265 2292
rect 12124 2252 12130 2264
rect 12253 2261 12265 2264
rect 12299 2261 12311 2295
rect 12544 2292 12572 2332
rect 12618 2320 12624 2372
rect 12676 2360 12682 2372
rect 12912 2360 12940 2391
rect 13078 2388 13084 2440
rect 13136 2428 13142 2440
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 13136 2400 13369 2428
rect 13136 2388 13142 2400
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 12989 2363 13047 2369
rect 12989 2360 13001 2363
rect 12676 2332 13001 2360
rect 12676 2320 12682 2332
rect 12989 2329 13001 2332
rect 13035 2329 13047 2363
rect 13372 2360 13400 2391
rect 13446 2388 13452 2440
rect 13504 2428 13510 2440
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 13504 2400 13737 2428
rect 13504 2388 13510 2400
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 13906 2388 13912 2440
rect 13964 2428 13970 2440
rect 14277 2431 14335 2437
rect 14277 2428 14289 2431
rect 13964 2400 14289 2428
rect 13964 2388 13970 2400
rect 14277 2397 14289 2400
rect 14323 2397 14335 2431
rect 14277 2391 14335 2397
rect 14366 2388 14372 2440
rect 14424 2428 14430 2440
rect 14645 2431 14703 2437
rect 14645 2428 14657 2431
rect 14424 2400 14657 2428
rect 14424 2388 14430 2400
rect 14645 2397 14657 2400
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 13817 2363 13875 2369
rect 13817 2360 13829 2363
rect 13372 2332 13829 2360
rect 12989 2323 13047 2329
rect 13817 2329 13829 2332
rect 13863 2329 13875 2363
rect 14660 2360 14688 2391
rect 14734 2388 14740 2440
rect 14792 2428 14798 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14792 2400 15025 2428
rect 14792 2388 14798 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 15194 2388 15200 2440
rect 15252 2428 15258 2440
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 15252 2400 15485 2428
rect 15252 2388 15258 2400
rect 15473 2397 15485 2400
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 15105 2363 15163 2369
rect 15105 2360 15117 2363
rect 13817 2323 13875 2329
rect 13924 2332 14504 2360
rect 14660 2332 15117 2360
rect 13924 2292 13952 2332
rect 14090 2292 14096 2304
rect 12544 2264 13952 2292
rect 14051 2264 14096 2292
rect 12253 2255 12311 2261
rect 14090 2252 14096 2264
rect 14148 2252 14154 2304
rect 14476 2301 14504 2332
rect 15105 2329 15117 2332
rect 15151 2329 15163 2363
rect 15105 2323 15163 2329
rect 14461 2295 14519 2301
rect 14461 2261 14473 2295
rect 14507 2261 14519 2295
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 14461 2255 14519 2261
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 15378 2252 15384 2304
rect 15436 2292 15442 2304
rect 15657 2295 15715 2301
rect 15657 2292 15669 2295
rect 15436 2264 15669 2292
rect 15436 2252 15442 2264
rect 15657 2261 15669 2264
rect 15703 2292 15715 2295
rect 16022 2292 16028 2304
rect 15703 2264 16028 2292
rect 15703 2261 15715 2264
rect 15657 2255 15715 2261
rect 16022 2252 16028 2264
rect 16080 2252 16086 2304
rect 1104 2202 16008 2224
rect 1104 2150 4698 2202
rect 4750 2150 4762 2202
rect 4814 2150 4826 2202
rect 4878 2150 4890 2202
rect 4942 2150 4954 2202
rect 5006 2150 8446 2202
rect 8498 2150 8510 2202
rect 8562 2150 8574 2202
rect 8626 2150 8638 2202
rect 8690 2150 8702 2202
rect 8754 2150 12194 2202
rect 12246 2150 12258 2202
rect 12310 2150 12322 2202
rect 12374 2150 12386 2202
rect 12438 2150 12450 2202
rect 12502 2150 16008 2202
rect 1104 2128 16008 2150
rect 6086 2048 6092 2100
rect 6144 2088 6150 2100
rect 6144 2060 6914 2088
rect 6144 2048 6150 2060
rect 6886 1952 6914 2060
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 11422 2088 11428 2100
rect 7340 2060 11428 2088
rect 7340 2048 7346 2060
rect 11422 2048 11428 2060
rect 11480 2048 11486 2100
rect 11974 2048 11980 2100
rect 12032 2088 12038 2100
rect 15286 2088 15292 2100
rect 12032 2060 15292 2088
rect 12032 2048 12038 2060
rect 15286 2048 15292 2060
rect 15344 2048 15350 2100
rect 9122 1980 9128 2032
rect 9180 2020 9186 2032
rect 12710 2020 12716 2032
rect 9180 1992 12716 2020
rect 9180 1980 9186 1992
rect 12710 1980 12716 1992
rect 12768 1980 12774 2032
rect 10134 1952 10140 1964
rect 6886 1924 10140 1952
rect 10134 1912 10140 1924
rect 10192 1912 10198 1964
rect 7742 1844 7748 1896
rect 7800 1884 7806 1896
rect 11514 1884 11520 1896
rect 7800 1856 11520 1884
rect 7800 1844 7806 1856
rect 11514 1844 11520 1856
rect 11572 1844 11578 1896
rect 9766 1776 9772 1828
rect 9824 1816 9830 1828
rect 14090 1816 14096 1828
rect 9824 1788 14096 1816
rect 9824 1776 9830 1788
rect 14090 1776 14096 1788
rect 14148 1776 14154 1828
rect 6270 1708 6276 1760
rect 6328 1748 6334 1760
rect 10962 1748 10968 1760
rect 6328 1720 10968 1748
rect 6328 1708 6334 1720
rect 10962 1708 10968 1720
rect 11020 1708 11026 1760
rect 4522 1640 4528 1692
rect 4580 1680 4586 1692
rect 9306 1680 9312 1692
rect 4580 1652 9312 1680
rect 4580 1640 4586 1652
rect 9306 1640 9312 1652
rect 9364 1640 9370 1692
rect 6914 1572 6920 1624
rect 6972 1612 6978 1624
rect 11882 1612 11888 1624
rect 6972 1584 11888 1612
rect 6972 1572 6978 1584
rect 11882 1572 11888 1584
rect 11940 1572 11946 1624
<< via1 >>
rect 6184 17620 6236 17672
rect 10876 17620 10928 17672
rect 9312 17552 9364 17604
rect 13084 17552 13136 17604
rect 9220 17484 9272 17536
rect 13636 17484 13688 17536
rect 4698 17382 4750 17434
rect 4762 17382 4814 17434
rect 4826 17382 4878 17434
rect 4890 17382 4942 17434
rect 4954 17382 5006 17434
rect 8446 17382 8498 17434
rect 8510 17382 8562 17434
rect 8574 17382 8626 17434
rect 8638 17382 8690 17434
rect 8702 17382 8754 17434
rect 12194 17382 12246 17434
rect 12258 17382 12310 17434
rect 12322 17382 12374 17434
rect 12386 17382 12438 17434
rect 12450 17382 12502 17434
rect 1400 17280 1452 17332
rect 1860 17280 1912 17332
rect 2228 17280 2280 17332
rect 2688 17323 2740 17332
rect 2688 17289 2697 17323
rect 2697 17289 2731 17323
rect 2731 17289 2740 17323
rect 2688 17280 2740 17289
rect 3056 17323 3108 17332
rect 3056 17289 3065 17323
rect 3065 17289 3099 17323
rect 3099 17289 3108 17323
rect 3056 17280 3108 17289
rect 3516 17280 3568 17332
rect 4160 17323 4212 17332
rect 4160 17289 4169 17323
rect 4169 17289 4203 17323
rect 4203 17289 4212 17323
rect 4160 17280 4212 17289
rect 4344 17280 4396 17332
rect 4620 17280 4672 17332
rect 5172 17280 5224 17332
rect 5632 17323 5684 17332
rect 5632 17289 5641 17323
rect 5641 17289 5675 17323
rect 5675 17289 5684 17323
rect 5632 17280 5684 17289
rect 6000 17323 6052 17332
rect 6000 17289 6009 17323
rect 6009 17289 6043 17323
rect 6043 17289 6052 17323
rect 6000 17280 6052 17289
rect 6460 17280 6512 17332
rect 6920 17280 6972 17332
rect 7288 17280 7340 17332
rect 7748 17280 7800 17332
rect 8300 17323 8352 17332
rect 8300 17289 8309 17323
rect 8309 17289 8343 17323
rect 8343 17289 8352 17323
rect 8300 17280 8352 17289
rect 8852 17280 8904 17332
rect 9404 17323 9456 17332
rect 9404 17289 9413 17323
rect 9413 17289 9447 17323
rect 9447 17289 9456 17323
rect 9404 17280 9456 17289
rect 10232 17280 10284 17332
rect 3884 17212 3936 17264
rect 2136 17187 2188 17196
rect 2136 17153 2145 17187
rect 2145 17153 2179 17187
rect 2179 17153 2188 17187
rect 2136 17144 2188 17153
rect 3148 17144 3200 17196
rect 3424 17144 3476 17196
rect 3608 17187 3660 17196
rect 3608 17153 3617 17187
rect 3617 17153 3651 17187
rect 3651 17153 3660 17187
rect 3608 17144 3660 17153
rect 4528 17144 4580 17196
rect 3792 17076 3844 17128
rect 4436 17076 4488 17128
rect 5540 17144 5592 17196
rect 5816 17187 5868 17196
rect 5816 17153 5825 17187
rect 5825 17153 5859 17187
rect 5859 17153 5868 17187
rect 5816 17144 5868 17153
rect 6184 17187 6236 17196
rect 6184 17153 6193 17187
rect 6193 17153 6227 17187
rect 6227 17153 6236 17187
rect 6184 17144 6236 17153
rect 6368 17144 6420 17196
rect 7104 17076 7156 17128
rect 7840 17076 7892 17128
rect 8208 17144 8260 17196
rect 9312 17212 9364 17264
rect 8944 17144 8996 17196
rect 9220 17187 9272 17196
rect 9220 17153 9229 17187
rect 9229 17153 9263 17187
rect 9263 17153 9272 17187
rect 9220 17144 9272 17153
rect 9772 17144 9824 17196
rect 14004 17280 14056 17332
rect 9404 17076 9456 17128
rect 9496 17076 9548 17128
rect 10692 17144 10744 17196
rect 11060 17144 11112 17196
rect 11520 17144 11572 17196
rect 11888 17144 11940 17196
rect 12532 17144 12584 17196
rect 12716 17144 12768 17196
rect 13176 17144 13228 17196
rect 13544 17144 13596 17196
rect 15568 17323 15620 17332
rect 15568 17289 15577 17323
rect 15577 17289 15611 17323
rect 15611 17289 15620 17323
rect 15568 17280 15620 17289
rect 11244 17076 11296 17128
rect 14464 17144 14516 17196
rect 14832 17144 14884 17196
rect 14556 17076 14608 17128
rect 9036 17008 9088 17060
rect 11704 17008 11756 17060
rect 8852 16940 8904 16992
rect 9312 16940 9364 16992
rect 10048 16983 10100 16992
rect 10048 16949 10057 16983
rect 10057 16949 10091 16983
rect 10091 16949 10100 16983
rect 10048 16940 10100 16949
rect 10784 16983 10836 16992
rect 10784 16949 10793 16983
rect 10793 16949 10827 16983
rect 10827 16949 10836 16983
rect 10784 16940 10836 16949
rect 11152 16983 11204 16992
rect 11152 16949 11161 16983
rect 11161 16949 11195 16983
rect 11195 16949 11204 16983
rect 11152 16940 11204 16949
rect 11612 16983 11664 16992
rect 11612 16949 11621 16983
rect 11621 16949 11655 16983
rect 11655 16949 11664 16983
rect 11612 16940 11664 16949
rect 11980 16983 12032 16992
rect 11980 16949 11989 16983
rect 11989 16949 12023 16983
rect 12023 16949 12032 16983
rect 11980 16940 12032 16949
rect 12624 16940 12676 16992
rect 12808 16983 12860 16992
rect 12808 16949 12817 16983
rect 12817 16949 12851 16983
rect 12851 16949 12860 16983
rect 12808 16940 12860 16949
rect 13544 16940 13596 16992
rect 13728 16940 13780 16992
rect 2824 16838 2876 16890
rect 2888 16838 2940 16890
rect 2952 16838 3004 16890
rect 3016 16838 3068 16890
rect 3080 16838 3132 16890
rect 6572 16838 6624 16890
rect 6636 16838 6688 16890
rect 6700 16838 6752 16890
rect 6764 16838 6816 16890
rect 6828 16838 6880 16890
rect 10320 16838 10372 16890
rect 10384 16838 10436 16890
rect 10448 16838 10500 16890
rect 10512 16838 10564 16890
rect 10576 16838 10628 16890
rect 14068 16838 14120 16890
rect 14132 16838 14184 16890
rect 14196 16838 14248 16890
rect 14260 16838 14312 16890
rect 14324 16838 14376 16890
rect 8944 16779 8996 16788
rect 8944 16745 8953 16779
rect 8953 16745 8987 16779
rect 8987 16745 8996 16779
rect 8944 16736 8996 16745
rect 10692 16779 10744 16788
rect 10692 16745 10701 16779
rect 10701 16745 10735 16779
rect 10735 16745 10744 16779
rect 10692 16736 10744 16745
rect 11060 16779 11112 16788
rect 11060 16745 11069 16779
rect 11069 16745 11103 16779
rect 11103 16745 11112 16779
rect 11060 16736 11112 16745
rect 11888 16779 11940 16788
rect 11888 16745 11897 16779
rect 11897 16745 11931 16779
rect 11931 16745 11940 16779
rect 11888 16736 11940 16745
rect 12716 16779 12768 16788
rect 12716 16745 12725 16779
rect 12725 16745 12759 16779
rect 12759 16745 12768 16779
rect 12716 16736 12768 16745
rect 13176 16779 13228 16788
rect 13176 16745 13185 16779
rect 13185 16745 13219 16779
rect 13219 16745 13228 16779
rect 13176 16736 13228 16745
rect 13452 16779 13504 16788
rect 13452 16745 13461 16779
rect 13461 16745 13495 16779
rect 13495 16745 13504 16779
rect 13452 16736 13504 16745
rect 14832 16736 14884 16788
rect 1952 16600 2004 16652
rect 1032 16464 1084 16516
rect 572 16396 624 16448
rect 5816 16668 5868 16720
rect 9956 16668 10008 16720
rect 15108 16668 15160 16720
rect 6184 16600 6236 16652
rect 11980 16600 12032 16652
rect 4252 16532 4304 16584
rect 3976 16464 4028 16516
rect 9220 16464 9272 16516
rect 15384 16532 15436 16584
rect 16120 16532 16172 16584
rect 4068 16396 4120 16448
rect 12624 16396 12676 16448
rect 15660 16464 15712 16516
rect 15384 16439 15436 16448
rect 15384 16405 15393 16439
rect 15393 16405 15427 16439
rect 15427 16405 15436 16439
rect 15384 16396 15436 16405
rect 15476 16396 15528 16448
rect 4698 16294 4750 16346
rect 4762 16294 4814 16346
rect 4826 16294 4878 16346
rect 4890 16294 4942 16346
rect 4954 16294 5006 16346
rect 8446 16294 8498 16346
rect 8510 16294 8562 16346
rect 8574 16294 8626 16346
rect 8638 16294 8690 16346
rect 8702 16294 8754 16346
rect 12194 16294 12246 16346
rect 12258 16294 12310 16346
rect 12322 16294 12374 16346
rect 12386 16294 12438 16346
rect 12450 16294 12502 16346
rect 204 16056 256 16108
rect 16948 16124 17000 16176
rect 16488 16056 16540 16108
rect 4620 15920 4672 15972
rect 15200 15895 15252 15904
rect 15200 15861 15209 15895
rect 15209 15861 15243 15895
rect 15243 15861 15252 15895
rect 15200 15852 15252 15861
rect 15292 15852 15344 15904
rect 2824 15750 2876 15802
rect 2888 15750 2940 15802
rect 2952 15750 3004 15802
rect 3016 15750 3068 15802
rect 3080 15750 3132 15802
rect 6572 15750 6624 15802
rect 6636 15750 6688 15802
rect 6700 15750 6752 15802
rect 6764 15750 6816 15802
rect 6828 15750 6880 15802
rect 10320 15750 10372 15802
rect 10384 15750 10436 15802
rect 10448 15750 10500 15802
rect 10512 15750 10564 15802
rect 10576 15750 10628 15802
rect 14068 15750 14120 15802
rect 14132 15750 14184 15802
rect 14196 15750 14248 15802
rect 14260 15750 14312 15802
rect 14324 15750 14376 15802
rect 15476 15691 15528 15700
rect 15476 15657 15485 15691
rect 15485 15657 15519 15691
rect 15519 15657 15528 15691
rect 15476 15648 15528 15657
rect 4698 15206 4750 15258
rect 4762 15206 4814 15258
rect 4826 15206 4878 15258
rect 4890 15206 4942 15258
rect 4954 15206 5006 15258
rect 8446 15206 8498 15258
rect 8510 15206 8562 15258
rect 8574 15206 8626 15258
rect 8638 15206 8690 15258
rect 8702 15206 8754 15258
rect 12194 15206 12246 15258
rect 12258 15206 12310 15258
rect 12322 15206 12374 15258
rect 12386 15206 12438 15258
rect 12450 15206 12502 15258
rect 2824 14662 2876 14714
rect 2888 14662 2940 14714
rect 2952 14662 3004 14714
rect 3016 14662 3068 14714
rect 3080 14662 3132 14714
rect 6572 14662 6624 14714
rect 6636 14662 6688 14714
rect 6700 14662 6752 14714
rect 6764 14662 6816 14714
rect 6828 14662 6880 14714
rect 10320 14662 10372 14714
rect 10384 14662 10436 14714
rect 10448 14662 10500 14714
rect 10512 14662 10564 14714
rect 10576 14662 10628 14714
rect 14068 14662 14120 14714
rect 14132 14662 14184 14714
rect 14196 14662 14248 14714
rect 14260 14662 14312 14714
rect 14324 14662 14376 14714
rect 4698 14118 4750 14170
rect 4762 14118 4814 14170
rect 4826 14118 4878 14170
rect 4890 14118 4942 14170
rect 4954 14118 5006 14170
rect 8446 14118 8498 14170
rect 8510 14118 8562 14170
rect 8574 14118 8626 14170
rect 8638 14118 8690 14170
rect 8702 14118 8754 14170
rect 12194 14118 12246 14170
rect 12258 14118 12310 14170
rect 12322 14118 12374 14170
rect 12386 14118 12438 14170
rect 12450 14118 12502 14170
rect 4620 13923 4672 13932
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 3332 13812 3384 13864
rect 8852 13676 8904 13728
rect 2824 13574 2876 13626
rect 2888 13574 2940 13626
rect 2952 13574 3004 13626
rect 3016 13574 3068 13626
rect 3080 13574 3132 13626
rect 6572 13574 6624 13626
rect 6636 13574 6688 13626
rect 6700 13574 6752 13626
rect 6764 13574 6816 13626
rect 6828 13574 6880 13626
rect 10320 13574 10372 13626
rect 10384 13574 10436 13626
rect 10448 13574 10500 13626
rect 10512 13574 10564 13626
rect 10576 13574 10628 13626
rect 14068 13574 14120 13626
rect 14132 13574 14184 13626
rect 14196 13574 14248 13626
rect 14260 13574 14312 13626
rect 14324 13574 14376 13626
rect 4160 13311 4212 13320
rect 4160 13277 4169 13311
rect 4169 13277 4203 13311
rect 4203 13277 4212 13311
rect 4160 13268 4212 13277
rect 4252 13268 4304 13320
rect 8024 13132 8076 13184
rect 4698 13030 4750 13082
rect 4762 13030 4814 13082
rect 4826 13030 4878 13082
rect 4890 13030 4942 13082
rect 4954 13030 5006 13082
rect 8446 13030 8498 13082
rect 8510 13030 8562 13082
rect 8574 13030 8626 13082
rect 8638 13030 8690 13082
rect 8702 13030 8754 13082
rect 12194 13030 12246 13082
rect 12258 13030 12310 13082
rect 12322 13030 12374 13082
rect 12386 13030 12438 13082
rect 12450 13030 12502 13082
rect 4068 12971 4120 12980
rect 4068 12937 4077 12971
rect 4077 12937 4111 12971
rect 4111 12937 4120 12971
rect 4068 12928 4120 12937
rect 3792 12860 3844 12912
rect 7104 12928 7156 12980
rect 9404 12971 9456 12980
rect 9404 12937 9413 12971
rect 9413 12937 9447 12971
rect 9447 12937 9456 12971
rect 9404 12928 9456 12937
rect 14556 12928 14608 12980
rect 10232 12860 10284 12912
rect 7380 12835 7432 12844
rect 6092 12724 6144 12776
rect 7380 12801 7389 12835
rect 7389 12801 7423 12835
rect 7423 12801 7432 12835
rect 7380 12792 7432 12801
rect 9588 12835 9640 12844
rect 9588 12801 9597 12835
rect 9597 12801 9631 12835
rect 9631 12801 9640 12835
rect 9588 12792 9640 12801
rect 8300 12724 8352 12776
rect 8852 12724 8904 12776
rect 3884 12656 3936 12708
rect 7656 12588 7708 12640
rect 15568 12631 15620 12640
rect 15568 12597 15577 12631
rect 15577 12597 15611 12631
rect 15611 12597 15620 12631
rect 15568 12588 15620 12597
rect 2824 12486 2876 12538
rect 2888 12486 2940 12538
rect 2952 12486 3004 12538
rect 3016 12486 3068 12538
rect 3080 12486 3132 12538
rect 6572 12486 6624 12538
rect 6636 12486 6688 12538
rect 6700 12486 6752 12538
rect 6764 12486 6816 12538
rect 6828 12486 6880 12538
rect 10320 12486 10372 12538
rect 10384 12486 10436 12538
rect 10448 12486 10500 12538
rect 10512 12486 10564 12538
rect 10576 12486 10628 12538
rect 14068 12486 14120 12538
rect 14132 12486 14184 12538
rect 14196 12486 14248 12538
rect 14260 12486 14312 12538
rect 14324 12486 14376 12538
rect 4698 11942 4750 11994
rect 4762 11942 4814 11994
rect 4826 11942 4878 11994
rect 4890 11942 4942 11994
rect 4954 11942 5006 11994
rect 8446 11942 8498 11994
rect 8510 11942 8562 11994
rect 8574 11942 8626 11994
rect 8638 11942 8690 11994
rect 8702 11942 8754 11994
rect 12194 11942 12246 11994
rect 12258 11942 12310 11994
rect 12322 11942 12374 11994
rect 12386 11942 12438 11994
rect 12450 11942 12502 11994
rect 4528 11840 4580 11892
rect 1400 11747 1452 11756
rect 1400 11713 1409 11747
rect 1409 11713 1443 11747
rect 1443 11713 1452 11747
rect 1400 11704 1452 11713
rect 7472 11747 7524 11756
rect 7472 11713 7481 11747
rect 7481 11713 7515 11747
rect 7515 11713 7524 11747
rect 7472 11704 7524 11713
rect 8116 11747 8168 11756
rect 8116 11713 8125 11747
rect 8125 11713 8159 11747
rect 8159 11713 8168 11747
rect 8116 11704 8168 11713
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 5448 11568 5500 11620
rect 5908 11500 5960 11552
rect 6920 11568 6972 11620
rect 2824 11398 2876 11450
rect 2888 11398 2940 11450
rect 2952 11398 3004 11450
rect 3016 11398 3068 11450
rect 3080 11398 3132 11450
rect 6572 11398 6624 11450
rect 6636 11398 6688 11450
rect 6700 11398 6752 11450
rect 6764 11398 6816 11450
rect 6828 11398 6880 11450
rect 10320 11398 10372 11450
rect 10384 11398 10436 11450
rect 10448 11398 10500 11450
rect 10512 11398 10564 11450
rect 10576 11398 10628 11450
rect 14068 11398 14120 11450
rect 14132 11398 14184 11450
rect 14196 11398 14248 11450
rect 14260 11398 14312 11450
rect 14324 11398 14376 11450
rect 6460 11296 6512 11348
rect 4344 11024 4396 11076
rect 5264 11024 5316 11076
rect 9128 11296 9180 11348
rect 9496 11296 9548 11348
rect 7932 11228 7984 11280
rect 9496 11203 9548 11212
rect 9496 11169 9505 11203
rect 9505 11169 9539 11203
rect 9539 11169 9548 11203
rect 9496 11160 9548 11169
rect 5632 10956 5684 11008
rect 7104 10956 7156 11008
rect 9680 11024 9732 11076
rect 9312 10956 9364 11008
rect 9404 10999 9456 11008
rect 9404 10965 9413 10999
rect 9413 10965 9447 10999
rect 9447 10965 9456 10999
rect 9404 10956 9456 10965
rect 12716 10956 12768 11008
rect 13728 10956 13780 11008
rect 4698 10854 4750 10906
rect 4762 10854 4814 10906
rect 4826 10854 4878 10906
rect 4890 10854 4942 10906
rect 4954 10854 5006 10906
rect 8446 10854 8498 10906
rect 8510 10854 8562 10906
rect 8574 10854 8626 10906
rect 8638 10854 8690 10906
rect 8702 10854 8754 10906
rect 12194 10854 12246 10906
rect 12258 10854 12310 10906
rect 12322 10854 12374 10906
rect 12386 10854 12438 10906
rect 12450 10854 12502 10906
rect 4160 10752 4212 10804
rect 4344 10727 4396 10736
rect 4344 10693 4353 10727
rect 4353 10693 4387 10727
rect 4387 10693 4396 10727
rect 4344 10684 4396 10693
rect 3424 10616 3476 10668
rect 7564 10752 7616 10804
rect 10232 10752 10284 10804
rect 10692 10752 10744 10804
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6276 10616 6328 10668
rect 3240 10548 3292 10600
rect 5540 10480 5592 10532
rect 6184 10480 6236 10532
rect 5080 10412 5132 10464
rect 5724 10455 5776 10464
rect 5724 10421 5733 10455
rect 5733 10421 5767 10455
rect 5767 10421 5776 10455
rect 5724 10412 5776 10421
rect 6000 10455 6052 10464
rect 6000 10421 6009 10455
rect 6009 10421 6043 10455
rect 6043 10421 6052 10455
rect 6000 10412 6052 10421
rect 7748 10684 7800 10736
rect 7840 10684 7892 10736
rect 11796 10684 11848 10736
rect 7288 10616 7340 10668
rect 9496 10616 9548 10668
rect 7012 10548 7064 10600
rect 9312 10548 9364 10600
rect 10140 10616 10192 10668
rect 10232 10548 10284 10600
rect 11152 10480 11204 10532
rect 8852 10412 8904 10464
rect 9864 10412 9916 10464
rect 10784 10412 10836 10464
rect 12900 10412 12952 10464
rect 15384 10412 15436 10464
rect 2824 10310 2876 10362
rect 2888 10310 2940 10362
rect 2952 10310 3004 10362
rect 3016 10310 3068 10362
rect 3080 10310 3132 10362
rect 6572 10310 6624 10362
rect 6636 10310 6688 10362
rect 6700 10310 6752 10362
rect 6764 10310 6816 10362
rect 6828 10310 6880 10362
rect 10320 10310 10372 10362
rect 10384 10310 10436 10362
rect 10448 10310 10500 10362
rect 10512 10310 10564 10362
rect 10576 10310 10628 10362
rect 14068 10310 14120 10362
rect 14132 10310 14184 10362
rect 14196 10310 14248 10362
rect 14260 10310 14312 10362
rect 14324 10310 14376 10362
rect 4712 10208 4764 10260
rect 6460 10208 6512 10260
rect 7104 10208 7156 10260
rect 9036 10208 9088 10260
rect 9956 10208 10008 10260
rect 10876 10251 10928 10260
rect 10876 10217 10885 10251
rect 10885 10217 10919 10251
rect 10919 10217 10928 10251
rect 10876 10208 10928 10217
rect 5448 10072 5500 10124
rect 5816 10072 5868 10124
rect 5908 10115 5960 10124
rect 5908 10081 5917 10115
rect 5917 10081 5951 10115
rect 5951 10081 5960 10115
rect 6184 10140 6236 10192
rect 5908 10072 5960 10081
rect 7564 10115 7616 10124
rect 7564 10081 7573 10115
rect 7573 10081 7607 10115
rect 7607 10081 7616 10115
rect 7564 10072 7616 10081
rect 8024 10072 8076 10124
rect 9864 10140 9916 10192
rect 10048 10140 10100 10192
rect 12716 10208 12768 10260
rect 13084 10251 13136 10260
rect 13084 10217 13093 10251
rect 13093 10217 13127 10251
rect 13127 10217 13136 10251
rect 13084 10208 13136 10217
rect 13360 10251 13412 10260
rect 13360 10217 13369 10251
rect 13369 10217 13403 10251
rect 13403 10217 13412 10251
rect 13360 10208 13412 10217
rect 13636 10251 13688 10260
rect 13636 10217 13645 10251
rect 13645 10217 13679 10251
rect 13679 10217 13688 10251
rect 13636 10208 13688 10217
rect 3332 10047 3384 10056
rect 3332 10013 3350 10047
rect 3350 10013 3384 10047
rect 3332 10004 3384 10013
rect 4712 10047 4764 10056
rect 4712 10013 4721 10047
rect 4721 10013 4755 10047
rect 4755 10013 4764 10047
rect 4712 10004 4764 10013
rect 4896 10004 4948 10056
rect 8300 10004 8352 10056
rect 9496 10072 9548 10124
rect 11888 10140 11940 10192
rect 12532 10183 12584 10192
rect 12532 10149 12541 10183
rect 12541 10149 12575 10183
rect 12575 10149 12584 10183
rect 12532 10140 12584 10149
rect 9128 10047 9180 10056
rect 9128 10013 9137 10047
rect 9137 10013 9171 10047
rect 9171 10013 9180 10047
rect 9128 10004 9180 10013
rect 9220 10004 9272 10056
rect 11244 10072 11296 10124
rect 11060 10047 11112 10056
rect 3976 9936 4028 9988
rect 2044 9868 2096 9920
rect 5172 9868 5224 9920
rect 9772 9936 9824 9988
rect 11060 10013 11069 10047
rect 11069 10013 11103 10047
rect 11103 10013 11112 10047
rect 11060 10004 11112 10013
rect 11704 10072 11756 10124
rect 12900 10072 12952 10124
rect 11980 10004 12032 10056
rect 12624 10004 12676 10056
rect 15292 10140 15344 10192
rect 15200 10072 15252 10124
rect 13820 10047 13872 10056
rect 13820 10013 13829 10047
rect 13829 10013 13863 10047
rect 13863 10013 13872 10047
rect 13820 10004 13872 10013
rect 7196 9868 7248 9920
rect 8208 9868 8260 9920
rect 9036 9868 9088 9920
rect 9220 9911 9272 9920
rect 9220 9877 9229 9911
rect 9229 9877 9263 9911
rect 9263 9877 9272 9911
rect 9220 9868 9272 9877
rect 9588 9911 9640 9920
rect 9588 9877 9597 9911
rect 9597 9877 9631 9911
rect 9631 9877 9640 9911
rect 9588 9868 9640 9877
rect 9956 9868 10008 9920
rect 11244 9868 11296 9920
rect 11428 9911 11480 9920
rect 11428 9877 11437 9911
rect 11437 9877 11471 9911
rect 11471 9877 11480 9911
rect 11428 9868 11480 9877
rect 11520 9868 11572 9920
rect 11796 9868 11848 9920
rect 12624 9868 12676 9920
rect 12716 9868 12768 9920
rect 14924 9936 14976 9988
rect 14740 9868 14792 9920
rect 4698 9766 4750 9818
rect 4762 9766 4814 9818
rect 4826 9766 4878 9818
rect 4890 9766 4942 9818
rect 4954 9766 5006 9818
rect 8446 9766 8498 9818
rect 8510 9766 8562 9818
rect 8574 9766 8626 9818
rect 8638 9766 8690 9818
rect 8702 9766 8754 9818
rect 12194 9766 12246 9818
rect 12258 9766 12310 9818
rect 12322 9766 12374 9818
rect 12386 9766 12438 9818
rect 12450 9766 12502 9818
rect 3424 9664 3476 9716
rect 5172 9664 5224 9716
rect 5448 9664 5500 9716
rect 3332 9596 3384 9648
rect 5816 9664 5868 9716
rect 6368 9664 6420 9716
rect 8300 9664 8352 9716
rect 9312 9707 9364 9716
rect 9312 9673 9321 9707
rect 9321 9673 9355 9707
rect 9355 9673 9364 9707
rect 9312 9664 9364 9673
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 7104 9528 7156 9580
rect 7380 9596 7432 9648
rect 8760 9596 8812 9648
rect 8852 9596 8904 9648
rect 9128 9596 9180 9648
rect 7656 9528 7708 9580
rect 8484 9528 8536 9580
rect 10232 9664 10284 9716
rect 12624 9664 12676 9716
rect 13636 9664 13688 9716
rect 13544 9596 13596 9648
rect 3240 9503 3292 9512
rect 3240 9469 3249 9503
rect 3249 9469 3283 9503
rect 3283 9469 3292 9503
rect 3240 9460 3292 9469
rect 4252 9460 4304 9512
rect 8208 9503 8260 9512
rect 3148 9392 3200 9444
rect 4160 9392 4212 9444
rect 2136 9324 2188 9376
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 12808 9528 12860 9580
rect 8852 9503 8904 9512
rect 6644 9392 6696 9444
rect 8852 9469 8861 9503
rect 8861 9469 8895 9503
rect 8895 9469 8904 9503
rect 8852 9460 8904 9469
rect 9312 9460 9364 9512
rect 11612 9460 11664 9512
rect 7840 9324 7892 9376
rect 8024 9324 8076 9376
rect 8760 9392 8812 9444
rect 9864 9392 9916 9444
rect 8300 9324 8352 9376
rect 10232 9324 10284 9376
rect 2824 9222 2876 9274
rect 2888 9222 2940 9274
rect 2952 9222 3004 9274
rect 3016 9222 3068 9274
rect 3080 9222 3132 9274
rect 6572 9222 6624 9274
rect 6636 9222 6688 9274
rect 6700 9222 6752 9274
rect 6764 9222 6816 9274
rect 6828 9222 6880 9274
rect 10320 9222 10372 9274
rect 10384 9222 10436 9274
rect 10448 9222 10500 9274
rect 10512 9222 10564 9274
rect 10576 9222 10628 9274
rect 14068 9222 14120 9274
rect 14132 9222 14184 9274
rect 14196 9222 14248 9274
rect 14260 9222 14312 9274
rect 14324 9222 14376 9274
rect 3608 9120 3660 9172
rect 7288 9120 7340 9172
rect 7472 9120 7524 9172
rect 8484 9095 8536 9104
rect 8484 9061 8493 9095
rect 8493 9061 8527 9095
rect 8527 9061 8536 9095
rect 8484 9052 8536 9061
rect 5816 8984 5868 9036
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 7012 8916 7064 8968
rect 9036 8984 9088 9036
rect 9496 9027 9548 9036
rect 9496 8993 9505 9027
rect 9505 8993 9539 9027
rect 9539 8993 9548 9027
rect 9496 8984 9548 8993
rect 6920 8848 6972 8900
rect 8024 8848 8076 8900
rect 12072 8916 12124 8968
rect 9404 8848 9456 8900
rect 4528 8780 4580 8832
rect 9864 8780 9916 8832
rect 10784 8780 10836 8832
rect 4698 8678 4750 8730
rect 4762 8678 4814 8730
rect 4826 8678 4878 8730
rect 4890 8678 4942 8730
rect 4954 8678 5006 8730
rect 8446 8678 8498 8730
rect 8510 8678 8562 8730
rect 8574 8678 8626 8730
rect 8638 8678 8690 8730
rect 8702 8678 8754 8730
rect 12194 8678 12246 8730
rect 12258 8678 12310 8730
rect 12322 8678 12374 8730
rect 12386 8678 12438 8730
rect 12450 8678 12502 8730
rect 6368 8576 6420 8628
rect 3332 8440 3384 8492
rect 3148 8372 3200 8424
rect 3424 8372 3476 8424
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 6092 8304 6144 8356
rect 8852 8576 8904 8628
rect 9864 8576 9916 8628
rect 10692 8576 10744 8628
rect 7840 8551 7892 8560
rect 7840 8517 7858 8551
rect 7858 8517 7892 8551
rect 7840 8508 7892 8517
rect 9680 8508 9732 8560
rect 7104 8440 7156 8492
rect 8208 8440 8260 8492
rect 12532 8372 12584 8424
rect 12808 8347 12860 8356
rect 12808 8313 12817 8347
rect 12817 8313 12851 8347
rect 12851 8313 12860 8347
rect 12808 8304 12860 8313
rect 7012 8236 7064 8288
rect 8208 8236 8260 8288
rect 2824 8134 2876 8186
rect 2888 8134 2940 8186
rect 2952 8134 3004 8186
rect 3016 8134 3068 8186
rect 3080 8134 3132 8186
rect 6572 8134 6624 8186
rect 6636 8134 6688 8186
rect 6700 8134 6752 8186
rect 6764 8134 6816 8186
rect 6828 8134 6880 8186
rect 10320 8134 10372 8186
rect 10384 8134 10436 8186
rect 10448 8134 10500 8186
rect 10512 8134 10564 8186
rect 10576 8134 10628 8186
rect 14068 8134 14120 8186
rect 14132 8134 14184 8186
rect 14196 8134 14248 8186
rect 14260 8134 14312 8186
rect 14324 8134 14376 8186
rect 7196 8075 7248 8084
rect 7196 8041 7205 8075
rect 7205 8041 7239 8075
rect 7239 8041 7248 8075
rect 7196 8032 7248 8041
rect 7564 8032 7616 8084
rect 8208 8032 8260 8084
rect 7012 7939 7064 7948
rect 7012 7905 7021 7939
rect 7021 7905 7055 7939
rect 7055 7905 7064 7939
rect 7012 7896 7064 7905
rect 7840 7939 7892 7948
rect 7840 7905 7849 7939
rect 7849 7905 7883 7939
rect 7883 7905 7892 7939
rect 7840 7896 7892 7905
rect 5264 7871 5316 7880
rect 5264 7837 5273 7871
rect 5273 7837 5307 7871
rect 5307 7837 5316 7871
rect 5264 7828 5316 7837
rect 9220 7828 9272 7880
rect 7932 7760 7984 7812
rect 4698 7590 4750 7642
rect 4762 7590 4814 7642
rect 4826 7590 4878 7642
rect 4890 7590 4942 7642
rect 4954 7590 5006 7642
rect 8446 7590 8498 7642
rect 8510 7590 8562 7642
rect 8574 7590 8626 7642
rect 8638 7590 8690 7642
rect 8702 7590 8754 7642
rect 12194 7590 12246 7642
rect 12258 7590 12310 7642
rect 12322 7590 12374 7642
rect 12386 7590 12438 7642
rect 12450 7590 12502 7642
rect 9128 7488 9180 7540
rect 10140 7420 10192 7472
rect 5448 7352 5500 7404
rect 8944 7352 8996 7404
rect 9312 7352 9364 7404
rect 3608 7216 3660 7268
rect 3976 7191 4028 7200
rect 3976 7157 3985 7191
rect 3985 7157 4019 7191
rect 4019 7157 4028 7191
rect 3976 7148 4028 7157
rect 4528 7191 4580 7200
rect 4528 7157 4537 7191
rect 4537 7157 4571 7191
rect 4571 7157 4580 7191
rect 4528 7148 4580 7157
rect 5632 7148 5684 7200
rect 9036 7148 9088 7200
rect 2824 7046 2876 7098
rect 2888 7046 2940 7098
rect 2952 7046 3004 7098
rect 3016 7046 3068 7098
rect 3080 7046 3132 7098
rect 6572 7046 6624 7098
rect 6636 7046 6688 7098
rect 6700 7046 6752 7098
rect 6764 7046 6816 7098
rect 6828 7046 6880 7098
rect 10320 7046 10372 7098
rect 10384 7046 10436 7098
rect 10448 7046 10500 7098
rect 10512 7046 10564 7098
rect 10576 7046 10628 7098
rect 14068 7046 14120 7098
rect 14132 7046 14184 7098
rect 14196 7046 14248 7098
rect 14260 7046 14312 7098
rect 14324 7046 14376 7098
rect 3148 6783 3200 6792
rect 3148 6749 3157 6783
rect 3157 6749 3191 6783
rect 3191 6749 3200 6783
rect 3148 6740 3200 6749
rect 3148 6604 3200 6656
rect 4698 6502 4750 6554
rect 4762 6502 4814 6554
rect 4826 6502 4878 6554
rect 4890 6502 4942 6554
rect 4954 6502 5006 6554
rect 8446 6502 8498 6554
rect 8510 6502 8562 6554
rect 8574 6502 8626 6554
rect 8638 6502 8690 6554
rect 8702 6502 8754 6554
rect 12194 6502 12246 6554
rect 12258 6502 12310 6554
rect 12322 6502 12374 6554
rect 12386 6502 12438 6554
rect 12450 6502 12502 6554
rect 2824 5958 2876 6010
rect 2888 5958 2940 6010
rect 2952 5958 3004 6010
rect 3016 5958 3068 6010
rect 3080 5958 3132 6010
rect 6572 5958 6624 6010
rect 6636 5958 6688 6010
rect 6700 5958 6752 6010
rect 6764 5958 6816 6010
rect 6828 5958 6880 6010
rect 10320 5958 10372 6010
rect 10384 5958 10436 6010
rect 10448 5958 10500 6010
rect 10512 5958 10564 6010
rect 10576 5958 10628 6010
rect 14068 5958 14120 6010
rect 14132 5958 14184 6010
rect 14196 5958 14248 6010
rect 14260 5958 14312 6010
rect 14324 5958 14376 6010
rect 4698 5414 4750 5466
rect 4762 5414 4814 5466
rect 4826 5414 4878 5466
rect 4890 5414 4942 5466
rect 4954 5414 5006 5466
rect 8446 5414 8498 5466
rect 8510 5414 8562 5466
rect 8574 5414 8626 5466
rect 8638 5414 8690 5466
rect 8702 5414 8754 5466
rect 12194 5414 12246 5466
rect 12258 5414 12310 5466
rect 12322 5414 12374 5466
rect 12386 5414 12438 5466
rect 12450 5414 12502 5466
rect 3148 5176 3200 5228
rect 1492 5015 1544 5024
rect 1492 4981 1501 5015
rect 1501 4981 1535 5015
rect 1535 4981 1544 5015
rect 1492 4972 1544 4981
rect 2824 4870 2876 4922
rect 2888 4870 2940 4922
rect 2952 4870 3004 4922
rect 3016 4870 3068 4922
rect 3080 4870 3132 4922
rect 6572 4870 6624 4922
rect 6636 4870 6688 4922
rect 6700 4870 6752 4922
rect 6764 4870 6816 4922
rect 6828 4870 6880 4922
rect 10320 4870 10372 4922
rect 10384 4870 10436 4922
rect 10448 4870 10500 4922
rect 10512 4870 10564 4922
rect 10576 4870 10628 4922
rect 14068 4870 14120 4922
rect 14132 4870 14184 4922
rect 14196 4870 14248 4922
rect 14260 4870 14312 4922
rect 14324 4870 14376 4922
rect 4698 4326 4750 4378
rect 4762 4326 4814 4378
rect 4826 4326 4878 4378
rect 4890 4326 4942 4378
rect 4954 4326 5006 4378
rect 8446 4326 8498 4378
rect 8510 4326 8562 4378
rect 8574 4326 8626 4378
rect 8638 4326 8690 4378
rect 8702 4326 8754 4378
rect 12194 4326 12246 4378
rect 12258 4326 12310 4378
rect 12322 4326 12374 4378
rect 12386 4326 12438 4378
rect 12450 4326 12502 4378
rect 2824 3782 2876 3834
rect 2888 3782 2940 3834
rect 2952 3782 3004 3834
rect 3016 3782 3068 3834
rect 3080 3782 3132 3834
rect 6572 3782 6624 3834
rect 6636 3782 6688 3834
rect 6700 3782 6752 3834
rect 6764 3782 6816 3834
rect 6828 3782 6880 3834
rect 10320 3782 10372 3834
rect 10384 3782 10436 3834
rect 10448 3782 10500 3834
rect 10512 3782 10564 3834
rect 10576 3782 10628 3834
rect 14068 3782 14120 3834
rect 14132 3782 14184 3834
rect 14196 3782 14248 3834
rect 14260 3782 14312 3834
rect 14324 3782 14376 3834
rect 13820 3680 13872 3732
rect 4528 3476 4580 3528
rect 16948 3476 17000 3528
rect 1032 3340 1084 3392
rect 15292 3383 15344 3392
rect 15292 3349 15301 3383
rect 15301 3349 15335 3383
rect 15335 3349 15344 3383
rect 15292 3340 15344 3349
rect 15660 3340 15712 3392
rect 4698 3238 4750 3290
rect 4762 3238 4814 3290
rect 4826 3238 4878 3290
rect 4890 3238 4942 3290
rect 4954 3238 5006 3290
rect 8446 3238 8498 3290
rect 8510 3238 8562 3290
rect 8574 3238 8626 3290
rect 8638 3238 8690 3290
rect 8702 3238 8754 3290
rect 12194 3238 12246 3290
rect 12258 3238 12310 3290
rect 12322 3238 12374 3290
rect 12386 3238 12438 3290
rect 12450 3238 12502 3290
rect 3240 3136 3292 3188
rect 14924 3179 14976 3188
rect 14924 3145 14933 3179
rect 14933 3145 14967 3179
rect 14967 3145 14976 3179
rect 14924 3136 14976 3145
rect 3976 3068 4028 3120
rect 14740 3068 14792 3120
rect 2044 3043 2096 3052
rect 2044 3009 2053 3043
rect 2053 3009 2087 3043
rect 2087 3009 2096 3043
rect 2044 3000 2096 3009
rect 2136 3043 2188 3052
rect 2136 3009 2145 3043
rect 2145 3009 2179 3043
rect 2179 3009 2188 3043
rect 2136 3000 2188 3009
rect 9588 2932 9640 2984
rect 572 2864 624 2916
rect 204 2796 256 2848
rect 8760 2839 8812 2848
rect 8760 2805 8769 2839
rect 8769 2805 8803 2839
rect 8803 2805 8812 2839
rect 8760 2796 8812 2805
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 10876 2839 10928 2848
rect 10876 2805 10885 2839
rect 10885 2805 10919 2839
rect 10919 2805 10928 2839
rect 10876 2796 10928 2805
rect 11336 2796 11388 2848
rect 12532 2796 12584 2848
rect 13452 2839 13504 2848
rect 13452 2805 13461 2839
rect 13461 2805 13495 2839
rect 13495 2805 13504 2839
rect 13452 2796 13504 2805
rect 13912 2839 13964 2848
rect 13912 2805 13921 2839
rect 13921 2805 13955 2839
rect 13955 2805 13964 2839
rect 13912 2796 13964 2805
rect 14740 2839 14792 2848
rect 14740 2805 14749 2839
rect 14749 2805 14783 2839
rect 14783 2805 14792 2839
rect 14740 2796 14792 2805
rect 15384 3043 15436 3052
rect 15384 3009 15393 3043
rect 15393 3009 15427 3043
rect 15427 3009 15436 3043
rect 15384 3000 15436 3009
rect 15660 3043 15712 3052
rect 15660 3009 15669 3043
rect 15669 3009 15703 3043
rect 15703 3009 15712 3043
rect 15660 3000 15712 3009
rect 15292 2932 15344 2984
rect 16488 2932 16540 2984
rect 15200 2864 15252 2916
rect 2824 2694 2876 2746
rect 2888 2694 2940 2746
rect 2952 2694 3004 2746
rect 3016 2694 3068 2746
rect 3080 2694 3132 2746
rect 6572 2694 6624 2746
rect 6636 2694 6688 2746
rect 6700 2694 6752 2746
rect 6764 2694 6816 2746
rect 6828 2694 6880 2746
rect 10320 2694 10372 2746
rect 10384 2694 10436 2746
rect 10448 2694 10500 2746
rect 10512 2694 10564 2746
rect 10576 2694 10628 2746
rect 14068 2694 14120 2746
rect 14132 2694 14184 2746
rect 14196 2694 14248 2746
rect 14260 2694 14312 2746
rect 14324 2694 14376 2746
rect 5080 2592 5132 2644
rect 5264 2592 5316 2644
rect 8300 2592 8352 2644
rect 8852 2592 8904 2644
rect 9864 2635 9916 2644
rect 9864 2601 9873 2635
rect 9873 2601 9907 2635
rect 9907 2601 9916 2635
rect 9864 2592 9916 2601
rect 12072 2592 12124 2644
rect 13636 2592 13688 2644
rect 3608 2524 3660 2576
rect 2688 2431 2740 2440
rect 2688 2397 2697 2431
rect 2697 2397 2731 2431
rect 2731 2397 2740 2431
rect 2688 2388 2740 2397
rect 4160 2456 4212 2508
rect 4252 2388 4304 2440
rect 4620 2388 4672 2440
rect 5632 2524 5684 2576
rect 5264 2431 5316 2440
rect 5264 2397 5266 2431
rect 5266 2397 5300 2431
rect 5300 2397 5316 2431
rect 5264 2388 5316 2397
rect 6092 2431 6144 2440
rect 6092 2397 6101 2431
rect 6101 2397 6135 2431
rect 6135 2397 6144 2431
rect 6092 2388 6144 2397
rect 6644 2431 6696 2440
rect 6644 2397 6653 2431
rect 6653 2397 6687 2431
rect 6687 2397 6696 2431
rect 6644 2388 6696 2397
rect 7288 2388 7340 2440
rect 9036 2456 9088 2508
rect 9404 2524 9456 2576
rect 10784 2524 10836 2576
rect 13268 2524 13320 2576
rect 9864 2456 9916 2508
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8668 2431 8720 2440
rect 6000 2320 6052 2372
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 8852 2388 8904 2440
rect 9220 2388 9272 2440
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 1492 2252 1544 2304
rect 1860 2252 1912 2304
rect 2320 2252 2372 2304
rect 2780 2252 2832 2304
rect 3148 2252 3200 2304
rect 3608 2252 3660 2304
rect 4068 2252 4120 2304
rect 4436 2252 4488 2304
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 5356 2252 5408 2304
rect 5724 2252 5776 2304
rect 6184 2252 6236 2304
rect 6644 2252 6696 2304
rect 7012 2252 7064 2304
rect 7472 2252 7524 2304
rect 7932 2252 7984 2304
rect 8300 2252 8352 2304
rect 8944 2320 8996 2372
rect 9128 2252 9180 2304
rect 9312 2295 9364 2304
rect 9312 2261 9321 2295
rect 9321 2261 9355 2295
rect 9355 2261 9364 2295
rect 9312 2252 9364 2261
rect 10048 2320 10100 2372
rect 10508 2388 10560 2440
rect 11060 2388 11112 2440
rect 11336 2388 11388 2440
rect 11796 2388 11848 2440
rect 12532 2388 12584 2440
rect 10968 2295 11020 2304
rect 10968 2261 10977 2295
rect 10977 2261 11011 2295
rect 11011 2261 11020 2295
rect 10968 2252 11020 2261
rect 11152 2252 11204 2304
rect 11520 2295 11572 2304
rect 11520 2261 11529 2295
rect 11529 2261 11563 2295
rect 11563 2261 11572 2295
rect 11888 2295 11940 2304
rect 11520 2252 11572 2261
rect 11888 2261 11897 2295
rect 11897 2261 11931 2295
rect 11931 2261 11940 2295
rect 11888 2252 11940 2261
rect 12072 2252 12124 2304
rect 12624 2320 12676 2372
rect 13084 2388 13136 2440
rect 13452 2388 13504 2440
rect 13912 2388 13964 2440
rect 14372 2388 14424 2440
rect 14740 2388 14792 2440
rect 15200 2388 15252 2440
rect 14096 2295 14148 2304
rect 14096 2261 14105 2295
rect 14105 2261 14139 2295
rect 14139 2261 14148 2295
rect 14096 2252 14148 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 15384 2252 15436 2304
rect 16028 2252 16080 2304
rect 4698 2150 4750 2202
rect 4762 2150 4814 2202
rect 4826 2150 4878 2202
rect 4890 2150 4942 2202
rect 4954 2150 5006 2202
rect 8446 2150 8498 2202
rect 8510 2150 8562 2202
rect 8574 2150 8626 2202
rect 8638 2150 8690 2202
rect 8702 2150 8754 2202
rect 12194 2150 12246 2202
rect 12258 2150 12310 2202
rect 12322 2150 12374 2202
rect 12386 2150 12438 2202
rect 12450 2150 12502 2202
rect 6092 2048 6144 2100
rect 7288 2048 7340 2100
rect 11428 2048 11480 2100
rect 11980 2048 12032 2100
rect 15292 2048 15344 2100
rect 9128 1980 9180 2032
rect 12716 1980 12768 2032
rect 10140 1912 10192 1964
rect 7748 1844 7800 1896
rect 11520 1844 11572 1896
rect 9772 1776 9824 1828
rect 14096 1776 14148 1828
rect 6276 1708 6328 1760
rect 10968 1708 11020 1760
rect 4528 1640 4580 1692
rect 9312 1640 9364 1692
rect 6920 1572 6972 1624
rect 11888 1572 11940 1624
<< metal2 >>
rect 202 19200 258 20000
rect 570 19200 626 20000
rect 1030 19200 1086 20000
rect 1398 19200 1454 20000
rect 1858 19200 1914 20000
rect 2226 19200 2282 20000
rect 2686 19200 2742 20000
rect 3054 19200 3110 20000
rect 3514 19200 3570 20000
rect 3974 19200 4030 20000
rect 4342 19200 4398 20000
rect 4802 19200 4858 20000
rect 5170 19200 5226 20000
rect 5630 19200 5686 20000
rect 5998 19200 6054 20000
rect 6458 19200 6514 20000
rect 6826 19200 6882 20000
rect 7286 19200 7342 20000
rect 7746 19200 7802 20000
rect 8114 19200 8170 20000
rect 8574 19200 8630 20000
rect 8680 19230 8892 19258
rect 216 16114 244 19200
rect 584 16454 612 19200
rect 1044 16522 1072 19200
rect 1412 17338 1440 19200
rect 1872 17338 1900 19200
rect 1950 18320 2006 18329
rect 1950 18255 2006 18264
rect 1400 17332 1452 17338
rect 1400 17274 1452 17280
rect 1860 17332 1912 17338
rect 1860 17274 1912 17280
rect 1964 16658 1992 18255
rect 2240 17338 2268 19200
rect 2700 17338 2728 19200
rect 3068 17338 3096 19200
rect 3528 17338 3556 19200
rect 2228 17332 2280 17338
rect 2228 17274 2280 17280
rect 2688 17332 2740 17338
rect 2688 17274 2740 17280
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3516 17332 3568 17338
rect 3988 17320 4016 19200
rect 4356 17338 4384 19200
rect 4816 17626 4844 19200
rect 4632 17598 4844 17626
rect 4632 17338 4660 17598
rect 4698 17436 5006 17456
rect 4698 17434 4704 17436
rect 4760 17434 4784 17436
rect 4840 17434 4864 17436
rect 4920 17434 4944 17436
rect 5000 17434 5006 17436
rect 4760 17382 4762 17434
rect 4942 17382 4944 17434
rect 4698 17380 4704 17382
rect 4760 17380 4784 17382
rect 4840 17380 4864 17382
rect 4920 17380 4944 17382
rect 5000 17380 5006 17382
rect 4698 17360 5006 17380
rect 5184 17338 5212 19200
rect 5644 17338 5672 19200
rect 6012 17338 6040 19200
rect 6184 17672 6236 17678
rect 6184 17614 6236 17620
rect 4160 17332 4212 17338
rect 3988 17292 4160 17320
rect 3516 17274 3568 17280
rect 4160 17274 4212 17280
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5632 17332 5684 17338
rect 5632 17274 5684 17280
rect 6000 17332 6052 17338
rect 6000 17274 6052 17280
rect 3884 17264 3936 17270
rect 3884 17206 3936 17212
rect 2136 17196 2188 17202
rect 2136 17138 2188 17144
rect 3148 17196 3200 17202
rect 3424 17196 3476 17202
rect 3200 17156 3280 17184
rect 3148 17138 3200 17144
rect 1952 16652 2004 16658
rect 1952 16594 2004 16600
rect 1032 16516 1084 16522
rect 1032 16458 1084 16464
rect 572 16448 624 16454
rect 572 16390 624 16396
rect 204 16108 256 16114
rect 204 16050 256 16056
rect 1400 11756 1452 11762
rect 1400 11698 1452 11704
rect 1412 11665 1440 11698
rect 1398 11656 1454 11665
rect 1398 11591 1454 11600
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 1490 8392 1546 8401
rect 1490 8327 1492 8336
rect 1544 8327 1546 8336
rect 1492 8298 1544 8304
rect 1492 5024 1544 5030
rect 1490 4992 1492 5001
rect 1544 4992 1546 5001
rect 1490 4927 1546 4936
rect 1032 3392 1084 3398
rect 1032 3334 1084 3340
rect 572 2916 624 2922
rect 572 2858 624 2864
rect 204 2848 256 2854
rect 204 2790 256 2796
rect 216 800 244 2790
rect 584 800 612 2858
rect 1044 800 1072 3334
rect 2056 3058 2084 9862
rect 2148 9382 2176 17138
rect 2824 16892 3132 16912
rect 2824 16890 2830 16892
rect 2886 16890 2910 16892
rect 2966 16890 2990 16892
rect 3046 16890 3070 16892
rect 3126 16890 3132 16892
rect 2886 16838 2888 16890
rect 3068 16838 3070 16890
rect 2824 16836 2830 16838
rect 2886 16836 2910 16838
rect 2966 16836 2990 16838
rect 3046 16836 3070 16838
rect 3126 16836 3132 16838
rect 2824 16816 3132 16836
rect 2824 15804 3132 15824
rect 2824 15802 2830 15804
rect 2886 15802 2910 15804
rect 2966 15802 2990 15804
rect 3046 15802 3070 15804
rect 3126 15802 3132 15804
rect 2886 15750 2888 15802
rect 3068 15750 3070 15802
rect 2824 15748 2830 15750
rect 2886 15748 2910 15750
rect 2966 15748 2990 15750
rect 3046 15748 3070 15750
rect 3126 15748 3132 15750
rect 2824 15728 3132 15748
rect 3146 15056 3202 15065
rect 3146 14991 3202 15000
rect 2824 14716 3132 14736
rect 2824 14714 2830 14716
rect 2886 14714 2910 14716
rect 2966 14714 2990 14716
rect 3046 14714 3070 14716
rect 3126 14714 3132 14716
rect 2886 14662 2888 14714
rect 3068 14662 3070 14714
rect 2824 14660 2830 14662
rect 2886 14660 2910 14662
rect 2966 14660 2990 14662
rect 3046 14660 3070 14662
rect 3126 14660 3132 14662
rect 2824 14640 3132 14660
rect 2824 13628 3132 13648
rect 2824 13626 2830 13628
rect 2886 13626 2910 13628
rect 2966 13626 2990 13628
rect 3046 13626 3070 13628
rect 3126 13626 3132 13628
rect 2886 13574 2888 13626
rect 3068 13574 3070 13626
rect 2824 13572 2830 13574
rect 2886 13572 2910 13574
rect 2966 13572 2990 13574
rect 3046 13572 3070 13574
rect 3126 13572 3132 13574
rect 2824 13552 3132 13572
rect 2824 12540 3132 12560
rect 2824 12538 2830 12540
rect 2886 12538 2910 12540
rect 2966 12538 2990 12540
rect 3046 12538 3070 12540
rect 3126 12538 3132 12540
rect 2886 12486 2888 12538
rect 3068 12486 3070 12538
rect 2824 12484 2830 12486
rect 2886 12484 2910 12486
rect 2966 12484 2990 12486
rect 3046 12484 3070 12486
rect 3126 12484 3132 12486
rect 2824 12464 3132 12484
rect 2824 11452 3132 11472
rect 2824 11450 2830 11452
rect 2886 11450 2910 11452
rect 2966 11450 2990 11452
rect 3046 11450 3070 11452
rect 3126 11450 3132 11452
rect 2886 11398 2888 11450
rect 3068 11398 3070 11450
rect 2824 11396 2830 11398
rect 2886 11396 2910 11398
rect 2966 11396 2990 11398
rect 3046 11396 3070 11398
rect 3126 11396 3132 11398
rect 2824 11376 3132 11396
rect 2824 10364 3132 10384
rect 2824 10362 2830 10364
rect 2886 10362 2910 10364
rect 2966 10362 2990 10364
rect 3046 10362 3070 10364
rect 3126 10362 3132 10364
rect 2886 10310 2888 10362
rect 3068 10310 3070 10362
rect 2824 10308 2830 10310
rect 2886 10308 2910 10310
rect 2966 10308 2990 10310
rect 3046 10308 3070 10310
rect 3126 10308 3132 10310
rect 2824 10288 3132 10308
rect 3160 9450 3188 14991
rect 3252 10606 3280 17156
rect 3424 17138 3476 17144
rect 3608 17196 3660 17202
rect 3608 17138 3660 17144
rect 3332 13864 3384 13870
rect 3332 13806 3384 13812
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3344 10062 3372 13806
rect 3436 10674 3464 17138
rect 3424 10668 3476 10674
rect 3424 10610 3476 10616
rect 3332 10056 3384 10062
rect 3332 9998 3384 10004
rect 3344 9654 3372 9998
rect 3424 9716 3476 9722
rect 3424 9658 3476 9664
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 3148 9444 3200 9450
rect 3148 9386 3200 9392
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 2824 9276 3132 9296
rect 2824 9274 2830 9276
rect 2886 9274 2910 9276
rect 2966 9274 2990 9276
rect 3046 9274 3070 9276
rect 3126 9274 3132 9276
rect 2886 9222 2888 9274
rect 3068 9222 3070 9274
rect 2824 9220 2830 9222
rect 2886 9220 2910 9222
rect 2966 9220 2990 9222
rect 3046 9220 3070 9222
rect 3126 9220 3132 9222
rect 2824 9200 3132 9220
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 2824 8188 3132 8208
rect 2824 8186 2830 8188
rect 2886 8186 2910 8188
rect 2966 8186 2990 8188
rect 3046 8186 3070 8188
rect 3126 8186 3132 8188
rect 2886 8134 2888 8186
rect 3068 8134 3070 8186
rect 2824 8132 2830 8134
rect 2886 8132 2910 8134
rect 2966 8132 2990 8134
rect 3046 8132 3070 8134
rect 3126 8132 3132 8134
rect 2824 8112 3132 8132
rect 2824 7100 3132 7120
rect 2824 7098 2830 7100
rect 2886 7098 2910 7100
rect 2966 7098 2990 7100
rect 3046 7098 3070 7100
rect 3126 7098 3132 7100
rect 2886 7046 2888 7098
rect 3068 7046 3070 7098
rect 2824 7044 2830 7046
rect 2886 7044 2910 7046
rect 2966 7044 2990 7046
rect 3046 7044 3070 7046
rect 3126 7044 3132 7046
rect 2824 7024 3132 7044
rect 3160 6798 3188 8366
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3148 6656 3200 6662
rect 3148 6598 3200 6604
rect 2824 6012 3132 6032
rect 2824 6010 2830 6012
rect 2886 6010 2910 6012
rect 2966 6010 2990 6012
rect 3046 6010 3070 6012
rect 3126 6010 3132 6012
rect 2886 5958 2888 6010
rect 3068 5958 3070 6010
rect 2824 5956 2830 5958
rect 2886 5956 2910 5958
rect 2966 5956 2990 5958
rect 3046 5956 3070 5958
rect 3126 5956 3132 5958
rect 2824 5936 3132 5956
rect 3160 5234 3188 6598
rect 3148 5228 3200 5234
rect 3148 5170 3200 5176
rect 2824 4924 3132 4944
rect 2824 4922 2830 4924
rect 2886 4922 2910 4924
rect 2966 4922 2990 4924
rect 3046 4922 3070 4924
rect 3126 4922 3132 4924
rect 2886 4870 2888 4922
rect 3068 4870 3070 4922
rect 2824 4868 2830 4870
rect 2886 4868 2910 4870
rect 2966 4868 2990 4870
rect 3046 4868 3070 4870
rect 3126 4868 3132 4870
rect 2824 4848 3132 4868
rect 2824 3836 3132 3856
rect 2824 3834 2830 3836
rect 2886 3834 2910 3836
rect 2966 3834 2990 3836
rect 3046 3834 3070 3836
rect 3126 3834 3132 3836
rect 2886 3782 2888 3834
rect 3068 3782 3070 3834
rect 2824 3780 2830 3782
rect 2886 3780 2910 3782
rect 2966 3780 2990 3782
rect 3046 3780 3070 3782
rect 3126 3780 3132 3782
rect 2824 3760 3132 3780
rect 3252 3194 3280 9454
rect 3344 8498 3372 9590
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3436 8430 3464 9658
rect 3620 9178 3648 17138
rect 3792 17128 3844 17134
rect 3792 17070 3844 17076
rect 3804 12918 3832 17070
rect 3792 12912 3844 12918
rect 3792 12854 3844 12860
rect 3896 12714 3924 17206
rect 6196 17202 6224 17614
rect 6472 17338 6500 19200
rect 6460 17332 6512 17338
rect 6840 17320 6868 19200
rect 7300 17338 7328 19200
rect 7760 17338 7788 19200
rect 6920 17332 6972 17338
rect 6840 17292 6920 17320
rect 6460 17274 6512 17280
rect 6920 17274 6972 17280
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7748 17332 7800 17338
rect 8128 17320 8156 19200
rect 8588 19122 8616 19200
rect 8680 19122 8708 19230
rect 8588 19094 8708 19122
rect 8446 17436 8754 17456
rect 8446 17434 8452 17436
rect 8508 17434 8532 17436
rect 8588 17434 8612 17436
rect 8668 17434 8692 17436
rect 8748 17434 8754 17436
rect 8508 17382 8510 17434
rect 8690 17382 8692 17434
rect 8446 17380 8452 17382
rect 8508 17380 8532 17382
rect 8588 17380 8612 17382
rect 8668 17380 8692 17382
rect 8748 17380 8754 17382
rect 8446 17360 8754 17380
rect 8864 17338 8892 19230
rect 8942 19200 8998 20000
rect 9402 19200 9458 20000
rect 9770 19200 9826 20000
rect 10230 19200 10286 20000
rect 10690 19200 10746 20000
rect 11058 19200 11114 20000
rect 11518 19200 11574 20000
rect 11886 19200 11942 20000
rect 12346 19200 12402 20000
rect 12714 19200 12770 20000
rect 13174 19200 13230 20000
rect 13542 19200 13598 20000
rect 14002 19200 14058 20000
rect 14462 19200 14518 20000
rect 14830 19200 14886 20000
rect 15290 19200 15346 20000
rect 15658 19200 15714 20000
rect 16118 19200 16174 20000
rect 16486 19200 16542 20000
rect 16946 19200 17002 20000
rect 8300 17332 8352 17338
rect 8128 17292 8300 17320
rect 7748 17274 7800 17280
rect 8300 17274 8352 17280
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8956 17202 8984 19200
rect 9312 17604 9364 17610
rect 9312 17546 9364 17552
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9232 17202 9260 17478
rect 9324 17270 9352 17546
rect 9416 17338 9444 19200
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9312 17264 9364 17270
rect 9312 17206 9364 17212
rect 9784 17202 9812 19200
rect 10244 17338 10272 19200
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10704 17202 10732 19200
rect 10876 17672 10928 17678
rect 10876 17614 10928 17620
rect 4528 17196 4580 17202
rect 4528 17138 4580 17144
rect 5540 17196 5592 17202
rect 5540 17138 5592 17144
rect 5816 17196 5868 17202
rect 5816 17138 5868 17144
rect 6184 17196 6236 17202
rect 6184 17138 6236 17144
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 8208 17196 8260 17202
rect 8208 17138 8260 17144
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 9220 17196 9272 17202
rect 9220 17138 9272 17144
rect 9772 17196 9824 17202
rect 9772 17138 9824 17144
rect 10692 17196 10744 17202
rect 10692 17138 10744 17144
rect 4436 17128 4488 17134
rect 4436 17070 4488 17076
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 3976 16516 4028 16522
rect 3976 16458 4028 16464
rect 3884 12708 3936 12714
rect 3884 12650 3936 12656
rect 3988 9994 4016 16458
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 4080 12986 4108 16390
rect 4264 13326 4292 16526
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 4252 13320 4304 13326
rect 4252 13262 4304 13268
rect 4068 12980 4120 12986
rect 4068 12922 4120 12928
rect 4172 10810 4200 13262
rect 4448 11778 4476 17070
rect 4540 11898 4568 17138
rect 4698 16348 5006 16368
rect 4698 16346 4704 16348
rect 4760 16346 4784 16348
rect 4840 16346 4864 16348
rect 4920 16346 4944 16348
rect 5000 16346 5006 16348
rect 4760 16294 4762 16346
rect 4942 16294 4944 16346
rect 4698 16292 4704 16294
rect 4760 16292 4784 16294
rect 4840 16292 4864 16294
rect 4920 16292 4944 16294
rect 5000 16292 5006 16294
rect 4698 16272 5006 16292
rect 4620 15972 4672 15978
rect 4620 15914 4672 15920
rect 4632 13938 4660 15914
rect 4698 15260 5006 15280
rect 4698 15258 4704 15260
rect 4760 15258 4784 15260
rect 4840 15258 4864 15260
rect 4920 15258 4944 15260
rect 5000 15258 5006 15260
rect 4760 15206 4762 15258
rect 4942 15206 4944 15258
rect 4698 15204 4704 15206
rect 4760 15204 4784 15206
rect 4840 15204 4864 15206
rect 4920 15204 4944 15206
rect 5000 15204 5006 15206
rect 4698 15184 5006 15204
rect 4698 14172 5006 14192
rect 4698 14170 4704 14172
rect 4760 14170 4784 14172
rect 4840 14170 4864 14172
rect 4920 14170 4944 14172
rect 5000 14170 5006 14172
rect 4760 14118 4762 14170
rect 4942 14118 4944 14170
rect 4698 14116 4704 14118
rect 4760 14116 4784 14118
rect 4840 14116 4864 14118
rect 4920 14116 4944 14118
rect 5000 14116 5006 14118
rect 4698 14096 5006 14116
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4698 13084 5006 13104
rect 4698 13082 4704 13084
rect 4760 13082 4784 13084
rect 4840 13082 4864 13084
rect 4920 13082 4944 13084
rect 5000 13082 5006 13084
rect 4760 13030 4762 13082
rect 4942 13030 4944 13082
rect 4698 13028 4704 13030
rect 4760 13028 4784 13030
rect 4840 13028 4864 13030
rect 4920 13028 4944 13030
rect 5000 13028 5006 13030
rect 4698 13008 5006 13028
rect 4698 11996 5006 12016
rect 4698 11994 4704 11996
rect 4760 11994 4784 11996
rect 4840 11994 4864 11996
rect 4920 11994 4944 11996
rect 5000 11994 5006 11996
rect 4760 11942 4762 11994
rect 4942 11942 4944 11994
rect 4698 11940 4704 11942
rect 4760 11940 4784 11942
rect 4840 11940 4864 11942
rect 4920 11940 4944 11942
rect 5000 11940 5006 11942
rect 4698 11920 5006 11940
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4448 11750 4568 11778
rect 4344 11076 4396 11082
rect 4344 11018 4396 11024
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4356 10742 4384 11018
rect 4344 10736 4396 10742
rect 4344 10678 4396 10684
rect 3976 9988 4028 9994
rect 3976 9930 4028 9936
rect 4252 9512 4304 9518
rect 4252 9454 4304 9460
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 3608 9172 3660 9178
rect 3608 9114 3660 9120
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3608 7268 3660 7274
rect 3608 7210 3660 7216
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 2044 3052 2096 3058
rect 2044 2994 2096 3000
rect 2136 3052 2188 3058
rect 2136 2994 2188 3000
rect 1492 2304 1544 2310
rect 1492 2246 1544 2252
rect 1860 2304 1912 2310
rect 1860 2246 1912 2252
rect 1504 800 1532 2246
rect 1872 800 1900 2246
rect 2148 1737 2176 2994
rect 2824 2748 3132 2768
rect 2824 2746 2830 2748
rect 2886 2746 2910 2748
rect 2966 2746 2990 2748
rect 3046 2746 3070 2748
rect 3126 2746 3132 2748
rect 2886 2694 2888 2746
rect 3068 2694 3070 2746
rect 2824 2692 2830 2694
rect 2886 2692 2910 2694
rect 2966 2692 2990 2694
rect 3046 2692 3070 2694
rect 3126 2692 3132 2694
rect 2824 2672 3132 2692
rect 3620 2582 3648 7210
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 3126 4016 7142
rect 3976 3120 4028 3126
rect 3976 3062 4028 3068
rect 3608 2576 3660 2582
rect 2686 2544 2742 2553
rect 3608 2518 3660 2524
rect 4172 2514 4200 9386
rect 2686 2479 2742 2488
rect 4160 2508 4212 2514
rect 2700 2446 2728 2479
rect 4160 2450 4212 2456
rect 4264 2446 4292 9454
rect 4540 8838 4568 11750
rect 5448 11620 5500 11626
rect 5448 11562 5500 11568
rect 5264 11076 5316 11082
rect 5264 11018 5316 11024
rect 4698 10908 5006 10928
rect 4698 10906 4704 10908
rect 4760 10906 4784 10908
rect 4840 10906 4864 10908
rect 4920 10906 4944 10908
rect 5000 10906 5006 10908
rect 4760 10854 4762 10906
rect 4942 10854 4944 10906
rect 4698 10852 4704 10854
rect 4760 10852 4784 10854
rect 4840 10852 4864 10854
rect 4920 10852 4944 10854
rect 5000 10852 5006 10854
rect 4698 10832 5006 10852
rect 5080 10464 5132 10470
rect 5080 10406 5132 10412
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4724 10062 4752 10202
rect 4712 10056 4764 10062
rect 4712 9998 4764 10004
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4908 9908 4936 9998
rect 4632 9880 4936 9908
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4632 8480 4660 9880
rect 4698 9820 5006 9840
rect 4698 9818 4704 9820
rect 4760 9818 4784 9820
rect 4840 9818 4864 9820
rect 4920 9818 4944 9820
rect 5000 9818 5006 9820
rect 4760 9766 4762 9818
rect 4942 9766 4944 9818
rect 4698 9764 4704 9766
rect 4760 9764 4784 9766
rect 4840 9764 4864 9766
rect 4920 9764 4944 9766
rect 5000 9764 5006 9766
rect 4698 9744 5006 9764
rect 4698 8732 5006 8752
rect 4698 8730 4704 8732
rect 4760 8730 4784 8732
rect 4840 8730 4864 8732
rect 4920 8730 4944 8732
rect 5000 8730 5006 8732
rect 4760 8678 4762 8730
rect 4942 8678 4944 8730
rect 4698 8676 4704 8678
rect 4760 8676 4784 8678
rect 4840 8676 4864 8678
rect 4920 8676 4944 8678
rect 5000 8676 5006 8678
rect 4698 8656 5006 8676
rect 4448 8452 4660 8480
rect 4448 3346 4476 8452
rect 4698 7644 5006 7664
rect 4698 7642 4704 7644
rect 4760 7642 4784 7644
rect 4840 7642 4864 7644
rect 4920 7642 4944 7644
rect 5000 7642 5006 7644
rect 4760 7590 4762 7642
rect 4942 7590 4944 7642
rect 4698 7588 4704 7590
rect 4760 7588 4784 7590
rect 4840 7588 4864 7590
rect 4920 7588 4944 7590
rect 5000 7588 5006 7590
rect 4698 7568 5006 7588
rect 4528 7200 4580 7206
rect 4528 7142 4580 7148
rect 4540 3534 4568 7142
rect 4698 6556 5006 6576
rect 4698 6554 4704 6556
rect 4760 6554 4784 6556
rect 4840 6554 4864 6556
rect 4920 6554 4944 6556
rect 5000 6554 5006 6556
rect 4760 6502 4762 6554
rect 4942 6502 4944 6554
rect 4698 6500 4704 6502
rect 4760 6500 4784 6502
rect 4840 6500 4864 6502
rect 4920 6500 4944 6502
rect 5000 6500 5006 6502
rect 4698 6480 5006 6500
rect 4698 5468 5006 5488
rect 4698 5466 4704 5468
rect 4760 5466 4784 5468
rect 4840 5466 4864 5468
rect 4920 5466 4944 5468
rect 5000 5466 5006 5468
rect 4760 5414 4762 5466
rect 4942 5414 4944 5466
rect 4698 5412 4704 5414
rect 4760 5412 4784 5414
rect 4840 5412 4864 5414
rect 4920 5412 4944 5414
rect 5000 5412 5006 5414
rect 4698 5392 5006 5412
rect 4698 4380 5006 4400
rect 4698 4378 4704 4380
rect 4760 4378 4784 4380
rect 4840 4378 4864 4380
rect 4920 4378 4944 4380
rect 5000 4378 5006 4380
rect 4760 4326 4762 4378
rect 4942 4326 4944 4378
rect 4698 4324 4704 4326
rect 4760 4324 4784 4326
rect 4840 4324 4864 4326
rect 4920 4324 4944 4326
rect 5000 4324 5006 4326
rect 4698 4304 5006 4324
rect 4528 3528 4580 3534
rect 4528 3470 4580 3476
rect 4448 3318 4568 3346
rect 2688 2440 2740 2446
rect 2688 2382 2740 2388
rect 4252 2440 4304 2446
rect 4252 2382 4304 2388
rect 2320 2304 2372 2310
rect 2320 2246 2372 2252
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 3148 2304 3200 2310
rect 3148 2246 3200 2252
rect 3608 2304 3660 2310
rect 3608 2246 3660 2252
rect 4068 2304 4120 2310
rect 4068 2246 4120 2252
rect 4436 2304 4488 2310
rect 4436 2246 4488 2252
rect 2134 1728 2190 1737
rect 2134 1663 2190 1672
rect 2332 800 2360 2246
rect 2792 800 2820 2246
rect 3160 800 3188 2246
rect 3620 800 3648 2246
rect 4080 800 4108 2246
rect 4448 800 4476 2246
rect 4540 1698 4568 3318
rect 4698 3292 5006 3312
rect 4698 3290 4704 3292
rect 4760 3290 4784 3292
rect 4840 3290 4864 3292
rect 4920 3290 4944 3292
rect 5000 3290 5006 3292
rect 4760 3238 4762 3290
rect 4942 3238 4944 3290
rect 4698 3236 4704 3238
rect 4760 3236 4784 3238
rect 4840 3236 4864 3238
rect 4920 3236 4944 3238
rect 5000 3236 5006 3238
rect 4698 3216 5006 3236
rect 5092 2650 5120 10406
rect 5172 9920 5224 9926
rect 5172 9862 5224 9868
rect 5184 9722 5212 9862
rect 5172 9716 5224 9722
rect 5172 9658 5224 9664
rect 5276 7886 5304 11018
rect 5460 10130 5488 11562
rect 5552 10538 5580 17138
rect 5828 16726 5856 17138
rect 5816 16720 5868 16726
rect 5816 16662 5868 16668
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6092 12776 6144 12782
rect 6092 12718 6144 12724
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5644 10674 5672 10950
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5540 10532 5592 10538
rect 5540 10474 5592 10480
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5448 10124 5500 10130
rect 5448 10066 5500 10072
rect 5736 9761 5764 10406
rect 5920 10130 5948 11494
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5722 9752 5778 9761
rect 5448 9716 5500 9722
rect 5828 9722 5856 10066
rect 5722 9687 5778 9696
rect 5816 9716 5868 9722
rect 5448 9658 5500 9664
rect 5816 9658 5868 9664
rect 5264 7880 5316 7886
rect 5264 7822 5316 7828
rect 5460 7410 5488 9658
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5828 9042 5856 9522
rect 5816 9036 5868 9042
rect 5816 8978 5868 8984
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5632 7200 5684 7206
rect 5632 7142 5684 7148
rect 5080 2644 5132 2650
rect 5080 2586 5132 2592
rect 5264 2644 5316 2650
rect 5264 2586 5316 2592
rect 5276 2446 5304 2586
rect 5644 2582 5672 7142
rect 5632 2576 5684 2582
rect 5632 2518 5684 2524
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 4632 1873 4660 2382
rect 6012 2378 6040 10406
rect 6104 8362 6132 12718
rect 6196 10674 6224 16594
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6196 10198 6224 10474
rect 6184 10192 6236 10198
rect 6184 10134 6236 10140
rect 6092 8356 6144 8362
rect 6092 8298 6144 8304
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6000 2372 6052 2378
rect 6000 2314 6052 2320
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 5356 2304 5408 2310
rect 5356 2246 5408 2252
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 4698 2204 5006 2224
rect 4698 2202 4704 2204
rect 4760 2202 4784 2204
rect 4840 2202 4864 2204
rect 4920 2202 4944 2204
rect 5000 2202 5006 2204
rect 4760 2150 4762 2202
rect 4942 2150 4944 2202
rect 4698 2148 4704 2150
rect 4760 2148 4784 2150
rect 4840 2148 4864 2150
rect 4920 2148 4944 2150
rect 5000 2148 5006 2150
rect 4698 2128 5006 2148
rect 4618 1864 4674 1873
rect 4618 1799 4674 1808
rect 4528 1692 4580 1698
rect 4528 1634 4580 1640
rect 5092 1170 5120 2246
rect 4908 1142 5120 1170
rect 4908 800 4936 1142
rect 5368 800 5396 2246
rect 5736 800 5764 2246
rect 6104 2106 6132 2382
rect 6184 2304 6236 2310
rect 6184 2246 6236 2252
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 6196 800 6224 2246
rect 6288 1766 6316 10610
rect 6380 10033 6408 17138
rect 7104 17128 7156 17134
rect 7104 17070 7156 17076
rect 7840 17128 7892 17134
rect 7840 17070 7892 17076
rect 6572 16892 6880 16912
rect 6572 16890 6578 16892
rect 6634 16890 6658 16892
rect 6714 16890 6738 16892
rect 6794 16890 6818 16892
rect 6874 16890 6880 16892
rect 6634 16838 6636 16890
rect 6816 16838 6818 16890
rect 6572 16836 6578 16838
rect 6634 16836 6658 16838
rect 6714 16836 6738 16838
rect 6794 16836 6818 16838
rect 6874 16836 6880 16838
rect 6572 16816 6880 16836
rect 6572 15804 6880 15824
rect 6572 15802 6578 15804
rect 6634 15802 6658 15804
rect 6714 15802 6738 15804
rect 6794 15802 6818 15804
rect 6874 15802 6880 15804
rect 6634 15750 6636 15802
rect 6816 15750 6818 15802
rect 6572 15748 6578 15750
rect 6634 15748 6658 15750
rect 6714 15748 6738 15750
rect 6794 15748 6818 15750
rect 6874 15748 6880 15750
rect 6572 15728 6880 15748
rect 6572 14716 6880 14736
rect 6572 14714 6578 14716
rect 6634 14714 6658 14716
rect 6714 14714 6738 14716
rect 6794 14714 6818 14716
rect 6874 14714 6880 14716
rect 6634 14662 6636 14714
rect 6816 14662 6818 14714
rect 6572 14660 6578 14662
rect 6634 14660 6658 14662
rect 6714 14660 6738 14662
rect 6794 14660 6818 14662
rect 6874 14660 6880 14662
rect 6572 14640 6880 14660
rect 6572 13628 6880 13648
rect 6572 13626 6578 13628
rect 6634 13626 6658 13628
rect 6714 13626 6738 13628
rect 6794 13626 6818 13628
rect 6874 13626 6880 13628
rect 6634 13574 6636 13626
rect 6816 13574 6818 13626
rect 6572 13572 6578 13574
rect 6634 13572 6658 13574
rect 6714 13572 6738 13574
rect 6794 13572 6818 13574
rect 6874 13572 6880 13574
rect 6572 13552 6880 13572
rect 7116 12986 7144 17070
rect 7104 12980 7156 12986
rect 7104 12922 7156 12928
rect 7380 12844 7432 12850
rect 7380 12786 7432 12792
rect 6572 12540 6880 12560
rect 6572 12538 6578 12540
rect 6634 12538 6658 12540
rect 6714 12538 6738 12540
rect 6794 12538 6818 12540
rect 6874 12538 6880 12540
rect 6634 12486 6636 12538
rect 6816 12486 6818 12538
rect 6572 12484 6578 12486
rect 6634 12484 6658 12486
rect 6714 12484 6738 12486
rect 6794 12484 6818 12486
rect 6874 12484 6880 12486
rect 6572 12464 6880 12484
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6572 11452 6880 11472
rect 6572 11450 6578 11452
rect 6634 11450 6658 11452
rect 6714 11450 6738 11452
rect 6794 11450 6818 11452
rect 6874 11450 6880 11452
rect 6634 11398 6636 11450
rect 6816 11398 6818 11450
rect 6572 11396 6578 11398
rect 6634 11396 6658 11398
rect 6714 11396 6738 11398
rect 6794 11396 6818 11398
rect 6874 11396 6880 11398
rect 6572 11376 6880 11396
rect 6460 11348 6512 11354
rect 6460 11290 6512 11296
rect 6472 10266 6500 11290
rect 6572 10364 6880 10384
rect 6572 10362 6578 10364
rect 6634 10362 6658 10364
rect 6714 10362 6738 10364
rect 6794 10362 6818 10364
rect 6874 10362 6880 10364
rect 6634 10310 6636 10362
rect 6816 10310 6818 10362
rect 6572 10308 6578 10310
rect 6634 10308 6658 10310
rect 6714 10308 6738 10310
rect 6794 10308 6818 10310
rect 6874 10308 6880 10310
rect 6572 10288 6880 10308
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6366 10024 6422 10033
rect 6366 9959 6422 9968
rect 6368 9716 6420 9722
rect 6932 9674 6960 11562
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6368 9658 6420 9664
rect 6380 8974 6408 9658
rect 6656 9646 6960 9674
rect 6656 9450 6684 9646
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6572 9276 6880 9296
rect 6572 9274 6578 9276
rect 6634 9274 6658 9276
rect 6714 9274 6738 9276
rect 6794 9274 6818 9276
rect 6874 9274 6880 9276
rect 6634 9222 6636 9274
rect 6816 9222 6818 9274
rect 6572 9220 6578 9222
rect 6634 9220 6658 9222
rect 6714 9220 6738 9222
rect 6794 9220 6818 9222
rect 6874 9220 6880 9222
rect 6572 9200 6880 9220
rect 7024 8974 7052 10542
rect 7116 10266 7144 10950
rect 7288 10668 7340 10674
rect 7288 10610 7340 10616
rect 7104 10260 7156 10266
rect 7104 10202 7156 10208
rect 7196 9920 7248 9926
rect 7196 9862 7248 9868
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 7012 8968 7064 8974
rect 7012 8910 7064 8916
rect 6380 8634 6408 8910
rect 6920 8900 6972 8906
rect 6920 8842 6972 8848
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6572 8188 6880 8208
rect 6572 8186 6578 8188
rect 6634 8186 6658 8188
rect 6714 8186 6738 8188
rect 6794 8186 6818 8188
rect 6874 8186 6880 8188
rect 6634 8134 6636 8186
rect 6816 8134 6818 8186
rect 6572 8132 6578 8134
rect 6634 8132 6658 8134
rect 6714 8132 6738 8134
rect 6794 8132 6818 8134
rect 6874 8132 6880 8134
rect 6572 8112 6880 8132
rect 6572 7100 6880 7120
rect 6572 7098 6578 7100
rect 6634 7098 6658 7100
rect 6714 7098 6738 7100
rect 6794 7098 6818 7100
rect 6874 7098 6880 7100
rect 6634 7046 6636 7098
rect 6816 7046 6818 7098
rect 6572 7044 6578 7046
rect 6634 7044 6658 7046
rect 6714 7044 6738 7046
rect 6794 7044 6818 7046
rect 6874 7044 6880 7046
rect 6572 7024 6880 7044
rect 6572 6012 6880 6032
rect 6572 6010 6578 6012
rect 6634 6010 6658 6012
rect 6714 6010 6738 6012
rect 6794 6010 6818 6012
rect 6874 6010 6880 6012
rect 6634 5958 6636 6010
rect 6816 5958 6818 6010
rect 6572 5956 6578 5958
rect 6634 5956 6658 5958
rect 6714 5956 6738 5958
rect 6794 5956 6818 5958
rect 6874 5956 6880 5958
rect 6572 5936 6880 5956
rect 6572 4924 6880 4944
rect 6572 4922 6578 4924
rect 6634 4922 6658 4924
rect 6714 4922 6738 4924
rect 6794 4922 6818 4924
rect 6874 4922 6880 4924
rect 6634 4870 6636 4922
rect 6816 4870 6818 4922
rect 6572 4868 6578 4870
rect 6634 4868 6658 4870
rect 6714 4868 6738 4870
rect 6794 4868 6818 4870
rect 6874 4868 6880 4870
rect 6572 4848 6880 4868
rect 6572 3836 6880 3856
rect 6572 3834 6578 3836
rect 6634 3834 6658 3836
rect 6714 3834 6738 3836
rect 6794 3834 6818 3836
rect 6874 3834 6880 3836
rect 6634 3782 6636 3834
rect 6816 3782 6818 3834
rect 6572 3780 6578 3782
rect 6634 3780 6658 3782
rect 6714 3780 6738 3782
rect 6794 3780 6818 3782
rect 6874 3780 6880 3782
rect 6572 3760 6880 3780
rect 6572 2748 6880 2768
rect 6572 2746 6578 2748
rect 6634 2746 6658 2748
rect 6714 2746 6738 2748
rect 6794 2746 6818 2748
rect 6874 2746 6880 2748
rect 6634 2694 6636 2746
rect 6816 2694 6818 2746
rect 6572 2692 6578 2694
rect 6634 2692 6658 2694
rect 6714 2692 6738 2694
rect 6794 2692 6818 2694
rect 6874 2692 6880 2694
rect 6572 2672 6880 2692
rect 6644 2440 6696 2446
rect 6642 2408 6644 2417
rect 6696 2408 6698 2417
rect 6642 2343 6698 2352
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6276 1760 6328 1766
rect 6276 1702 6328 1708
rect 6656 800 6684 2246
rect 6932 1630 6960 8842
rect 7024 8294 7052 8910
rect 7116 8498 7144 9522
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 7024 7954 7052 8230
rect 7208 8090 7236 9862
rect 7300 9178 7328 10610
rect 7392 9654 7420 12786
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7472 11756 7524 11762
rect 7472 11698 7524 11704
rect 7380 9648 7432 9654
rect 7380 9590 7432 9596
rect 7484 9178 7512 11698
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7576 10810 7604 11630
rect 7564 10804 7616 10810
rect 7564 10746 7616 10752
rect 7668 10690 7696 12582
rect 7852 10742 7880 17070
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 7932 11280 7984 11286
rect 7932 11222 7984 11228
rect 7576 10662 7696 10690
rect 7748 10736 7800 10742
rect 7748 10678 7800 10684
rect 7840 10736 7892 10742
rect 7840 10678 7892 10684
rect 7576 10130 7604 10662
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7472 9172 7524 9178
rect 7472 9114 7524 9120
rect 7576 8090 7604 10066
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7668 9489 7696 9522
rect 7654 9480 7710 9489
rect 7654 9415 7710 9424
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7564 8084 7616 8090
rect 7564 8026 7616 8032
rect 7012 7948 7064 7954
rect 7012 7890 7064 7896
rect 7288 2440 7340 2446
rect 7288 2382 7340 2388
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6920 1624 6972 1630
rect 6920 1566 6972 1572
rect 7024 800 7052 2246
rect 7300 2106 7328 2382
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7484 800 7512 2246
rect 7760 1902 7788 10678
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 7852 8566 7880 9318
rect 7840 8560 7892 8566
rect 7840 8502 7892 8508
rect 7852 7954 7880 8502
rect 7840 7948 7892 7954
rect 7840 7890 7892 7896
rect 7944 7818 7972 11222
rect 8036 10130 8064 13126
rect 8116 11756 8168 11762
rect 8116 11698 8168 11704
rect 8024 10124 8076 10130
rect 8024 10066 8076 10072
rect 8036 9382 8064 10066
rect 8024 9376 8076 9382
rect 8024 9318 8076 9324
rect 8036 8906 8064 9318
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7932 7812 7984 7818
rect 7932 7754 7984 7760
rect 7838 2544 7894 2553
rect 7838 2479 7894 2488
rect 7852 2446 7880 2479
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 7932 2304 7984 2310
rect 7932 2246 7984 2252
rect 7748 1896 7800 1902
rect 7748 1838 7800 1844
rect 7944 800 7972 2246
rect 8128 1601 8156 11698
rect 8220 10577 8248 17138
rect 8852 16992 8904 16998
rect 8852 16934 8904 16940
rect 8446 16348 8754 16368
rect 8446 16346 8452 16348
rect 8508 16346 8532 16348
rect 8588 16346 8612 16348
rect 8668 16346 8692 16348
rect 8748 16346 8754 16348
rect 8508 16294 8510 16346
rect 8690 16294 8692 16346
rect 8446 16292 8452 16294
rect 8508 16292 8532 16294
rect 8588 16292 8612 16294
rect 8668 16292 8692 16294
rect 8748 16292 8754 16294
rect 8446 16272 8754 16292
rect 8446 15260 8754 15280
rect 8446 15258 8452 15260
rect 8508 15258 8532 15260
rect 8588 15258 8612 15260
rect 8668 15258 8692 15260
rect 8748 15258 8754 15260
rect 8508 15206 8510 15258
rect 8690 15206 8692 15258
rect 8446 15204 8452 15206
rect 8508 15204 8532 15206
rect 8588 15204 8612 15206
rect 8668 15204 8692 15206
rect 8748 15204 8754 15206
rect 8446 15184 8754 15204
rect 8864 14770 8892 16934
rect 8956 16794 8984 17138
rect 9404 17128 9456 17134
rect 9404 17070 9456 17076
rect 9496 17128 9548 17134
rect 9496 17070 9548 17076
rect 9036 17060 9088 17066
rect 9036 17002 9088 17008
rect 8944 16788 8996 16794
rect 8944 16730 8996 16736
rect 8864 14742 8984 14770
rect 8446 14172 8754 14192
rect 8446 14170 8452 14172
rect 8508 14170 8532 14172
rect 8588 14170 8612 14172
rect 8668 14170 8692 14172
rect 8748 14170 8754 14172
rect 8508 14118 8510 14170
rect 8690 14118 8692 14170
rect 8446 14116 8452 14118
rect 8508 14116 8532 14118
rect 8588 14116 8612 14118
rect 8668 14116 8692 14118
rect 8748 14116 8754 14118
rect 8446 14096 8754 14116
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8446 13084 8754 13104
rect 8446 13082 8452 13084
rect 8508 13082 8532 13084
rect 8588 13082 8612 13084
rect 8668 13082 8692 13084
rect 8748 13082 8754 13084
rect 8508 13030 8510 13082
rect 8690 13030 8692 13082
rect 8446 13028 8452 13030
rect 8508 13028 8532 13030
rect 8588 13028 8612 13030
rect 8668 13028 8692 13030
rect 8748 13028 8754 13030
rect 8446 13008 8754 13028
rect 8864 12782 8892 13670
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8852 12776 8904 12782
rect 8852 12718 8904 12724
rect 8206 10568 8262 10577
rect 8206 10503 8262 10512
rect 8312 10146 8340 12718
rect 8446 11996 8754 12016
rect 8446 11994 8452 11996
rect 8508 11994 8532 11996
rect 8588 11994 8612 11996
rect 8668 11994 8692 11996
rect 8748 11994 8754 11996
rect 8508 11942 8510 11994
rect 8690 11942 8692 11994
rect 8446 11940 8452 11942
rect 8508 11940 8532 11942
rect 8588 11940 8612 11942
rect 8668 11940 8692 11942
rect 8748 11940 8754 11942
rect 8446 11920 8754 11940
rect 8446 10908 8754 10928
rect 8446 10906 8452 10908
rect 8508 10906 8532 10908
rect 8588 10906 8612 10908
rect 8668 10906 8692 10908
rect 8748 10906 8754 10908
rect 8508 10854 8510 10906
rect 8690 10854 8692 10906
rect 8446 10852 8452 10854
rect 8508 10852 8532 10854
rect 8588 10852 8612 10854
rect 8668 10852 8692 10854
rect 8748 10852 8754 10854
rect 8446 10832 8754 10852
rect 8864 10470 8892 12718
rect 8852 10464 8904 10470
rect 8852 10406 8904 10412
rect 8956 10248 8984 14742
rect 9048 10266 9076 17002
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9128 11348 9180 11354
rect 9128 11290 9180 11296
rect 8220 10118 8340 10146
rect 8864 10220 8984 10248
rect 9036 10260 9088 10266
rect 8220 9926 8248 10118
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8208 9920 8260 9926
rect 8208 9862 8260 9868
rect 8220 9602 8248 9862
rect 8312 9722 8340 9998
rect 8446 9820 8754 9840
rect 8446 9818 8452 9820
rect 8508 9818 8532 9820
rect 8588 9818 8612 9820
rect 8668 9818 8692 9820
rect 8748 9818 8754 9820
rect 8508 9766 8510 9818
rect 8690 9766 8692 9818
rect 8446 9764 8452 9766
rect 8508 9764 8532 9766
rect 8588 9764 8612 9766
rect 8668 9764 8692 9766
rect 8748 9764 8754 9766
rect 8446 9744 8754 9764
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8864 9654 8892 10220
rect 9036 10202 9088 10208
rect 9140 10146 9168 11290
rect 9232 10826 9260 16458
rect 9324 11014 9352 16934
rect 9416 12986 9444 17070
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9508 11354 9536 17070
rect 10048 16992 10100 16998
rect 10048 16934 10100 16940
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9588 12844 9640 12850
rect 9588 12786 9640 12792
rect 9496 11348 9548 11354
rect 9496 11290 9548 11296
rect 9496 11212 9548 11218
rect 9496 11154 9548 11160
rect 9312 11008 9364 11014
rect 9312 10950 9364 10956
rect 9404 11008 9456 11014
rect 9404 10950 9456 10956
rect 9416 10826 9444 10950
rect 9232 10798 9444 10826
rect 9312 10600 9364 10606
rect 9312 10542 9364 10548
rect 8956 10118 9260 10146
rect 8760 9648 8812 9654
rect 8220 9574 8340 9602
rect 8760 9590 8812 9596
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8312 9466 8340 9574
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8220 8498 8248 9454
rect 8312 9438 8432 9466
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8208 8492 8260 8498
rect 8208 8434 8260 8440
rect 8220 8294 8248 8434
rect 8208 8288 8260 8294
rect 8208 8230 8260 8236
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8220 2009 8248 8026
rect 8312 2650 8340 9318
rect 8404 8945 8432 9438
rect 8496 9110 8524 9522
rect 8772 9450 8800 9590
rect 8852 9512 8904 9518
rect 8852 9454 8904 9460
rect 8760 9444 8812 9450
rect 8760 9386 8812 9392
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8390 8936 8446 8945
rect 8390 8871 8446 8880
rect 8446 8732 8754 8752
rect 8446 8730 8452 8732
rect 8508 8730 8532 8732
rect 8588 8730 8612 8732
rect 8668 8730 8692 8732
rect 8748 8730 8754 8732
rect 8508 8678 8510 8730
rect 8690 8678 8692 8730
rect 8446 8676 8452 8678
rect 8508 8676 8532 8678
rect 8588 8676 8612 8678
rect 8668 8676 8692 8678
rect 8748 8676 8754 8678
rect 8446 8656 8754 8676
rect 8864 8634 8892 9454
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 8446 7644 8754 7664
rect 8446 7642 8452 7644
rect 8508 7642 8532 7644
rect 8588 7642 8612 7644
rect 8668 7642 8692 7644
rect 8748 7642 8754 7644
rect 8508 7590 8510 7642
rect 8690 7590 8692 7642
rect 8446 7588 8452 7590
rect 8508 7588 8532 7590
rect 8588 7588 8612 7590
rect 8668 7588 8692 7590
rect 8748 7588 8754 7590
rect 8446 7568 8754 7588
rect 8446 6556 8754 6576
rect 8446 6554 8452 6556
rect 8508 6554 8532 6556
rect 8588 6554 8612 6556
rect 8668 6554 8692 6556
rect 8748 6554 8754 6556
rect 8508 6502 8510 6554
rect 8690 6502 8692 6554
rect 8446 6500 8452 6502
rect 8508 6500 8532 6502
rect 8588 6500 8612 6502
rect 8668 6500 8692 6502
rect 8748 6500 8754 6502
rect 8446 6480 8754 6500
rect 8446 5468 8754 5488
rect 8446 5466 8452 5468
rect 8508 5466 8532 5468
rect 8588 5466 8612 5468
rect 8668 5466 8692 5468
rect 8748 5466 8754 5468
rect 8508 5414 8510 5466
rect 8690 5414 8692 5466
rect 8446 5412 8452 5414
rect 8508 5412 8532 5414
rect 8588 5412 8612 5414
rect 8668 5412 8692 5414
rect 8748 5412 8754 5414
rect 8446 5392 8754 5412
rect 8446 4380 8754 4400
rect 8446 4378 8452 4380
rect 8508 4378 8532 4380
rect 8588 4378 8612 4380
rect 8668 4378 8692 4380
rect 8748 4378 8754 4380
rect 8508 4326 8510 4378
rect 8690 4326 8692 4378
rect 8446 4324 8452 4326
rect 8508 4324 8532 4326
rect 8588 4324 8612 4326
rect 8668 4324 8692 4326
rect 8748 4324 8754 4326
rect 8446 4304 8754 4324
rect 8446 3292 8754 3312
rect 8446 3290 8452 3292
rect 8508 3290 8532 3292
rect 8588 3290 8612 3292
rect 8668 3290 8692 3292
rect 8748 3290 8754 3292
rect 8508 3238 8510 3290
rect 8690 3238 8692 3290
rect 8446 3236 8452 3238
rect 8508 3236 8532 3238
rect 8588 3236 8612 3238
rect 8668 3236 8692 3238
rect 8748 3236 8754 3238
rect 8446 3216 8754 3236
rect 8760 2848 8812 2854
rect 8760 2790 8812 2796
rect 8666 2680 8722 2689
rect 8300 2644 8352 2650
rect 8666 2615 8722 2624
rect 8300 2586 8352 2592
rect 8680 2446 8708 2615
rect 8668 2440 8720 2446
rect 8772 2428 8800 2790
rect 8864 2650 8892 8570
rect 8956 7410 8984 10118
rect 9232 10062 9260 10118
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9220 10056 9272 10062
rect 9220 9998 9272 10004
rect 9036 9920 9088 9926
rect 9036 9862 9088 9868
rect 9048 9042 9076 9862
rect 9140 9761 9168 9998
rect 9220 9920 9272 9926
rect 9220 9862 9272 9868
rect 9126 9752 9182 9761
rect 9126 9687 9182 9696
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9036 9036 9088 9042
rect 9036 8978 9088 8984
rect 9034 8936 9090 8945
rect 9034 8871 9090 8880
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 9048 7290 9076 8871
rect 9140 7546 9168 9590
rect 9232 7886 9260 9862
rect 9324 9722 9352 10542
rect 9312 9716 9364 9722
rect 9312 9658 9364 9664
rect 9312 9512 9364 9518
rect 9310 9480 9312 9489
rect 9364 9480 9366 9489
rect 9310 9415 9366 9424
rect 9416 9058 9444 10798
rect 9508 10674 9536 11154
rect 9496 10668 9548 10674
rect 9496 10610 9548 10616
rect 9508 10130 9536 10610
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9324 9030 9444 9058
rect 9508 9042 9536 10066
rect 9600 9926 9628 12786
rect 9680 11076 9732 11082
rect 9680 11018 9732 11024
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9496 9036 9548 9042
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 9324 7410 9352 9030
rect 9496 8978 9548 8984
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9312 7404 9364 7410
rect 9312 7346 9364 7352
rect 8956 7262 9076 7290
rect 8852 2644 8904 2650
rect 8852 2586 8904 2592
rect 8852 2440 8904 2446
rect 8772 2400 8852 2428
rect 8668 2382 8720 2388
rect 8852 2382 8904 2388
rect 8300 2304 8352 2310
rect 8300 2246 8352 2252
rect 8206 2000 8262 2009
rect 8206 1935 8262 1944
rect 8114 1592 8170 1601
rect 8114 1527 8170 1536
rect 8312 800 8340 2246
rect 8446 2204 8754 2224
rect 8446 2202 8452 2204
rect 8508 2202 8532 2204
rect 8588 2202 8612 2204
rect 8668 2202 8692 2204
rect 8748 2202 8754 2204
rect 8508 2150 8510 2202
rect 8690 2150 8692 2202
rect 8446 2148 8452 2150
rect 8508 2148 8532 2150
rect 8588 2148 8612 2150
rect 8668 2148 8692 2150
rect 8748 2148 8754 2150
rect 8446 2128 8754 2148
rect 8864 1850 8892 2382
rect 8956 2378 8984 7262
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9048 2514 9076 7142
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9036 2508 9088 2514
rect 9036 2450 9088 2456
rect 9232 2446 9260 2790
rect 9416 2582 9444 8842
rect 9600 2990 9628 9862
rect 9692 8566 9720 11018
rect 9864 10464 9916 10470
rect 9864 10406 9916 10412
rect 9876 10198 9904 10406
rect 9968 10266 9996 16662
rect 10060 12434 10088 16934
rect 10320 16892 10628 16912
rect 10320 16890 10326 16892
rect 10382 16890 10406 16892
rect 10462 16890 10486 16892
rect 10542 16890 10566 16892
rect 10622 16890 10628 16892
rect 10382 16838 10384 16890
rect 10564 16838 10566 16890
rect 10320 16836 10326 16838
rect 10382 16836 10406 16838
rect 10462 16836 10486 16838
rect 10542 16836 10566 16838
rect 10622 16836 10628 16838
rect 10320 16816 10628 16836
rect 10704 16794 10732 17138
rect 10784 16992 10836 16998
rect 10784 16934 10836 16940
rect 10692 16788 10744 16794
rect 10692 16730 10744 16736
rect 10320 15804 10628 15824
rect 10320 15802 10326 15804
rect 10382 15802 10406 15804
rect 10462 15802 10486 15804
rect 10542 15802 10566 15804
rect 10622 15802 10628 15804
rect 10382 15750 10384 15802
rect 10564 15750 10566 15802
rect 10320 15748 10326 15750
rect 10382 15748 10406 15750
rect 10462 15748 10486 15750
rect 10542 15748 10566 15750
rect 10622 15748 10628 15750
rect 10320 15728 10628 15748
rect 10320 14716 10628 14736
rect 10320 14714 10326 14716
rect 10382 14714 10406 14716
rect 10462 14714 10486 14716
rect 10542 14714 10566 14716
rect 10622 14714 10628 14716
rect 10382 14662 10384 14714
rect 10564 14662 10566 14714
rect 10320 14660 10326 14662
rect 10382 14660 10406 14662
rect 10462 14660 10486 14662
rect 10542 14660 10566 14662
rect 10622 14660 10628 14662
rect 10320 14640 10628 14660
rect 10320 13628 10628 13648
rect 10320 13626 10326 13628
rect 10382 13626 10406 13628
rect 10462 13626 10486 13628
rect 10542 13626 10566 13628
rect 10622 13626 10628 13628
rect 10382 13574 10384 13626
rect 10564 13574 10566 13626
rect 10320 13572 10326 13574
rect 10382 13572 10406 13574
rect 10462 13572 10486 13574
rect 10542 13572 10566 13574
rect 10622 13572 10628 13574
rect 10320 13552 10628 13572
rect 10232 12912 10284 12918
rect 10232 12854 10284 12860
rect 10060 12406 10180 12434
rect 10152 10674 10180 12406
rect 10244 10810 10272 12854
rect 10320 12540 10628 12560
rect 10320 12538 10326 12540
rect 10382 12538 10406 12540
rect 10462 12538 10486 12540
rect 10542 12538 10566 12540
rect 10622 12538 10628 12540
rect 10382 12486 10384 12538
rect 10564 12486 10566 12538
rect 10320 12484 10326 12486
rect 10382 12484 10406 12486
rect 10462 12484 10486 12486
rect 10542 12484 10566 12486
rect 10622 12484 10628 12486
rect 10320 12464 10628 12484
rect 10320 11452 10628 11472
rect 10320 11450 10326 11452
rect 10382 11450 10406 11452
rect 10462 11450 10486 11452
rect 10542 11450 10566 11452
rect 10622 11450 10628 11452
rect 10382 11398 10384 11450
rect 10564 11398 10566 11450
rect 10320 11396 10326 11398
rect 10382 11396 10406 11398
rect 10462 11396 10486 11398
rect 10542 11396 10566 11398
rect 10622 11396 10628 11398
rect 10320 11376 10628 11396
rect 10232 10804 10284 10810
rect 10232 10746 10284 10752
rect 10692 10804 10744 10810
rect 10692 10746 10744 10752
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9864 10192 9916 10198
rect 9864 10134 9916 10140
rect 10048 10192 10100 10198
rect 10048 10134 10100 10140
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9680 8560 9732 8566
rect 9680 8502 9732 8508
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9494 2680 9550 2689
rect 9494 2615 9550 2624
rect 9404 2576 9456 2582
rect 9404 2518 9456 2524
rect 9220 2440 9272 2446
rect 9220 2382 9272 2388
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 9128 2304 9180 2310
rect 9128 2246 9180 2252
rect 9140 2038 9168 2246
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 8772 1822 8892 1850
rect 8772 800 8800 1822
rect 9232 800 9260 2382
rect 9312 2304 9364 2310
rect 9508 2281 9536 2615
rect 9680 2440 9732 2446
rect 9600 2400 9680 2428
rect 9312 2246 9364 2252
rect 9494 2272 9550 2281
rect 9324 1698 9352 2246
rect 9494 2207 9550 2216
rect 9312 1692 9364 1698
rect 9312 1634 9364 1640
rect 9600 800 9628 2400
rect 9680 2382 9732 2388
rect 9784 1834 9812 9930
rect 9956 9920 10008 9926
rect 9956 9862 10008 9868
rect 9864 9444 9916 9450
rect 9864 9386 9916 9392
rect 9876 8838 9904 9386
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9876 2650 9904 8570
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9968 2530 9996 9862
rect 9876 2514 9996 2530
rect 9864 2508 9996 2514
rect 9916 2502 9996 2508
rect 10060 2530 10088 10134
rect 10152 7478 10180 10610
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 10244 9722 10272 10542
rect 10320 10364 10628 10384
rect 10320 10362 10326 10364
rect 10382 10362 10406 10364
rect 10462 10362 10486 10364
rect 10542 10362 10566 10364
rect 10622 10362 10628 10364
rect 10382 10310 10384 10362
rect 10564 10310 10566 10362
rect 10320 10308 10326 10310
rect 10382 10308 10406 10310
rect 10462 10308 10486 10310
rect 10542 10308 10566 10310
rect 10622 10308 10628 10310
rect 10320 10288 10628 10308
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10232 9376 10284 9382
rect 10232 9318 10284 9324
rect 10140 7472 10192 7478
rect 10140 7414 10192 7420
rect 10060 2502 10180 2530
rect 9864 2450 9916 2456
rect 10048 2372 10100 2378
rect 10048 2314 10100 2320
rect 9772 1828 9824 1834
rect 9772 1770 9824 1776
rect 10060 800 10088 2314
rect 10152 1970 10180 2502
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 10244 1873 10272 9318
rect 10320 9276 10628 9296
rect 10320 9274 10326 9276
rect 10382 9274 10406 9276
rect 10462 9274 10486 9276
rect 10542 9274 10566 9276
rect 10622 9274 10628 9276
rect 10382 9222 10384 9274
rect 10564 9222 10566 9274
rect 10320 9220 10326 9222
rect 10382 9220 10406 9222
rect 10462 9220 10486 9222
rect 10542 9220 10566 9222
rect 10622 9220 10628 9222
rect 10320 9200 10628 9220
rect 10704 8634 10732 10746
rect 10796 10470 10824 16934
rect 10784 10464 10836 10470
rect 10784 10406 10836 10412
rect 10888 10266 10916 17614
rect 11072 17202 11100 19200
rect 11532 17202 11560 19200
rect 11900 17202 11928 19200
rect 12360 17626 12388 19200
rect 12360 17598 12572 17626
rect 12194 17436 12502 17456
rect 12194 17434 12200 17436
rect 12256 17434 12280 17436
rect 12336 17434 12360 17436
rect 12416 17434 12440 17436
rect 12496 17434 12502 17436
rect 12256 17382 12258 17434
rect 12438 17382 12440 17434
rect 12194 17380 12200 17382
rect 12256 17380 12280 17382
rect 12336 17380 12360 17382
rect 12416 17380 12440 17382
rect 12496 17380 12502 17382
rect 12194 17360 12502 17380
rect 12544 17202 12572 17598
rect 12728 17202 12756 19200
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 11060 17196 11112 17202
rect 11060 17138 11112 17144
rect 11520 17196 11572 17202
rect 11520 17138 11572 17144
rect 11888 17196 11940 17202
rect 11888 17138 11940 17144
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12716 17196 12768 17202
rect 12716 17138 12768 17144
rect 11072 16794 11100 17138
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 11164 10538 11192 16934
rect 11152 10532 11204 10538
rect 11152 10474 11204 10480
rect 10876 10260 10928 10266
rect 10876 10202 10928 10208
rect 11256 10130 11284 17070
rect 11704 17060 11756 17066
rect 11704 17002 11756 17008
rect 11612 16992 11664 16998
rect 11612 16934 11664 16940
rect 11244 10124 11296 10130
rect 11244 10066 11296 10072
rect 11060 10056 11112 10062
rect 11060 9998 11112 10004
rect 11426 10024 11482 10033
rect 10784 8832 10836 8838
rect 10784 8774 10836 8780
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 10320 8188 10628 8208
rect 10320 8186 10326 8188
rect 10382 8186 10406 8188
rect 10462 8186 10486 8188
rect 10542 8186 10566 8188
rect 10622 8186 10628 8188
rect 10382 8134 10384 8186
rect 10564 8134 10566 8186
rect 10320 8132 10326 8134
rect 10382 8132 10406 8134
rect 10462 8132 10486 8134
rect 10542 8132 10566 8134
rect 10622 8132 10628 8134
rect 10320 8112 10628 8132
rect 10320 7100 10628 7120
rect 10320 7098 10326 7100
rect 10382 7098 10406 7100
rect 10462 7098 10486 7100
rect 10542 7098 10566 7100
rect 10622 7098 10628 7100
rect 10382 7046 10384 7098
rect 10564 7046 10566 7098
rect 10320 7044 10326 7046
rect 10382 7044 10406 7046
rect 10462 7044 10486 7046
rect 10542 7044 10566 7046
rect 10622 7044 10628 7046
rect 10320 7024 10628 7044
rect 10320 6012 10628 6032
rect 10320 6010 10326 6012
rect 10382 6010 10406 6012
rect 10462 6010 10486 6012
rect 10542 6010 10566 6012
rect 10622 6010 10628 6012
rect 10382 5958 10384 6010
rect 10564 5958 10566 6010
rect 10320 5956 10326 5958
rect 10382 5956 10406 5958
rect 10462 5956 10486 5958
rect 10542 5956 10566 5958
rect 10622 5956 10628 5958
rect 10320 5936 10628 5956
rect 10320 4924 10628 4944
rect 10320 4922 10326 4924
rect 10382 4922 10406 4924
rect 10462 4922 10486 4924
rect 10542 4922 10566 4924
rect 10622 4922 10628 4924
rect 10382 4870 10384 4922
rect 10564 4870 10566 4922
rect 10320 4868 10326 4870
rect 10382 4868 10406 4870
rect 10462 4868 10486 4870
rect 10542 4868 10566 4870
rect 10622 4868 10628 4870
rect 10320 4848 10628 4868
rect 10320 3836 10628 3856
rect 10320 3834 10326 3836
rect 10382 3834 10406 3836
rect 10462 3834 10486 3836
rect 10542 3834 10566 3836
rect 10622 3834 10628 3836
rect 10382 3782 10384 3834
rect 10564 3782 10566 3834
rect 10320 3780 10326 3782
rect 10382 3780 10406 3782
rect 10462 3780 10486 3782
rect 10542 3780 10566 3782
rect 10622 3780 10628 3782
rect 10320 3760 10628 3780
rect 10320 2748 10628 2768
rect 10320 2746 10326 2748
rect 10382 2746 10406 2748
rect 10462 2746 10486 2748
rect 10542 2746 10566 2748
rect 10622 2746 10628 2748
rect 10382 2694 10384 2746
rect 10564 2694 10566 2746
rect 10320 2692 10326 2694
rect 10382 2692 10406 2694
rect 10462 2692 10486 2694
rect 10542 2692 10566 2694
rect 10622 2692 10628 2694
rect 10320 2672 10628 2692
rect 10796 2582 10824 8774
rect 10876 2848 10928 2854
rect 10876 2790 10928 2796
rect 10784 2576 10836 2582
rect 10784 2518 10836 2524
rect 10508 2440 10560 2446
rect 10508 2382 10560 2388
rect 10888 2428 10916 2790
rect 11072 2530 11100 9998
rect 11426 9959 11482 9968
rect 11440 9926 11468 9959
rect 11244 9920 11296 9926
rect 11244 9862 11296 9868
rect 11428 9920 11480 9926
rect 11428 9862 11480 9868
rect 11520 9920 11572 9926
rect 11520 9862 11572 9868
rect 11072 2502 11192 2530
rect 11060 2440 11112 2446
rect 10888 2400 11060 2428
rect 10230 1864 10286 1873
rect 10230 1799 10286 1808
rect 10520 800 10548 2382
rect 10888 800 10916 2400
rect 11060 2382 11112 2388
rect 11164 2310 11192 2502
rect 11256 2417 11284 9862
rect 11532 6914 11560 9862
rect 11624 9518 11652 16934
rect 11716 10130 11744 17002
rect 11900 16794 11928 17138
rect 11980 16992 12032 16998
rect 11980 16934 12032 16940
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 11888 16788 11940 16794
rect 11888 16730 11940 16736
rect 11992 16658 12020 16934
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12636 16574 12664 16934
rect 12728 16794 12756 17138
rect 12808 16992 12860 16998
rect 12808 16934 12860 16940
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12544 16546 12664 16574
rect 12194 16348 12502 16368
rect 12194 16346 12200 16348
rect 12256 16346 12280 16348
rect 12336 16346 12360 16348
rect 12416 16346 12440 16348
rect 12496 16346 12502 16348
rect 12256 16294 12258 16346
rect 12438 16294 12440 16346
rect 12194 16292 12200 16294
rect 12256 16292 12280 16294
rect 12336 16292 12360 16294
rect 12416 16292 12440 16294
rect 12496 16292 12502 16294
rect 12194 16272 12502 16292
rect 12194 15260 12502 15280
rect 12194 15258 12200 15260
rect 12256 15258 12280 15260
rect 12336 15258 12360 15260
rect 12416 15258 12440 15260
rect 12496 15258 12502 15260
rect 12256 15206 12258 15258
rect 12438 15206 12440 15258
rect 12194 15204 12200 15206
rect 12256 15204 12280 15206
rect 12336 15204 12360 15206
rect 12416 15204 12440 15206
rect 12496 15204 12502 15206
rect 12194 15184 12502 15204
rect 12194 14172 12502 14192
rect 12194 14170 12200 14172
rect 12256 14170 12280 14172
rect 12336 14170 12360 14172
rect 12416 14170 12440 14172
rect 12496 14170 12502 14172
rect 12256 14118 12258 14170
rect 12438 14118 12440 14170
rect 12194 14116 12200 14118
rect 12256 14116 12280 14118
rect 12336 14116 12360 14118
rect 12416 14116 12440 14118
rect 12496 14116 12502 14118
rect 12194 14096 12502 14116
rect 12194 13084 12502 13104
rect 12194 13082 12200 13084
rect 12256 13082 12280 13084
rect 12336 13082 12360 13084
rect 12416 13082 12440 13084
rect 12496 13082 12502 13084
rect 12256 13030 12258 13082
rect 12438 13030 12440 13082
rect 12194 13028 12200 13030
rect 12256 13028 12280 13030
rect 12336 13028 12360 13030
rect 12416 13028 12440 13030
rect 12496 13028 12502 13030
rect 12194 13008 12502 13028
rect 12194 11996 12502 12016
rect 12194 11994 12200 11996
rect 12256 11994 12280 11996
rect 12336 11994 12360 11996
rect 12416 11994 12440 11996
rect 12496 11994 12502 11996
rect 12256 11942 12258 11994
rect 12438 11942 12440 11994
rect 12194 11940 12200 11942
rect 12256 11940 12280 11942
rect 12336 11940 12360 11942
rect 12416 11940 12440 11942
rect 12496 11940 12502 11942
rect 12194 11920 12502 11940
rect 12194 10908 12502 10928
rect 12194 10906 12200 10908
rect 12256 10906 12280 10908
rect 12336 10906 12360 10908
rect 12416 10906 12440 10908
rect 12496 10906 12502 10908
rect 12256 10854 12258 10906
rect 12438 10854 12440 10906
rect 12194 10852 12200 10854
rect 12256 10852 12280 10854
rect 12336 10852 12360 10854
rect 12416 10852 12440 10854
rect 12496 10852 12502 10854
rect 12194 10832 12502 10852
rect 11796 10736 11848 10742
rect 12544 10690 12572 16546
rect 12624 16448 12676 16454
rect 12624 16390 12676 16396
rect 11796 10678 11848 10684
rect 11704 10124 11756 10130
rect 11704 10066 11756 10072
rect 11808 9926 11836 10678
rect 12452 10662 12572 10690
rect 11888 10192 11940 10198
rect 11888 10134 11940 10140
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11612 9512 11664 9518
rect 11612 9454 11664 9460
rect 11440 6886 11560 6914
rect 11336 2848 11388 2854
rect 11336 2790 11388 2796
rect 11348 2446 11376 2790
rect 11336 2440 11388 2446
rect 11242 2408 11298 2417
rect 11336 2382 11388 2388
rect 11242 2343 11298 2352
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 11152 2304 11204 2310
rect 11152 2246 11204 2252
rect 10980 1766 11008 2246
rect 10968 1760 11020 1766
rect 10968 1702 11020 1708
rect 11348 800 11376 2382
rect 11440 2106 11468 6886
rect 11900 2553 11928 10134
rect 11980 10056 12032 10062
rect 11980 9998 12032 10004
rect 12452 10010 12480 10662
rect 12530 10568 12586 10577
rect 12530 10503 12586 10512
rect 12544 10198 12572 10503
rect 12532 10192 12584 10198
rect 12532 10134 12584 10140
rect 12636 10062 12664 16390
rect 12716 11008 12768 11014
rect 12716 10950 12768 10956
rect 12728 10266 12756 10950
rect 12716 10260 12768 10266
rect 12716 10202 12768 10208
rect 12624 10056 12676 10062
rect 11886 2544 11942 2553
rect 11886 2479 11942 2488
rect 11796 2440 11848 2446
rect 11796 2382 11848 2388
rect 11520 2304 11572 2310
rect 11520 2246 11572 2252
rect 11428 2100 11480 2106
rect 11428 2042 11480 2048
rect 11532 1902 11560 2246
rect 11520 1896 11572 1902
rect 11520 1838 11572 1844
rect 11808 800 11836 2382
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 1630 11928 2246
rect 11992 2106 12020 9998
rect 12452 9982 12572 10010
rect 12624 9998 12676 10004
rect 12194 9820 12502 9840
rect 12194 9818 12200 9820
rect 12256 9818 12280 9820
rect 12336 9818 12360 9820
rect 12416 9818 12440 9820
rect 12496 9818 12502 9820
rect 12256 9766 12258 9818
rect 12438 9766 12440 9818
rect 12194 9764 12200 9766
rect 12256 9764 12280 9766
rect 12336 9764 12360 9766
rect 12416 9764 12440 9766
rect 12496 9764 12502 9766
rect 12194 9744 12502 9764
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12084 2650 12112 8910
rect 12194 8732 12502 8752
rect 12194 8730 12200 8732
rect 12256 8730 12280 8732
rect 12336 8730 12360 8732
rect 12416 8730 12440 8732
rect 12496 8730 12502 8732
rect 12256 8678 12258 8730
rect 12438 8678 12440 8730
rect 12194 8676 12200 8678
rect 12256 8676 12280 8678
rect 12336 8676 12360 8678
rect 12416 8676 12440 8678
rect 12496 8676 12502 8678
rect 12194 8656 12502 8676
rect 12544 8430 12572 9982
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12716 9920 12768 9926
rect 12716 9862 12768 9868
rect 12636 9722 12664 9862
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12194 7644 12502 7664
rect 12194 7642 12200 7644
rect 12256 7642 12280 7644
rect 12336 7642 12360 7644
rect 12416 7642 12440 7644
rect 12496 7642 12502 7644
rect 12256 7590 12258 7642
rect 12438 7590 12440 7642
rect 12194 7588 12200 7590
rect 12256 7588 12280 7590
rect 12336 7588 12360 7590
rect 12416 7588 12440 7590
rect 12496 7588 12502 7590
rect 12194 7568 12502 7588
rect 12194 6556 12502 6576
rect 12194 6554 12200 6556
rect 12256 6554 12280 6556
rect 12336 6554 12360 6556
rect 12416 6554 12440 6556
rect 12496 6554 12502 6556
rect 12256 6502 12258 6554
rect 12438 6502 12440 6554
rect 12194 6500 12200 6502
rect 12256 6500 12280 6502
rect 12336 6500 12360 6502
rect 12416 6500 12440 6502
rect 12496 6500 12502 6502
rect 12194 6480 12502 6500
rect 12194 5468 12502 5488
rect 12194 5466 12200 5468
rect 12256 5466 12280 5468
rect 12336 5466 12360 5468
rect 12416 5466 12440 5468
rect 12496 5466 12502 5468
rect 12256 5414 12258 5466
rect 12438 5414 12440 5466
rect 12194 5412 12200 5414
rect 12256 5412 12280 5414
rect 12336 5412 12360 5414
rect 12416 5412 12440 5414
rect 12496 5412 12502 5414
rect 12194 5392 12502 5412
rect 12194 4380 12502 4400
rect 12194 4378 12200 4380
rect 12256 4378 12280 4380
rect 12336 4378 12360 4380
rect 12416 4378 12440 4380
rect 12496 4378 12502 4380
rect 12256 4326 12258 4378
rect 12438 4326 12440 4378
rect 12194 4324 12200 4326
rect 12256 4324 12280 4326
rect 12336 4324 12360 4326
rect 12416 4324 12440 4326
rect 12496 4324 12502 4326
rect 12194 4304 12502 4324
rect 12194 3292 12502 3312
rect 12194 3290 12200 3292
rect 12256 3290 12280 3292
rect 12336 3290 12360 3292
rect 12416 3290 12440 3292
rect 12496 3290 12502 3292
rect 12256 3238 12258 3290
rect 12438 3238 12440 3290
rect 12194 3236 12200 3238
rect 12256 3236 12280 3238
rect 12336 3236 12360 3238
rect 12416 3236 12440 3238
rect 12496 3236 12502 3238
rect 12194 3216 12502 3236
rect 12532 2848 12584 2854
rect 12532 2790 12584 2796
rect 12072 2644 12124 2650
rect 12072 2586 12124 2592
rect 12544 2446 12572 2790
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12072 2304 12124 2310
rect 12072 2246 12124 2252
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 11888 1624 11940 1630
rect 12084 1601 12112 2246
rect 12194 2204 12502 2224
rect 12194 2202 12200 2204
rect 12256 2202 12280 2204
rect 12336 2202 12360 2204
rect 12416 2202 12440 2204
rect 12496 2202 12502 2204
rect 12256 2150 12258 2202
rect 12438 2150 12440 2202
rect 12194 2148 12200 2150
rect 12256 2148 12280 2150
rect 12336 2148 12360 2150
rect 12416 2148 12440 2150
rect 12496 2148 12502 2150
rect 12194 2128 12502 2148
rect 12544 1850 12572 2382
rect 12624 2372 12676 2378
rect 12624 2314 12676 2320
rect 12176 1822 12572 1850
rect 11888 1566 11940 1572
rect 12070 1592 12126 1601
rect 12070 1527 12126 1536
rect 12176 800 12204 1822
rect 12636 800 12664 2314
rect 12728 2038 12756 9862
rect 12820 9586 12848 16934
rect 12900 10464 12952 10470
rect 12900 10406 12952 10412
rect 12912 10130 12940 10406
rect 13096 10266 13124 17546
rect 13188 17202 13216 19200
rect 13556 17202 13584 19200
rect 13636 17536 13688 17542
rect 13636 17478 13688 17484
rect 13176 17196 13228 17202
rect 13176 17138 13228 17144
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13188 16794 13216 17138
rect 13556 17082 13584 17138
rect 13464 17054 13584 17082
rect 13464 16794 13492 17054
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13176 16788 13228 16794
rect 13176 16730 13228 16736
rect 13452 16788 13504 16794
rect 13452 16730 13504 16736
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13360 10260 13412 10266
rect 13360 10202 13412 10208
rect 12900 10124 12952 10130
rect 12900 10066 12952 10072
rect 12808 9580 12860 9586
rect 12808 9522 12860 9528
rect 12808 8356 12860 8362
rect 12808 8298 12860 8304
rect 12820 7449 12848 8298
rect 12806 7440 12862 7449
rect 12806 7375 12862 7384
rect 13268 2576 13320 2582
rect 13268 2518 13320 2524
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 12716 2032 12768 2038
rect 12716 1974 12768 1980
rect 13096 800 13124 2382
rect 13280 1737 13308 2518
rect 13372 2417 13400 10202
rect 13556 9654 13584 16934
rect 13648 10266 13676 17478
rect 14016 17338 14044 19200
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 14476 17202 14504 19200
rect 14844 17202 14872 19200
rect 14464 17196 14516 17202
rect 14464 17138 14516 17144
rect 14832 17196 14884 17202
rect 14832 17138 14884 17144
rect 14556 17128 14608 17134
rect 14556 17070 14608 17076
rect 13728 16992 13780 16998
rect 13728 16934 13780 16940
rect 13740 11014 13768 16934
rect 14068 16892 14376 16912
rect 14068 16890 14074 16892
rect 14130 16890 14154 16892
rect 14210 16890 14234 16892
rect 14290 16890 14314 16892
rect 14370 16890 14376 16892
rect 14130 16838 14132 16890
rect 14312 16838 14314 16890
rect 14068 16836 14074 16838
rect 14130 16836 14154 16838
rect 14210 16836 14234 16838
rect 14290 16836 14314 16838
rect 14370 16836 14376 16838
rect 14068 16816 14376 16836
rect 14068 15804 14376 15824
rect 14068 15802 14074 15804
rect 14130 15802 14154 15804
rect 14210 15802 14234 15804
rect 14290 15802 14314 15804
rect 14370 15802 14376 15804
rect 14130 15750 14132 15802
rect 14312 15750 14314 15802
rect 14068 15748 14074 15750
rect 14130 15748 14154 15750
rect 14210 15748 14234 15750
rect 14290 15748 14314 15750
rect 14370 15748 14376 15750
rect 14068 15728 14376 15748
rect 14068 14716 14376 14736
rect 14068 14714 14074 14716
rect 14130 14714 14154 14716
rect 14210 14714 14234 14716
rect 14290 14714 14314 14716
rect 14370 14714 14376 14716
rect 14130 14662 14132 14714
rect 14312 14662 14314 14714
rect 14068 14660 14074 14662
rect 14130 14660 14154 14662
rect 14210 14660 14234 14662
rect 14290 14660 14314 14662
rect 14370 14660 14376 14662
rect 14068 14640 14376 14660
rect 14068 13628 14376 13648
rect 14068 13626 14074 13628
rect 14130 13626 14154 13628
rect 14210 13626 14234 13628
rect 14290 13626 14314 13628
rect 14370 13626 14376 13628
rect 14130 13574 14132 13626
rect 14312 13574 14314 13626
rect 14068 13572 14074 13574
rect 14130 13572 14154 13574
rect 14210 13572 14234 13574
rect 14290 13572 14314 13574
rect 14370 13572 14376 13574
rect 14068 13552 14376 13572
rect 14568 12986 14596 17070
rect 14844 16794 14872 17138
rect 14832 16788 14884 16794
rect 14832 16730 14884 16736
rect 15108 16720 15160 16726
rect 15304 16674 15332 19200
rect 15566 17504 15622 17513
rect 15566 17439 15622 17448
rect 15580 17338 15608 17439
rect 15568 17332 15620 17338
rect 15568 17274 15620 17280
rect 15160 16668 15332 16674
rect 15108 16662 15332 16668
rect 15120 16646 15332 16662
rect 15304 16574 15332 16646
rect 15384 16584 15436 16590
rect 15304 16546 15384 16574
rect 15384 16526 15436 16532
rect 15672 16522 15700 19200
rect 16132 16590 16160 19200
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15476 16448 15528 16454
rect 15476 16390 15528 16396
rect 15200 15904 15252 15910
rect 15200 15846 15252 15852
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 14556 12980 14608 12986
rect 14556 12922 14608 12928
rect 14068 12540 14376 12560
rect 14068 12538 14074 12540
rect 14130 12538 14154 12540
rect 14210 12538 14234 12540
rect 14290 12538 14314 12540
rect 14370 12538 14376 12540
rect 14130 12486 14132 12538
rect 14312 12486 14314 12538
rect 14068 12484 14074 12486
rect 14130 12484 14154 12486
rect 14210 12484 14234 12486
rect 14290 12484 14314 12486
rect 14370 12484 14376 12486
rect 14068 12464 14376 12484
rect 14068 11452 14376 11472
rect 14068 11450 14074 11452
rect 14130 11450 14154 11452
rect 14210 11450 14234 11452
rect 14290 11450 14314 11452
rect 14370 11450 14376 11452
rect 14130 11398 14132 11450
rect 14312 11398 14314 11450
rect 14068 11396 14074 11398
rect 14130 11396 14154 11398
rect 14210 11396 14234 11398
rect 14290 11396 14314 11398
rect 14370 11396 14376 11398
rect 14068 11376 14376 11396
rect 13728 11008 13780 11014
rect 13728 10950 13780 10956
rect 14068 10364 14376 10384
rect 14068 10362 14074 10364
rect 14130 10362 14154 10364
rect 14210 10362 14234 10364
rect 14290 10362 14314 10364
rect 14370 10362 14376 10364
rect 14130 10310 14132 10362
rect 14312 10310 14314 10362
rect 14068 10308 14074 10310
rect 14130 10308 14154 10310
rect 14210 10308 14234 10310
rect 14290 10308 14314 10310
rect 14370 10308 14376 10310
rect 14068 10288 14376 10308
rect 13636 10260 13688 10266
rect 13636 10202 13688 10208
rect 15212 10130 15240 15846
rect 15304 10198 15332 15846
rect 15396 10470 15424 16390
rect 15488 15706 15516 16390
rect 16500 16114 16528 19200
rect 16960 16182 16988 19200
rect 16948 16176 17000 16182
rect 16948 16118 17000 16124
rect 16488 16108 16540 16114
rect 16488 16050 16540 16056
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15568 12640 15620 12646
rect 15568 12582 15620 12588
rect 15580 12481 15608 12582
rect 15566 12472 15622 12481
rect 15566 12407 15622 12416
rect 15384 10464 15436 10470
rect 15384 10406 15436 10412
rect 15292 10192 15344 10198
rect 15292 10134 15344 10140
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 13820 10056 13872 10062
rect 13820 9998 13872 10004
rect 13636 9716 13688 9722
rect 13636 9658 13688 9664
rect 13544 9648 13596 9654
rect 13544 9590 13596 9596
rect 13452 2848 13504 2854
rect 13452 2790 13504 2796
rect 13464 2446 13492 2790
rect 13648 2650 13676 9658
rect 13832 3738 13860 9998
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14740 9920 14792 9926
rect 14740 9862 14792 9868
rect 14068 9276 14376 9296
rect 14068 9274 14074 9276
rect 14130 9274 14154 9276
rect 14210 9274 14234 9276
rect 14290 9274 14314 9276
rect 14370 9274 14376 9276
rect 14130 9222 14132 9274
rect 14312 9222 14314 9274
rect 14068 9220 14074 9222
rect 14130 9220 14154 9222
rect 14210 9220 14234 9222
rect 14290 9220 14314 9222
rect 14370 9220 14376 9222
rect 14068 9200 14376 9220
rect 14068 8188 14376 8208
rect 14068 8186 14074 8188
rect 14130 8186 14154 8188
rect 14210 8186 14234 8188
rect 14290 8186 14314 8188
rect 14370 8186 14376 8188
rect 14130 8134 14132 8186
rect 14312 8134 14314 8186
rect 14068 8132 14074 8134
rect 14130 8132 14154 8134
rect 14210 8132 14234 8134
rect 14290 8132 14314 8134
rect 14370 8132 14376 8134
rect 14068 8112 14376 8132
rect 14068 7100 14376 7120
rect 14068 7098 14074 7100
rect 14130 7098 14154 7100
rect 14210 7098 14234 7100
rect 14290 7098 14314 7100
rect 14370 7098 14376 7100
rect 14130 7046 14132 7098
rect 14312 7046 14314 7098
rect 14068 7044 14074 7046
rect 14130 7044 14154 7046
rect 14210 7044 14234 7046
rect 14290 7044 14314 7046
rect 14370 7044 14376 7046
rect 14068 7024 14376 7044
rect 14068 6012 14376 6032
rect 14068 6010 14074 6012
rect 14130 6010 14154 6012
rect 14210 6010 14234 6012
rect 14290 6010 14314 6012
rect 14370 6010 14376 6012
rect 14130 5958 14132 6010
rect 14312 5958 14314 6010
rect 14068 5956 14074 5958
rect 14130 5956 14154 5958
rect 14210 5956 14234 5958
rect 14290 5956 14314 5958
rect 14370 5956 14376 5958
rect 14068 5936 14376 5956
rect 14068 4924 14376 4944
rect 14068 4922 14074 4924
rect 14130 4922 14154 4924
rect 14210 4922 14234 4924
rect 14290 4922 14314 4924
rect 14370 4922 14376 4924
rect 14130 4870 14132 4922
rect 14312 4870 14314 4922
rect 14068 4868 14074 4870
rect 14130 4868 14154 4870
rect 14210 4868 14234 4870
rect 14290 4868 14314 4870
rect 14370 4868 14376 4870
rect 14068 4848 14376 4868
rect 14068 3836 14376 3856
rect 14068 3834 14074 3836
rect 14130 3834 14154 3836
rect 14210 3834 14234 3836
rect 14290 3834 14314 3836
rect 14370 3834 14376 3836
rect 14130 3782 14132 3834
rect 14312 3782 14314 3834
rect 14068 3780 14074 3782
rect 14130 3780 14154 3782
rect 14210 3780 14234 3782
rect 14290 3780 14314 3782
rect 14370 3780 14376 3782
rect 14068 3760 14376 3780
rect 13820 3732 13872 3738
rect 13820 3674 13872 3680
rect 14752 3126 14780 9862
rect 14936 3194 14964 9930
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 15660 3392 15712 3398
rect 15660 3334 15712 3340
rect 14924 3188 14976 3194
rect 14924 3130 14976 3136
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 15304 2990 15332 3334
rect 15672 3058 15700 3334
rect 15384 3052 15436 3058
rect 15384 2994 15436 3000
rect 15660 3052 15712 3058
rect 15660 2994 15712 3000
rect 15292 2984 15344 2990
rect 15292 2926 15344 2932
rect 15200 2916 15252 2922
rect 15200 2858 15252 2864
rect 13912 2848 13964 2854
rect 13912 2790 13964 2796
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13924 2446 13952 2790
rect 14068 2748 14376 2768
rect 14068 2746 14074 2748
rect 14130 2746 14154 2748
rect 14210 2746 14234 2748
rect 14290 2746 14314 2748
rect 14370 2746 14376 2748
rect 14130 2694 14132 2746
rect 14312 2694 14314 2746
rect 14068 2692 14074 2694
rect 14130 2692 14154 2694
rect 14210 2692 14234 2694
rect 14290 2692 14314 2694
rect 14370 2692 14376 2694
rect 14068 2672 14376 2692
rect 14752 2446 14780 2790
rect 15212 2446 15240 2858
rect 13452 2440 13504 2446
rect 13358 2408 13414 2417
rect 13452 2382 13504 2388
rect 13912 2440 13964 2446
rect 13912 2382 13964 2388
rect 14372 2440 14424 2446
rect 14372 2382 14424 2388
rect 14740 2440 14792 2446
rect 14740 2382 14792 2388
rect 15200 2440 15252 2446
rect 15200 2382 15252 2388
rect 13358 2343 13414 2352
rect 13266 1728 13322 1737
rect 13266 1663 13322 1672
rect 13464 800 13492 2382
rect 13924 800 13952 2382
rect 14096 2304 14148 2310
rect 14096 2246 14148 2252
rect 14108 1834 14136 2246
rect 14096 1828 14148 1834
rect 14096 1770 14148 1776
rect 14384 800 14412 2382
rect 14752 800 14780 2382
rect 15212 800 15240 2382
rect 15396 2310 15424 2994
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15384 2304 15436 2310
rect 15384 2246 15436 2252
rect 15304 2106 15332 2246
rect 15292 2100 15344 2106
rect 15292 2042 15344 2048
rect 15672 800 15700 2994
rect 16488 2984 16540 2990
rect 16488 2926 16540 2932
rect 16028 2304 16080 2310
rect 16028 2246 16080 2252
rect 16040 800 16068 2246
rect 16500 800 16528 2926
rect 16960 800 16988 3470
rect 202 0 258 800
rect 570 0 626 800
rect 1030 0 1086 800
rect 1490 0 1546 800
rect 1858 0 1914 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3146 0 3202 800
rect 3606 0 3662 800
rect 4066 0 4122 800
rect 4434 0 4490 800
rect 4894 0 4950 800
rect 5354 0 5410 800
rect 5722 0 5778 800
rect 6182 0 6238 800
rect 6642 0 6698 800
rect 7010 0 7066 800
rect 7470 0 7526 800
rect 7930 0 7986 800
rect 8298 0 8354 800
rect 8758 0 8814 800
rect 9218 0 9274 800
rect 9586 0 9642 800
rect 10046 0 10102 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11334 0 11390 800
rect 11794 0 11850 800
rect 12162 0 12218 800
rect 12622 0 12678 800
rect 13082 0 13138 800
rect 13450 0 13506 800
rect 13910 0 13966 800
rect 14370 0 14426 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 15658 0 15714 800
rect 16026 0 16082 800
rect 16486 0 16542 800
rect 16946 0 17002 800
<< via2 >>
rect 1950 18264 2006 18320
rect 4704 17434 4760 17436
rect 4784 17434 4840 17436
rect 4864 17434 4920 17436
rect 4944 17434 5000 17436
rect 4704 17382 4750 17434
rect 4750 17382 4760 17434
rect 4784 17382 4814 17434
rect 4814 17382 4826 17434
rect 4826 17382 4840 17434
rect 4864 17382 4878 17434
rect 4878 17382 4890 17434
rect 4890 17382 4920 17434
rect 4944 17382 4954 17434
rect 4954 17382 5000 17434
rect 4704 17380 4760 17382
rect 4784 17380 4840 17382
rect 4864 17380 4920 17382
rect 4944 17380 5000 17382
rect 1398 11600 1454 11656
rect 1490 8356 1546 8392
rect 1490 8336 1492 8356
rect 1492 8336 1544 8356
rect 1544 8336 1546 8356
rect 1490 4972 1492 4992
rect 1492 4972 1544 4992
rect 1544 4972 1546 4992
rect 1490 4936 1546 4972
rect 2830 16890 2886 16892
rect 2910 16890 2966 16892
rect 2990 16890 3046 16892
rect 3070 16890 3126 16892
rect 2830 16838 2876 16890
rect 2876 16838 2886 16890
rect 2910 16838 2940 16890
rect 2940 16838 2952 16890
rect 2952 16838 2966 16890
rect 2990 16838 3004 16890
rect 3004 16838 3016 16890
rect 3016 16838 3046 16890
rect 3070 16838 3080 16890
rect 3080 16838 3126 16890
rect 2830 16836 2886 16838
rect 2910 16836 2966 16838
rect 2990 16836 3046 16838
rect 3070 16836 3126 16838
rect 2830 15802 2886 15804
rect 2910 15802 2966 15804
rect 2990 15802 3046 15804
rect 3070 15802 3126 15804
rect 2830 15750 2876 15802
rect 2876 15750 2886 15802
rect 2910 15750 2940 15802
rect 2940 15750 2952 15802
rect 2952 15750 2966 15802
rect 2990 15750 3004 15802
rect 3004 15750 3016 15802
rect 3016 15750 3046 15802
rect 3070 15750 3080 15802
rect 3080 15750 3126 15802
rect 2830 15748 2886 15750
rect 2910 15748 2966 15750
rect 2990 15748 3046 15750
rect 3070 15748 3126 15750
rect 3146 15000 3202 15056
rect 2830 14714 2886 14716
rect 2910 14714 2966 14716
rect 2990 14714 3046 14716
rect 3070 14714 3126 14716
rect 2830 14662 2876 14714
rect 2876 14662 2886 14714
rect 2910 14662 2940 14714
rect 2940 14662 2952 14714
rect 2952 14662 2966 14714
rect 2990 14662 3004 14714
rect 3004 14662 3016 14714
rect 3016 14662 3046 14714
rect 3070 14662 3080 14714
rect 3080 14662 3126 14714
rect 2830 14660 2886 14662
rect 2910 14660 2966 14662
rect 2990 14660 3046 14662
rect 3070 14660 3126 14662
rect 2830 13626 2886 13628
rect 2910 13626 2966 13628
rect 2990 13626 3046 13628
rect 3070 13626 3126 13628
rect 2830 13574 2876 13626
rect 2876 13574 2886 13626
rect 2910 13574 2940 13626
rect 2940 13574 2952 13626
rect 2952 13574 2966 13626
rect 2990 13574 3004 13626
rect 3004 13574 3016 13626
rect 3016 13574 3046 13626
rect 3070 13574 3080 13626
rect 3080 13574 3126 13626
rect 2830 13572 2886 13574
rect 2910 13572 2966 13574
rect 2990 13572 3046 13574
rect 3070 13572 3126 13574
rect 2830 12538 2886 12540
rect 2910 12538 2966 12540
rect 2990 12538 3046 12540
rect 3070 12538 3126 12540
rect 2830 12486 2876 12538
rect 2876 12486 2886 12538
rect 2910 12486 2940 12538
rect 2940 12486 2952 12538
rect 2952 12486 2966 12538
rect 2990 12486 3004 12538
rect 3004 12486 3016 12538
rect 3016 12486 3046 12538
rect 3070 12486 3080 12538
rect 3080 12486 3126 12538
rect 2830 12484 2886 12486
rect 2910 12484 2966 12486
rect 2990 12484 3046 12486
rect 3070 12484 3126 12486
rect 2830 11450 2886 11452
rect 2910 11450 2966 11452
rect 2990 11450 3046 11452
rect 3070 11450 3126 11452
rect 2830 11398 2876 11450
rect 2876 11398 2886 11450
rect 2910 11398 2940 11450
rect 2940 11398 2952 11450
rect 2952 11398 2966 11450
rect 2990 11398 3004 11450
rect 3004 11398 3016 11450
rect 3016 11398 3046 11450
rect 3070 11398 3080 11450
rect 3080 11398 3126 11450
rect 2830 11396 2886 11398
rect 2910 11396 2966 11398
rect 2990 11396 3046 11398
rect 3070 11396 3126 11398
rect 2830 10362 2886 10364
rect 2910 10362 2966 10364
rect 2990 10362 3046 10364
rect 3070 10362 3126 10364
rect 2830 10310 2876 10362
rect 2876 10310 2886 10362
rect 2910 10310 2940 10362
rect 2940 10310 2952 10362
rect 2952 10310 2966 10362
rect 2990 10310 3004 10362
rect 3004 10310 3016 10362
rect 3016 10310 3046 10362
rect 3070 10310 3080 10362
rect 3080 10310 3126 10362
rect 2830 10308 2886 10310
rect 2910 10308 2966 10310
rect 2990 10308 3046 10310
rect 3070 10308 3126 10310
rect 2830 9274 2886 9276
rect 2910 9274 2966 9276
rect 2990 9274 3046 9276
rect 3070 9274 3126 9276
rect 2830 9222 2876 9274
rect 2876 9222 2886 9274
rect 2910 9222 2940 9274
rect 2940 9222 2952 9274
rect 2952 9222 2966 9274
rect 2990 9222 3004 9274
rect 3004 9222 3016 9274
rect 3016 9222 3046 9274
rect 3070 9222 3080 9274
rect 3080 9222 3126 9274
rect 2830 9220 2886 9222
rect 2910 9220 2966 9222
rect 2990 9220 3046 9222
rect 3070 9220 3126 9222
rect 2830 8186 2886 8188
rect 2910 8186 2966 8188
rect 2990 8186 3046 8188
rect 3070 8186 3126 8188
rect 2830 8134 2876 8186
rect 2876 8134 2886 8186
rect 2910 8134 2940 8186
rect 2940 8134 2952 8186
rect 2952 8134 2966 8186
rect 2990 8134 3004 8186
rect 3004 8134 3016 8186
rect 3016 8134 3046 8186
rect 3070 8134 3080 8186
rect 3080 8134 3126 8186
rect 2830 8132 2886 8134
rect 2910 8132 2966 8134
rect 2990 8132 3046 8134
rect 3070 8132 3126 8134
rect 2830 7098 2886 7100
rect 2910 7098 2966 7100
rect 2990 7098 3046 7100
rect 3070 7098 3126 7100
rect 2830 7046 2876 7098
rect 2876 7046 2886 7098
rect 2910 7046 2940 7098
rect 2940 7046 2952 7098
rect 2952 7046 2966 7098
rect 2990 7046 3004 7098
rect 3004 7046 3016 7098
rect 3016 7046 3046 7098
rect 3070 7046 3080 7098
rect 3080 7046 3126 7098
rect 2830 7044 2886 7046
rect 2910 7044 2966 7046
rect 2990 7044 3046 7046
rect 3070 7044 3126 7046
rect 2830 6010 2886 6012
rect 2910 6010 2966 6012
rect 2990 6010 3046 6012
rect 3070 6010 3126 6012
rect 2830 5958 2876 6010
rect 2876 5958 2886 6010
rect 2910 5958 2940 6010
rect 2940 5958 2952 6010
rect 2952 5958 2966 6010
rect 2990 5958 3004 6010
rect 3004 5958 3016 6010
rect 3016 5958 3046 6010
rect 3070 5958 3080 6010
rect 3080 5958 3126 6010
rect 2830 5956 2886 5958
rect 2910 5956 2966 5958
rect 2990 5956 3046 5958
rect 3070 5956 3126 5958
rect 2830 4922 2886 4924
rect 2910 4922 2966 4924
rect 2990 4922 3046 4924
rect 3070 4922 3126 4924
rect 2830 4870 2876 4922
rect 2876 4870 2886 4922
rect 2910 4870 2940 4922
rect 2940 4870 2952 4922
rect 2952 4870 2966 4922
rect 2990 4870 3004 4922
rect 3004 4870 3016 4922
rect 3016 4870 3046 4922
rect 3070 4870 3080 4922
rect 3080 4870 3126 4922
rect 2830 4868 2886 4870
rect 2910 4868 2966 4870
rect 2990 4868 3046 4870
rect 3070 4868 3126 4870
rect 2830 3834 2886 3836
rect 2910 3834 2966 3836
rect 2990 3834 3046 3836
rect 3070 3834 3126 3836
rect 2830 3782 2876 3834
rect 2876 3782 2886 3834
rect 2910 3782 2940 3834
rect 2940 3782 2952 3834
rect 2952 3782 2966 3834
rect 2990 3782 3004 3834
rect 3004 3782 3016 3834
rect 3016 3782 3046 3834
rect 3070 3782 3080 3834
rect 3080 3782 3126 3834
rect 2830 3780 2886 3782
rect 2910 3780 2966 3782
rect 2990 3780 3046 3782
rect 3070 3780 3126 3782
rect 8452 17434 8508 17436
rect 8532 17434 8588 17436
rect 8612 17434 8668 17436
rect 8692 17434 8748 17436
rect 8452 17382 8498 17434
rect 8498 17382 8508 17434
rect 8532 17382 8562 17434
rect 8562 17382 8574 17434
rect 8574 17382 8588 17434
rect 8612 17382 8626 17434
rect 8626 17382 8638 17434
rect 8638 17382 8668 17434
rect 8692 17382 8702 17434
rect 8702 17382 8748 17434
rect 8452 17380 8508 17382
rect 8532 17380 8588 17382
rect 8612 17380 8668 17382
rect 8692 17380 8748 17382
rect 4704 16346 4760 16348
rect 4784 16346 4840 16348
rect 4864 16346 4920 16348
rect 4944 16346 5000 16348
rect 4704 16294 4750 16346
rect 4750 16294 4760 16346
rect 4784 16294 4814 16346
rect 4814 16294 4826 16346
rect 4826 16294 4840 16346
rect 4864 16294 4878 16346
rect 4878 16294 4890 16346
rect 4890 16294 4920 16346
rect 4944 16294 4954 16346
rect 4954 16294 5000 16346
rect 4704 16292 4760 16294
rect 4784 16292 4840 16294
rect 4864 16292 4920 16294
rect 4944 16292 5000 16294
rect 4704 15258 4760 15260
rect 4784 15258 4840 15260
rect 4864 15258 4920 15260
rect 4944 15258 5000 15260
rect 4704 15206 4750 15258
rect 4750 15206 4760 15258
rect 4784 15206 4814 15258
rect 4814 15206 4826 15258
rect 4826 15206 4840 15258
rect 4864 15206 4878 15258
rect 4878 15206 4890 15258
rect 4890 15206 4920 15258
rect 4944 15206 4954 15258
rect 4954 15206 5000 15258
rect 4704 15204 4760 15206
rect 4784 15204 4840 15206
rect 4864 15204 4920 15206
rect 4944 15204 5000 15206
rect 4704 14170 4760 14172
rect 4784 14170 4840 14172
rect 4864 14170 4920 14172
rect 4944 14170 5000 14172
rect 4704 14118 4750 14170
rect 4750 14118 4760 14170
rect 4784 14118 4814 14170
rect 4814 14118 4826 14170
rect 4826 14118 4840 14170
rect 4864 14118 4878 14170
rect 4878 14118 4890 14170
rect 4890 14118 4920 14170
rect 4944 14118 4954 14170
rect 4954 14118 5000 14170
rect 4704 14116 4760 14118
rect 4784 14116 4840 14118
rect 4864 14116 4920 14118
rect 4944 14116 5000 14118
rect 4704 13082 4760 13084
rect 4784 13082 4840 13084
rect 4864 13082 4920 13084
rect 4944 13082 5000 13084
rect 4704 13030 4750 13082
rect 4750 13030 4760 13082
rect 4784 13030 4814 13082
rect 4814 13030 4826 13082
rect 4826 13030 4840 13082
rect 4864 13030 4878 13082
rect 4878 13030 4890 13082
rect 4890 13030 4920 13082
rect 4944 13030 4954 13082
rect 4954 13030 5000 13082
rect 4704 13028 4760 13030
rect 4784 13028 4840 13030
rect 4864 13028 4920 13030
rect 4944 13028 5000 13030
rect 4704 11994 4760 11996
rect 4784 11994 4840 11996
rect 4864 11994 4920 11996
rect 4944 11994 5000 11996
rect 4704 11942 4750 11994
rect 4750 11942 4760 11994
rect 4784 11942 4814 11994
rect 4814 11942 4826 11994
rect 4826 11942 4840 11994
rect 4864 11942 4878 11994
rect 4878 11942 4890 11994
rect 4890 11942 4920 11994
rect 4944 11942 4954 11994
rect 4954 11942 5000 11994
rect 4704 11940 4760 11942
rect 4784 11940 4840 11942
rect 4864 11940 4920 11942
rect 4944 11940 5000 11942
rect 2830 2746 2886 2748
rect 2910 2746 2966 2748
rect 2990 2746 3046 2748
rect 3070 2746 3126 2748
rect 2830 2694 2876 2746
rect 2876 2694 2886 2746
rect 2910 2694 2940 2746
rect 2940 2694 2952 2746
rect 2952 2694 2966 2746
rect 2990 2694 3004 2746
rect 3004 2694 3016 2746
rect 3016 2694 3046 2746
rect 3070 2694 3080 2746
rect 3080 2694 3126 2746
rect 2830 2692 2886 2694
rect 2910 2692 2966 2694
rect 2990 2692 3046 2694
rect 3070 2692 3126 2694
rect 2686 2488 2742 2544
rect 4704 10906 4760 10908
rect 4784 10906 4840 10908
rect 4864 10906 4920 10908
rect 4944 10906 5000 10908
rect 4704 10854 4750 10906
rect 4750 10854 4760 10906
rect 4784 10854 4814 10906
rect 4814 10854 4826 10906
rect 4826 10854 4840 10906
rect 4864 10854 4878 10906
rect 4878 10854 4890 10906
rect 4890 10854 4920 10906
rect 4944 10854 4954 10906
rect 4954 10854 5000 10906
rect 4704 10852 4760 10854
rect 4784 10852 4840 10854
rect 4864 10852 4920 10854
rect 4944 10852 5000 10854
rect 4704 9818 4760 9820
rect 4784 9818 4840 9820
rect 4864 9818 4920 9820
rect 4944 9818 5000 9820
rect 4704 9766 4750 9818
rect 4750 9766 4760 9818
rect 4784 9766 4814 9818
rect 4814 9766 4826 9818
rect 4826 9766 4840 9818
rect 4864 9766 4878 9818
rect 4878 9766 4890 9818
rect 4890 9766 4920 9818
rect 4944 9766 4954 9818
rect 4954 9766 5000 9818
rect 4704 9764 4760 9766
rect 4784 9764 4840 9766
rect 4864 9764 4920 9766
rect 4944 9764 5000 9766
rect 4704 8730 4760 8732
rect 4784 8730 4840 8732
rect 4864 8730 4920 8732
rect 4944 8730 5000 8732
rect 4704 8678 4750 8730
rect 4750 8678 4760 8730
rect 4784 8678 4814 8730
rect 4814 8678 4826 8730
rect 4826 8678 4840 8730
rect 4864 8678 4878 8730
rect 4878 8678 4890 8730
rect 4890 8678 4920 8730
rect 4944 8678 4954 8730
rect 4954 8678 5000 8730
rect 4704 8676 4760 8678
rect 4784 8676 4840 8678
rect 4864 8676 4920 8678
rect 4944 8676 5000 8678
rect 4704 7642 4760 7644
rect 4784 7642 4840 7644
rect 4864 7642 4920 7644
rect 4944 7642 5000 7644
rect 4704 7590 4750 7642
rect 4750 7590 4760 7642
rect 4784 7590 4814 7642
rect 4814 7590 4826 7642
rect 4826 7590 4840 7642
rect 4864 7590 4878 7642
rect 4878 7590 4890 7642
rect 4890 7590 4920 7642
rect 4944 7590 4954 7642
rect 4954 7590 5000 7642
rect 4704 7588 4760 7590
rect 4784 7588 4840 7590
rect 4864 7588 4920 7590
rect 4944 7588 5000 7590
rect 4704 6554 4760 6556
rect 4784 6554 4840 6556
rect 4864 6554 4920 6556
rect 4944 6554 5000 6556
rect 4704 6502 4750 6554
rect 4750 6502 4760 6554
rect 4784 6502 4814 6554
rect 4814 6502 4826 6554
rect 4826 6502 4840 6554
rect 4864 6502 4878 6554
rect 4878 6502 4890 6554
rect 4890 6502 4920 6554
rect 4944 6502 4954 6554
rect 4954 6502 5000 6554
rect 4704 6500 4760 6502
rect 4784 6500 4840 6502
rect 4864 6500 4920 6502
rect 4944 6500 5000 6502
rect 4704 5466 4760 5468
rect 4784 5466 4840 5468
rect 4864 5466 4920 5468
rect 4944 5466 5000 5468
rect 4704 5414 4750 5466
rect 4750 5414 4760 5466
rect 4784 5414 4814 5466
rect 4814 5414 4826 5466
rect 4826 5414 4840 5466
rect 4864 5414 4878 5466
rect 4878 5414 4890 5466
rect 4890 5414 4920 5466
rect 4944 5414 4954 5466
rect 4954 5414 5000 5466
rect 4704 5412 4760 5414
rect 4784 5412 4840 5414
rect 4864 5412 4920 5414
rect 4944 5412 5000 5414
rect 4704 4378 4760 4380
rect 4784 4378 4840 4380
rect 4864 4378 4920 4380
rect 4944 4378 5000 4380
rect 4704 4326 4750 4378
rect 4750 4326 4760 4378
rect 4784 4326 4814 4378
rect 4814 4326 4826 4378
rect 4826 4326 4840 4378
rect 4864 4326 4878 4378
rect 4878 4326 4890 4378
rect 4890 4326 4920 4378
rect 4944 4326 4954 4378
rect 4954 4326 5000 4378
rect 4704 4324 4760 4326
rect 4784 4324 4840 4326
rect 4864 4324 4920 4326
rect 4944 4324 5000 4326
rect 2134 1672 2190 1728
rect 4704 3290 4760 3292
rect 4784 3290 4840 3292
rect 4864 3290 4920 3292
rect 4944 3290 5000 3292
rect 4704 3238 4750 3290
rect 4750 3238 4760 3290
rect 4784 3238 4814 3290
rect 4814 3238 4826 3290
rect 4826 3238 4840 3290
rect 4864 3238 4878 3290
rect 4878 3238 4890 3290
rect 4890 3238 4920 3290
rect 4944 3238 4954 3290
rect 4954 3238 5000 3290
rect 4704 3236 4760 3238
rect 4784 3236 4840 3238
rect 4864 3236 4920 3238
rect 4944 3236 5000 3238
rect 5722 9696 5778 9752
rect 4704 2202 4760 2204
rect 4784 2202 4840 2204
rect 4864 2202 4920 2204
rect 4944 2202 5000 2204
rect 4704 2150 4750 2202
rect 4750 2150 4760 2202
rect 4784 2150 4814 2202
rect 4814 2150 4826 2202
rect 4826 2150 4840 2202
rect 4864 2150 4878 2202
rect 4878 2150 4890 2202
rect 4890 2150 4920 2202
rect 4944 2150 4954 2202
rect 4954 2150 5000 2202
rect 4704 2148 4760 2150
rect 4784 2148 4840 2150
rect 4864 2148 4920 2150
rect 4944 2148 5000 2150
rect 4618 1808 4674 1864
rect 6578 16890 6634 16892
rect 6658 16890 6714 16892
rect 6738 16890 6794 16892
rect 6818 16890 6874 16892
rect 6578 16838 6624 16890
rect 6624 16838 6634 16890
rect 6658 16838 6688 16890
rect 6688 16838 6700 16890
rect 6700 16838 6714 16890
rect 6738 16838 6752 16890
rect 6752 16838 6764 16890
rect 6764 16838 6794 16890
rect 6818 16838 6828 16890
rect 6828 16838 6874 16890
rect 6578 16836 6634 16838
rect 6658 16836 6714 16838
rect 6738 16836 6794 16838
rect 6818 16836 6874 16838
rect 6578 15802 6634 15804
rect 6658 15802 6714 15804
rect 6738 15802 6794 15804
rect 6818 15802 6874 15804
rect 6578 15750 6624 15802
rect 6624 15750 6634 15802
rect 6658 15750 6688 15802
rect 6688 15750 6700 15802
rect 6700 15750 6714 15802
rect 6738 15750 6752 15802
rect 6752 15750 6764 15802
rect 6764 15750 6794 15802
rect 6818 15750 6828 15802
rect 6828 15750 6874 15802
rect 6578 15748 6634 15750
rect 6658 15748 6714 15750
rect 6738 15748 6794 15750
rect 6818 15748 6874 15750
rect 6578 14714 6634 14716
rect 6658 14714 6714 14716
rect 6738 14714 6794 14716
rect 6818 14714 6874 14716
rect 6578 14662 6624 14714
rect 6624 14662 6634 14714
rect 6658 14662 6688 14714
rect 6688 14662 6700 14714
rect 6700 14662 6714 14714
rect 6738 14662 6752 14714
rect 6752 14662 6764 14714
rect 6764 14662 6794 14714
rect 6818 14662 6828 14714
rect 6828 14662 6874 14714
rect 6578 14660 6634 14662
rect 6658 14660 6714 14662
rect 6738 14660 6794 14662
rect 6818 14660 6874 14662
rect 6578 13626 6634 13628
rect 6658 13626 6714 13628
rect 6738 13626 6794 13628
rect 6818 13626 6874 13628
rect 6578 13574 6624 13626
rect 6624 13574 6634 13626
rect 6658 13574 6688 13626
rect 6688 13574 6700 13626
rect 6700 13574 6714 13626
rect 6738 13574 6752 13626
rect 6752 13574 6764 13626
rect 6764 13574 6794 13626
rect 6818 13574 6828 13626
rect 6828 13574 6874 13626
rect 6578 13572 6634 13574
rect 6658 13572 6714 13574
rect 6738 13572 6794 13574
rect 6818 13572 6874 13574
rect 6578 12538 6634 12540
rect 6658 12538 6714 12540
rect 6738 12538 6794 12540
rect 6818 12538 6874 12540
rect 6578 12486 6624 12538
rect 6624 12486 6634 12538
rect 6658 12486 6688 12538
rect 6688 12486 6700 12538
rect 6700 12486 6714 12538
rect 6738 12486 6752 12538
rect 6752 12486 6764 12538
rect 6764 12486 6794 12538
rect 6818 12486 6828 12538
rect 6828 12486 6874 12538
rect 6578 12484 6634 12486
rect 6658 12484 6714 12486
rect 6738 12484 6794 12486
rect 6818 12484 6874 12486
rect 6578 11450 6634 11452
rect 6658 11450 6714 11452
rect 6738 11450 6794 11452
rect 6818 11450 6874 11452
rect 6578 11398 6624 11450
rect 6624 11398 6634 11450
rect 6658 11398 6688 11450
rect 6688 11398 6700 11450
rect 6700 11398 6714 11450
rect 6738 11398 6752 11450
rect 6752 11398 6764 11450
rect 6764 11398 6794 11450
rect 6818 11398 6828 11450
rect 6828 11398 6874 11450
rect 6578 11396 6634 11398
rect 6658 11396 6714 11398
rect 6738 11396 6794 11398
rect 6818 11396 6874 11398
rect 6578 10362 6634 10364
rect 6658 10362 6714 10364
rect 6738 10362 6794 10364
rect 6818 10362 6874 10364
rect 6578 10310 6624 10362
rect 6624 10310 6634 10362
rect 6658 10310 6688 10362
rect 6688 10310 6700 10362
rect 6700 10310 6714 10362
rect 6738 10310 6752 10362
rect 6752 10310 6764 10362
rect 6764 10310 6794 10362
rect 6818 10310 6828 10362
rect 6828 10310 6874 10362
rect 6578 10308 6634 10310
rect 6658 10308 6714 10310
rect 6738 10308 6794 10310
rect 6818 10308 6874 10310
rect 6366 9968 6422 10024
rect 6578 9274 6634 9276
rect 6658 9274 6714 9276
rect 6738 9274 6794 9276
rect 6818 9274 6874 9276
rect 6578 9222 6624 9274
rect 6624 9222 6634 9274
rect 6658 9222 6688 9274
rect 6688 9222 6700 9274
rect 6700 9222 6714 9274
rect 6738 9222 6752 9274
rect 6752 9222 6764 9274
rect 6764 9222 6794 9274
rect 6818 9222 6828 9274
rect 6828 9222 6874 9274
rect 6578 9220 6634 9222
rect 6658 9220 6714 9222
rect 6738 9220 6794 9222
rect 6818 9220 6874 9222
rect 6578 8186 6634 8188
rect 6658 8186 6714 8188
rect 6738 8186 6794 8188
rect 6818 8186 6874 8188
rect 6578 8134 6624 8186
rect 6624 8134 6634 8186
rect 6658 8134 6688 8186
rect 6688 8134 6700 8186
rect 6700 8134 6714 8186
rect 6738 8134 6752 8186
rect 6752 8134 6764 8186
rect 6764 8134 6794 8186
rect 6818 8134 6828 8186
rect 6828 8134 6874 8186
rect 6578 8132 6634 8134
rect 6658 8132 6714 8134
rect 6738 8132 6794 8134
rect 6818 8132 6874 8134
rect 6578 7098 6634 7100
rect 6658 7098 6714 7100
rect 6738 7098 6794 7100
rect 6818 7098 6874 7100
rect 6578 7046 6624 7098
rect 6624 7046 6634 7098
rect 6658 7046 6688 7098
rect 6688 7046 6700 7098
rect 6700 7046 6714 7098
rect 6738 7046 6752 7098
rect 6752 7046 6764 7098
rect 6764 7046 6794 7098
rect 6818 7046 6828 7098
rect 6828 7046 6874 7098
rect 6578 7044 6634 7046
rect 6658 7044 6714 7046
rect 6738 7044 6794 7046
rect 6818 7044 6874 7046
rect 6578 6010 6634 6012
rect 6658 6010 6714 6012
rect 6738 6010 6794 6012
rect 6818 6010 6874 6012
rect 6578 5958 6624 6010
rect 6624 5958 6634 6010
rect 6658 5958 6688 6010
rect 6688 5958 6700 6010
rect 6700 5958 6714 6010
rect 6738 5958 6752 6010
rect 6752 5958 6764 6010
rect 6764 5958 6794 6010
rect 6818 5958 6828 6010
rect 6828 5958 6874 6010
rect 6578 5956 6634 5958
rect 6658 5956 6714 5958
rect 6738 5956 6794 5958
rect 6818 5956 6874 5958
rect 6578 4922 6634 4924
rect 6658 4922 6714 4924
rect 6738 4922 6794 4924
rect 6818 4922 6874 4924
rect 6578 4870 6624 4922
rect 6624 4870 6634 4922
rect 6658 4870 6688 4922
rect 6688 4870 6700 4922
rect 6700 4870 6714 4922
rect 6738 4870 6752 4922
rect 6752 4870 6764 4922
rect 6764 4870 6794 4922
rect 6818 4870 6828 4922
rect 6828 4870 6874 4922
rect 6578 4868 6634 4870
rect 6658 4868 6714 4870
rect 6738 4868 6794 4870
rect 6818 4868 6874 4870
rect 6578 3834 6634 3836
rect 6658 3834 6714 3836
rect 6738 3834 6794 3836
rect 6818 3834 6874 3836
rect 6578 3782 6624 3834
rect 6624 3782 6634 3834
rect 6658 3782 6688 3834
rect 6688 3782 6700 3834
rect 6700 3782 6714 3834
rect 6738 3782 6752 3834
rect 6752 3782 6764 3834
rect 6764 3782 6794 3834
rect 6818 3782 6828 3834
rect 6828 3782 6874 3834
rect 6578 3780 6634 3782
rect 6658 3780 6714 3782
rect 6738 3780 6794 3782
rect 6818 3780 6874 3782
rect 6578 2746 6634 2748
rect 6658 2746 6714 2748
rect 6738 2746 6794 2748
rect 6818 2746 6874 2748
rect 6578 2694 6624 2746
rect 6624 2694 6634 2746
rect 6658 2694 6688 2746
rect 6688 2694 6700 2746
rect 6700 2694 6714 2746
rect 6738 2694 6752 2746
rect 6752 2694 6764 2746
rect 6764 2694 6794 2746
rect 6818 2694 6828 2746
rect 6828 2694 6874 2746
rect 6578 2692 6634 2694
rect 6658 2692 6714 2694
rect 6738 2692 6794 2694
rect 6818 2692 6874 2694
rect 6642 2388 6644 2408
rect 6644 2388 6696 2408
rect 6696 2388 6698 2408
rect 6642 2352 6698 2388
rect 7654 9424 7710 9480
rect 7838 2488 7894 2544
rect 8452 16346 8508 16348
rect 8532 16346 8588 16348
rect 8612 16346 8668 16348
rect 8692 16346 8748 16348
rect 8452 16294 8498 16346
rect 8498 16294 8508 16346
rect 8532 16294 8562 16346
rect 8562 16294 8574 16346
rect 8574 16294 8588 16346
rect 8612 16294 8626 16346
rect 8626 16294 8638 16346
rect 8638 16294 8668 16346
rect 8692 16294 8702 16346
rect 8702 16294 8748 16346
rect 8452 16292 8508 16294
rect 8532 16292 8588 16294
rect 8612 16292 8668 16294
rect 8692 16292 8748 16294
rect 8452 15258 8508 15260
rect 8532 15258 8588 15260
rect 8612 15258 8668 15260
rect 8692 15258 8748 15260
rect 8452 15206 8498 15258
rect 8498 15206 8508 15258
rect 8532 15206 8562 15258
rect 8562 15206 8574 15258
rect 8574 15206 8588 15258
rect 8612 15206 8626 15258
rect 8626 15206 8638 15258
rect 8638 15206 8668 15258
rect 8692 15206 8702 15258
rect 8702 15206 8748 15258
rect 8452 15204 8508 15206
rect 8532 15204 8588 15206
rect 8612 15204 8668 15206
rect 8692 15204 8748 15206
rect 8452 14170 8508 14172
rect 8532 14170 8588 14172
rect 8612 14170 8668 14172
rect 8692 14170 8748 14172
rect 8452 14118 8498 14170
rect 8498 14118 8508 14170
rect 8532 14118 8562 14170
rect 8562 14118 8574 14170
rect 8574 14118 8588 14170
rect 8612 14118 8626 14170
rect 8626 14118 8638 14170
rect 8638 14118 8668 14170
rect 8692 14118 8702 14170
rect 8702 14118 8748 14170
rect 8452 14116 8508 14118
rect 8532 14116 8588 14118
rect 8612 14116 8668 14118
rect 8692 14116 8748 14118
rect 8452 13082 8508 13084
rect 8532 13082 8588 13084
rect 8612 13082 8668 13084
rect 8692 13082 8748 13084
rect 8452 13030 8498 13082
rect 8498 13030 8508 13082
rect 8532 13030 8562 13082
rect 8562 13030 8574 13082
rect 8574 13030 8588 13082
rect 8612 13030 8626 13082
rect 8626 13030 8638 13082
rect 8638 13030 8668 13082
rect 8692 13030 8702 13082
rect 8702 13030 8748 13082
rect 8452 13028 8508 13030
rect 8532 13028 8588 13030
rect 8612 13028 8668 13030
rect 8692 13028 8748 13030
rect 8206 10512 8262 10568
rect 8452 11994 8508 11996
rect 8532 11994 8588 11996
rect 8612 11994 8668 11996
rect 8692 11994 8748 11996
rect 8452 11942 8498 11994
rect 8498 11942 8508 11994
rect 8532 11942 8562 11994
rect 8562 11942 8574 11994
rect 8574 11942 8588 11994
rect 8612 11942 8626 11994
rect 8626 11942 8638 11994
rect 8638 11942 8668 11994
rect 8692 11942 8702 11994
rect 8702 11942 8748 11994
rect 8452 11940 8508 11942
rect 8532 11940 8588 11942
rect 8612 11940 8668 11942
rect 8692 11940 8748 11942
rect 8452 10906 8508 10908
rect 8532 10906 8588 10908
rect 8612 10906 8668 10908
rect 8692 10906 8748 10908
rect 8452 10854 8498 10906
rect 8498 10854 8508 10906
rect 8532 10854 8562 10906
rect 8562 10854 8574 10906
rect 8574 10854 8588 10906
rect 8612 10854 8626 10906
rect 8626 10854 8638 10906
rect 8638 10854 8668 10906
rect 8692 10854 8702 10906
rect 8702 10854 8748 10906
rect 8452 10852 8508 10854
rect 8532 10852 8588 10854
rect 8612 10852 8668 10854
rect 8692 10852 8748 10854
rect 8452 9818 8508 9820
rect 8532 9818 8588 9820
rect 8612 9818 8668 9820
rect 8692 9818 8748 9820
rect 8452 9766 8498 9818
rect 8498 9766 8508 9818
rect 8532 9766 8562 9818
rect 8562 9766 8574 9818
rect 8574 9766 8588 9818
rect 8612 9766 8626 9818
rect 8626 9766 8638 9818
rect 8638 9766 8668 9818
rect 8692 9766 8702 9818
rect 8702 9766 8748 9818
rect 8452 9764 8508 9766
rect 8532 9764 8588 9766
rect 8612 9764 8668 9766
rect 8692 9764 8748 9766
rect 8390 8880 8446 8936
rect 8452 8730 8508 8732
rect 8532 8730 8588 8732
rect 8612 8730 8668 8732
rect 8692 8730 8748 8732
rect 8452 8678 8498 8730
rect 8498 8678 8508 8730
rect 8532 8678 8562 8730
rect 8562 8678 8574 8730
rect 8574 8678 8588 8730
rect 8612 8678 8626 8730
rect 8626 8678 8638 8730
rect 8638 8678 8668 8730
rect 8692 8678 8702 8730
rect 8702 8678 8748 8730
rect 8452 8676 8508 8678
rect 8532 8676 8588 8678
rect 8612 8676 8668 8678
rect 8692 8676 8748 8678
rect 8452 7642 8508 7644
rect 8532 7642 8588 7644
rect 8612 7642 8668 7644
rect 8692 7642 8748 7644
rect 8452 7590 8498 7642
rect 8498 7590 8508 7642
rect 8532 7590 8562 7642
rect 8562 7590 8574 7642
rect 8574 7590 8588 7642
rect 8612 7590 8626 7642
rect 8626 7590 8638 7642
rect 8638 7590 8668 7642
rect 8692 7590 8702 7642
rect 8702 7590 8748 7642
rect 8452 7588 8508 7590
rect 8532 7588 8588 7590
rect 8612 7588 8668 7590
rect 8692 7588 8748 7590
rect 8452 6554 8508 6556
rect 8532 6554 8588 6556
rect 8612 6554 8668 6556
rect 8692 6554 8748 6556
rect 8452 6502 8498 6554
rect 8498 6502 8508 6554
rect 8532 6502 8562 6554
rect 8562 6502 8574 6554
rect 8574 6502 8588 6554
rect 8612 6502 8626 6554
rect 8626 6502 8638 6554
rect 8638 6502 8668 6554
rect 8692 6502 8702 6554
rect 8702 6502 8748 6554
rect 8452 6500 8508 6502
rect 8532 6500 8588 6502
rect 8612 6500 8668 6502
rect 8692 6500 8748 6502
rect 8452 5466 8508 5468
rect 8532 5466 8588 5468
rect 8612 5466 8668 5468
rect 8692 5466 8748 5468
rect 8452 5414 8498 5466
rect 8498 5414 8508 5466
rect 8532 5414 8562 5466
rect 8562 5414 8574 5466
rect 8574 5414 8588 5466
rect 8612 5414 8626 5466
rect 8626 5414 8638 5466
rect 8638 5414 8668 5466
rect 8692 5414 8702 5466
rect 8702 5414 8748 5466
rect 8452 5412 8508 5414
rect 8532 5412 8588 5414
rect 8612 5412 8668 5414
rect 8692 5412 8748 5414
rect 8452 4378 8508 4380
rect 8532 4378 8588 4380
rect 8612 4378 8668 4380
rect 8692 4378 8748 4380
rect 8452 4326 8498 4378
rect 8498 4326 8508 4378
rect 8532 4326 8562 4378
rect 8562 4326 8574 4378
rect 8574 4326 8588 4378
rect 8612 4326 8626 4378
rect 8626 4326 8638 4378
rect 8638 4326 8668 4378
rect 8692 4326 8702 4378
rect 8702 4326 8748 4378
rect 8452 4324 8508 4326
rect 8532 4324 8588 4326
rect 8612 4324 8668 4326
rect 8692 4324 8748 4326
rect 8452 3290 8508 3292
rect 8532 3290 8588 3292
rect 8612 3290 8668 3292
rect 8692 3290 8748 3292
rect 8452 3238 8498 3290
rect 8498 3238 8508 3290
rect 8532 3238 8562 3290
rect 8562 3238 8574 3290
rect 8574 3238 8588 3290
rect 8612 3238 8626 3290
rect 8626 3238 8638 3290
rect 8638 3238 8668 3290
rect 8692 3238 8702 3290
rect 8702 3238 8748 3290
rect 8452 3236 8508 3238
rect 8532 3236 8588 3238
rect 8612 3236 8668 3238
rect 8692 3236 8748 3238
rect 8666 2624 8722 2680
rect 9126 9696 9182 9752
rect 9034 8880 9090 8936
rect 9310 9460 9312 9480
rect 9312 9460 9364 9480
rect 9364 9460 9366 9480
rect 9310 9424 9366 9460
rect 8206 1944 8262 2000
rect 8114 1536 8170 1592
rect 8452 2202 8508 2204
rect 8532 2202 8588 2204
rect 8612 2202 8668 2204
rect 8692 2202 8748 2204
rect 8452 2150 8498 2202
rect 8498 2150 8508 2202
rect 8532 2150 8562 2202
rect 8562 2150 8574 2202
rect 8574 2150 8588 2202
rect 8612 2150 8626 2202
rect 8626 2150 8638 2202
rect 8638 2150 8668 2202
rect 8692 2150 8702 2202
rect 8702 2150 8748 2202
rect 8452 2148 8508 2150
rect 8532 2148 8588 2150
rect 8612 2148 8668 2150
rect 8692 2148 8748 2150
rect 10326 16890 10382 16892
rect 10406 16890 10462 16892
rect 10486 16890 10542 16892
rect 10566 16890 10622 16892
rect 10326 16838 10372 16890
rect 10372 16838 10382 16890
rect 10406 16838 10436 16890
rect 10436 16838 10448 16890
rect 10448 16838 10462 16890
rect 10486 16838 10500 16890
rect 10500 16838 10512 16890
rect 10512 16838 10542 16890
rect 10566 16838 10576 16890
rect 10576 16838 10622 16890
rect 10326 16836 10382 16838
rect 10406 16836 10462 16838
rect 10486 16836 10542 16838
rect 10566 16836 10622 16838
rect 10326 15802 10382 15804
rect 10406 15802 10462 15804
rect 10486 15802 10542 15804
rect 10566 15802 10622 15804
rect 10326 15750 10372 15802
rect 10372 15750 10382 15802
rect 10406 15750 10436 15802
rect 10436 15750 10448 15802
rect 10448 15750 10462 15802
rect 10486 15750 10500 15802
rect 10500 15750 10512 15802
rect 10512 15750 10542 15802
rect 10566 15750 10576 15802
rect 10576 15750 10622 15802
rect 10326 15748 10382 15750
rect 10406 15748 10462 15750
rect 10486 15748 10542 15750
rect 10566 15748 10622 15750
rect 10326 14714 10382 14716
rect 10406 14714 10462 14716
rect 10486 14714 10542 14716
rect 10566 14714 10622 14716
rect 10326 14662 10372 14714
rect 10372 14662 10382 14714
rect 10406 14662 10436 14714
rect 10436 14662 10448 14714
rect 10448 14662 10462 14714
rect 10486 14662 10500 14714
rect 10500 14662 10512 14714
rect 10512 14662 10542 14714
rect 10566 14662 10576 14714
rect 10576 14662 10622 14714
rect 10326 14660 10382 14662
rect 10406 14660 10462 14662
rect 10486 14660 10542 14662
rect 10566 14660 10622 14662
rect 10326 13626 10382 13628
rect 10406 13626 10462 13628
rect 10486 13626 10542 13628
rect 10566 13626 10622 13628
rect 10326 13574 10372 13626
rect 10372 13574 10382 13626
rect 10406 13574 10436 13626
rect 10436 13574 10448 13626
rect 10448 13574 10462 13626
rect 10486 13574 10500 13626
rect 10500 13574 10512 13626
rect 10512 13574 10542 13626
rect 10566 13574 10576 13626
rect 10576 13574 10622 13626
rect 10326 13572 10382 13574
rect 10406 13572 10462 13574
rect 10486 13572 10542 13574
rect 10566 13572 10622 13574
rect 10326 12538 10382 12540
rect 10406 12538 10462 12540
rect 10486 12538 10542 12540
rect 10566 12538 10622 12540
rect 10326 12486 10372 12538
rect 10372 12486 10382 12538
rect 10406 12486 10436 12538
rect 10436 12486 10448 12538
rect 10448 12486 10462 12538
rect 10486 12486 10500 12538
rect 10500 12486 10512 12538
rect 10512 12486 10542 12538
rect 10566 12486 10576 12538
rect 10576 12486 10622 12538
rect 10326 12484 10382 12486
rect 10406 12484 10462 12486
rect 10486 12484 10542 12486
rect 10566 12484 10622 12486
rect 10326 11450 10382 11452
rect 10406 11450 10462 11452
rect 10486 11450 10542 11452
rect 10566 11450 10622 11452
rect 10326 11398 10372 11450
rect 10372 11398 10382 11450
rect 10406 11398 10436 11450
rect 10436 11398 10448 11450
rect 10448 11398 10462 11450
rect 10486 11398 10500 11450
rect 10500 11398 10512 11450
rect 10512 11398 10542 11450
rect 10566 11398 10576 11450
rect 10576 11398 10622 11450
rect 10326 11396 10382 11398
rect 10406 11396 10462 11398
rect 10486 11396 10542 11398
rect 10566 11396 10622 11398
rect 9494 2624 9550 2680
rect 9494 2216 9550 2272
rect 10326 10362 10382 10364
rect 10406 10362 10462 10364
rect 10486 10362 10542 10364
rect 10566 10362 10622 10364
rect 10326 10310 10372 10362
rect 10372 10310 10382 10362
rect 10406 10310 10436 10362
rect 10436 10310 10448 10362
rect 10448 10310 10462 10362
rect 10486 10310 10500 10362
rect 10500 10310 10512 10362
rect 10512 10310 10542 10362
rect 10566 10310 10576 10362
rect 10576 10310 10622 10362
rect 10326 10308 10382 10310
rect 10406 10308 10462 10310
rect 10486 10308 10542 10310
rect 10566 10308 10622 10310
rect 10326 9274 10382 9276
rect 10406 9274 10462 9276
rect 10486 9274 10542 9276
rect 10566 9274 10622 9276
rect 10326 9222 10372 9274
rect 10372 9222 10382 9274
rect 10406 9222 10436 9274
rect 10436 9222 10448 9274
rect 10448 9222 10462 9274
rect 10486 9222 10500 9274
rect 10500 9222 10512 9274
rect 10512 9222 10542 9274
rect 10566 9222 10576 9274
rect 10576 9222 10622 9274
rect 10326 9220 10382 9222
rect 10406 9220 10462 9222
rect 10486 9220 10542 9222
rect 10566 9220 10622 9222
rect 12200 17434 12256 17436
rect 12280 17434 12336 17436
rect 12360 17434 12416 17436
rect 12440 17434 12496 17436
rect 12200 17382 12246 17434
rect 12246 17382 12256 17434
rect 12280 17382 12310 17434
rect 12310 17382 12322 17434
rect 12322 17382 12336 17434
rect 12360 17382 12374 17434
rect 12374 17382 12386 17434
rect 12386 17382 12416 17434
rect 12440 17382 12450 17434
rect 12450 17382 12496 17434
rect 12200 17380 12256 17382
rect 12280 17380 12336 17382
rect 12360 17380 12416 17382
rect 12440 17380 12496 17382
rect 10326 8186 10382 8188
rect 10406 8186 10462 8188
rect 10486 8186 10542 8188
rect 10566 8186 10622 8188
rect 10326 8134 10372 8186
rect 10372 8134 10382 8186
rect 10406 8134 10436 8186
rect 10436 8134 10448 8186
rect 10448 8134 10462 8186
rect 10486 8134 10500 8186
rect 10500 8134 10512 8186
rect 10512 8134 10542 8186
rect 10566 8134 10576 8186
rect 10576 8134 10622 8186
rect 10326 8132 10382 8134
rect 10406 8132 10462 8134
rect 10486 8132 10542 8134
rect 10566 8132 10622 8134
rect 10326 7098 10382 7100
rect 10406 7098 10462 7100
rect 10486 7098 10542 7100
rect 10566 7098 10622 7100
rect 10326 7046 10372 7098
rect 10372 7046 10382 7098
rect 10406 7046 10436 7098
rect 10436 7046 10448 7098
rect 10448 7046 10462 7098
rect 10486 7046 10500 7098
rect 10500 7046 10512 7098
rect 10512 7046 10542 7098
rect 10566 7046 10576 7098
rect 10576 7046 10622 7098
rect 10326 7044 10382 7046
rect 10406 7044 10462 7046
rect 10486 7044 10542 7046
rect 10566 7044 10622 7046
rect 10326 6010 10382 6012
rect 10406 6010 10462 6012
rect 10486 6010 10542 6012
rect 10566 6010 10622 6012
rect 10326 5958 10372 6010
rect 10372 5958 10382 6010
rect 10406 5958 10436 6010
rect 10436 5958 10448 6010
rect 10448 5958 10462 6010
rect 10486 5958 10500 6010
rect 10500 5958 10512 6010
rect 10512 5958 10542 6010
rect 10566 5958 10576 6010
rect 10576 5958 10622 6010
rect 10326 5956 10382 5958
rect 10406 5956 10462 5958
rect 10486 5956 10542 5958
rect 10566 5956 10622 5958
rect 10326 4922 10382 4924
rect 10406 4922 10462 4924
rect 10486 4922 10542 4924
rect 10566 4922 10622 4924
rect 10326 4870 10372 4922
rect 10372 4870 10382 4922
rect 10406 4870 10436 4922
rect 10436 4870 10448 4922
rect 10448 4870 10462 4922
rect 10486 4870 10500 4922
rect 10500 4870 10512 4922
rect 10512 4870 10542 4922
rect 10566 4870 10576 4922
rect 10576 4870 10622 4922
rect 10326 4868 10382 4870
rect 10406 4868 10462 4870
rect 10486 4868 10542 4870
rect 10566 4868 10622 4870
rect 10326 3834 10382 3836
rect 10406 3834 10462 3836
rect 10486 3834 10542 3836
rect 10566 3834 10622 3836
rect 10326 3782 10372 3834
rect 10372 3782 10382 3834
rect 10406 3782 10436 3834
rect 10436 3782 10448 3834
rect 10448 3782 10462 3834
rect 10486 3782 10500 3834
rect 10500 3782 10512 3834
rect 10512 3782 10542 3834
rect 10566 3782 10576 3834
rect 10576 3782 10622 3834
rect 10326 3780 10382 3782
rect 10406 3780 10462 3782
rect 10486 3780 10542 3782
rect 10566 3780 10622 3782
rect 10326 2746 10382 2748
rect 10406 2746 10462 2748
rect 10486 2746 10542 2748
rect 10566 2746 10622 2748
rect 10326 2694 10372 2746
rect 10372 2694 10382 2746
rect 10406 2694 10436 2746
rect 10436 2694 10448 2746
rect 10448 2694 10462 2746
rect 10486 2694 10500 2746
rect 10500 2694 10512 2746
rect 10512 2694 10542 2746
rect 10566 2694 10576 2746
rect 10576 2694 10622 2746
rect 10326 2692 10382 2694
rect 10406 2692 10462 2694
rect 10486 2692 10542 2694
rect 10566 2692 10622 2694
rect 11426 9968 11482 10024
rect 10230 1808 10286 1864
rect 12200 16346 12256 16348
rect 12280 16346 12336 16348
rect 12360 16346 12416 16348
rect 12440 16346 12496 16348
rect 12200 16294 12246 16346
rect 12246 16294 12256 16346
rect 12280 16294 12310 16346
rect 12310 16294 12322 16346
rect 12322 16294 12336 16346
rect 12360 16294 12374 16346
rect 12374 16294 12386 16346
rect 12386 16294 12416 16346
rect 12440 16294 12450 16346
rect 12450 16294 12496 16346
rect 12200 16292 12256 16294
rect 12280 16292 12336 16294
rect 12360 16292 12416 16294
rect 12440 16292 12496 16294
rect 12200 15258 12256 15260
rect 12280 15258 12336 15260
rect 12360 15258 12416 15260
rect 12440 15258 12496 15260
rect 12200 15206 12246 15258
rect 12246 15206 12256 15258
rect 12280 15206 12310 15258
rect 12310 15206 12322 15258
rect 12322 15206 12336 15258
rect 12360 15206 12374 15258
rect 12374 15206 12386 15258
rect 12386 15206 12416 15258
rect 12440 15206 12450 15258
rect 12450 15206 12496 15258
rect 12200 15204 12256 15206
rect 12280 15204 12336 15206
rect 12360 15204 12416 15206
rect 12440 15204 12496 15206
rect 12200 14170 12256 14172
rect 12280 14170 12336 14172
rect 12360 14170 12416 14172
rect 12440 14170 12496 14172
rect 12200 14118 12246 14170
rect 12246 14118 12256 14170
rect 12280 14118 12310 14170
rect 12310 14118 12322 14170
rect 12322 14118 12336 14170
rect 12360 14118 12374 14170
rect 12374 14118 12386 14170
rect 12386 14118 12416 14170
rect 12440 14118 12450 14170
rect 12450 14118 12496 14170
rect 12200 14116 12256 14118
rect 12280 14116 12336 14118
rect 12360 14116 12416 14118
rect 12440 14116 12496 14118
rect 12200 13082 12256 13084
rect 12280 13082 12336 13084
rect 12360 13082 12416 13084
rect 12440 13082 12496 13084
rect 12200 13030 12246 13082
rect 12246 13030 12256 13082
rect 12280 13030 12310 13082
rect 12310 13030 12322 13082
rect 12322 13030 12336 13082
rect 12360 13030 12374 13082
rect 12374 13030 12386 13082
rect 12386 13030 12416 13082
rect 12440 13030 12450 13082
rect 12450 13030 12496 13082
rect 12200 13028 12256 13030
rect 12280 13028 12336 13030
rect 12360 13028 12416 13030
rect 12440 13028 12496 13030
rect 12200 11994 12256 11996
rect 12280 11994 12336 11996
rect 12360 11994 12416 11996
rect 12440 11994 12496 11996
rect 12200 11942 12246 11994
rect 12246 11942 12256 11994
rect 12280 11942 12310 11994
rect 12310 11942 12322 11994
rect 12322 11942 12336 11994
rect 12360 11942 12374 11994
rect 12374 11942 12386 11994
rect 12386 11942 12416 11994
rect 12440 11942 12450 11994
rect 12450 11942 12496 11994
rect 12200 11940 12256 11942
rect 12280 11940 12336 11942
rect 12360 11940 12416 11942
rect 12440 11940 12496 11942
rect 12200 10906 12256 10908
rect 12280 10906 12336 10908
rect 12360 10906 12416 10908
rect 12440 10906 12496 10908
rect 12200 10854 12246 10906
rect 12246 10854 12256 10906
rect 12280 10854 12310 10906
rect 12310 10854 12322 10906
rect 12322 10854 12336 10906
rect 12360 10854 12374 10906
rect 12374 10854 12386 10906
rect 12386 10854 12416 10906
rect 12440 10854 12450 10906
rect 12450 10854 12496 10906
rect 12200 10852 12256 10854
rect 12280 10852 12336 10854
rect 12360 10852 12416 10854
rect 12440 10852 12496 10854
rect 11242 2352 11298 2408
rect 12530 10512 12586 10568
rect 11886 2488 11942 2544
rect 12200 9818 12256 9820
rect 12280 9818 12336 9820
rect 12360 9818 12416 9820
rect 12440 9818 12496 9820
rect 12200 9766 12246 9818
rect 12246 9766 12256 9818
rect 12280 9766 12310 9818
rect 12310 9766 12322 9818
rect 12322 9766 12336 9818
rect 12360 9766 12374 9818
rect 12374 9766 12386 9818
rect 12386 9766 12416 9818
rect 12440 9766 12450 9818
rect 12450 9766 12496 9818
rect 12200 9764 12256 9766
rect 12280 9764 12336 9766
rect 12360 9764 12416 9766
rect 12440 9764 12496 9766
rect 12200 8730 12256 8732
rect 12280 8730 12336 8732
rect 12360 8730 12416 8732
rect 12440 8730 12496 8732
rect 12200 8678 12246 8730
rect 12246 8678 12256 8730
rect 12280 8678 12310 8730
rect 12310 8678 12322 8730
rect 12322 8678 12336 8730
rect 12360 8678 12374 8730
rect 12374 8678 12386 8730
rect 12386 8678 12416 8730
rect 12440 8678 12450 8730
rect 12450 8678 12496 8730
rect 12200 8676 12256 8678
rect 12280 8676 12336 8678
rect 12360 8676 12416 8678
rect 12440 8676 12496 8678
rect 12200 7642 12256 7644
rect 12280 7642 12336 7644
rect 12360 7642 12416 7644
rect 12440 7642 12496 7644
rect 12200 7590 12246 7642
rect 12246 7590 12256 7642
rect 12280 7590 12310 7642
rect 12310 7590 12322 7642
rect 12322 7590 12336 7642
rect 12360 7590 12374 7642
rect 12374 7590 12386 7642
rect 12386 7590 12416 7642
rect 12440 7590 12450 7642
rect 12450 7590 12496 7642
rect 12200 7588 12256 7590
rect 12280 7588 12336 7590
rect 12360 7588 12416 7590
rect 12440 7588 12496 7590
rect 12200 6554 12256 6556
rect 12280 6554 12336 6556
rect 12360 6554 12416 6556
rect 12440 6554 12496 6556
rect 12200 6502 12246 6554
rect 12246 6502 12256 6554
rect 12280 6502 12310 6554
rect 12310 6502 12322 6554
rect 12322 6502 12336 6554
rect 12360 6502 12374 6554
rect 12374 6502 12386 6554
rect 12386 6502 12416 6554
rect 12440 6502 12450 6554
rect 12450 6502 12496 6554
rect 12200 6500 12256 6502
rect 12280 6500 12336 6502
rect 12360 6500 12416 6502
rect 12440 6500 12496 6502
rect 12200 5466 12256 5468
rect 12280 5466 12336 5468
rect 12360 5466 12416 5468
rect 12440 5466 12496 5468
rect 12200 5414 12246 5466
rect 12246 5414 12256 5466
rect 12280 5414 12310 5466
rect 12310 5414 12322 5466
rect 12322 5414 12336 5466
rect 12360 5414 12374 5466
rect 12374 5414 12386 5466
rect 12386 5414 12416 5466
rect 12440 5414 12450 5466
rect 12450 5414 12496 5466
rect 12200 5412 12256 5414
rect 12280 5412 12336 5414
rect 12360 5412 12416 5414
rect 12440 5412 12496 5414
rect 12200 4378 12256 4380
rect 12280 4378 12336 4380
rect 12360 4378 12416 4380
rect 12440 4378 12496 4380
rect 12200 4326 12246 4378
rect 12246 4326 12256 4378
rect 12280 4326 12310 4378
rect 12310 4326 12322 4378
rect 12322 4326 12336 4378
rect 12360 4326 12374 4378
rect 12374 4326 12386 4378
rect 12386 4326 12416 4378
rect 12440 4326 12450 4378
rect 12450 4326 12496 4378
rect 12200 4324 12256 4326
rect 12280 4324 12336 4326
rect 12360 4324 12416 4326
rect 12440 4324 12496 4326
rect 12200 3290 12256 3292
rect 12280 3290 12336 3292
rect 12360 3290 12416 3292
rect 12440 3290 12496 3292
rect 12200 3238 12246 3290
rect 12246 3238 12256 3290
rect 12280 3238 12310 3290
rect 12310 3238 12322 3290
rect 12322 3238 12336 3290
rect 12360 3238 12374 3290
rect 12374 3238 12386 3290
rect 12386 3238 12416 3290
rect 12440 3238 12450 3290
rect 12450 3238 12496 3290
rect 12200 3236 12256 3238
rect 12280 3236 12336 3238
rect 12360 3236 12416 3238
rect 12440 3236 12496 3238
rect 12200 2202 12256 2204
rect 12280 2202 12336 2204
rect 12360 2202 12416 2204
rect 12440 2202 12496 2204
rect 12200 2150 12246 2202
rect 12246 2150 12256 2202
rect 12280 2150 12310 2202
rect 12310 2150 12322 2202
rect 12322 2150 12336 2202
rect 12360 2150 12374 2202
rect 12374 2150 12386 2202
rect 12386 2150 12416 2202
rect 12440 2150 12450 2202
rect 12450 2150 12496 2202
rect 12200 2148 12256 2150
rect 12280 2148 12336 2150
rect 12360 2148 12416 2150
rect 12440 2148 12496 2150
rect 12070 1536 12126 1592
rect 12806 7384 12862 7440
rect 14074 16890 14130 16892
rect 14154 16890 14210 16892
rect 14234 16890 14290 16892
rect 14314 16890 14370 16892
rect 14074 16838 14120 16890
rect 14120 16838 14130 16890
rect 14154 16838 14184 16890
rect 14184 16838 14196 16890
rect 14196 16838 14210 16890
rect 14234 16838 14248 16890
rect 14248 16838 14260 16890
rect 14260 16838 14290 16890
rect 14314 16838 14324 16890
rect 14324 16838 14370 16890
rect 14074 16836 14130 16838
rect 14154 16836 14210 16838
rect 14234 16836 14290 16838
rect 14314 16836 14370 16838
rect 14074 15802 14130 15804
rect 14154 15802 14210 15804
rect 14234 15802 14290 15804
rect 14314 15802 14370 15804
rect 14074 15750 14120 15802
rect 14120 15750 14130 15802
rect 14154 15750 14184 15802
rect 14184 15750 14196 15802
rect 14196 15750 14210 15802
rect 14234 15750 14248 15802
rect 14248 15750 14260 15802
rect 14260 15750 14290 15802
rect 14314 15750 14324 15802
rect 14324 15750 14370 15802
rect 14074 15748 14130 15750
rect 14154 15748 14210 15750
rect 14234 15748 14290 15750
rect 14314 15748 14370 15750
rect 14074 14714 14130 14716
rect 14154 14714 14210 14716
rect 14234 14714 14290 14716
rect 14314 14714 14370 14716
rect 14074 14662 14120 14714
rect 14120 14662 14130 14714
rect 14154 14662 14184 14714
rect 14184 14662 14196 14714
rect 14196 14662 14210 14714
rect 14234 14662 14248 14714
rect 14248 14662 14260 14714
rect 14260 14662 14290 14714
rect 14314 14662 14324 14714
rect 14324 14662 14370 14714
rect 14074 14660 14130 14662
rect 14154 14660 14210 14662
rect 14234 14660 14290 14662
rect 14314 14660 14370 14662
rect 14074 13626 14130 13628
rect 14154 13626 14210 13628
rect 14234 13626 14290 13628
rect 14314 13626 14370 13628
rect 14074 13574 14120 13626
rect 14120 13574 14130 13626
rect 14154 13574 14184 13626
rect 14184 13574 14196 13626
rect 14196 13574 14210 13626
rect 14234 13574 14248 13626
rect 14248 13574 14260 13626
rect 14260 13574 14290 13626
rect 14314 13574 14324 13626
rect 14324 13574 14370 13626
rect 14074 13572 14130 13574
rect 14154 13572 14210 13574
rect 14234 13572 14290 13574
rect 14314 13572 14370 13574
rect 15566 17448 15622 17504
rect 14074 12538 14130 12540
rect 14154 12538 14210 12540
rect 14234 12538 14290 12540
rect 14314 12538 14370 12540
rect 14074 12486 14120 12538
rect 14120 12486 14130 12538
rect 14154 12486 14184 12538
rect 14184 12486 14196 12538
rect 14196 12486 14210 12538
rect 14234 12486 14248 12538
rect 14248 12486 14260 12538
rect 14260 12486 14290 12538
rect 14314 12486 14324 12538
rect 14324 12486 14370 12538
rect 14074 12484 14130 12486
rect 14154 12484 14210 12486
rect 14234 12484 14290 12486
rect 14314 12484 14370 12486
rect 14074 11450 14130 11452
rect 14154 11450 14210 11452
rect 14234 11450 14290 11452
rect 14314 11450 14370 11452
rect 14074 11398 14120 11450
rect 14120 11398 14130 11450
rect 14154 11398 14184 11450
rect 14184 11398 14196 11450
rect 14196 11398 14210 11450
rect 14234 11398 14248 11450
rect 14248 11398 14260 11450
rect 14260 11398 14290 11450
rect 14314 11398 14324 11450
rect 14324 11398 14370 11450
rect 14074 11396 14130 11398
rect 14154 11396 14210 11398
rect 14234 11396 14290 11398
rect 14314 11396 14370 11398
rect 14074 10362 14130 10364
rect 14154 10362 14210 10364
rect 14234 10362 14290 10364
rect 14314 10362 14370 10364
rect 14074 10310 14120 10362
rect 14120 10310 14130 10362
rect 14154 10310 14184 10362
rect 14184 10310 14196 10362
rect 14196 10310 14210 10362
rect 14234 10310 14248 10362
rect 14248 10310 14260 10362
rect 14260 10310 14290 10362
rect 14314 10310 14324 10362
rect 14324 10310 14370 10362
rect 14074 10308 14130 10310
rect 14154 10308 14210 10310
rect 14234 10308 14290 10310
rect 14314 10308 14370 10310
rect 15566 12416 15622 12472
rect 14074 9274 14130 9276
rect 14154 9274 14210 9276
rect 14234 9274 14290 9276
rect 14314 9274 14370 9276
rect 14074 9222 14120 9274
rect 14120 9222 14130 9274
rect 14154 9222 14184 9274
rect 14184 9222 14196 9274
rect 14196 9222 14210 9274
rect 14234 9222 14248 9274
rect 14248 9222 14260 9274
rect 14260 9222 14290 9274
rect 14314 9222 14324 9274
rect 14324 9222 14370 9274
rect 14074 9220 14130 9222
rect 14154 9220 14210 9222
rect 14234 9220 14290 9222
rect 14314 9220 14370 9222
rect 14074 8186 14130 8188
rect 14154 8186 14210 8188
rect 14234 8186 14290 8188
rect 14314 8186 14370 8188
rect 14074 8134 14120 8186
rect 14120 8134 14130 8186
rect 14154 8134 14184 8186
rect 14184 8134 14196 8186
rect 14196 8134 14210 8186
rect 14234 8134 14248 8186
rect 14248 8134 14260 8186
rect 14260 8134 14290 8186
rect 14314 8134 14324 8186
rect 14324 8134 14370 8186
rect 14074 8132 14130 8134
rect 14154 8132 14210 8134
rect 14234 8132 14290 8134
rect 14314 8132 14370 8134
rect 14074 7098 14130 7100
rect 14154 7098 14210 7100
rect 14234 7098 14290 7100
rect 14314 7098 14370 7100
rect 14074 7046 14120 7098
rect 14120 7046 14130 7098
rect 14154 7046 14184 7098
rect 14184 7046 14196 7098
rect 14196 7046 14210 7098
rect 14234 7046 14248 7098
rect 14248 7046 14260 7098
rect 14260 7046 14290 7098
rect 14314 7046 14324 7098
rect 14324 7046 14370 7098
rect 14074 7044 14130 7046
rect 14154 7044 14210 7046
rect 14234 7044 14290 7046
rect 14314 7044 14370 7046
rect 14074 6010 14130 6012
rect 14154 6010 14210 6012
rect 14234 6010 14290 6012
rect 14314 6010 14370 6012
rect 14074 5958 14120 6010
rect 14120 5958 14130 6010
rect 14154 5958 14184 6010
rect 14184 5958 14196 6010
rect 14196 5958 14210 6010
rect 14234 5958 14248 6010
rect 14248 5958 14260 6010
rect 14260 5958 14290 6010
rect 14314 5958 14324 6010
rect 14324 5958 14370 6010
rect 14074 5956 14130 5958
rect 14154 5956 14210 5958
rect 14234 5956 14290 5958
rect 14314 5956 14370 5958
rect 14074 4922 14130 4924
rect 14154 4922 14210 4924
rect 14234 4922 14290 4924
rect 14314 4922 14370 4924
rect 14074 4870 14120 4922
rect 14120 4870 14130 4922
rect 14154 4870 14184 4922
rect 14184 4870 14196 4922
rect 14196 4870 14210 4922
rect 14234 4870 14248 4922
rect 14248 4870 14260 4922
rect 14260 4870 14290 4922
rect 14314 4870 14324 4922
rect 14324 4870 14370 4922
rect 14074 4868 14130 4870
rect 14154 4868 14210 4870
rect 14234 4868 14290 4870
rect 14314 4868 14370 4870
rect 14074 3834 14130 3836
rect 14154 3834 14210 3836
rect 14234 3834 14290 3836
rect 14314 3834 14370 3836
rect 14074 3782 14120 3834
rect 14120 3782 14130 3834
rect 14154 3782 14184 3834
rect 14184 3782 14196 3834
rect 14196 3782 14210 3834
rect 14234 3782 14248 3834
rect 14248 3782 14260 3834
rect 14260 3782 14290 3834
rect 14314 3782 14324 3834
rect 14324 3782 14370 3834
rect 14074 3780 14130 3782
rect 14154 3780 14210 3782
rect 14234 3780 14290 3782
rect 14314 3780 14370 3782
rect 14074 2746 14130 2748
rect 14154 2746 14210 2748
rect 14234 2746 14290 2748
rect 14314 2746 14370 2748
rect 14074 2694 14120 2746
rect 14120 2694 14130 2746
rect 14154 2694 14184 2746
rect 14184 2694 14196 2746
rect 14196 2694 14210 2746
rect 14234 2694 14248 2746
rect 14248 2694 14260 2746
rect 14260 2694 14290 2746
rect 14314 2694 14324 2746
rect 14324 2694 14370 2746
rect 14074 2692 14130 2694
rect 14154 2692 14210 2694
rect 14234 2692 14290 2694
rect 14314 2692 14370 2694
rect 13358 2352 13414 2408
rect 13266 1672 13322 1728
<< metal3 >>
rect 0 18322 800 18352
rect 1945 18322 2011 18325
rect 0 18320 2011 18322
rect 0 18264 1950 18320
rect 2006 18264 2011 18320
rect 0 18262 2011 18264
rect 0 18232 800 18262
rect 1945 18259 2011 18262
rect 15561 17506 15627 17509
rect 16400 17506 17200 17536
rect 15561 17504 17200 17506
rect 15561 17448 15566 17504
rect 15622 17448 17200 17504
rect 15561 17446 17200 17448
rect 15561 17443 15627 17446
rect 4692 17440 5012 17441
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 17375 5012 17376
rect 8440 17440 8760 17441
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 17375 8760 17376
rect 12188 17440 12508 17441
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 16400 17416 17200 17446
rect 12188 17375 12508 17376
rect 2818 16896 3138 16897
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 16831 3138 16832
rect 6566 16896 6886 16897
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 16831 6886 16832
rect 10314 16896 10634 16897
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 16831 10634 16832
rect 14062 16896 14382 16897
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 16831 14382 16832
rect 4692 16352 5012 16353
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 16287 5012 16288
rect 8440 16352 8760 16353
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 16287 8760 16288
rect 12188 16352 12508 16353
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 16287 12508 16288
rect 2818 15808 3138 15809
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 15743 3138 15744
rect 6566 15808 6886 15809
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 15743 6886 15744
rect 10314 15808 10634 15809
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 15743 10634 15744
rect 14062 15808 14382 15809
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 15743 14382 15744
rect 4692 15264 5012 15265
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 15199 5012 15200
rect 8440 15264 8760 15265
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 15199 8760 15200
rect 12188 15264 12508 15265
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 15199 12508 15200
rect 0 15058 800 15088
rect 3141 15058 3207 15061
rect 0 15056 3207 15058
rect 0 15000 3146 15056
rect 3202 15000 3207 15056
rect 0 14998 3207 15000
rect 0 14968 800 14998
rect 3141 14995 3207 14998
rect 2818 14720 3138 14721
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 14655 3138 14656
rect 6566 14720 6886 14721
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 14655 6886 14656
rect 10314 14720 10634 14721
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 14655 10634 14656
rect 14062 14720 14382 14721
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 14655 14382 14656
rect 4692 14176 5012 14177
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 14111 5012 14112
rect 8440 14176 8760 14177
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 14111 8760 14112
rect 12188 14176 12508 14177
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 14111 12508 14112
rect 2818 13632 3138 13633
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 13567 3138 13568
rect 6566 13632 6886 13633
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 13567 6886 13568
rect 10314 13632 10634 13633
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 13567 10634 13568
rect 14062 13632 14382 13633
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 13567 14382 13568
rect 4692 13088 5012 13089
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 13023 5012 13024
rect 8440 13088 8760 13089
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 13023 8760 13024
rect 12188 13088 12508 13089
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 13023 12508 13024
rect 2818 12544 3138 12545
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 12479 3138 12480
rect 6566 12544 6886 12545
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 12479 6886 12480
rect 10314 12544 10634 12545
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 12479 10634 12480
rect 14062 12544 14382 12545
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 12479 14382 12480
rect 15561 12474 15627 12477
rect 16400 12474 17200 12504
rect 15561 12472 17200 12474
rect 15561 12416 15566 12472
rect 15622 12416 17200 12472
rect 15561 12414 17200 12416
rect 15561 12411 15627 12414
rect 16400 12384 17200 12414
rect 4692 12000 5012 12001
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 11935 5012 11936
rect 8440 12000 8760 12001
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 11935 8760 11936
rect 12188 12000 12508 12001
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 11935 12508 11936
rect 0 11658 800 11688
rect 1393 11658 1459 11661
rect 0 11656 1459 11658
rect 0 11600 1398 11656
rect 1454 11600 1459 11656
rect 0 11598 1459 11600
rect 0 11568 800 11598
rect 1393 11595 1459 11598
rect 2818 11456 3138 11457
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 11391 3138 11392
rect 6566 11456 6886 11457
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 11391 6886 11392
rect 10314 11456 10634 11457
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 11391 10634 11392
rect 14062 11456 14382 11457
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 11391 14382 11392
rect 4692 10912 5012 10913
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 10847 5012 10848
rect 8440 10912 8760 10913
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 10847 8760 10848
rect 12188 10912 12508 10913
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 10847 12508 10848
rect 8201 10570 8267 10573
rect 12525 10570 12591 10573
rect 8201 10568 12591 10570
rect 8201 10512 8206 10568
rect 8262 10512 12530 10568
rect 12586 10512 12591 10568
rect 8201 10510 12591 10512
rect 8201 10507 8267 10510
rect 12525 10507 12591 10510
rect 2818 10368 3138 10369
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 10303 3138 10304
rect 6566 10368 6886 10369
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 6566 10303 6886 10304
rect 10314 10368 10634 10369
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 10314 10303 10634 10304
rect 14062 10368 14382 10369
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 10303 14382 10304
rect 6361 10026 6427 10029
rect 11421 10026 11487 10029
rect 6361 10024 11487 10026
rect 6361 9968 6366 10024
rect 6422 9968 11426 10024
rect 11482 9968 11487 10024
rect 6361 9966 11487 9968
rect 6361 9963 6427 9966
rect 11421 9963 11487 9966
rect 4692 9824 5012 9825
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 9759 5012 9760
rect 8440 9824 8760 9825
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 9759 8760 9760
rect 12188 9824 12508 9825
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 9759 12508 9760
rect 5717 9756 5783 9757
rect 5717 9752 5764 9756
rect 5828 9754 5834 9756
rect 9121 9754 9187 9757
rect 9254 9754 9260 9756
rect 5717 9696 5722 9752
rect 5717 9692 5764 9696
rect 5828 9694 5874 9754
rect 9121 9752 9260 9754
rect 9121 9696 9126 9752
rect 9182 9696 9260 9752
rect 9121 9694 9260 9696
rect 5828 9692 5834 9694
rect 5717 9691 5783 9692
rect 9121 9691 9187 9694
rect 9254 9692 9260 9694
rect 9324 9692 9330 9756
rect 7649 9482 7715 9485
rect 9305 9482 9371 9485
rect 7649 9480 9371 9482
rect 7649 9424 7654 9480
rect 7710 9424 9310 9480
rect 9366 9424 9371 9480
rect 7649 9422 9371 9424
rect 7649 9419 7715 9422
rect 9305 9419 9371 9422
rect 2818 9280 3138 9281
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 9215 3138 9216
rect 6566 9280 6886 9281
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 9215 6886 9216
rect 10314 9280 10634 9281
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 9215 10634 9216
rect 14062 9280 14382 9281
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 9215 14382 9216
rect 8385 8938 8451 8941
rect 9029 8938 9095 8941
rect 8385 8936 9095 8938
rect 8385 8880 8390 8936
rect 8446 8880 9034 8936
rect 9090 8880 9095 8936
rect 8385 8878 9095 8880
rect 8385 8875 8451 8878
rect 9029 8875 9095 8878
rect 4692 8736 5012 8737
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 8671 5012 8672
rect 8440 8736 8760 8737
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 8671 8760 8672
rect 12188 8736 12508 8737
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 8671 12508 8672
rect 0 8394 800 8424
rect 1485 8394 1551 8397
rect 0 8392 1551 8394
rect 0 8336 1490 8392
rect 1546 8336 1551 8392
rect 0 8334 1551 8336
rect 0 8304 800 8334
rect 1485 8331 1551 8334
rect 2818 8192 3138 8193
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 8127 3138 8128
rect 6566 8192 6886 8193
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 8127 6886 8128
rect 10314 8192 10634 8193
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 8127 10634 8128
rect 14062 8192 14382 8193
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 8127 14382 8128
rect 4692 7648 5012 7649
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 7583 5012 7584
rect 8440 7648 8760 7649
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 7583 8760 7584
rect 12188 7648 12508 7649
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 7583 12508 7584
rect 12801 7442 12867 7445
rect 16400 7442 17200 7472
rect 12801 7440 17200 7442
rect 12801 7384 12806 7440
rect 12862 7384 17200 7440
rect 12801 7382 17200 7384
rect 12801 7379 12867 7382
rect 16400 7352 17200 7382
rect 2818 7104 3138 7105
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 7039 3138 7040
rect 6566 7104 6886 7105
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 7039 6886 7040
rect 10314 7104 10634 7105
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 7039 10634 7040
rect 14062 7104 14382 7105
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 7039 14382 7040
rect 4692 6560 5012 6561
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 6495 5012 6496
rect 8440 6560 8760 6561
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 6495 8760 6496
rect 12188 6560 12508 6561
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 6495 12508 6496
rect 2818 6016 3138 6017
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 5951 3138 5952
rect 6566 6016 6886 6017
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 5951 6886 5952
rect 10314 6016 10634 6017
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 5951 10634 5952
rect 14062 6016 14382 6017
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 5951 14382 5952
rect 4692 5472 5012 5473
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 5407 5012 5408
rect 8440 5472 8760 5473
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 5407 8760 5408
rect 12188 5472 12508 5473
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 5407 12508 5408
rect 0 4994 800 5024
rect 1485 4994 1551 4997
rect 0 4992 1551 4994
rect 0 4936 1490 4992
rect 1546 4936 1551 4992
rect 0 4934 1551 4936
rect 0 4904 800 4934
rect 1485 4931 1551 4934
rect 2818 4928 3138 4929
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 4863 3138 4864
rect 6566 4928 6886 4929
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 4863 6886 4864
rect 10314 4928 10634 4929
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 4863 10634 4864
rect 14062 4928 14382 4929
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 4863 14382 4864
rect 4692 4384 5012 4385
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 4319 5012 4320
rect 8440 4384 8760 4385
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 4319 8760 4320
rect 12188 4384 12508 4385
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 4319 12508 4320
rect 2818 3840 3138 3841
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 3775 3138 3776
rect 6566 3840 6886 3841
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 3775 6886 3776
rect 10314 3840 10634 3841
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10314 3775 10634 3776
rect 14062 3840 14382 3841
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 3775 14382 3776
rect 4692 3296 5012 3297
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 3231 5012 3232
rect 8440 3296 8760 3297
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 3231 8760 3232
rect 12188 3296 12508 3297
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 3231 12508 3232
rect 2818 2752 3138 2753
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2687 3138 2688
rect 6566 2752 6886 2753
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 6566 2687 6886 2688
rect 10314 2752 10634 2753
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2687 10634 2688
rect 14062 2752 14382 2753
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2687 14382 2688
rect 8661 2682 8727 2685
rect 9489 2682 9555 2685
rect 8661 2680 9555 2682
rect 8661 2624 8666 2680
rect 8722 2624 9494 2680
rect 9550 2624 9555 2680
rect 8661 2622 9555 2624
rect 8661 2619 8727 2622
rect 9489 2619 9555 2622
rect 2681 2546 2747 2549
rect 5758 2546 5764 2548
rect 2681 2544 5764 2546
rect 2681 2488 2686 2544
rect 2742 2488 5764 2544
rect 2681 2486 5764 2488
rect 2681 2483 2747 2486
rect 5758 2484 5764 2486
rect 5828 2484 5834 2548
rect 7833 2546 7899 2549
rect 11881 2546 11947 2549
rect 16400 2546 17200 2576
rect 7833 2544 11947 2546
rect 7833 2488 7838 2544
rect 7894 2488 11886 2544
rect 11942 2488 11947 2544
rect 7833 2486 11947 2488
rect 7833 2483 7899 2486
rect 11881 2483 11947 2486
rect 16254 2486 17200 2546
rect 6637 2410 6703 2413
rect 11237 2410 11303 2413
rect 13353 2410 13419 2413
rect 6637 2408 11303 2410
rect 6637 2352 6642 2408
rect 6698 2352 11242 2408
rect 11298 2352 11303 2408
rect 6637 2350 11303 2352
rect 6637 2347 6703 2350
rect 11237 2347 11303 2350
rect 12022 2408 13419 2410
rect 12022 2352 13358 2408
rect 13414 2352 13419 2408
rect 12022 2350 13419 2352
rect 9489 2274 9555 2277
rect 12022 2274 12082 2350
rect 13353 2347 13419 2350
rect 9489 2272 12082 2274
rect 9489 2216 9494 2272
rect 9550 2216 12082 2272
rect 9489 2214 12082 2216
rect 16254 2274 16314 2486
rect 16400 2456 17200 2486
rect 16254 2214 16498 2274
rect 9489 2211 9555 2214
rect 4692 2208 5012 2209
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2143 5012 2144
rect 8440 2208 8760 2209
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2143 8760 2144
rect 12188 2208 12508 2209
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2143 12508 2144
rect 8201 2002 8267 2005
rect 16438 2002 16498 2214
rect 8201 2000 16498 2002
rect 8201 1944 8206 2000
rect 8262 1944 16498 2000
rect 8201 1942 16498 1944
rect 8201 1939 8267 1942
rect 4613 1866 4679 1869
rect 10225 1866 10291 1869
rect 4613 1864 10291 1866
rect 4613 1808 4618 1864
rect 4674 1808 10230 1864
rect 10286 1808 10291 1864
rect 4613 1806 10291 1808
rect 4613 1803 4679 1806
rect 10225 1803 10291 1806
rect 0 1730 800 1760
rect 2129 1730 2195 1733
rect 0 1728 2195 1730
rect 0 1672 2134 1728
rect 2190 1672 2195 1728
rect 0 1670 2195 1672
rect 0 1640 800 1670
rect 2129 1667 2195 1670
rect 9254 1668 9260 1732
rect 9324 1730 9330 1732
rect 13261 1730 13327 1733
rect 9324 1728 13327 1730
rect 9324 1672 13266 1728
rect 13322 1672 13327 1728
rect 9324 1670 13327 1672
rect 9324 1668 9330 1670
rect 13261 1667 13327 1670
rect 8109 1594 8175 1597
rect 12065 1594 12131 1597
rect 8109 1592 12131 1594
rect 8109 1536 8114 1592
rect 8170 1536 12070 1592
rect 12126 1536 12131 1592
rect 8109 1534 12131 1536
rect 8109 1531 8175 1534
rect 12065 1531 12131 1534
<< via3 >>
rect 4700 17436 4764 17440
rect 4700 17380 4704 17436
rect 4704 17380 4760 17436
rect 4760 17380 4764 17436
rect 4700 17376 4764 17380
rect 4780 17436 4844 17440
rect 4780 17380 4784 17436
rect 4784 17380 4840 17436
rect 4840 17380 4844 17436
rect 4780 17376 4844 17380
rect 4860 17436 4924 17440
rect 4860 17380 4864 17436
rect 4864 17380 4920 17436
rect 4920 17380 4924 17436
rect 4860 17376 4924 17380
rect 4940 17436 5004 17440
rect 4940 17380 4944 17436
rect 4944 17380 5000 17436
rect 5000 17380 5004 17436
rect 4940 17376 5004 17380
rect 8448 17436 8512 17440
rect 8448 17380 8452 17436
rect 8452 17380 8508 17436
rect 8508 17380 8512 17436
rect 8448 17376 8512 17380
rect 8528 17436 8592 17440
rect 8528 17380 8532 17436
rect 8532 17380 8588 17436
rect 8588 17380 8592 17436
rect 8528 17376 8592 17380
rect 8608 17436 8672 17440
rect 8608 17380 8612 17436
rect 8612 17380 8668 17436
rect 8668 17380 8672 17436
rect 8608 17376 8672 17380
rect 8688 17436 8752 17440
rect 8688 17380 8692 17436
rect 8692 17380 8748 17436
rect 8748 17380 8752 17436
rect 8688 17376 8752 17380
rect 12196 17436 12260 17440
rect 12196 17380 12200 17436
rect 12200 17380 12256 17436
rect 12256 17380 12260 17436
rect 12196 17376 12260 17380
rect 12276 17436 12340 17440
rect 12276 17380 12280 17436
rect 12280 17380 12336 17436
rect 12336 17380 12340 17436
rect 12276 17376 12340 17380
rect 12356 17436 12420 17440
rect 12356 17380 12360 17436
rect 12360 17380 12416 17436
rect 12416 17380 12420 17436
rect 12356 17376 12420 17380
rect 12436 17436 12500 17440
rect 12436 17380 12440 17436
rect 12440 17380 12496 17436
rect 12496 17380 12500 17436
rect 12436 17376 12500 17380
rect 2826 16892 2890 16896
rect 2826 16836 2830 16892
rect 2830 16836 2886 16892
rect 2886 16836 2890 16892
rect 2826 16832 2890 16836
rect 2906 16892 2970 16896
rect 2906 16836 2910 16892
rect 2910 16836 2966 16892
rect 2966 16836 2970 16892
rect 2906 16832 2970 16836
rect 2986 16892 3050 16896
rect 2986 16836 2990 16892
rect 2990 16836 3046 16892
rect 3046 16836 3050 16892
rect 2986 16832 3050 16836
rect 3066 16892 3130 16896
rect 3066 16836 3070 16892
rect 3070 16836 3126 16892
rect 3126 16836 3130 16892
rect 3066 16832 3130 16836
rect 6574 16892 6638 16896
rect 6574 16836 6578 16892
rect 6578 16836 6634 16892
rect 6634 16836 6638 16892
rect 6574 16832 6638 16836
rect 6654 16892 6718 16896
rect 6654 16836 6658 16892
rect 6658 16836 6714 16892
rect 6714 16836 6718 16892
rect 6654 16832 6718 16836
rect 6734 16892 6798 16896
rect 6734 16836 6738 16892
rect 6738 16836 6794 16892
rect 6794 16836 6798 16892
rect 6734 16832 6798 16836
rect 6814 16892 6878 16896
rect 6814 16836 6818 16892
rect 6818 16836 6874 16892
rect 6874 16836 6878 16892
rect 6814 16832 6878 16836
rect 10322 16892 10386 16896
rect 10322 16836 10326 16892
rect 10326 16836 10382 16892
rect 10382 16836 10386 16892
rect 10322 16832 10386 16836
rect 10402 16892 10466 16896
rect 10402 16836 10406 16892
rect 10406 16836 10462 16892
rect 10462 16836 10466 16892
rect 10402 16832 10466 16836
rect 10482 16892 10546 16896
rect 10482 16836 10486 16892
rect 10486 16836 10542 16892
rect 10542 16836 10546 16892
rect 10482 16832 10546 16836
rect 10562 16892 10626 16896
rect 10562 16836 10566 16892
rect 10566 16836 10622 16892
rect 10622 16836 10626 16892
rect 10562 16832 10626 16836
rect 14070 16892 14134 16896
rect 14070 16836 14074 16892
rect 14074 16836 14130 16892
rect 14130 16836 14134 16892
rect 14070 16832 14134 16836
rect 14150 16892 14214 16896
rect 14150 16836 14154 16892
rect 14154 16836 14210 16892
rect 14210 16836 14214 16892
rect 14150 16832 14214 16836
rect 14230 16892 14294 16896
rect 14230 16836 14234 16892
rect 14234 16836 14290 16892
rect 14290 16836 14294 16892
rect 14230 16832 14294 16836
rect 14310 16892 14374 16896
rect 14310 16836 14314 16892
rect 14314 16836 14370 16892
rect 14370 16836 14374 16892
rect 14310 16832 14374 16836
rect 4700 16348 4764 16352
rect 4700 16292 4704 16348
rect 4704 16292 4760 16348
rect 4760 16292 4764 16348
rect 4700 16288 4764 16292
rect 4780 16348 4844 16352
rect 4780 16292 4784 16348
rect 4784 16292 4840 16348
rect 4840 16292 4844 16348
rect 4780 16288 4844 16292
rect 4860 16348 4924 16352
rect 4860 16292 4864 16348
rect 4864 16292 4920 16348
rect 4920 16292 4924 16348
rect 4860 16288 4924 16292
rect 4940 16348 5004 16352
rect 4940 16292 4944 16348
rect 4944 16292 5000 16348
rect 5000 16292 5004 16348
rect 4940 16288 5004 16292
rect 8448 16348 8512 16352
rect 8448 16292 8452 16348
rect 8452 16292 8508 16348
rect 8508 16292 8512 16348
rect 8448 16288 8512 16292
rect 8528 16348 8592 16352
rect 8528 16292 8532 16348
rect 8532 16292 8588 16348
rect 8588 16292 8592 16348
rect 8528 16288 8592 16292
rect 8608 16348 8672 16352
rect 8608 16292 8612 16348
rect 8612 16292 8668 16348
rect 8668 16292 8672 16348
rect 8608 16288 8672 16292
rect 8688 16348 8752 16352
rect 8688 16292 8692 16348
rect 8692 16292 8748 16348
rect 8748 16292 8752 16348
rect 8688 16288 8752 16292
rect 12196 16348 12260 16352
rect 12196 16292 12200 16348
rect 12200 16292 12256 16348
rect 12256 16292 12260 16348
rect 12196 16288 12260 16292
rect 12276 16348 12340 16352
rect 12276 16292 12280 16348
rect 12280 16292 12336 16348
rect 12336 16292 12340 16348
rect 12276 16288 12340 16292
rect 12356 16348 12420 16352
rect 12356 16292 12360 16348
rect 12360 16292 12416 16348
rect 12416 16292 12420 16348
rect 12356 16288 12420 16292
rect 12436 16348 12500 16352
rect 12436 16292 12440 16348
rect 12440 16292 12496 16348
rect 12496 16292 12500 16348
rect 12436 16288 12500 16292
rect 2826 15804 2890 15808
rect 2826 15748 2830 15804
rect 2830 15748 2886 15804
rect 2886 15748 2890 15804
rect 2826 15744 2890 15748
rect 2906 15804 2970 15808
rect 2906 15748 2910 15804
rect 2910 15748 2966 15804
rect 2966 15748 2970 15804
rect 2906 15744 2970 15748
rect 2986 15804 3050 15808
rect 2986 15748 2990 15804
rect 2990 15748 3046 15804
rect 3046 15748 3050 15804
rect 2986 15744 3050 15748
rect 3066 15804 3130 15808
rect 3066 15748 3070 15804
rect 3070 15748 3126 15804
rect 3126 15748 3130 15804
rect 3066 15744 3130 15748
rect 6574 15804 6638 15808
rect 6574 15748 6578 15804
rect 6578 15748 6634 15804
rect 6634 15748 6638 15804
rect 6574 15744 6638 15748
rect 6654 15804 6718 15808
rect 6654 15748 6658 15804
rect 6658 15748 6714 15804
rect 6714 15748 6718 15804
rect 6654 15744 6718 15748
rect 6734 15804 6798 15808
rect 6734 15748 6738 15804
rect 6738 15748 6794 15804
rect 6794 15748 6798 15804
rect 6734 15744 6798 15748
rect 6814 15804 6878 15808
rect 6814 15748 6818 15804
rect 6818 15748 6874 15804
rect 6874 15748 6878 15804
rect 6814 15744 6878 15748
rect 10322 15804 10386 15808
rect 10322 15748 10326 15804
rect 10326 15748 10382 15804
rect 10382 15748 10386 15804
rect 10322 15744 10386 15748
rect 10402 15804 10466 15808
rect 10402 15748 10406 15804
rect 10406 15748 10462 15804
rect 10462 15748 10466 15804
rect 10402 15744 10466 15748
rect 10482 15804 10546 15808
rect 10482 15748 10486 15804
rect 10486 15748 10542 15804
rect 10542 15748 10546 15804
rect 10482 15744 10546 15748
rect 10562 15804 10626 15808
rect 10562 15748 10566 15804
rect 10566 15748 10622 15804
rect 10622 15748 10626 15804
rect 10562 15744 10626 15748
rect 14070 15804 14134 15808
rect 14070 15748 14074 15804
rect 14074 15748 14130 15804
rect 14130 15748 14134 15804
rect 14070 15744 14134 15748
rect 14150 15804 14214 15808
rect 14150 15748 14154 15804
rect 14154 15748 14210 15804
rect 14210 15748 14214 15804
rect 14150 15744 14214 15748
rect 14230 15804 14294 15808
rect 14230 15748 14234 15804
rect 14234 15748 14290 15804
rect 14290 15748 14294 15804
rect 14230 15744 14294 15748
rect 14310 15804 14374 15808
rect 14310 15748 14314 15804
rect 14314 15748 14370 15804
rect 14370 15748 14374 15804
rect 14310 15744 14374 15748
rect 4700 15260 4764 15264
rect 4700 15204 4704 15260
rect 4704 15204 4760 15260
rect 4760 15204 4764 15260
rect 4700 15200 4764 15204
rect 4780 15260 4844 15264
rect 4780 15204 4784 15260
rect 4784 15204 4840 15260
rect 4840 15204 4844 15260
rect 4780 15200 4844 15204
rect 4860 15260 4924 15264
rect 4860 15204 4864 15260
rect 4864 15204 4920 15260
rect 4920 15204 4924 15260
rect 4860 15200 4924 15204
rect 4940 15260 5004 15264
rect 4940 15204 4944 15260
rect 4944 15204 5000 15260
rect 5000 15204 5004 15260
rect 4940 15200 5004 15204
rect 8448 15260 8512 15264
rect 8448 15204 8452 15260
rect 8452 15204 8508 15260
rect 8508 15204 8512 15260
rect 8448 15200 8512 15204
rect 8528 15260 8592 15264
rect 8528 15204 8532 15260
rect 8532 15204 8588 15260
rect 8588 15204 8592 15260
rect 8528 15200 8592 15204
rect 8608 15260 8672 15264
rect 8608 15204 8612 15260
rect 8612 15204 8668 15260
rect 8668 15204 8672 15260
rect 8608 15200 8672 15204
rect 8688 15260 8752 15264
rect 8688 15204 8692 15260
rect 8692 15204 8748 15260
rect 8748 15204 8752 15260
rect 8688 15200 8752 15204
rect 12196 15260 12260 15264
rect 12196 15204 12200 15260
rect 12200 15204 12256 15260
rect 12256 15204 12260 15260
rect 12196 15200 12260 15204
rect 12276 15260 12340 15264
rect 12276 15204 12280 15260
rect 12280 15204 12336 15260
rect 12336 15204 12340 15260
rect 12276 15200 12340 15204
rect 12356 15260 12420 15264
rect 12356 15204 12360 15260
rect 12360 15204 12416 15260
rect 12416 15204 12420 15260
rect 12356 15200 12420 15204
rect 12436 15260 12500 15264
rect 12436 15204 12440 15260
rect 12440 15204 12496 15260
rect 12496 15204 12500 15260
rect 12436 15200 12500 15204
rect 2826 14716 2890 14720
rect 2826 14660 2830 14716
rect 2830 14660 2886 14716
rect 2886 14660 2890 14716
rect 2826 14656 2890 14660
rect 2906 14716 2970 14720
rect 2906 14660 2910 14716
rect 2910 14660 2966 14716
rect 2966 14660 2970 14716
rect 2906 14656 2970 14660
rect 2986 14716 3050 14720
rect 2986 14660 2990 14716
rect 2990 14660 3046 14716
rect 3046 14660 3050 14716
rect 2986 14656 3050 14660
rect 3066 14716 3130 14720
rect 3066 14660 3070 14716
rect 3070 14660 3126 14716
rect 3126 14660 3130 14716
rect 3066 14656 3130 14660
rect 6574 14716 6638 14720
rect 6574 14660 6578 14716
rect 6578 14660 6634 14716
rect 6634 14660 6638 14716
rect 6574 14656 6638 14660
rect 6654 14716 6718 14720
rect 6654 14660 6658 14716
rect 6658 14660 6714 14716
rect 6714 14660 6718 14716
rect 6654 14656 6718 14660
rect 6734 14716 6798 14720
rect 6734 14660 6738 14716
rect 6738 14660 6794 14716
rect 6794 14660 6798 14716
rect 6734 14656 6798 14660
rect 6814 14716 6878 14720
rect 6814 14660 6818 14716
rect 6818 14660 6874 14716
rect 6874 14660 6878 14716
rect 6814 14656 6878 14660
rect 10322 14716 10386 14720
rect 10322 14660 10326 14716
rect 10326 14660 10382 14716
rect 10382 14660 10386 14716
rect 10322 14656 10386 14660
rect 10402 14716 10466 14720
rect 10402 14660 10406 14716
rect 10406 14660 10462 14716
rect 10462 14660 10466 14716
rect 10402 14656 10466 14660
rect 10482 14716 10546 14720
rect 10482 14660 10486 14716
rect 10486 14660 10542 14716
rect 10542 14660 10546 14716
rect 10482 14656 10546 14660
rect 10562 14716 10626 14720
rect 10562 14660 10566 14716
rect 10566 14660 10622 14716
rect 10622 14660 10626 14716
rect 10562 14656 10626 14660
rect 14070 14716 14134 14720
rect 14070 14660 14074 14716
rect 14074 14660 14130 14716
rect 14130 14660 14134 14716
rect 14070 14656 14134 14660
rect 14150 14716 14214 14720
rect 14150 14660 14154 14716
rect 14154 14660 14210 14716
rect 14210 14660 14214 14716
rect 14150 14656 14214 14660
rect 14230 14716 14294 14720
rect 14230 14660 14234 14716
rect 14234 14660 14290 14716
rect 14290 14660 14294 14716
rect 14230 14656 14294 14660
rect 14310 14716 14374 14720
rect 14310 14660 14314 14716
rect 14314 14660 14370 14716
rect 14370 14660 14374 14716
rect 14310 14656 14374 14660
rect 4700 14172 4764 14176
rect 4700 14116 4704 14172
rect 4704 14116 4760 14172
rect 4760 14116 4764 14172
rect 4700 14112 4764 14116
rect 4780 14172 4844 14176
rect 4780 14116 4784 14172
rect 4784 14116 4840 14172
rect 4840 14116 4844 14172
rect 4780 14112 4844 14116
rect 4860 14172 4924 14176
rect 4860 14116 4864 14172
rect 4864 14116 4920 14172
rect 4920 14116 4924 14172
rect 4860 14112 4924 14116
rect 4940 14172 5004 14176
rect 4940 14116 4944 14172
rect 4944 14116 5000 14172
rect 5000 14116 5004 14172
rect 4940 14112 5004 14116
rect 8448 14172 8512 14176
rect 8448 14116 8452 14172
rect 8452 14116 8508 14172
rect 8508 14116 8512 14172
rect 8448 14112 8512 14116
rect 8528 14172 8592 14176
rect 8528 14116 8532 14172
rect 8532 14116 8588 14172
rect 8588 14116 8592 14172
rect 8528 14112 8592 14116
rect 8608 14172 8672 14176
rect 8608 14116 8612 14172
rect 8612 14116 8668 14172
rect 8668 14116 8672 14172
rect 8608 14112 8672 14116
rect 8688 14172 8752 14176
rect 8688 14116 8692 14172
rect 8692 14116 8748 14172
rect 8748 14116 8752 14172
rect 8688 14112 8752 14116
rect 12196 14172 12260 14176
rect 12196 14116 12200 14172
rect 12200 14116 12256 14172
rect 12256 14116 12260 14172
rect 12196 14112 12260 14116
rect 12276 14172 12340 14176
rect 12276 14116 12280 14172
rect 12280 14116 12336 14172
rect 12336 14116 12340 14172
rect 12276 14112 12340 14116
rect 12356 14172 12420 14176
rect 12356 14116 12360 14172
rect 12360 14116 12416 14172
rect 12416 14116 12420 14172
rect 12356 14112 12420 14116
rect 12436 14172 12500 14176
rect 12436 14116 12440 14172
rect 12440 14116 12496 14172
rect 12496 14116 12500 14172
rect 12436 14112 12500 14116
rect 2826 13628 2890 13632
rect 2826 13572 2830 13628
rect 2830 13572 2886 13628
rect 2886 13572 2890 13628
rect 2826 13568 2890 13572
rect 2906 13628 2970 13632
rect 2906 13572 2910 13628
rect 2910 13572 2966 13628
rect 2966 13572 2970 13628
rect 2906 13568 2970 13572
rect 2986 13628 3050 13632
rect 2986 13572 2990 13628
rect 2990 13572 3046 13628
rect 3046 13572 3050 13628
rect 2986 13568 3050 13572
rect 3066 13628 3130 13632
rect 3066 13572 3070 13628
rect 3070 13572 3126 13628
rect 3126 13572 3130 13628
rect 3066 13568 3130 13572
rect 6574 13628 6638 13632
rect 6574 13572 6578 13628
rect 6578 13572 6634 13628
rect 6634 13572 6638 13628
rect 6574 13568 6638 13572
rect 6654 13628 6718 13632
rect 6654 13572 6658 13628
rect 6658 13572 6714 13628
rect 6714 13572 6718 13628
rect 6654 13568 6718 13572
rect 6734 13628 6798 13632
rect 6734 13572 6738 13628
rect 6738 13572 6794 13628
rect 6794 13572 6798 13628
rect 6734 13568 6798 13572
rect 6814 13628 6878 13632
rect 6814 13572 6818 13628
rect 6818 13572 6874 13628
rect 6874 13572 6878 13628
rect 6814 13568 6878 13572
rect 10322 13628 10386 13632
rect 10322 13572 10326 13628
rect 10326 13572 10382 13628
rect 10382 13572 10386 13628
rect 10322 13568 10386 13572
rect 10402 13628 10466 13632
rect 10402 13572 10406 13628
rect 10406 13572 10462 13628
rect 10462 13572 10466 13628
rect 10402 13568 10466 13572
rect 10482 13628 10546 13632
rect 10482 13572 10486 13628
rect 10486 13572 10542 13628
rect 10542 13572 10546 13628
rect 10482 13568 10546 13572
rect 10562 13628 10626 13632
rect 10562 13572 10566 13628
rect 10566 13572 10622 13628
rect 10622 13572 10626 13628
rect 10562 13568 10626 13572
rect 14070 13628 14134 13632
rect 14070 13572 14074 13628
rect 14074 13572 14130 13628
rect 14130 13572 14134 13628
rect 14070 13568 14134 13572
rect 14150 13628 14214 13632
rect 14150 13572 14154 13628
rect 14154 13572 14210 13628
rect 14210 13572 14214 13628
rect 14150 13568 14214 13572
rect 14230 13628 14294 13632
rect 14230 13572 14234 13628
rect 14234 13572 14290 13628
rect 14290 13572 14294 13628
rect 14230 13568 14294 13572
rect 14310 13628 14374 13632
rect 14310 13572 14314 13628
rect 14314 13572 14370 13628
rect 14370 13572 14374 13628
rect 14310 13568 14374 13572
rect 4700 13084 4764 13088
rect 4700 13028 4704 13084
rect 4704 13028 4760 13084
rect 4760 13028 4764 13084
rect 4700 13024 4764 13028
rect 4780 13084 4844 13088
rect 4780 13028 4784 13084
rect 4784 13028 4840 13084
rect 4840 13028 4844 13084
rect 4780 13024 4844 13028
rect 4860 13084 4924 13088
rect 4860 13028 4864 13084
rect 4864 13028 4920 13084
rect 4920 13028 4924 13084
rect 4860 13024 4924 13028
rect 4940 13084 5004 13088
rect 4940 13028 4944 13084
rect 4944 13028 5000 13084
rect 5000 13028 5004 13084
rect 4940 13024 5004 13028
rect 8448 13084 8512 13088
rect 8448 13028 8452 13084
rect 8452 13028 8508 13084
rect 8508 13028 8512 13084
rect 8448 13024 8512 13028
rect 8528 13084 8592 13088
rect 8528 13028 8532 13084
rect 8532 13028 8588 13084
rect 8588 13028 8592 13084
rect 8528 13024 8592 13028
rect 8608 13084 8672 13088
rect 8608 13028 8612 13084
rect 8612 13028 8668 13084
rect 8668 13028 8672 13084
rect 8608 13024 8672 13028
rect 8688 13084 8752 13088
rect 8688 13028 8692 13084
rect 8692 13028 8748 13084
rect 8748 13028 8752 13084
rect 8688 13024 8752 13028
rect 12196 13084 12260 13088
rect 12196 13028 12200 13084
rect 12200 13028 12256 13084
rect 12256 13028 12260 13084
rect 12196 13024 12260 13028
rect 12276 13084 12340 13088
rect 12276 13028 12280 13084
rect 12280 13028 12336 13084
rect 12336 13028 12340 13084
rect 12276 13024 12340 13028
rect 12356 13084 12420 13088
rect 12356 13028 12360 13084
rect 12360 13028 12416 13084
rect 12416 13028 12420 13084
rect 12356 13024 12420 13028
rect 12436 13084 12500 13088
rect 12436 13028 12440 13084
rect 12440 13028 12496 13084
rect 12496 13028 12500 13084
rect 12436 13024 12500 13028
rect 2826 12540 2890 12544
rect 2826 12484 2830 12540
rect 2830 12484 2886 12540
rect 2886 12484 2890 12540
rect 2826 12480 2890 12484
rect 2906 12540 2970 12544
rect 2906 12484 2910 12540
rect 2910 12484 2966 12540
rect 2966 12484 2970 12540
rect 2906 12480 2970 12484
rect 2986 12540 3050 12544
rect 2986 12484 2990 12540
rect 2990 12484 3046 12540
rect 3046 12484 3050 12540
rect 2986 12480 3050 12484
rect 3066 12540 3130 12544
rect 3066 12484 3070 12540
rect 3070 12484 3126 12540
rect 3126 12484 3130 12540
rect 3066 12480 3130 12484
rect 6574 12540 6638 12544
rect 6574 12484 6578 12540
rect 6578 12484 6634 12540
rect 6634 12484 6638 12540
rect 6574 12480 6638 12484
rect 6654 12540 6718 12544
rect 6654 12484 6658 12540
rect 6658 12484 6714 12540
rect 6714 12484 6718 12540
rect 6654 12480 6718 12484
rect 6734 12540 6798 12544
rect 6734 12484 6738 12540
rect 6738 12484 6794 12540
rect 6794 12484 6798 12540
rect 6734 12480 6798 12484
rect 6814 12540 6878 12544
rect 6814 12484 6818 12540
rect 6818 12484 6874 12540
rect 6874 12484 6878 12540
rect 6814 12480 6878 12484
rect 10322 12540 10386 12544
rect 10322 12484 10326 12540
rect 10326 12484 10382 12540
rect 10382 12484 10386 12540
rect 10322 12480 10386 12484
rect 10402 12540 10466 12544
rect 10402 12484 10406 12540
rect 10406 12484 10462 12540
rect 10462 12484 10466 12540
rect 10402 12480 10466 12484
rect 10482 12540 10546 12544
rect 10482 12484 10486 12540
rect 10486 12484 10542 12540
rect 10542 12484 10546 12540
rect 10482 12480 10546 12484
rect 10562 12540 10626 12544
rect 10562 12484 10566 12540
rect 10566 12484 10622 12540
rect 10622 12484 10626 12540
rect 10562 12480 10626 12484
rect 14070 12540 14134 12544
rect 14070 12484 14074 12540
rect 14074 12484 14130 12540
rect 14130 12484 14134 12540
rect 14070 12480 14134 12484
rect 14150 12540 14214 12544
rect 14150 12484 14154 12540
rect 14154 12484 14210 12540
rect 14210 12484 14214 12540
rect 14150 12480 14214 12484
rect 14230 12540 14294 12544
rect 14230 12484 14234 12540
rect 14234 12484 14290 12540
rect 14290 12484 14294 12540
rect 14230 12480 14294 12484
rect 14310 12540 14374 12544
rect 14310 12484 14314 12540
rect 14314 12484 14370 12540
rect 14370 12484 14374 12540
rect 14310 12480 14374 12484
rect 4700 11996 4764 12000
rect 4700 11940 4704 11996
rect 4704 11940 4760 11996
rect 4760 11940 4764 11996
rect 4700 11936 4764 11940
rect 4780 11996 4844 12000
rect 4780 11940 4784 11996
rect 4784 11940 4840 11996
rect 4840 11940 4844 11996
rect 4780 11936 4844 11940
rect 4860 11996 4924 12000
rect 4860 11940 4864 11996
rect 4864 11940 4920 11996
rect 4920 11940 4924 11996
rect 4860 11936 4924 11940
rect 4940 11996 5004 12000
rect 4940 11940 4944 11996
rect 4944 11940 5000 11996
rect 5000 11940 5004 11996
rect 4940 11936 5004 11940
rect 8448 11996 8512 12000
rect 8448 11940 8452 11996
rect 8452 11940 8508 11996
rect 8508 11940 8512 11996
rect 8448 11936 8512 11940
rect 8528 11996 8592 12000
rect 8528 11940 8532 11996
rect 8532 11940 8588 11996
rect 8588 11940 8592 11996
rect 8528 11936 8592 11940
rect 8608 11996 8672 12000
rect 8608 11940 8612 11996
rect 8612 11940 8668 11996
rect 8668 11940 8672 11996
rect 8608 11936 8672 11940
rect 8688 11996 8752 12000
rect 8688 11940 8692 11996
rect 8692 11940 8748 11996
rect 8748 11940 8752 11996
rect 8688 11936 8752 11940
rect 12196 11996 12260 12000
rect 12196 11940 12200 11996
rect 12200 11940 12256 11996
rect 12256 11940 12260 11996
rect 12196 11936 12260 11940
rect 12276 11996 12340 12000
rect 12276 11940 12280 11996
rect 12280 11940 12336 11996
rect 12336 11940 12340 11996
rect 12276 11936 12340 11940
rect 12356 11996 12420 12000
rect 12356 11940 12360 11996
rect 12360 11940 12416 11996
rect 12416 11940 12420 11996
rect 12356 11936 12420 11940
rect 12436 11996 12500 12000
rect 12436 11940 12440 11996
rect 12440 11940 12496 11996
rect 12496 11940 12500 11996
rect 12436 11936 12500 11940
rect 2826 11452 2890 11456
rect 2826 11396 2830 11452
rect 2830 11396 2886 11452
rect 2886 11396 2890 11452
rect 2826 11392 2890 11396
rect 2906 11452 2970 11456
rect 2906 11396 2910 11452
rect 2910 11396 2966 11452
rect 2966 11396 2970 11452
rect 2906 11392 2970 11396
rect 2986 11452 3050 11456
rect 2986 11396 2990 11452
rect 2990 11396 3046 11452
rect 3046 11396 3050 11452
rect 2986 11392 3050 11396
rect 3066 11452 3130 11456
rect 3066 11396 3070 11452
rect 3070 11396 3126 11452
rect 3126 11396 3130 11452
rect 3066 11392 3130 11396
rect 6574 11452 6638 11456
rect 6574 11396 6578 11452
rect 6578 11396 6634 11452
rect 6634 11396 6638 11452
rect 6574 11392 6638 11396
rect 6654 11452 6718 11456
rect 6654 11396 6658 11452
rect 6658 11396 6714 11452
rect 6714 11396 6718 11452
rect 6654 11392 6718 11396
rect 6734 11452 6798 11456
rect 6734 11396 6738 11452
rect 6738 11396 6794 11452
rect 6794 11396 6798 11452
rect 6734 11392 6798 11396
rect 6814 11452 6878 11456
rect 6814 11396 6818 11452
rect 6818 11396 6874 11452
rect 6874 11396 6878 11452
rect 6814 11392 6878 11396
rect 10322 11452 10386 11456
rect 10322 11396 10326 11452
rect 10326 11396 10382 11452
rect 10382 11396 10386 11452
rect 10322 11392 10386 11396
rect 10402 11452 10466 11456
rect 10402 11396 10406 11452
rect 10406 11396 10462 11452
rect 10462 11396 10466 11452
rect 10402 11392 10466 11396
rect 10482 11452 10546 11456
rect 10482 11396 10486 11452
rect 10486 11396 10542 11452
rect 10542 11396 10546 11452
rect 10482 11392 10546 11396
rect 10562 11452 10626 11456
rect 10562 11396 10566 11452
rect 10566 11396 10622 11452
rect 10622 11396 10626 11452
rect 10562 11392 10626 11396
rect 14070 11452 14134 11456
rect 14070 11396 14074 11452
rect 14074 11396 14130 11452
rect 14130 11396 14134 11452
rect 14070 11392 14134 11396
rect 14150 11452 14214 11456
rect 14150 11396 14154 11452
rect 14154 11396 14210 11452
rect 14210 11396 14214 11452
rect 14150 11392 14214 11396
rect 14230 11452 14294 11456
rect 14230 11396 14234 11452
rect 14234 11396 14290 11452
rect 14290 11396 14294 11452
rect 14230 11392 14294 11396
rect 14310 11452 14374 11456
rect 14310 11396 14314 11452
rect 14314 11396 14370 11452
rect 14370 11396 14374 11452
rect 14310 11392 14374 11396
rect 4700 10908 4764 10912
rect 4700 10852 4704 10908
rect 4704 10852 4760 10908
rect 4760 10852 4764 10908
rect 4700 10848 4764 10852
rect 4780 10908 4844 10912
rect 4780 10852 4784 10908
rect 4784 10852 4840 10908
rect 4840 10852 4844 10908
rect 4780 10848 4844 10852
rect 4860 10908 4924 10912
rect 4860 10852 4864 10908
rect 4864 10852 4920 10908
rect 4920 10852 4924 10908
rect 4860 10848 4924 10852
rect 4940 10908 5004 10912
rect 4940 10852 4944 10908
rect 4944 10852 5000 10908
rect 5000 10852 5004 10908
rect 4940 10848 5004 10852
rect 8448 10908 8512 10912
rect 8448 10852 8452 10908
rect 8452 10852 8508 10908
rect 8508 10852 8512 10908
rect 8448 10848 8512 10852
rect 8528 10908 8592 10912
rect 8528 10852 8532 10908
rect 8532 10852 8588 10908
rect 8588 10852 8592 10908
rect 8528 10848 8592 10852
rect 8608 10908 8672 10912
rect 8608 10852 8612 10908
rect 8612 10852 8668 10908
rect 8668 10852 8672 10908
rect 8608 10848 8672 10852
rect 8688 10908 8752 10912
rect 8688 10852 8692 10908
rect 8692 10852 8748 10908
rect 8748 10852 8752 10908
rect 8688 10848 8752 10852
rect 12196 10908 12260 10912
rect 12196 10852 12200 10908
rect 12200 10852 12256 10908
rect 12256 10852 12260 10908
rect 12196 10848 12260 10852
rect 12276 10908 12340 10912
rect 12276 10852 12280 10908
rect 12280 10852 12336 10908
rect 12336 10852 12340 10908
rect 12276 10848 12340 10852
rect 12356 10908 12420 10912
rect 12356 10852 12360 10908
rect 12360 10852 12416 10908
rect 12416 10852 12420 10908
rect 12356 10848 12420 10852
rect 12436 10908 12500 10912
rect 12436 10852 12440 10908
rect 12440 10852 12496 10908
rect 12496 10852 12500 10908
rect 12436 10848 12500 10852
rect 2826 10364 2890 10368
rect 2826 10308 2830 10364
rect 2830 10308 2886 10364
rect 2886 10308 2890 10364
rect 2826 10304 2890 10308
rect 2906 10364 2970 10368
rect 2906 10308 2910 10364
rect 2910 10308 2966 10364
rect 2966 10308 2970 10364
rect 2906 10304 2970 10308
rect 2986 10364 3050 10368
rect 2986 10308 2990 10364
rect 2990 10308 3046 10364
rect 3046 10308 3050 10364
rect 2986 10304 3050 10308
rect 3066 10364 3130 10368
rect 3066 10308 3070 10364
rect 3070 10308 3126 10364
rect 3126 10308 3130 10364
rect 3066 10304 3130 10308
rect 6574 10364 6638 10368
rect 6574 10308 6578 10364
rect 6578 10308 6634 10364
rect 6634 10308 6638 10364
rect 6574 10304 6638 10308
rect 6654 10364 6718 10368
rect 6654 10308 6658 10364
rect 6658 10308 6714 10364
rect 6714 10308 6718 10364
rect 6654 10304 6718 10308
rect 6734 10364 6798 10368
rect 6734 10308 6738 10364
rect 6738 10308 6794 10364
rect 6794 10308 6798 10364
rect 6734 10304 6798 10308
rect 6814 10364 6878 10368
rect 6814 10308 6818 10364
rect 6818 10308 6874 10364
rect 6874 10308 6878 10364
rect 6814 10304 6878 10308
rect 10322 10364 10386 10368
rect 10322 10308 10326 10364
rect 10326 10308 10382 10364
rect 10382 10308 10386 10364
rect 10322 10304 10386 10308
rect 10402 10364 10466 10368
rect 10402 10308 10406 10364
rect 10406 10308 10462 10364
rect 10462 10308 10466 10364
rect 10402 10304 10466 10308
rect 10482 10364 10546 10368
rect 10482 10308 10486 10364
rect 10486 10308 10542 10364
rect 10542 10308 10546 10364
rect 10482 10304 10546 10308
rect 10562 10364 10626 10368
rect 10562 10308 10566 10364
rect 10566 10308 10622 10364
rect 10622 10308 10626 10364
rect 10562 10304 10626 10308
rect 14070 10364 14134 10368
rect 14070 10308 14074 10364
rect 14074 10308 14130 10364
rect 14130 10308 14134 10364
rect 14070 10304 14134 10308
rect 14150 10364 14214 10368
rect 14150 10308 14154 10364
rect 14154 10308 14210 10364
rect 14210 10308 14214 10364
rect 14150 10304 14214 10308
rect 14230 10364 14294 10368
rect 14230 10308 14234 10364
rect 14234 10308 14290 10364
rect 14290 10308 14294 10364
rect 14230 10304 14294 10308
rect 14310 10364 14374 10368
rect 14310 10308 14314 10364
rect 14314 10308 14370 10364
rect 14370 10308 14374 10364
rect 14310 10304 14374 10308
rect 4700 9820 4764 9824
rect 4700 9764 4704 9820
rect 4704 9764 4760 9820
rect 4760 9764 4764 9820
rect 4700 9760 4764 9764
rect 4780 9820 4844 9824
rect 4780 9764 4784 9820
rect 4784 9764 4840 9820
rect 4840 9764 4844 9820
rect 4780 9760 4844 9764
rect 4860 9820 4924 9824
rect 4860 9764 4864 9820
rect 4864 9764 4920 9820
rect 4920 9764 4924 9820
rect 4860 9760 4924 9764
rect 4940 9820 5004 9824
rect 4940 9764 4944 9820
rect 4944 9764 5000 9820
rect 5000 9764 5004 9820
rect 4940 9760 5004 9764
rect 8448 9820 8512 9824
rect 8448 9764 8452 9820
rect 8452 9764 8508 9820
rect 8508 9764 8512 9820
rect 8448 9760 8512 9764
rect 8528 9820 8592 9824
rect 8528 9764 8532 9820
rect 8532 9764 8588 9820
rect 8588 9764 8592 9820
rect 8528 9760 8592 9764
rect 8608 9820 8672 9824
rect 8608 9764 8612 9820
rect 8612 9764 8668 9820
rect 8668 9764 8672 9820
rect 8608 9760 8672 9764
rect 8688 9820 8752 9824
rect 8688 9764 8692 9820
rect 8692 9764 8748 9820
rect 8748 9764 8752 9820
rect 8688 9760 8752 9764
rect 12196 9820 12260 9824
rect 12196 9764 12200 9820
rect 12200 9764 12256 9820
rect 12256 9764 12260 9820
rect 12196 9760 12260 9764
rect 12276 9820 12340 9824
rect 12276 9764 12280 9820
rect 12280 9764 12336 9820
rect 12336 9764 12340 9820
rect 12276 9760 12340 9764
rect 12356 9820 12420 9824
rect 12356 9764 12360 9820
rect 12360 9764 12416 9820
rect 12416 9764 12420 9820
rect 12356 9760 12420 9764
rect 12436 9820 12500 9824
rect 12436 9764 12440 9820
rect 12440 9764 12496 9820
rect 12496 9764 12500 9820
rect 12436 9760 12500 9764
rect 5764 9752 5828 9756
rect 5764 9696 5778 9752
rect 5778 9696 5828 9752
rect 5764 9692 5828 9696
rect 9260 9692 9324 9756
rect 2826 9276 2890 9280
rect 2826 9220 2830 9276
rect 2830 9220 2886 9276
rect 2886 9220 2890 9276
rect 2826 9216 2890 9220
rect 2906 9276 2970 9280
rect 2906 9220 2910 9276
rect 2910 9220 2966 9276
rect 2966 9220 2970 9276
rect 2906 9216 2970 9220
rect 2986 9276 3050 9280
rect 2986 9220 2990 9276
rect 2990 9220 3046 9276
rect 3046 9220 3050 9276
rect 2986 9216 3050 9220
rect 3066 9276 3130 9280
rect 3066 9220 3070 9276
rect 3070 9220 3126 9276
rect 3126 9220 3130 9276
rect 3066 9216 3130 9220
rect 6574 9276 6638 9280
rect 6574 9220 6578 9276
rect 6578 9220 6634 9276
rect 6634 9220 6638 9276
rect 6574 9216 6638 9220
rect 6654 9276 6718 9280
rect 6654 9220 6658 9276
rect 6658 9220 6714 9276
rect 6714 9220 6718 9276
rect 6654 9216 6718 9220
rect 6734 9276 6798 9280
rect 6734 9220 6738 9276
rect 6738 9220 6794 9276
rect 6794 9220 6798 9276
rect 6734 9216 6798 9220
rect 6814 9276 6878 9280
rect 6814 9220 6818 9276
rect 6818 9220 6874 9276
rect 6874 9220 6878 9276
rect 6814 9216 6878 9220
rect 10322 9276 10386 9280
rect 10322 9220 10326 9276
rect 10326 9220 10382 9276
rect 10382 9220 10386 9276
rect 10322 9216 10386 9220
rect 10402 9276 10466 9280
rect 10402 9220 10406 9276
rect 10406 9220 10462 9276
rect 10462 9220 10466 9276
rect 10402 9216 10466 9220
rect 10482 9276 10546 9280
rect 10482 9220 10486 9276
rect 10486 9220 10542 9276
rect 10542 9220 10546 9276
rect 10482 9216 10546 9220
rect 10562 9276 10626 9280
rect 10562 9220 10566 9276
rect 10566 9220 10622 9276
rect 10622 9220 10626 9276
rect 10562 9216 10626 9220
rect 14070 9276 14134 9280
rect 14070 9220 14074 9276
rect 14074 9220 14130 9276
rect 14130 9220 14134 9276
rect 14070 9216 14134 9220
rect 14150 9276 14214 9280
rect 14150 9220 14154 9276
rect 14154 9220 14210 9276
rect 14210 9220 14214 9276
rect 14150 9216 14214 9220
rect 14230 9276 14294 9280
rect 14230 9220 14234 9276
rect 14234 9220 14290 9276
rect 14290 9220 14294 9276
rect 14230 9216 14294 9220
rect 14310 9276 14374 9280
rect 14310 9220 14314 9276
rect 14314 9220 14370 9276
rect 14370 9220 14374 9276
rect 14310 9216 14374 9220
rect 4700 8732 4764 8736
rect 4700 8676 4704 8732
rect 4704 8676 4760 8732
rect 4760 8676 4764 8732
rect 4700 8672 4764 8676
rect 4780 8732 4844 8736
rect 4780 8676 4784 8732
rect 4784 8676 4840 8732
rect 4840 8676 4844 8732
rect 4780 8672 4844 8676
rect 4860 8732 4924 8736
rect 4860 8676 4864 8732
rect 4864 8676 4920 8732
rect 4920 8676 4924 8732
rect 4860 8672 4924 8676
rect 4940 8732 5004 8736
rect 4940 8676 4944 8732
rect 4944 8676 5000 8732
rect 5000 8676 5004 8732
rect 4940 8672 5004 8676
rect 8448 8732 8512 8736
rect 8448 8676 8452 8732
rect 8452 8676 8508 8732
rect 8508 8676 8512 8732
rect 8448 8672 8512 8676
rect 8528 8732 8592 8736
rect 8528 8676 8532 8732
rect 8532 8676 8588 8732
rect 8588 8676 8592 8732
rect 8528 8672 8592 8676
rect 8608 8732 8672 8736
rect 8608 8676 8612 8732
rect 8612 8676 8668 8732
rect 8668 8676 8672 8732
rect 8608 8672 8672 8676
rect 8688 8732 8752 8736
rect 8688 8676 8692 8732
rect 8692 8676 8748 8732
rect 8748 8676 8752 8732
rect 8688 8672 8752 8676
rect 12196 8732 12260 8736
rect 12196 8676 12200 8732
rect 12200 8676 12256 8732
rect 12256 8676 12260 8732
rect 12196 8672 12260 8676
rect 12276 8732 12340 8736
rect 12276 8676 12280 8732
rect 12280 8676 12336 8732
rect 12336 8676 12340 8732
rect 12276 8672 12340 8676
rect 12356 8732 12420 8736
rect 12356 8676 12360 8732
rect 12360 8676 12416 8732
rect 12416 8676 12420 8732
rect 12356 8672 12420 8676
rect 12436 8732 12500 8736
rect 12436 8676 12440 8732
rect 12440 8676 12496 8732
rect 12496 8676 12500 8732
rect 12436 8672 12500 8676
rect 2826 8188 2890 8192
rect 2826 8132 2830 8188
rect 2830 8132 2886 8188
rect 2886 8132 2890 8188
rect 2826 8128 2890 8132
rect 2906 8188 2970 8192
rect 2906 8132 2910 8188
rect 2910 8132 2966 8188
rect 2966 8132 2970 8188
rect 2906 8128 2970 8132
rect 2986 8188 3050 8192
rect 2986 8132 2990 8188
rect 2990 8132 3046 8188
rect 3046 8132 3050 8188
rect 2986 8128 3050 8132
rect 3066 8188 3130 8192
rect 3066 8132 3070 8188
rect 3070 8132 3126 8188
rect 3126 8132 3130 8188
rect 3066 8128 3130 8132
rect 6574 8188 6638 8192
rect 6574 8132 6578 8188
rect 6578 8132 6634 8188
rect 6634 8132 6638 8188
rect 6574 8128 6638 8132
rect 6654 8188 6718 8192
rect 6654 8132 6658 8188
rect 6658 8132 6714 8188
rect 6714 8132 6718 8188
rect 6654 8128 6718 8132
rect 6734 8188 6798 8192
rect 6734 8132 6738 8188
rect 6738 8132 6794 8188
rect 6794 8132 6798 8188
rect 6734 8128 6798 8132
rect 6814 8188 6878 8192
rect 6814 8132 6818 8188
rect 6818 8132 6874 8188
rect 6874 8132 6878 8188
rect 6814 8128 6878 8132
rect 10322 8188 10386 8192
rect 10322 8132 10326 8188
rect 10326 8132 10382 8188
rect 10382 8132 10386 8188
rect 10322 8128 10386 8132
rect 10402 8188 10466 8192
rect 10402 8132 10406 8188
rect 10406 8132 10462 8188
rect 10462 8132 10466 8188
rect 10402 8128 10466 8132
rect 10482 8188 10546 8192
rect 10482 8132 10486 8188
rect 10486 8132 10542 8188
rect 10542 8132 10546 8188
rect 10482 8128 10546 8132
rect 10562 8188 10626 8192
rect 10562 8132 10566 8188
rect 10566 8132 10622 8188
rect 10622 8132 10626 8188
rect 10562 8128 10626 8132
rect 14070 8188 14134 8192
rect 14070 8132 14074 8188
rect 14074 8132 14130 8188
rect 14130 8132 14134 8188
rect 14070 8128 14134 8132
rect 14150 8188 14214 8192
rect 14150 8132 14154 8188
rect 14154 8132 14210 8188
rect 14210 8132 14214 8188
rect 14150 8128 14214 8132
rect 14230 8188 14294 8192
rect 14230 8132 14234 8188
rect 14234 8132 14290 8188
rect 14290 8132 14294 8188
rect 14230 8128 14294 8132
rect 14310 8188 14374 8192
rect 14310 8132 14314 8188
rect 14314 8132 14370 8188
rect 14370 8132 14374 8188
rect 14310 8128 14374 8132
rect 4700 7644 4764 7648
rect 4700 7588 4704 7644
rect 4704 7588 4760 7644
rect 4760 7588 4764 7644
rect 4700 7584 4764 7588
rect 4780 7644 4844 7648
rect 4780 7588 4784 7644
rect 4784 7588 4840 7644
rect 4840 7588 4844 7644
rect 4780 7584 4844 7588
rect 4860 7644 4924 7648
rect 4860 7588 4864 7644
rect 4864 7588 4920 7644
rect 4920 7588 4924 7644
rect 4860 7584 4924 7588
rect 4940 7644 5004 7648
rect 4940 7588 4944 7644
rect 4944 7588 5000 7644
rect 5000 7588 5004 7644
rect 4940 7584 5004 7588
rect 8448 7644 8512 7648
rect 8448 7588 8452 7644
rect 8452 7588 8508 7644
rect 8508 7588 8512 7644
rect 8448 7584 8512 7588
rect 8528 7644 8592 7648
rect 8528 7588 8532 7644
rect 8532 7588 8588 7644
rect 8588 7588 8592 7644
rect 8528 7584 8592 7588
rect 8608 7644 8672 7648
rect 8608 7588 8612 7644
rect 8612 7588 8668 7644
rect 8668 7588 8672 7644
rect 8608 7584 8672 7588
rect 8688 7644 8752 7648
rect 8688 7588 8692 7644
rect 8692 7588 8748 7644
rect 8748 7588 8752 7644
rect 8688 7584 8752 7588
rect 12196 7644 12260 7648
rect 12196 7588 12200 7644
rect 12200 7588 12256 7644
rect 12256 7588 12260 7644
rect 12196 7584 12260 7588
rect 12276 7644 12340 7648
rect 12276 7588 12280 7644
rect 12280 7588 12336 7644
rect 12336 7588 12340 7644
rect 12276 7584 12340 7588
rect 12356 7644 12420 7648
rect 12356 7588 12360 7644
rect 12360 7588 12416 7644
rect 12416 7588 12420 7644
rect 12356 7584 12420 7588
rect 12436 7644 12500 7648
rect 12436 7588 12440 7644
rect 12440 7588 12496 7644
rect 12496 7588 12500 7644
rect 12436 7584 12500 7588
rect 2826 7100 2890 7104
rect 2826 7044 2830 7100
rect 2830 7044 2886 7100
rect 2886 7044 2890 7100
rect 2826 7040 2890 7044
rect 2906 7100 2970 7104
rect 2906 7044 2910 7100
rect 2910 7044 2966 7100
rect 2966 7044 2970 7100
rect 2906 7040 2970 7044
rect 2986 7100 3050 7104
rect 2986 7044 2990 7100
rect 2990 7044 3046 7100
rect 3046 7044 3050 7100
rect 2986 7040 3050 7044
rect 3066 7100 3130 7104
rect 3066 7044 3070 7100
rect 3070 7044 3126 7100
rect 3126 7044 3130 7100
rect 3066 7040 3130 7044
rect 6574 7100 6638 7104
rect 6574 7044 6578 7100
rect 6578 7044 6634 7100
rect 6634 7044 6638 7100
rect 6574 7040 6638 7044
rect 6654 7100 6718 7104
rect 6654 7044 6658 7100
rect 6658 7044 6714 7100
rect 6714 7044 6718 7100
rect 6654 7040 6718 7044
rect 6734 7100 6798 7104
rect 6734 7044 6738 7100
rect 6738 7044 6794 7100
rect 6794 7044 6798 7100
rect 6734 7040 6798 7044
rect 6814 7100 6878 7104
rect 6814 7044 6818 7100
rect 6818 7044 6874 7100
rect 6874 7044 6878 7100
rect 6814 7040 6878 7044
rect 10322 7100 10386 7104
rect 10322 7044 10326 7100
rect 10326 7044 10382 7100
rect 10382 7044 10386 7100
rect 10322 7040 10386 7044
rect 10402 7100 10466 7104
rect 10402 7044 10406 7100
rect 10406 7044 10462 7100
rect 10462 7044 10466 7100
rect 10402 7040 10466 7044
rect 10482 7100 10546 7104
rect 10482 7044 10486 7100
rect 10486 7044 10542 7100
rect 10542 7044 10546 7100
rect 10482 7040 10546 7044
rect 10562 7100 10626 7104
rect 10562 7044 10566 7100
rect 10566 7044 10622 7100
rect 10622 7044 10626 7100
rect 10562 7040 10626 7044
rect 14070 7100 14134 7104
rect 14070 7044 14074 7100
rect 14074 7044 14130 7100
rect 14130 7044 14134 7100
rect 14070 7040 14134 7044
rect 14150 7100 14214 7104
rect 14150 7044 14154 7100
rect 14154 7044 14210 7100
rect 14210 7044 14214 7100
rect 14150 7040 14214 7044
rect 14230 7100 14294 7104
rect 14230 7044 14234 7100
rect 14234 7044 14290 7100
rect 14290 7044 14294 7100
rect 14230 7040 14294 7044
rect 14310 7100 14374 7104
rect 14310 7044 14314 7100
rect 14314 7044 14370 7100
rect 14370 7044 14374 7100
rect 14310 7040 14374 7044
rect 4700 6556 4764 6560
rect 4700 6500 4704 6556
rect 4704 6500 4760 6556
rect 4760 6500 4764 6556
rect 4700 6496 4764 6500
rect 4780 6556 4844 6560
rect 4780 6500 4784 6556
rect 4784 6500 4840 6556
rect 4840 6500 4844 6556
rect 4780 6496 4844 6500
rect 4860 6556 4924 6560
rect 4860 6500 4864 6556
rect 4864 6500 4920 6556
rect 4920 6500 4924 6556
rect 4860 6496 4924 6500
rect 4940 6556 5004 6560
rect 4940 6500 4944 6556
rect 4944 6500 5000 6556
rect 5000 6500 5004 6556
rect 4940 6496 5004 6500
rect 8448 6556 8512 6560
rect 8448 6500 8452 6556
rect 8452 6500 8508 6556
rect 8508 6500 8512 6556
rect 8448 6496 8512 6500
rect 8528 6556 8592 6560
rect 8528 6500 8532 6556
rect 8532 6500 8588 6556
rect 8588 6500 8592 6556
rect 8528 6496 8592 6500
rect 8608 6556 8672 6560
rect 8608 6500 8612 6556
rect 8612 6500 8668 6556
rect 8668 6500 8672 6556
rect 8608 6496 8672 6500
rect 8688 6556 8752 6560
rect 8688 6500 8692 6556
rect 8692 6500 8748 6556
rect 8748 6500 8752 6556
rect 8688 6496 8752 6500
rect 12196 6556 12260 6560
rect 12196 6500 12200 6556
rect 12200 6500 12256 6556
rect 12256 6500 12260 6556
rect 12196 6496 12260 6500
rect 12276 6556 12340 6560
rect 12276 6500 12280 6556
rect 12280 6500 12336 6556
rect 12336 6500 12340 6556
rect 12276 6496 12340 6500
rect 12356 6556 12420 6560
rect 12356 6500 12360 6556
rect 12360 6500 12416 6556
rect 12416 6500 12420 6556
rect 12356 6496 12420 6500
rect 12436 6556 12500 6560
rect 12436 6500 12440 6556
rect 12440 6500 12496 6556
rect 12496 6500 12500 6556
rect 12436 6496 12500 6500
rect 2826 6012 2890 6016
rect 2826 5956 2830 6012
rect 2830 5956 2886 6012
rect 2886 5956 2890 6012
rect 2826 5952 2890 5956
rect 2906 6012 2970 6016
rect 2906 5956 2910 6012
rect 2910 5956 2966 6012
rect 2966 5956 2970 6012
rect 2906 5952 2970 5956
rect 2986 6012 3050 6016
rect 2986 5956 2990 6012
rect 2990 5956 3046 6012
rect 3046 5956 3050 6012
rect 2986 5952 3050 5956
rect 3066 6012 3130 6016
rect 3066 5956 3070 6012
rect 3070 5956 3126 6012
rect 3126 5956 3130 6012
rect 3066 5952 3130 5956
rect 6574 6012 6638 6016
rect 6574 5956 6578 6012
rect 6578 5956 6634 6012
rect 6634 5956 6638 6012
rect 6574 5952 6638 5956
rect 6654 6012 6718 6016
rect 6654 5956 6658 6012
rect 6658 5956 6714 6012
rect 6714 5956 6718 6012
rect 6654 5952 6718 5956
rect 6734 6012 6798 6016
rect 6734 5956 6738 6012
rect 6738 5956 6794 6012
rect 6794 5956 6798 6012
rect 6734 5952 6798 5956
rect 6814 6012 6878 6016
rect 6814 5956 6818 6012
rect 6818 5956 6874 6012
rect 6874 5956 6878 6012
rect 6814 5952 6878 5956
rect 10322 6012 10386 6016
rect 10322 5956 10326 6012
rect 10326 5956 10382 6012
rect 10382 5956 10386 6012
rect 10322 5952 10386 5956
rect 10402 6012 10466 6016
rect 10402 5956 10406 6012
rect 10406 5956 10462 6012
rect 10462 5956 10466 6012
rect 10402 5952 10466 5956
rect 10482 6012 10546 6016
rect 10482 5956 10486 6012
rect 10486 5956 10542 6012
rect 10542 5956 10546 6012
rect 10482 5952 10546 5956
rect 10562 6012 10626 6016
rect 10562 5956 10566 6012
rect 10566 5956 10622 6012
rect 10622 5956 10626 6012
rect 10562 5952 10626 5956
rect 14070 6012 14134 6016
rect 14070 5956 14074 6012
rect 14074 5956 14130 6012
rect 14130 5956 14134 6012
rect 14070 5952 14134 5956
rect 14150 6012 14214 6016
rect 14150 5956 14154 6012
rect 14154 5956 14210 6012
rect 14210 5956 14214 6012
rect 14150 5952 14214 5956
rect 14230 6012 14294 6016
rect 14230 5956 14234 6012
rect 14234 5956 14290 6012
rect 14290 5956 14294 6012
rect 14230 5952 14294 5956
rect 14310 6012 14374 6016
rect 14310 5956 14314 6012
rect 14314 5956 14370 6012
rect 14370 5956 14374 6012
rect 14310 5952 14374 5956
rect 4700 5468 4764 5472
rect 4700 5412 4704 5468
rect 4704 5412 4760 5468
rect 4760 5412 4764 5468
rect 4700 5408 4764 5412
rect 4780 5468 4844 5472
rect 4780 5412 4784 5468
rect 4784 5412 4840 5468
rect 4840 5412 4844 5468
rect 4780 5408 4844 5412
rect 4860 5468 4924 5472
rect 4860 5412 4864 5468
rect 4864 5412 4920 5468
rect 4920 5412 4924 5468
rect 4860 5408 4924 5412
rect 4940 5468 5004 5472
rect 4940 5412 4944 5468
rect 4944 5412 5000 5468
rect 5000 5412 5004 5468
rect 4940 5408 5004 5412
rect 8448 5468 8512 5472
rect 8448 5412 8452 5468
rect 8452 5412 8508 5468
rect 8508 5412 8512 5468
rect 8448 5408 8512 5412
rect 8528 5468 8592 5472
rect 8528 5412 8532 5468
rect 8532 5412 8588 5468
rect 8588 5412 8592 5468
rect 8528 5408 8592 5412
rect 8608 5468 8672 5472
rect 8608 5412 8612 5468
rect 8612 5412 8668 5468
rect 8668 5412 8672 5468
rect 8608 5408 8672 5412
rect 8688 5468 8752 5472
rect 8688 5412 8692 5468
rect 8692 5412 8748 5468
rect 8748 5412 8752 5468
rect 8688 5408 8752 5412
rect 12196 5468 12260 5472
rect 12196 5412 12200 5468
rect 12200 5412 12256 5468
rect 12256 5412 12260 5468
rect 12196 5408 12260 5412
rect 12276 5468 12340 5472
rect 12276 5412 12280 5468
rect 12280 5412 12336 5468
rect 12336 5412 12340 5468
rect 12276 5408 12340 5412
rect 12356 5468 12420 5472
rect 12356 5412 12360 5468
rect 12360 5412 12416 5468
rect 12416 5412 12420 5468
rect 12356 5408 12420 5412
rect 12436 5468 12500 5472
rect 12436 5412 12440 5468
rect 12440 5412 12496 5468
rect 12496 5412 12500 5468
rect 12436 5408 12500 5412
rect 2826 4924 2890 4928
rect 2826 4868 2830 4924
rect 2830 4868 2886 4924
rect 2886 4868 2890 4924
rect 2826 4864 2890 4868
rect 2906 4924 2970 4928
rect 2906 4868 2910 4924
rect 2910 4868 2966 4924
rect 2966 4868 2970 4924
rect 2906 4864 2970 4868
rect 2986 4924 3050 4928
rect 2986 4868 2990 4924
rect 2990 4868 3046 4924
rect 3046 4868 3050 4924
rect 2986 4864 3050 4868
rect 3066 4924 3130 4928
rect 3066 4868 3070 4924
rect 3070 4868 3126 4924
rect 3126 4868 3130 4924
rect 3066 4864 3130 4868
rect 6574 4924 6638 4928
rect 6574 4868 6578 4924
rect 6578 4868 6634 4924
rect 6634 4868 6638 4924
rect 6574 4864 6638 4868
rect 6654 4924 6718 4928
rect 6654 4868 6658 4924
rect 6658 4868 6714 4924
rect 6714 4868 6718 4924
rect 6654 4864 6718 4868
rect 6734 4924 6798 4928
rect 6734 4868 6738 4924
rect 6738 4868 6794 4924
rect 6794 4868 6798 4924
rect 6734 4864 6798 4868
rect 6814 4924 6878 4928
rect 6814 4868 6818 4924
rect 6818 4868 6874 4924
rect 6874 4868 6878 4924
rect 6814 4864 6878 4868
rect 10322 4924 10386 4928
rect 10322 4868 10326 4924
rect 10326 4868 10382 4924
rect 10382 4868 10386 4924
rect 10322 4864 10386 4868
rect 10402 4924 10466 4928
rect 10402 4868 10406 4924
rect 10406 4868 10462 4924
rect 10462 4868 10466 4924
rect 10402 4864 10466 4868
rect 10482 4924 10546 4928
rect 10482 4868 10486 4924
rect 10486 4868 10542 4924
rect 10542 4868 10546 4924
rect 10482 4864 10546 4868
rect 10562 4924 10626 4928
rect 10562 4868 10566 4924
rect 10566 4868 10622 4924
rect 10622 4868 10626 4924
rect 10562 4864 10626 4868
rect 14070 4924 14134 4928
rect 14070 4868 14074 4924
rect 14074 4868 14130 4924
rect 14130 4868 14134 4924
rect 14070 4864 14134 4868
rect 14150 4924 14214 4928
rect 14150 4868 14154 4924
rect 14154 4868 14210 4924
rect 14210 4868 14214 4924
rect 14150 4864 14214 4868
rect 14230 4924 14294 4928
rect 14230 4868 14234 4924
rect 14234 4868 14290 4924
rect 14290 4868 14294 4924
rect 14230 4864 14294 4868
rect 14310 4924 14374 4928
rect 14310 4868 14314 4924
rect 14314 4868 14370 4924
rect 14370 4868 14374 4924
rect 14310 4864 14374 4868
rect 4700 4380 4764 4384
rect 4700 4324 4704 4380
rect 4704 4324 4760 4380
rect 4760 4324 4764 4380
rect 4700 4320 4764 4324
rect 4780 4380 4844 4384
rect 4780 4324 4784 4380
rect 4784 4324 4840 4380
rect 4840 4324 4844 4380
rect 4780 4320 4844 4324
rect 4860 4380 4924 4384
rect 4860 4324 4864 4380
rect 4864 4324 4920 4380
rect 4920 4324 4924 4380
rect 4860 4320 4924 4324
rect 4940 4380 5004 4384
rect 4940 4324 4944 4380
rect 4944 4324 5000 4380
rect 5000 4324 5004 4380
rect 4940 4320 5004 4324
rect 8448 4380 8512 4384
rect 8448 4324 8452 4380
rect 8452 4324 8508 4380
rect 8508 4324 8512 4380
rect 8448 4320 8512 4324
rect 8528 4380 8592 4384
rect 8528 4324 8532 4380
rect 8532 4324 8588 4380
rect 8588 4324 8592 4380
rect 8528 4320 8592 4324
rect 8608 4380 8672 4384
rect 8608 4324 8612 4380
rect 8612 4324 8668 4380
rect 8668 4324 8672 4380
rect 8608 4320 8672 4324
rect 8688 4380 8752 4384
rect 8688 4324 8692 4380
rect 8692 4324 8748 4380
rect 8748 4324 8752 4380
rect 8688 4320 8752 4324
rect 12196 4380 12260 4384
rect 12196 4324 12200 4380
rect 12200 4324 12256 4380
rect 12256 4324 12260 4380
rect 12196 4320 12260 4324
rect 12276 4380 12340 4384
rect 12276 4324 12280 4380
rect 12280 4324 12336 4380
rect 12336 4324 12340 4380
rect 12276 4320 12340 4324
rect 12356 4380 12420 4384
rect 12356 4324 12360 4380
rect 12360 4324 12416 4380
rect 12416 4324 12420 4380
rect 12356 4320 12420 4324
rect 12436 4380 12500 4384
rect 12436 4324 12440 4380
rect 12440 4324 12496 4380
rect 12496 4324 12500 4380
rect 12436 4320 12500 4324
rect 2826 3836 2890 3840
rect 2826 3780 2830 3836
rect 2830 3780 2886 3836
rect 2886 3780 2890 3836
rect 2826 3776 2890 3780
rect 2906 3836 2970 3840
rect 2906 3780 2910 3836
rect 2910 3780 2966 3836
rect 2966 3780 2970 3836
rect 2906 3776 2970 3780
rect 2986 3836 3050 3840
rect 2986 3780 2990 3836
rect 2990 3780 3046 3836
rect 3046 3780 3050 3836
rect 2986 3776 3050 3780
rect 3066 3836 3130 3840
rect 3066 3780 3070 3836
rect 3070 3780 3126 3836
rect 3126 3780 3130 3836
rect 3066 3776 3130 3780
rect 6574 3836 6638 3840
rect 6574 3780 6578 3836
rect 6578 3780 6634 3836
rect 6634 3780 6638 3836
rect 6574 3776 6638 3780
rect 6654 3836 6718 3840
rect 6654 3780 6658 3836
rect 6658 3780 6714 3836
rect 6714 3780 6718 3836
rect 6654 3776 6718 3780
rect 6734 3836 6798 3840
rect 6734 3780 6738 3836
rect 6738 3780 6794 3836
rect 6794 3780 6798 3836
rect 6734 3776 6798 3780
rect 6814 3836 6878 3840
rect 6814 3780 6818 3836
rect 6818 3780 6874 3836
rect 6874 3780 6878 3836
rect 6814 3776 6878 3780
rect 10322 3836 10386 3840
rect 10322 3780 10326 3836
rect 10326 3780 10382 3836
rect 10382 3780 10386 3836
rect 10322 3776 10386 3780
rect 10402 3836 10466 3840
rect 10402 3780 10406 3836
rect 10406 3780 10462 3836
rect 10462 3780 10466 3836
rect 10402 3776 10466 3780
rect 10482 3836 10546 3840
rect 10482 3780 10486 3836
rect 10486 3780 10542 3836
rect 10542 3780 10546 3836
rect 10482 3776 10546 3780
rect 10562 3836 10626 3840
rect 10562 3780 10566 3836
rect 10566 3780 10622 3836
rect 10622 3780 10626 3836
rect 10562 3776 10626 3780
rect 14070 3836 14134 3840
rect 14070 3780 14074 3836
rect 14074 3780 14130 3836
rect 14130 3780 14134 3836
rect 14070 3776 14134 3780
rect 14150 3836 14214 3840
rect 14150 3780 14154 3836
rect 14154 3780 14210 3836
rect 14210 3780 14214 3836
rect 14150 3776 14214 3780
rect 14230 3836 14294 3840
rect 14230 3780 14234 3836
rect 14234 3780 14290 3836
rect 14290 3780 14294 3836
rect 14230 3776 14294 3780
rect 14310 3836 14374 3840
rect 14310 3780 14314 3836
rect 14314 3780 14370 3836
rect 14370 3780 14374 3836
rect 14310 3776 14374 3780
rect 4700 3292 4764 3296
rect 4700 3236 4704 3292
rect 4704 3236 4760 3292
rect 4760 3236 4764 3292
rect 4700 3232 4764 3236
rect 4780 3292 4844 3296
rect 4780 3236 4784 3292
rect 4784 3236 4840 3292
rect 4840 3236 4844 3292
rect 4780 3232 4844 3236
rect 4860 3292 4924 3296
rect 4860 3236 4864 3292
rect 4864 3236 4920 3292
rect 4920 3236 4924 3292
rect 4860 3232 4924 3236
rect 4940 3292 5004 3296
rect 4940 3236 4944 3292
rect 4944 3236 5000 3292
rect 5000 3236 5004 3292
rect 4940 3232 5004 3236
rect 8448 3292 8512 3296
rect 8448 3236 8452 3292
rect 8452 3236 8508 3292
rect 8508 3236 8512 3292
rect 8448 3232 8512 3236
rect 8528 3292 8592 3296
rect 8528 3236 8532 3292
rect 8532 3236 8588 3292
rect 8588 3236 8592 3292
rect 8528 3232 8592 3236
rect 8608 3292 8672 3296
rect 8608 3236 8612 3292
rect 8612 3236 8668 3292
rect 8668 3236 8672 3292
rect 8608 3232 8672 3236
rect 8688 3292 8752 3296
rect 8688 3236 8692 3292
rect 8692 3236 8748 3292
rect 8748 3236 8752 3292
rect 8688 3232 8752 3236
rect 12196 3292 12260 3296
rect 12196 3236 12200 3292
rect 12200 3236 12256 3292
rect 12256 3236 12260 3292
rect 12196 3232 12260 3236
rect 12276 3292 12340 3296
rect 12276 3236 12280 3292
rect 12280 3236 12336 3292
rect 12336 3236 12340 3292
rect 12276 3232 12340 3236
rect 12356 3292 12420 3296
rect 12356 3236 12360 3292
rect 12360 3236 12416 3292
rect 12416 3236 12420 3292
rect 12356 3232 12420 3236
rect 12436 3292 12500 3296
rect 12436 3236 12440 3292
rect 12440 3236 12496 3292
rect 12496 3236 12500 3292
rect 12436 3232 12500 3236
rect 2826 2748 2890 2752
rect 2826 2692 2830 2748
rect 2830 2692 2886 2748
rect 2886 2692 2890 2748
rect 2826 2688 2890 2692
rect 2906 2748 2970 2752
rect 2906 2692 2910 2748
rect 2910 2692 2966 2748
rect 2966 2692 2970 2748
rect 2906 2688 2970 2692
rect 2986 2748 3050 2752
rect 2986 2692 2990 2748
rect 2990 2692 3046 2748
rect 3046 2692 3050 2748
rect 2986 2688 3050 2692
rect 3066 2748 3130 2752
rect 3066 2692 3070 2748
rect 3070 2692 3126 2748
rect 3126 2692 3130 2748
rect 3066 2688 3130 2692
rect 6574 2748 6638 2752
rect 6574 2692 6578 2748
rect 6578 2692 6634 2748
rect 6634 2692 6638 2748
rect 6574 2688 6638 2692
rect 6654 2748 6718 2752
rect 6654 2692 6658 2748
rect 6658 2692 6714 2748
rect 6714 2692 6718 2748
rect 6654 2688 6718 2692
rect 6734 2748 6798 2752
rect 6734 2692 6738 2748
rect 6738 2692 6794 2748
rect 6794 2692 6798 2748
rect 6734 2688 6798 2692
rect 6814 2748 6878 2752
rect 6814 2692 6818 2748
rect 6818 2692 6874 2748
rect 6874 2692 6878 2748
rect 6814 2688 6878 2692
rect 10322 2748 10386 2752
rect 10322 2692 10326 2748
rect 10326 2692 10382 2748
rect 10382 2692 10386 2748
rect 10322 2688 10386 2692
rect 10402 2748 10466 2752
rect 10402 2692 10406 2748
rect 10406 2692 10462 2748
rect 10462 2692 10466 2748
rect 10402 2688 10466 2692
rect 10482 2748 10546 2752
rect 10482 2692 10486 2748
rect 10486 2692 10542 2748
rect 10542 2692 10546 2748
rect 10482 2688 10546 2692
rect 10562 2748 10626 2752
rect 10562 2692 10566 2748
rect 10566 2692 10622 2748
rect 10622 2692 10626 2748
rect 10562 2688 10626 2692
rect 14070 2748 14134 2752
rect 14070 2692 14074 2748
rect 14074 2692 14130 2748
rect 14130 2692 14134 2748
rect 14070 2688 14134 2692
rect 14150 2748 14214 2752
rect 14150 2692 14154 2748
rect 14154 2692 14210 2748
rect 14210 2692 14214 2748
rect 14150 2688 14214 2692
rect 14230 2748 14294 2752
rect 14230 2692 14234 2748
rect 14234 2692 14290 2748
rect 14290 2692 14294 2748
rect 14230 2688 14294 2692
rect 14310 2748 14374 2752
rect 14310 2692 14314 2748
rect 14314 2692 14370 2748
rect 14370 2692 14374 2748
rect 14310 2688 14374 2692
rect 5764 2484 5828 2548
rect 4700 2204 4764 2208
rect 4700 2148 4704 2204
rect 4704 2148 4760 2204
rect 4760 2148 4764 2204
rect 4700 2144 4764 2148
rect 4780 2204 4844 2208
rect 4780 2148 4784 2204
rect 4784 2148 4840 2204
rect 4840 2148 4844 2204
rect 4780 2144 4844 2148
rect 4860 2204 4924 2208
rect 4860 2148 4864 2204
rect 4864 2148 4920 2204
rect 4920 2148 4924 2204
rect 4860 2144 4924 2148
rect 4940 2204 5004 2208
rect 4940 2148 4944 2204
rect 4944 2148 5000 2204
rect 5000 2148 5004 2204
rect 4940 2144 5004 2148
rect 8448 2204 8512 2208
rect 8448 2148 8452 2204
rect 8452 2148 8508 2204
rect 8508 2148 8512 2204
rect 8448 2144 8512 2148
rect 8528 2204 8592 2208
rect 8528 2148 8532 2204
rect 8532 2148 8588 2204
rect 8588 2148 8592 2204
rect 8528 2144 8592 2148
rect 8608 2204 8672 2208
rect 8608 2148 8612 2204
rect 8612 2148 8668 2204
rect 8668 2148 8672 2204
rect 8608 2144 8672 2148
rect 8688 2204 8752 2208
rect 8688 2148 8692 2204
rect 8692 2148 8748 2204
rect 8748 2148 8752 2204
rect 8688 2144 8752 2148
rect 12196 2204 12260 2208
rect 12196 2148 12200 2204
rect 12200 2148 12256 2204
rect 12256 2148 12260 2204
rect 12196 2144 12260 2148
rect 12276 2204 12340 2208
rect 12276 2148 12280 2204
rect 12280 2148 12336 2204
rect 12336 2148 12340 2204
rect 12276 2144 12340 2148
rect 12356 2204 12420 2208
rect 12356 2148 12360 2204
rect 12360 2148 12416 2204
rect 12416 2148 12420 2204
rect 12356 2144 12420 2148
rect 12436 2204 12500 2208
rect 12436 2148 12440 2204
rect 12440 2148 12496 2204
rect 12496 2148 12500 2204
rect 12436 2144 12500 2148
rect 9260 1668 9324 1732
<< metal4 >>
rect 2818 16896 3138 17456
rect 2818 16832 2826 16896
rect 2890 16832 2906 16896
rect 2970 16832 2986 16896
rect 3050 16832 3066 16896
rect 3130 16832 3138 16896
rect 2818 15808 3138 16832
rect 2818 15744 2826 15808
rect 2890 15744 2906 15808
rect 2970 15744 2986 15808
rect 3050 15744 3066 15808
rect 3130 15744 3138 15808
rect 2818 14720 3138 15744
rect 2818 14656 2826 14720
rect 2890 14656 2906 14720
rect 2970 14656 2986 14720
rect 3050 14656 3066 14720
rect 3130 14656 3138 14720
rect 2818 13632 3138 14656
rect 2818 13568 2826 13632
rect 2890 13568 2906 13632
rect 2970 13568 2986 13632
rect 3050 13568 3066 13632
rect 3130 13568 3138 13632
rect 2818 12544 3138 13568
rect 2818 12480 2826 12544
rect 2890 12480 2906 12544
rect 2970 12480 2986 12544
rect 3050 12480 3066 12544
rect 3130 12480 3138 12544
rect 2818 11456 3138 12480
rect 2818 11392 2826 11456
rect 2890 11392 2906 11456
rect 2970 11392 2986 11456
rect 3050 11392 3066 11456
rect 3130 11392 3138 11456
rect 2818 10368 3138 11392
rect 2818 10304 2826 10368
rect 2890 10304 2906 10368
rect 2970 10304 2986 10368
rect 3050 10304 3066 10368
rect 3130 10304 3138 10368
rect 2818 9280 3138 10304
rect 2818 9216 2826 9280
rect 2890 9216 2906 9280
rect 2970 9216 2986 9280
rect 3050 9216 3066 9280
rect 3130 9216 3138 9280
rect 2818 8192 3138 9216
rect 2818 8128 2826 8192
rect 2890 8128 2906 8192
rect 2970 8128 2986 8192
rect 3050 8128 3066 8192
rect 3130 8128 3138 8192
rect 2818 7104 3138 8128
rect 2818 7040 2826 7104
rect 2890 7040 2906 7104
rect 2970 7040 2986 7104
rect 3050 7040 3066 7104
rect 3130 7040 3138 7104
rect 2818 6016 3138 7040
rect 2818 5952 2826 6016
rect 2890 5952 2906 6016
rect 2970 5952 2986 6016
rect 3050 5952 3066 6016
rect 3130 5952 3138 6016
rect 2818 4928 3138 5952
rect 2818 4864 2826 4928
rect 2890 4864 2906 4928
rect 2970 4864 2986 4928
rect 3050 4864 3066 4928
rect 3130 4864 3138 4928
rect 2818 3840 3138 4864
rect 2818 3776 2826 3840
rect 2890 3776 2906 3840
rect 2970 3776 2986 3840
rect 3050 3776 3066 3840
rect 3130 3776 3138 3840
rect 2818 2752 3138 3776
rect 2818 2688 2826 2752
rect 2890 2688 2906 2752
rect 2970 2688 2986 2752
rect 3050 2688 3066 2752
rect 3130 2688 3138 2752
rect 2818 2128 3138 2688
rect 4692 17440 5012 17456
rect 4692 17376 4700 17440
rect 4764 17376 4780 17440
rect 4844 17376 4860 17440
rect 4924 17376 4940 17440
rect 5004 17376 5012 17440
rect 4692 16352 5012 17376
rect 4692 16288 4700 16352
rect 4764 16288 4780 16352
rect 4844 16288 4860 16352
rect 4924 16288 4940 16352
rect 5004 16288 5012 16352
rect 4692 15264 5012 16288
rect 4692 15200 4700 15264
rect 4764 15200 4780 15264
rect 4844 15200 4860 15264
rect 4924 15200 4940 15264
rect 5004 15200 5012 15264
rect 4692 14176 5012 15200
rect 4692 14112 4700 14176
rect 4764 14112 4780 14176
rect 4844 14112 4860 14176
rect 4924 14112 4940 14176
rect 5004 14112 5012 14176
rect 4692 13088 5012 14112
rect 4692 13024 4700 13088
rect 4764 13024 4780 13088
rect 4844 13024 4860 13088
rect 4924 13024 4940 13088
rect 5004 13024 5012 13088
rect 4692 12000 5012 13024
rect 4692 11936 4700 12000
rect 4764 11936 4780 12000
rect 4844 11936 4860 12000
rect 4924 11936 4940 12000
rect 5004 11936 5012 12000
rect 4692 10912 5012 11936
rect 4692 10848 4700 10912
rect 4764 10848 4780 10912
rect 4844 10848 4860 10912
rect 4924 10848 4940 10912
rect 5004 10848 5012 10912
rect 4692 9824 5012 10848
rect 4692 9760 4700 9824
rect 4764 9760 4780 9824
rect 4844 9760 4860 9824
rect 4924 9760 4940 9824
rect 5004 9760 5012 9824
rect 4692 8736 5012 9760
rect 6566 16896 6886 17456
rect 6566 16832 6574 16896
rect 6638 16832 6654 16896
rect 6718 16832 6734 16896
rect 6798 16832 6814 16896
rect 6878 16832 6886 16896
rect 6566 15808 6886 16832
rect 6566 15744 6574 15808
rect 6638 15744 6654 15808
rect 6718 15744 6734 15808
rect 6798 15744 6814 15808
rect 6878 15744 6886 15808
rect 6566 14720 6886 15744
rect 6566 14656 6574 14720
rect 6638 14656 6654 14720
rect 6718 14656 6734 14720
rect 6798 14656 6814 14720
rect 6878 14656 6886 14720
rect 6566 13632 6886 14656
rect 6566 13568 6574 13632
rect 6638 13568 6654 13632
rect 6718 13568 6734 13632
rect 6798 13568 6814 13632
rect 6878 13568 6886 13632
rect 6566 12544 6886 13568
rect 6566 12480 6574 12544
rect 6638 12480 6654 12544
rect 6718 12480 6734 12544
rect 6798 12480 6814 12544
rect 6878 12480 6886 12544
rect 6566 11456 6886 12480
rect 6566 11392 6574 11456
rect 6638 11392 6654 11456
rect 6718 11392 6734 11456
rect 6798 11392 6814 11456
rect 6878 11392 6886 11456
rect 6566 10368 6886 11392
rect 6566 10304 6574 10368
rect 6638 10304 6654 10368
rect 6718 10304 6734 10368
rect 6798 10304 6814 10368
rect 6878 10304 6886 10368
rect 5763 9756 5829 9757
rect 5763 9692 5764 9756
rect 5828 9692 5829 9756
rect 5763 9691 5829 9692
rect 4692 8672 4700 8736
rect 4764 8672 4780 8736
rect 4844 8672 4860 8736
rect 4924 8672 4940 8736
rect 5004 8672 5012 8736
rect 4692 7648 5012 8672
rect 4692 7584 4700 7648
rect 4764 7584 4780 7648
rect 4844 7584 4860 7648
rect 4924 7584 4940 7648
rect 5004 7584 5012 7648
rect 4692 6560 5012 7584
rect 4692 6496 4700 6560
rect 4764 6496 4780 6560
rect 4844 6496 4860 6560
rect 4924 6496 4940 6560
rect 5004 6496 5012 6560
rect 4692 5472 5012 6496
rect 4692 5408 4700 5472
rect 4764 5408 4780 5472
rect 4844 5408 4860 5472
rect 4924 5408 4940 5472
rect 5004 5408 5012 5472
rect 4692 4384 5012 5408
rect 4692 4320 4700 4384
rect 4764 4320 4780 4384
rect 4844 4320 4860 4384
rect 4924 4320 4940 4384
rect 5004 4320 5012 4384
rect 4692 3296 5012 4320
rect 4692 3232 4700 3296
rect 4764 3232 4780 3296
rect 4844 3232 4860 3296
rect 4924 3232 4940 3296
rect 5004 3232 5012 3296
rect 4692 2208 5012 3232
rect 5766 2549 5826 9691
rect 6566 9280 6886 10304
rect 6566 9216 6574 9280
rect 6638 9216 6654 9280
rect 6718 9216 6734 9280
rect 6798 9216 6814 9280
rect 6878 9216 6886 9280
rect 6566 8192 6886 9216
rect 6566 8128 6574 8192
rect 6638 8128 6654 8192
rect 6718 8128 6734 8192
rect 6798 8128 6814 8192
rect 6878 8128 6886 8192
rect 6566 7104 6886 8128
rect 6566 7040 6574 7104
rect 6638 7040 6654 7104
rect 6718 7040 6734 7104
rect 6798 7040 6814 7104
rect 6878 7040 6886 7104
rect 6566 6016 6886 7040
rect 6566 5952 6574 6016
rect 6638 5952 6654 6016
rect 6718 5952 6734 6016
rect 6798 5952 6814 6016
rect 6878 5952 6886 6016
rect 6566 4928 6886 5952
rect 6566 4864 6574 4928
rect 6638 4864 6654 4928
rect 6718 4864 6734 4928
rect 6798 4864 6814 4928
rect 6878 4864 6886 4928
rect 6566 3840 6886 4864
rect 6566 3776 6574 3840
rect 6638 3776 6654 3840
rect 6718 3776 6734 3840
rect 6798 3776 6814 3840
rect 6878 3776 6886 3840
rect 6566 2752 6886 3776
rect 6566 2688 6574 2752
rect 6638 2688 6654 2752
rect 6718 2688 6734 2752
rect 6798 2688 6814 2752
rect 6878 2688 6886 2752
rect 5763 2548 5829 2549
rect 5763 2484 5764 2548
rect 5828 2484 5829 2548
rect 5763 2483 5829 2484
rect 4692 2144 4700 2208
rect 4764 2144 4780 2208
rect 4844 2144 4860 2208
rect 4924 2144 4940 2208
rect 5004 2144 5012 2208
rect 4692 2128 5012 2144
rect 6566 2128 6886 2688
rect 8440 17440 8760 17456
rect 8440 17376 8448 17440
rect 8512 17376 8528 17440
rect 8592 17376 8608 17440
rect 8672 17376 8688 17440
rect 8752 17376 8760 17440
rect 8440 16352 8760 17376
rect 8440 16288 8448 16352
rect 8512 16288 8528 16352
rect 8592 16288 8608 16352
rect 8672 16288 8688 16352
rect 8752 16288 8760 16352
rect 8440 15264 8760 16288
rect 8440 15200 8448 15264
rect 8512 15200 8528 15264
rect 8592 15200 8608 15264
rect 8672 15200 8688 15264
rect 8752 15200 8760 15264
rect 8440 14176 8760 15200
rect 8440 14112 8448 14176
rect 8512 14112 8528 14176
rect 8592 14112 8608 14176
rect 8672 14112 8688 14176
rect 8752 14112 8760 14176
rect 8440 13088 8760 14112
rect 8440 13024 8448 13088
rect 8512 13024 8528 13088
rect 8592 13024 8608 13088
rect 8672 13024 8688 13088
rect 8752 13024 8760 13088
rect 8440 12000 8760 13024
rect 8440 11936 8448 12000
rect 8512 11936 8528 12000
rect 8592 11936 8608 12000
rect 8672 11936 8688 12000
rect 8752 11936 8760 12000
rect 8440 10912 8760 11936
rect 8440 10848 8448 10912
rect 8512 10848 8528 10912
rect 8592 10848 8608 10912
rect 8672 10848 8688 10912
rect 8752 10848 8760 10912
rect 8440 9824 8760 10848
rect 8440 9760 8448 9824
rect 8512 9760 8528 9824
rect 8592 9760 8608 9824
rect 8672 9760 8688 9824
rect 8752 9760 8760 9824
rect 8440 8736 8760 9760
rect 10314 16896 10634 17456
rect 10314 16832 10322 16896
rect 10386 16832 10402 16896
rect 10466 16832 10482 16896
rect 10546 16832 10562 16896
rect 10626 16832 10634 16896
rect 10314 15808 10634 16832
rect 10314 15744 10322 15808
rect 10386 15744 10402 15808
rect 10466 15744 10482 15808
rect 10546 15744 10562 15808
rect 10626 15744 10634 15808
rect 10314 14720 10634 15744
rect 10314 14656 10322 14720
rect 10386 14656 10402 14720
rect 10466 14656 10482 14720
rect 10546 14656 10562 14720
rect 10626 14656 10634 14720
rect 10314 13632 10634 14656
rect 10314 13568 10322 13632
rect 10386 13568 10402 13632
rect 10466 13568 10482 13632
rect 10546 13568 10562 13632
rect 10626 13568 10634 13632
rect 10314 12544 10634 13568
rect 10314 12480 10322 12544
rect 10386 12480 10402 12544
rect 10466 12480 10482 12544
rect 10546 12480 10562 12544
rect 10626 12480 10634 12544
rect 10314 11456 10634 12480
rect 10314 11392 10322 11456
rect 10386 11392 10402 11456
rect 10466 11392 10482 11456
rect 10546 11392 10562 11456
rect 10626 11392 10634 11456
rect 10314 10368 10634 11392
rect 10314 10304 10322 10368
rect 10386 10304 10402 10368
rect 10466 10304 10482 10368
rect 10546 10304 10562 10368
rect 10626 10304 10634 10368
rect 9259 9756 9325 9757
rect 9259 9692 9260 9756
rect 9324 9692 9325 9756
rect 9259 9691 9325 9692
rect 8440 8672 8448 8736
rect 8512 8672 8528 8736
rect 8592 8672 8608 8736
rect 8672 8672 8688 8736
rect 8752 8672 8760 8736
rect 8440 7648 8760 8672
rect 8440 7584 8448 7648
rect 8512 7584 8528 7648
rect 8592 7584 8608 7648
rect 8672 7584 8688 7648
rect 8752 7584 8760 7648
rect 8440 6560 8760 7584
rect 8440 6496 8448 6560
rect 8512 6496 8528 6560
rect 8592 6496 8608 6560
rect 8672 6496 8688 6560
rect 8752 6496 8760 6560
rect 8440 5472 8760 6496
rect 8440 5408 8448 5472
rect 8512 5408 8528 5472
rect 8592 5408 8608 5472
rect 8672 5408 8688 5472
rect 8752 5408 8760 5472
rect 8440 4384 8760 5408
rect 8440 4320 8448 4384
rect 8512 4320 8528 4384
rect 8592 4320 8608 4384
rect 8672 4320 8688 4384
rect 8752 4320 8760 4384
rect 8440 3296 8760 4320
rect 8440 3232 8448 3296
rect 8512 3232 8528 3296
rect 8592 3232 8608 3296
rect 8672 3232 8688 3296
rect 8752 3232 8760 3296
rect 8440 2208 8760 3232
rect 8440 2144 8448 2208
rect 8512 2144 8528 2208
rect 8592 2144 8608 2208
rect 8672 2144 8688 2208
rect 8752 2144 8760 2208
rect 8440 2128 8760 2144
rect 9262 1733 9322 9691
rect 10314 9280 10634 10304
rect 10314 9216 10322 9280
rect 10386 9216 10402 9280
rect 10466 9216 10482 9280
rect 10546 9216 10562 9280
rect 10626 9216 10634 9280
rect 10314 8192 10634 9216
rect 10314 8128 10322 8192
rect 10386 8128 10402 8192
rect 10466 8128 10482 8192
rect 10546 8128 10562 8192
rect 10626 8128 10634 8192
rect 10314 7104 10634 8128
rect 10314 7040 10322 7104
rect 10386 7040 10402 7104
rect 10466 7040 10482 7104
rect 10546 7040 10562 7104
rect 10626 7040 10634 7104
rect 10314 6016 10634 7040
rect 10314 5952 10322 6016
rect 10386 5952 10402 6016
rect 10466 5952 10482 6016
rect 10546 5952 10562 6016
rect 10626 5952 10634 6016
rect 10314 4928 10634 5952
rect 10314 4864 10322 4928
rect 10386 4864 10402 4928
rect 10466 4864 10482 4928
rect 10546 4864 10562 4928
rect 10626 4864 10634 4928
rect 10314 3840 10634 4864
rect 10314 3776 10322 3840
rect 10386 3776 10402 3840
rect 10466 3776 10482 3840
rect 10546 3776 10562 3840
rect 10626 3776 10634 3840
rect 10314 2752 10634 3776
rect 10314 2688 10322 2752
rect 10386 2688 10402 2752
rect 10466 2688 10482 2752
rect 10546 2688 10562 2752
rect 10626 2688 10634 2752
rect 10314 2128 10634 2688
rect 12188 17440 12508 17456
rect 12188 17376 12196 17440
rect 12260 17376 12276 17440
rect 12340 17376 12356 17440
rect 12420 17376 12436 17440
rect 12500 17376 12508 17440
rect 12188 16352 12508 17376
rect 12188 16288 12196 16352
rect 12260 16288 12276 16352
rect 12340 16288 12356 16352
rect 12420 16288 12436 16352
rect 12500 16288 12508 16352
rect 12188 15264 12508 16288
rect 12188 15200 12196 15264
rect 12260 15200 12276 15264
rect 12340 15200 12356 15264
rect 12420 15200 12436 15264
rect 12500 15200 12508 15264
rect 12188 14176 12508 15200
rect 12188 14112 12196 14176
rect 12260 14112 12276 14176
rect 12340 14112 12356 14176
rect 12420 14112 12436 14176
rect 12500 14112 12508 14176
rect 12188 13088 12508 14112
rect 12188 13024 12196 13088
rect 12260 13024 12276 13088
rect 12340 13024 12356 13088
rect 12420 13024 12436 13088
rect 12500 13024 12508 13088
rect 12188 12000 12508 13024
rect 12188 11936 12196 12000
rect 12260 11936 12276 12000
rect 12340 11936 12356 12000
rect 12420 11936 12436 12000
rect 12500 11936 12508 12000
rect 12188 10912 12508 11936
rect 12188 10848 12196 10912
rect 12260 10848 12276 10912
rect 12340 10848 12356 10912
rect 12420 10848 12436 10912
rect 12500 10848 12508 10912
rect 12188 9824 12508 10848
rect 12188 9760 12196 9824
rect 12260 9760 12276 9824
rect 12340 9760 12356 9824
rect 12420 9760 12436 9824
rect 12500 9760 12508 9824
rect 12188 8736 12508 9760
rect 12188 8672 12196 8736
rect 12260 8672 12276 8736
rect 12340 8672 12356 8736
rect 12420 8672 12436 8736
rect 12500 8672 12508 8736
rect 12188 7648 12508 8672
rect 12188 7584 12196 7648
rect 12260 7584 12276 7648
rect 12340 7584 12356 7648
rect 12420 7584 12436 7648
rect 12500 7584 12508 7648
rect 12188 6560 12508 7584
rect 12188 6496 12196 6560
rect 12260 6496 12276 6560
rect 12340 6496 12356 6560
rect 12420 6496 12436 6560
rect 12500 6496 12508 6560
rect 12188 5472 12508 6496
rect 12188 5408 12196 5472
rect 12260 5408 12276 5472
rect 12340 5408 12356 5472
rect 12420 5408 12436 5472
rect 12500 5408 12508 5472
rect 12188 4384 12508 5408
rect 12188 4320 12196 4384
rect 12260 4320 12276 4384
rect 12340 4320 12356 4384
rect 12420 4320 12436 4384
rect 12500 4320 12508 4384
rect 12188 3296 12508 4320
rect 12188 3232 12196 3296
rect 12260 3232 12276 3296
rect 12340 3232 12356 3296
rect 12420 3232 12436 3296
rect 12500 3232 12508 3296
rect 12188 2208 12508 3232
rect 12188 2144 12196 2208
rect 12260 2144 12276 2208
rect 12340 2144 12356 2208
rect 12420 2144 12436 2208
rect 12500 2144 12508 2208
rect 12188 2128 12508 2144
rect 14062 16896 14382 17456
rect 14062 16832 14070 16896
rect 14134 16832 14150 16896
rect 14214 16832 14230 16896
rect 14294 16832 14310 16896
rect 14374 16832 14382 16896
rect 14062 15808 14382 16832
rect 14062 15744 14070 15808
rect 14134 15744 14150 15808
rect 14214 15744 14230 15808
rect 14294 15744 14310 15808
rect 14374 15744 14382 15808
rect 14062 14720 14382 15744
rect 14062 14656 14070 14720
rect 14134 14656 14150 14720
rect 14214 14656 14230 14720
rect 14294 14656 14310 14720
rect 14374 14656 14382 14720
rect 14062 13632 14382 14656
rect 14062 13568 14070 13632
rect 14134 13568 14150 13632
rect 14214 13568 14230 13632
rect 14294 13568 14310 13632
rect 14374 13568 14382 13632
rect 14062 12544 14382 13568
rect 14062 12480 14070 12544
rect 14134 12480 14150 12544
rect 14214 12480 14230 12544
rect 14294 12480 14310 12544
rect 14374 12480 14382 12544
rect 14062 11456 14382 12480
rect 14062 11392 14070 11456
rect 14134 11392 14150 11456
rect 14214 11392 14230 11456
rect 14294 11392 14310 11456
rect 14374 11392 14382 11456
rect 14062 10368 14382 11392
rect 14062 10304 14070 10368
rect 14134 10304 14150 10368
rect 14214 10304 14230 10368
rect 14294 10304 14310 10368
rect 14374 10304 14382 10368
rect 14062 9280 14382 10304
rect 14062 9216 14070 9280
rect 14134 9216 14150 9280
rect 14214 9216 14230 9280
rect 14294 9216 14310 9280
rect 14374 9216 14382 9280
rect 14062 8192 14382 9216
rect 14062 8128 14070 8192
rect 14134 8128 14150 8192
rect 14214 8128 14230 8192
rect 14294 8128 14310 8192
rect 14374 8128 14382 8192
rect 14062 7104 14382 8128
rect 14062 7040 14070 7104
rect 14134 7040 14150 7104
rect 14214 7040 14230 7104
rect 14294 7040 14310 7104
rect 14374 7040 14382 7104
rect 14062 6016 14382 7040
rect 14062 5952 14070 6016
rect 14134 5952 14150 6016
rect 14214 5952 14230 6016
rect 14294 5952 14310 6016
rect 14374 5952 14382 6016
rect 14062 4928 14382 5952
rect 14062 4864 14070 4928
rect 14134 4864 14150 4928
rect 14214 4864 14230 4928
rect 14294 4864 14310 4928
rect 14374 4864 14382 4928
rect 14062 3840 14382 4864
rect 14062 3776 14070 3840
rect 14134 3776 14150 3840
rect 14214 3776 14230 3840
rect 14294 3776 14310 3840
rect 14374 3776 14382 3840
rect 14062 2752 14382 3776
rect 14062 2688 14070 2752
rect 14134 2688 14150 2752
rect 14214 2688 14230 2752
rect 14294 2688 14310 2752
rect 14374 2688 14382 2752
rect 14062 2128 14382 2688
rect 9259 1732 9325 1733
rect 9259 1668 9260 1732
rect 9324 1668 9325 1732
rect 9259 1667 9325 1668
use sky130_fd_sc_hd__diode_2  ANTENNA__21__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 2576 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 13984 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 14076 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 15272 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 14812 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 14628 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 15364 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 15180 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 10580 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 11408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 10948 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 11684 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 12236 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 13156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 9108 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 13248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 14536 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 15364 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 14628 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 14812 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 9476 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 10304 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 10764 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 11132 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 12420 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 11960 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 13248 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 12788 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 1840 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18
timestamp 1649977179
transform 1 0 2760 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 1649977179
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46
timestamp 1649977179
transform 1 0 5336 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 1649977179
transform 1 0 7912 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88
timestamp 1649977179
transform 1 0 9200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1649977179
transform 1 0 9568 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_106
timestamp 1649977179
transform 1 0 10856 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_116
timestamp 1649977179
transform 1 0 11776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_120
timestamp 1649977179
transform 1 0 12144 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_134
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_144
timestamp 1649977179
transform 1 0 14352 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_148
timestamp 1649977179
transform 1 0 14720 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_16 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_28
timestamp 1649977179
transform 1 0 3680 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_40
timestamp 1649977179
transform 1 0 4784 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_85
timestamp 1649977179
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_101
timestamp 1649977179
transform 1 0 10396 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_107
timestamp 1649977179
transform 1 0 10948 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_115
timestamp 1649977179
transform 1 0 11684 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_121
timestamp 1649977179
transform 1 0 12236 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_141
timestamp 1649977179
transform 1 0 14076 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_7
timestamp 1649977179
transform 1 0 1748 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_19 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_155
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_157
timestamp 1649977179
transform 1 0 15548 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_7
timestamp 1649977179
transform 1 0 1748 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_19
timestamp 1649977179
transform 1 0 2852 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_31
timestamp 1649977179
transform 1 0 3956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_157
timestamp 1649977179
transform 1 0 15548 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_157
timestamp 1649977179
transform 1 0 15548 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_19
timestamp 1649977179
transform 1 0 2852 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_23
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_40
timestamp 1649977179
transform 1 0 4784 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_46
timestamp 1649977179
transform 1 0 5336 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1649977179
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_68
timestamp 1649977179
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_80
timestamp 1649977179
transform 1 0 8464 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_91
timestamp 1649977179
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_157
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_75
timestamp 1649977179
transform 1 0 8004 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_7
timestamp 1649977179
transform 1 0 1748 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_89
timestamp 1649977179
transform 1 0 9292 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1649977179
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_128
timestamp 1649977179
transform 1 0 12880 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_140
timestamp 1649977179
transform 1 0 13984 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_152
timestamp 1649977179
transform 1 0 15088 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_158
timestamp 1649977179
transform 1 0 15640 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_94
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_106
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_118
timestamp 1649977179
transform 1 0 11960 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_130
timestamp 1649977179
transform 1 0 13064 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_24
timestamp 1649977179
transform 1 0 3312 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_36
timestamp 1649977179
transform 1 0 4416 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_48
timestamp 1649977179
transform 1 0 5520 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_52
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_78
timestamp 1649977179
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_13_96
timestamp 1649977179
transform 1 0 9936 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_26
timestamp 1649977179
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_73
timestamp 1649977179
transform 1 0 7820 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_44
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_62
timestamp 1649977179
transform 1 0 6808 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_67
timestamp 1649977179
transform 1 0 7268 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_84
timestamp 1649977179
transform 1 0 8832 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_157
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_76
timestamp 1649977179
transform 1 0 8096 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_8
timestamp 1649977179
transform 1 0 1840 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_20
timestamp 1649977179
transform 1 0 2944 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_32
timestamp 1649977179
transform 1 0 4048 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_77
timestamp 1649977179
transform 1 0 8188 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_89
timestamp 1649977179
transform 1 0 9292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_101
timestamp 1649977179
transform 1 0 10396 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_109
timestamp 1649977179
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_157
timestamp 1649977179
transform 1 0 15548 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_35
timestamp 1649977179
transform 1 0 4324 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_41
timestamp 1649977179
transform 1 0 4876 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_48
timestamp 1649977179
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_89
timestamp 1649977179
transform 1 0 9292 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_145
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_49
timestamp 1649977179
transform 1 0 5612 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_61
timestamp 1649977179
transform 1 0 6716 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_73
timestamp 1649977179
transform 1 0 7820 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_81
timestamp 1649977179
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_31
timestamp 1649977179
transform 1 0 3956 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_157
timestamp 1649977179
transform 1 0 15548 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_157
timestamp 1649977179
transform 1 0 15548 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_8
timestamp 1649977179
transform 1 0 1840 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_20
timestamp 1649977179
transform 1 0 2944 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_32
timestamp 1649977179
transform 1 0 4048 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_44
timestamp 1649977179
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_16
timestamp 1649977179
transform 1 0 2576 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_87
timestamp 1649977179
transform 1 0 9108 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_99
timestamp 1649977179
transform 1 0 10212 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1649977179
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_115
timestamp 1649977179
transform 1 0 11684 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_118
timestamp 1649977179
transform 1 0 11960 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_124
timestamp 1649977179
transform 1 0 12512 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_127
timestamp 1649977179
transform 1 0 12788 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_132
timestamp 1649977179
transform 1 0 13248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1649977179
transform 1 0 15640 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_29
timestamp 1649977179
transform 1 0 3772 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_67
timestamp 1649977179
transform 1 0 7268 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_72
timestamp 1649977179
transform 1 0 7728 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_94
timestamp 1649977179
transform 1 0 9752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_108
timestamp 1649977179
transform 1 0 11040 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_117
timestamp 1649977179
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_126
timestamp 1649977179
transform 1 0 12696 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_135
timestamp 1649977179
transform 1 0 13524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_139
timestamp 1649977179
transform 1 0 13892 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 16008 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 16008 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 16008 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 16008 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 16008 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 16008 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 16008 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 16008 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 16008 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 16008 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 16008 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 16008 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 16008 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 16008 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 16008 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 16008 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 3680 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _02_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _03_
timestamp 1649977179
transform 1 0 4600 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _04_
timestamp 1649977179
transform 1 0 5612 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _05_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _06_
timestamp 1649977179
transform 1 0 6532 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _07_
timestamp 1649977179
transform 1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _08_
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _09_
timestamp 1649977179
transform 1 0 7912 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _10_
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _11_
timestamp 1649977179
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _12_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _13_
timestamp 1649977179
transform 1 0 10304 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _14_
timestamp 1649977179
transform 1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _15_
timestamp 1649977179
transform 1 0 11408 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _16_
timestamp 1649977179
transform 1 0 11960 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _17_
timestamp 1649977179
transform 1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _18_
timestamp 1649977179
transform 1 0 12512 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _19_
timestamp 1649977179
transform 1 0 13064 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _20_
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _21_
timestamp 1649977179
transform -1 0 14444 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _22_
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1649977179
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _24_
timestamp 1649977179
transform 1 0 4508 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _25_
timestamp 1649977179
transform 1 0 5428 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _26_
timestamp 1649977179
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1649977179
transform 1 0 5704 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _28_
timestamp 1649977179
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _29_
timestamp 1649977179
transform 1 0 5980 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _30_
timestamp 1649977179
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _31_
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _32_
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _33_
timestamp 1649977179
transform 1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _34_
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _35_
timestamp 1649977179
transform 1 0 10580 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _36_
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _37_
timestamp 1649977179
transform 1 0 11684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _38_
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _39_
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _40_
timestamp 1649977179
transform 1 0 12788 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _41_
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _42_
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 8096 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.prog_clk
timestamp 1649977179
transform -1 0 4416 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 2392 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 13524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform 1 0 15272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 15456 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 10120 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 10580 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 10948 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform 1 0 12696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform 1 0 13248 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform 1 0 13616 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 14076 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 14536 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 14904 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 15364 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 15088 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 14812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 15456 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 9476 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 10120 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 11592 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 11960 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 12420 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 1656 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform -1 0 2392 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.INV_SOC_DIR .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.IN_PROTECT_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5888 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_2  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.ISOL_EN_GATE .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 4692 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_8  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_0_.OUT_PROTECT_GATE
timestamp 1649977179
transform -1 0 3312 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfxtp_1  logical_tile_io_mode_io__0.ltile_phy_iopad_0.EMBEDDED_IO_HD_sky130_fd_sc_hd__dfxtp_1_mem.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 7360 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 8280 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_ipin_0.sky130_fd_sc_hd__dfxtp_1_3_
timestamp 1649977179
transform -1 0 8188 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9384 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 8832 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9108 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_2_
timestamp 1649977179
transform 1 0 9200 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_ipin_0.mux_l2_in_3__89 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l2_in_3_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 7084 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l3_in_1_
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_ipin_0.mux_l4_in_0_
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_ipin_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2944 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output45 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15364 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output46
timestamp 1649977179
transform -1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output47
timestamp 1649977179
transform -1 0 4876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output48
timestamp 1649977179
transform -1 0 5336 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output49
timestamp 1649977179
transform -1 0 5796 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output50
timestamp 1649977179
transform -1 0 6164 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output51
timestamp 1649977179
transform -1 0 6716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output52
timestamp 1649977179
transform -1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output53
timestamp 1649977179
transform -1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 7912 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform -1 0 8372 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform -1 0 8740 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform -1 0 1748 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform -1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform -1 0 2760 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 3220 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 3588 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform -1 0 4140 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform -1 0 4508 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform -1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform -1 0 5152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 5520 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform -1 0 6256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform -1 0 6900 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 7268 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform -1 0 8188 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform -1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform -1 0 9292 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 1840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform -1 0 2576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 2944 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 3680 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 4416 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 4784 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform -1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 15364 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12696 0 -1 8704
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 202 19200 258 20000 6 IO_ISOL_N
port 0 nsew signal input
rlabel metal4 s 4692 2128 5012 17456 6 VGND
port 1 nsew ground input
rlabel metal4 s 8440 2128 8760 17456 6 VGND
port 1 nsew ground input
rlabel metal4 s 12188 2128 12508 17456 6 VGND
port 1 nsew ground input
rlabel metal4 s 2818 2128 3138 17456 6 VPWR
port 2 nsew power input
rlabel metal4 s 6566 2128 6886 17456 6 VPWR
port 2 nsew power input
rlabel metal4 s 10314 2128 10634 17456 6 VPWR
port 2 nsew power input
rlabel metal4 s 14062 2128 14382 17456 6 VPWR
port 2 nsew power input
rlabel metal3 s 0 18232 800 18352 6 ccff_head
port 3 nsew signal input
rlabel metal3 s 16400 12384 17200 12504 6 ccff_tail
port 4 nsew signal tristate
rlabel metal2 s 8758 0 8814 800 6 chany_bottom_in[0]
port 5 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 chany_bottom_in[10]
port 6 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 chany_bottom_in[11]
port 7 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 chany_bottom_in[12]
port 8 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_in[13]
port 9 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 chany_bottom_in[14]
port 10 nsew signal input
rlabel metal2 s 15198 0 15254 800 6 chany_bottom_in[15]
port 11 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 chany_bottom_in[16]
port 12 nsew signal input
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_in[17]
port 13 nsew signal input
rlabel metal2 s 16486 0 16542 800 6 chany_bottom_in[18]
port 14 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 chany_bottom_in[19]
port 15 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 chany_bottom_in[1]
port 16 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 chany_bottom_in[2]
port 17 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[3]
port 18 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 chany_bottom_in[4]
port 19 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 chany_bottom_in[5]
port 20 nsew signal input
rlabel metal2 s 11334 0 11390 800 6 chany_bottom_in[6]
port 21 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 chany_bottom_in[7]
port 22 nsew signal input
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_in[8]
port 23 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 chany_bottom_in[9]
port 24 nsew signal input
rlabel metal2 s 202 0 258 800 6 chany_bottom_out[0]
port 25 nsew signal tristate
rlabel metal2 s 4434 0 4490 800 6 chany_bottom_out[10]
port 26 nsew signal tristate
rlabel metal2 s 4894 0 4950 800 6 chany_bottom_out[11]
port 27 nsew signal tristate
rlabel metal2 s 5354 0 5410 800 6 chany_bottom_out[12]
port 28 nsew signal tristate
rlabel metal2 s 5722 0 5778 800 6 chany_bottom_out[13]
port 29 nsew signal tristate
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_out[14]
port 30 nsew signal tristate
rlabel metal2 s 6642 0 6698 800 6 chany_bottom_out[15]
port 31 nsew signal tristate
rlabel metal2 s 7010 0 7066 800 6 chany_bottom_out[16]
port 32 nsew signal tristate
rlabel metal2 s 7470 0 7526 800 6 chany_bottom_out[17]
port 33 nsew signal tristate
rlabel metal2 s 7930 0 7986 800 6 chany_bottom_out[18]
port 34 nsew signal tristate
rlabel metal2 s 8298 0 8354 800 6 chany_bottom_out[19]
port 35 nsew signal tristate
rlabel metal2 s 570 0 626 800 6 chany_bottom_out[1]
port 36 nsew signal tristate
rlabel metal2 s 1030 0 1086 800 6 chany_bottom_out[2]
port 37 nsew signal tristate
rlabel metal2 s 1490 0 1546 800 6 chany_bottom_out[3]
port 38 nsew signal tristate
rlabel metal2 s 1858 0 1914 800 6 chany_bottom_out[4]
port 39 nsew signal tristate
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_out[5]
port 40 nsew signal tristate
rlabel metal2 s 2778 0 2834 800 6 chany_bottom_out[6]
port 41 nsew signal tristate
rlabel metal2 s 3146 0 3202 800 6 chany_bottom_out[7]
port 42 nsew signal tristate
rlabel metal2 s 3606 0 3662 800 6 chany_bottom_out[8]
port 43 nsew signal tristate
rlabel metal2 s 4066 0 4122 800 6 chany_bottom_out[9]
port 44 nsew signal tristate
rlabel metal2 s 8942 19200 8998 20000 6 chany_top_in[0]
port 45 nsew signal input
rlabel metal2 s 13174 19200 13230 20000 6 chany_top_in[10]
port 46 nsew signal input
rlabel metal2 s 13542 19200 13598 20000 6 chany_top_in[11]
port 47 nsew signal input
rlabel metal2 s 14002 19200 14058 20000 6 chany_top_in[12]
port 48 nsew signal input
rlabel metal2 s 14462 19200 14518 20000 6 chany_top_in[13]
port 49 nsew signal input
rlabel metal2 s 14830 19200 14886 20000 6 chany_top_in[14]
port 50 nsew signal input
rlabel metal2 s 15290 19200 15346 20000 6 chany_top_in[15]
port 51 nsew signal input
rlabel metal2 s 15658 19200 15714 20000 6 chany_top_in[16]
port 52 nsew signal input
rlabel metal2 s 16118 19200 16174 20000 6 chany_top_in[17]
port 53 nsew signal input
rlabel metal2 s 16486 19200 16542 20000 6 chany_top_in[18]
port 54 nsew signal input
rlabel metal2 s 16946 19200 17002 20000 6 chany_top_in[19]
port 55 nsew signal input
rlabel metal2 s 9402 19200 9458 20000 6 chany_top_in[1]
port 56 nsew signal input
rlabel metal2 s 9770 19200 9826 20000 6 chany_top_in[2]
port 57 nsew signal input
rlabel metal2 s 10230 19200 10286 20000 6 chany_top_in[3]
port 58 nsew signal input
rlabel metal2 s 10690 19200 10746 20000 6 chany_top_in[4]
port 59 nsew signal input
rlabel metal2 s 11058 19200 11114 20000 6 chany_top_in[5]
port 60 nsew signal input
rlabel metal2 s 11518 19200 11574 20000 6 chany_top_in[6]
port 61 nsew signal input
rlabel metal2 s 11886 19200 11942 20000 6 chany_top_in[7]
port 62 nsew signal input
rlabel metal2 s 12346 19200 12402 20000 6 chany_top_in[8]
port 63 nsew signal input
rlabel metal2 s 12714 19200 12770 20000 6 chany_top_in[9]
port 64 nsew signal input
rlabel metal2 s 570 19200 626 20000 6 chany_top_out[0]
port 65 nsew signal tristate
rlabel metal2 s 4802 19200 4858 20000 6 chany_top_out[10]
port 66 nsew signal tristate
rlabel metal2 s 5170 19200 5226 20000 6 chany_top_out[11]
port 67 nsew signal tristate
rlabel metal2 s 5630 19200 5686 20000 6 chany_top_out[12]
port 68 nsew signal tristate
rlabel metal2 s 5998 19200 6054 20000 6 chany_top_out[13]
port 69 nsew signal tristate
rlabel metal2 s 6458 19200 6514 20000 6 chany_top_out[14]
port 70 nsew signal tristate
rlabel metal2 s 6826 19200 6882 20000 6 chany_top_out[15]
port 71 nsew signal tristate
rlabel metal2 s 7286 19200 7342 20000 6 chany_top_out[16]
port 72 nsew signal tristate
rlabel metal2 s 7746 19200 7802 20000 6 chany_top_out[17]
port 73 nsew signal tristate
rlabel metal2 s 8114 19200 8170 20000 6 chany_top_out[18]
port 74 nsew signal tristate
rlabel metal2 s 8574 19200 8630 20000 6 chany_top_out[19]
port 75 nsew signal tristate
rlabel metal2 s 1030 19200 1086 20000 6 chany_top_out[1]
port 76 nsew signal tristate
rlabel metal2 s 1398 19200 1454 20000 6 chany_top_out[2]
port 77 nsew signal tristate
rlabel metal2 s 1858 19200 1914 20000 6 chany_top_out[3]
port 78 nsew signal tristate
rlabel metal2 s 2226 19200 2282 20000 6 chany_top_out[4]
port 79 nsew signal tristate
rlabel metal2 s 2686 19200 2742 20000 6 chany_top_out[5]
port 80 nsew signal tristate
rlabel metal2 s 3054 19200 3110 20000 6 chany_top_out[6]
port 81 nsew signal tristate
rlabel metal2 s 3514 19200 3570 20000 6 chany_top_out[7]
port 82 nsew signal tristate
rlabel metal2 s 3974 19200 4030 20000 6 chany_top_out[8]
port 83 nsew signal tristate
rlabel metal2 s 4342 19200 4398 20000 6 chany_top_out[9]
port 84 nsew signal tristate
rlabel metal3 s 0 8304 800 8424 6 gfpga_pad_EMBEDDED_IO_HD_SOC_DIR
port 85 nsew signal tristate
rlabel metal3 s 0 11568 800 11688 6 gfpga_pad_EMBEDDED_IO_HD_SOC_IN
port 86 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 gfpga_pad_EMBEDDED_IO_HD_SOC_OUT
port 87 nsew signal tristate
rlabel metal3 s 0 4904 800 5024 6 left_grid_pin_0_
port 88 nsew signal tristate
rlabel metal3 s 16400 7352 17200 7472 6 prog_clk_0_E_in
port 89 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 right_width_0_height_0__pin_0_
port 90 nsew signal input
rlabel metal3 s 16400 2456 17200 2576 6 right_width_0_height_0__pin_1_lower
port 91 nsew signal tristate
rlabel metal3 s 16400 17416 17200 17536 6 right_width_0_height_0__pin_1_upper
port 92 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 17200 20000
<< end >>
