module tie_array (VGND,
    VPWR,
    x);
 inout VGND;
 inout VPWR;
 output [7:0] x;

 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;

 sky130_fd_sc_hd__decap_3 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_0_88 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_10_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_102 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_11_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_12_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_102 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_13_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_14_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_102 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_15_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_100 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_59 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_83 ();
 sky130_fd_sc_hd__decap_12 FILLER_16_88 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_28 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_57 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_2_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_99 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_20 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_31 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_12 FILLER_3_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_95 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_4_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_99 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_100 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_82 ();
 sky130_fd_sc_hd__decap_12 FILLER_5_88 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_6_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_102 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_7_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_94 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_30 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_42 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_54 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_78 ();
 sky130_fd_sc_hd__decap_12 FILLER_8_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_102 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_51 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_58 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_70 ();
 sky130_fd_sc_hd__decap_12 FILLER_9_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_94 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__conb_1 \conb_1[0]  (.LO(net1));
 sky130_fd_sc_hd__conb_1 \conb_1[1]  (.LO(net2));
 sky130_fd_sc_hd__conb_1 \conb_1[2]  (.LO(net3));
 sky130_fd_sc_hd__conb_1 \conb_1[3]  (.LO(net4));
 sky130_fd_sc_hd__conb_1 \conb_1[4]  (.LO(net5));
 sky130_fd_sc_hd__conb_1 \conb_1[5]  (.LO(net6));
 sky130_fd_sc_hd__conb_1 \conb_1[6]  (.LO(net7));
 sky130_fd_sc_hd__conb_1 \conb_1[7]  (.LO(net8));
 sky130_fd_sc_hd__clkbuf_2 output1 (.A(net1),
    .X(x[0]));
 sky130_fd_sc_hd__clkbuf_2 output2 (.A(net2),
    .X(x[1]));
 sky130_fd_sc_hd__clkbuf_2 output3 (.A(net3),
    .X(x[2]));
 sky130_fd_sc_hd__clkbuf_2 output4 (.A(net4),
    .X(x[3]));
 sky130_fd_sc_hd__clkbuf_2 output5 (.A(net5),
    .X(x[4]));
 sky130_fd_sc_hd__clkbuf_2 output6 (.A(net6),
    .X(x[5]));
 sky130_fd_sc_hd__clkbuf_2 output7 (.A(net7),
    .X(x[6]));
 sky130_fd_sc_hd__clkbuf_2 output8 (.A(net8),
    .X(x[7]));
endmodule
