magic
tech sky130A
magscale 1 2
timestamp 1650625444
<< viali >>
rect 19625 20553 19659 20587
rect 18797 20485 18831 20519
rect 20177 20485 20211 20519
rect 5825 20417 5859 20451
rect 6377 20417 6411 20451
rect 17509 20417 17543 20451
rect 17785 20417 17819 20451
rect 19441 20417 19475 20451
rect 20545 20417 20579 20451
rect 21097 20417 21131 20451
rect 6009 20213 6043 20247
rect 17325 20213 17359 20247
rect 20085 20213 20119 20247
rect 20729 20213 20763 20247
rect 21281 20213 21315 20247
rect 18889 20009 18923 20043
rect 20177 20009 20211 20043
rect 20729 20009 20763 20043
rect 13093 19941 13127 19975
rect 6377 19805 6411 19839
rect 12909 19805 12943 19839
rect 18705 19805 18739 19839
rect 19533 19805 19567 19839
rect 19993 19805 20027 19839
rect 20545 19805 20579 19839
rect 21097 19805 21131 19839
rect 6561 19737 6595 19771
rect 19717 19669 19751 19703
rect 21281 19669 21315 19703
rect 19717 19465 19751 19499
rect 19993 19465 20027 19499
rect 21281 19465 21315 19499
rect 18429 19329 18463 19363
rect 19073 19329 19107 19363
rect 19533 19329 19567 19363
rect 20177 19329 20211 19363
rect 20545 19329 20579 19363
rect 21097 19329 21131 19363
rect 18613 19193 18647 19227
rect 19257 19193 19291 19227
rect 20729 19193 20763 19227
rect 12173 18921 12207 18955
rect 20361 18921 20395 18955
rect 20821 18921 20855 18955
rect 9505 18717 9539 18751
rect 11989 18717 12023 18751
rect 20177 18717 20211 18751
rect 20637 18717 20671 18751
rect 21097 18717 21131 18751
rect 9689 18581 9723 18615
rect 21281 18581 21315 18615
rect 12449 18377 12483 18411
rect 8401 18241 8435 18275
rect 12265 18241 12299 18275
rect 20821 18241 20855 18275
rect 21097 18241 21131 18275
rect 8585 18105 8619 18139
rect 20637 18037 20671 18071
rect 21281 18037 21315 18071
rect 11621 17833 11655 17867
rect 20269 17833 20303 17867
rect 11437 17629 11471 17663
rect 20085 17629 20119 17663
rect 20545 17629 20579 17663
rect 21097 17629 21131 17663
rect 20729 17493 20763 17527
rect 21281 17493 21315 17527
rect 20085 17289 20119 17323
rect 20821 17289 20855 17323
rect 19901 17153 19935 17187
rect 20637 17153 20671 17187
rect 21097 17153 21131 17187
rect 21281 16949 21315 16983
rect 20821 16745 20855 16779
rect 18245 16541 18279 16575
rect 20177 16541 20211 16575
rect 20637 16541 20671 16575
rect 21097 16541 21131 16575
rect 18429 16405 18463 16439
rect 20361 16405 20395 16439
rect 21281 16405 21315 16439
rect 14749 16201 14783 16235
rect 20177 16201 20211 16235
rect 20821 16201 20855 16235
rect 14565 16065 14599 16099
rect 19993 16065 20027 16099
rect 20637 16065 20671 16099
rect 21097 16065 21131 16099
rect 19717 15861 19751 15895
rect 21281 15861 21315 15895
rect 20361 15657 20395 15691
rect 18889 15453 18923 15487
rect 19717 15453 19751 15487
rect 20177 15453 20211 15487
rect 20637 15453 20671 15487
rect 21097 15453 21131 15487
rect 19441 15317 19475 15351
rect 19901 15317 19935 15351
rect 20821 15317 20855 15351
rect 21281 15317 21315 15351
rect 9505 15113 9539 15147
rect 20361 15113 20395 15147
rect 20821 15113 20855 15147
rect 9321 14977 9355 15011
rect 11621 14977 11655 15011
rect 19257 14977 19291 15011
rect 19717 14977 19751 15011
rect 20177 14977 20211 15011
rect 20637 14977 20671 15011
rect 21097 14977 21131 15011
rect 18889 14909 18923 14943
rect 11805 14841 11839 14875
rect 19901 14841 19935 14875
rect 18245 14773 18279 14807
rect 19441 14773 19475 14807
rect 21281 14773 21315 14807
rect 20085 14569 20119 14603
rect 17969 14501 18003 14535
rect 20361 14501 20395 14535
rect 8953 14365 8987 14399
rect 17509 14365 17543 14399
rect 17785 14365 17819 14399
rect 18429 14365 18463 14399
rect 18705 14365 18739 14399
rect 19625 14365 19659 14399
rect 19901 14365 19935 14399
rect 20545 14365 20579 14399
rect 21097 14365 21131 14399
rect 9137 14229 9171 14263
rect 18245 14229 18279 14263
rect 18889 14229 18923 14263
rect 19441 14229 19475 14263
rect 21281 14229 21315 14263
rect 11713 14025 11747 14059
rect 18153 14025 18187 14059
rect 19073 14025 19107 14059
rect 20453 13957 20487 13991
rect 11529 13889 11563 13923
rect 17141 13889 17175 13923
rect 17969 13889 18003 13923
rect 18889 13889 18923 13923
rect 19349 13889 19383 13923
rect 19993 13889 20027 13923
rect 21097 13889 21131 13923
rect 16681 13821 16715 13855
rect 17417 13821 17451 13855
rect 18613 13821 18647 13855
rect 13737 13481 13771 13515
rect 20361 13481 20395 13515
rect 16129 13413 16163 13447
rect 13553 13277 13587 13311
rect 17242 13277 17276 13311
rect 17509 13277 17543 13311
rect 17969 13277 18003 13311
rect 18429 13277 18463 13311
rect 19257 13277 19291 13311
rect 20177 13277 20211 13311
rect 20729 13277 20763 13311
rect 15761 13141 15795 13175
rect 17785 13141 17819 13175
rect 18245 13141 18279 13175
rect 18705 13141 18739 13175
rect 19901 13141 19935 13175
rect 21373 13141 21407 13175
rect 18061 12937 18095 12971
rect 15853 12869 15887 12903
rect 17417 12801 17451 12835
rect 17969 12801 18003 12835
rect 18797 12801 18831 12835
rect 20361 12801 20395 12835
rect 20637 12801 20671 12835
rect 16313 12733 16347 12767
rect 17877 12733 17911 12767
rect 18429 12665 18463 12699
rect 15209 12597 15243 12631
rect 16773 12597 16807 12631
rect 19441 12597 19475 12631
rect 19717 12597 19751 12631
rect 21281 12597 21315 12631
rect 15485 12393 15519 12427
rect 18797 12393 18831 12427
rect 21281 12393 21315 12427
rect 15025 12189 15059 12223
rect 15301 12189 15335 12223
rect 15761 12189 15795 12223
rect 17417 12189 17451 12223
rect 19257 12189 19291 12223
rect 19524 12189 19558 12223
rect 21097 12189 21131 12223
rect 16028 12121 16062 12155
rect 17684 12121 17718 12155
rect 14197 12053 14231 12087
rect 14473 12053 14507 12087
rect 14841 12053 14875 12087
rect 17141 12053 17175 12087
rect 20637 12053 20671 12087
rect 15025 11849 15059 11883
rect 16221 11849 16255 11883
rect 17785 11849 17819 11883
rect 20453 11849 20487 11883
rect 18328 11781 18362 11815
rect 1685 11713 1719 11747
rect 13921 11713 13955 11747
rect 15209 11713 15243 11747
rect 15853 11713 15887 11747
rect 16681 11713 16715 11747
rect 17141 11713 17175 11747
rect 20361 11713 20395 11747
rect 21097 11713 21131 11747
rect 15577 11645 15611 11679
rect 15761 11645 15795 11679
rect 18061 11645 18095 11679
rect 20545 11645 20579 11679
rect 2053 11577 2087 11611
rect 13645 11577 13679 11611
rect 19441 11577 19475 11611
rect 1501 11509 1535 11543
rect 13277 11509 13311 11543
rect 14565 11509 14599 11543
rect 19993 11509 20027 11543
rect 21281 11509 21315 11543
rect 12449 11305 12483 11339
rect 16681 11305 16715 11339
rect 19809 11305 19843 11339
rect 13277 11237 13311 11271
rect 16129 11237 16163 11271
rect 18613 11237 18647 11271
rect 19257 11237 19291 11271
rect 13737 11169 13771 11203
rect 17141 11169 17175 11203
rect 13093 11101 13127 11135
rect 14749 11101 14783 11135
rect 16497 11101 16531 11135
rect 17969 11101 18003 11135
rect 19441 11101 19475 11135
rect 21189 11101 21223 11135
rect 12817 11033 12851 11067
rect 15016 11033 15050 11067
rect 20922 11033 20956 11067
rect 14289 10965 14323 10999
rect 17233 10965 17267 10999
rect 17325 10965 17359 10999
rect 17693 10965 17727 10999
rect 13921 10761 13955 10795
rect 19441 10761 19475 10795
rect 19809 10761 19843 10795
rect 19901 10761 19935 10795
rect 20913 10761 20947 10795
rect 14464 10693 14498 10727
rect 19073 10693 19107 10727
rect 20821 10693 20855 10727
rect 12265 10625 12299 10659
rect 12808 10625 12842 10659
rect 14197 10625 14231 10659
rect 16313 10625 16347 10659
rect 18081 10625 18115 10659
rect 12541 10557 12575 10591
rect 18337 10557 18371 10591
rect 18613 10557 18647 10591
rect 19993 10557 20027 10591
rect 21005 10557 21039 10591
rect 12081 10489 12115 10523
rect 11805 10421 11839 10455
rect 15577 10421 15611 10455
rect 16129 10421 16163 10455
rect 16957 10421 16991 10455
rect 20453 10421 20487 10455
rect 14841 10217 14875 10251
rect 15853 10217 15887 10251
rect 16773 10217 16807 10251
rect 17049 10217 17083 10251
rect 20361 10217 20395 10251
rect 18889 10149 18923 10183
rect 14197 10081 14231 10115
rect 15301 10081 15335 10115
rect 19809 10081 19843 10115
rect 19901 10081 19935 10115
rect 11161 10013 11195 10047
rect 13553 10013 13587 10047
rect 14473 10013 14507 10047
rect 16129 10013 16163 10047
rect 17233 10013 17267 10047
rect 17509 10013 17543 10047
rect 19717 10013 19751 10047
rect 21005 10013 21039 10047
rect 15485 9945 15519 9979
rect 17754 9945 17788 9979
rect 11805 9877 11839 9911
rect 12081 9877 12115 9911
rect 12541 9877 12575 9911
rect 12909 9877 12943 9911
rect 14381 9877 14415 9911
rect 15393 9877 15427 9911
rect 19349 9877 19383 9911
rect 21373 9877 21407 9911
rect 11161 9673 11195 9707
rect 12909 9673 12943 9707
rect 18061 9673 18095 9707
rect 9045 9605 9079 9639
rect 14197 9605 14231 9639
rect 15761 9605 15795 9639
rect 17049 9605 17083 9639
rect 18153 9605 18187 9639
rect 19840 9605 19874 9639
rect 21005 9605 21039 9639
rect 9137 9537 9171 9571
rect 9781 9537 9815 9571
rect 10048 9537 10082 9571
rect 11529 9537 11563 9571
rect 11796 9537 11830 9571
rect 13553 9537 13587 9571
rect 14841 9537 14875 9571
rect 20361 9537 20395 9571
rect 8861 9469 8895 9503
rect 14013 9469 14047 9503
rect 14105 9469 14139 9503
rect 16221 9469 16255 9503
rect 16773 9469 16807 9503
rect 16957 9469 16991 9503
rect 18245 9469 18279 9503
rect 20085 9469 20119 9503
rect 9505 9401 9539 9435
rect 13369 9401 13403 9435
rect 14565 9401 14599 9435
rect 17693 9401 17727 9435
rect 18705 9401 18739 9435
rect 15485 9333 15519 9367
rect 17417 9333 17451 9367
rect 21281 9333 21315 9367
rect 13737 9129 13771 9163
rect 18153 9129 18187 9163
rect 20913 9129 20947 9163
rect 10701 9061 10735 9095
rect 17785 9061 17819 9095
rect 7665 8993 7699 9027
rect 11161 8993 11195 9027
rect 18613 8993 18647 9027
rect 18797 8993 18831 9027
rect 7941 8925 7975 8959
rect 8953 8925 8987 8959
rect 11345 8925 11379 8959
rect 12357 8925 12391 8959
rect 12624 8925 12658 8959
rect 14105 8925 14139 8959
rect 15761 8925 15795 8959
rect 17601 8925 17635 8959
rect 19533 8925 19567 8959
rect 21373 8925 21407 8959
rect 8585 8857 8619 8891
rect 9198 8857 9232 8891
rect 14372 8857 14406 8891
rect 16028 8857 16062 8891
rect 19800 8857 19834 8891
rect 10333 8789 10367 8823
rect 11253 8789 11287 8823
rect 11713 8789 11747 8823
rect 12081 8789 12115 8823
rect 15485 8789 15519 8823
rect 17141 8789 17175 8823
rect 18521 8789 18555 8823
rect 21189 8789 21223 8823
rect 8125 8585 8159 8619
rect 11161 8585 11195 8619
rect 12173 8585 12207 8619
rect 13645 8585 13679 8619
rect 14841 8585 14875 8619
rect 16037 8585 16071 8619
rect 18337 8585 18371 8619
rect 19533 8585 19567 8619
rect 19993 8585 20027 8619
rect 10793 8517 10827 8551
rect 13277 8517 13311 8551
rect 14473 8517 14507 8551
rect 18705 8517 18739 8551
rect 21106 8517 21140 8551
rect 9238 8449 9272 8483
rect 9505 8449 9539 8483
rect 9965 8449 9999 8483
rect 11529 8449 11563 8483
rect 13185 8449 13219 8483
rect 14381 8449 14415 8483
rect 15669 8449 15703 8483
rect 16681 8449 16715 8483
rect 16948 8449 16982 8483
rect 19349 8449 19383 8483
rect 21373 8449 21407 8483
rect 10517 8381 10551 8415
rect 10701 8381 10735 8415
rect 12633 8381 12667 8415
rect 13001 8381 13035 8415
rect 14197 8381 14231 8415
rect 15485 8381 15519 8415
rect 15577 8381 15611 8415
rect 18797 8381 18831 8415
rect 18889 8381 18923 8415
rect 18061 8313 18095 8347
rect 10149 8245 10183 8279
rect 10885 8041 10919 8075
rect 13093 8041 13127 8075
rect 17877 8041 17911 8075
rect 19717 7973 19751 8007
rect 9597 7905 9631 7939
rect 19257 7905 19291 7939
rect 20269 7905 20303 7939
rect 7481 7837 7515 7871
rect 8585 7837 8619 7871
rect 9689 7837 9723 7871
rect 12817 7837 12851 7871
rect 13737 7837 13771 7871
rect 16129 7837 16163 7871
rect 18613 7837 18647 7871
rect 20085 7837 20119 7871
rect 20729 7837 20763 7871
rect 6929 7769 6963 7803
rect 12173 7769 12207 7803
rect 14381 7769 14415 7803
rect 16405 7769 16439 7803
rect 7665 7701 7699 7735
rect 7941 7701 7975 7735
rect 9137 7701 9171 7735
rect 9781 7701 9815 7735
rect 10149 7701 10183 7735
rect 12633 7701 12667 7735
rect 18797 7701 18831 7735
rect 20177 7701 20211 7735
rect 21373 7701 21407 7735
rect 10609 7497 10643 7531
rect 11161 7497 11195 7531
rect 13645 7497 13679 7531
rect 16221 7497 16255 7531
rect 18337 7497 18371 7531
rect 19993 7497 20027 7531
rect 20545 7497 20579 7531
rect 20913 7497 20947 7531
rect 6653 7429 6687 7463
rect 8309 7429 8343 7463
rect 9485 7429 9519 7463
rect 14188 7429 14222 7463
rect 17224 7429 17258 7463
rect 7389 7361 7423 7395
rect 7849 7361 7883 7395
rect 8953 7361 8987 7395
rect 10977 7361 11011 7395
rect 11989 7361 12023 7395
rect 12265 7361 12299 7395
rect 12532 7361 12566 7395
rect 13921 7361 13955 7395
rect 15577 7361 15611 7395
rect 18613 7361 18647 7395
rect 19901 7361 19935 7395
rect 21005 7361 21039 7395
rect 7113 7293 7147 7327
rect 9229 7293 9263 7327
rect 16957 7293 16991 7327
rect 19257 7293 19291 7327
rect 20177 7293 20211 7327
rect 21097 7293 21131 7327
rect 8033 7225 8067 7259
rect 7573 7157 7607 7191
rect 11805 7157 11839 7191
rect 15301 7157 15335 7191
rect 19533 7157 19567 7191
rect 7941 6885 7975 6919
rect 9689 6885 9723 6919
rect 11897 6885 11931 6919
rect 5825 6817 5859 6851
rect 9045 6817 9079 6851
rect 10517 6817 10551 6851
rect 12725 6817 12759 6851
rect 15393 6817 15427 6851
rect 16773 6817 16807 6851
rect 17417 6817 17451 6851
rect 18245 6817 18279 6851
rect 6561 6749 6595 6783
rect 7021 6749 7055 6783
rect 8585 6749 8619 6783
rect 9321 6749 9355 6783
rect 10057 6749 10091 6783
rect 12541 6749 12575 6783
rect 13461 6749 13495 6783
rect 14933 6749 14967 6783
rect 15577 6749 15611 6783
rect 17601 6749 17635 6783
rect 18889 6749 18923 6783
rect 19257 6749 19291 6783
rect 19809 6749 19843 6783
rect 6285 6681 6319 6715
rect 10762 6681 10796 6715
rect 12633 6681 12667 6715
rect 16589 6681 16623 6715
rect 20076 6681 20110 6715
rect 6745 6613 6779 6647
rect 7205 6613 7239 6647
rect 7665 6613 7699 6647
rect 9229 6613 9263 6647
rect 10241 6613 10275 6647
rect 12173 6613 12207 6647
rect 13645 6613 13679 6647
rect 14289 6613 14323 6647
rect 15485 6613 15519 6647
rect 15945 6613 15979 6647
rect 16221 6613 16255 6647
rect 16681 6613 16715 6647
rect 17509 6613 17543 6647
rect 17969 6613 18003 6647
rect 19441 6613 19475 6647
rect 21189 6613 21223 6647
rect 9597 6409 9631 6443
rect 11529 6409 11563 6443
rect 13829 6409 13863 6443
rect 20453 6409 20487 6443
rect 21281 6409 21315 6443
rect 7297 6341 7331 6375
rect 8462 6341 8496 6375
rect 11897 6341 11931 6375
rect 6377 6273 6411 6307
rect 6837 6273 6871 6307
rect 7941 6273 7975 6307
rect 10241 6273 10275 6307
rect 10517 6273 10551 6307
rect 12541 6273 12575 6307
rect 13461 6273 13495 6307
rect 14105 6273 14139 6307
rect 14924 6273 14958 6307
rect 16773 6273 16807 6307
rect 17029 6273 17063 6307
rect 18429 6273 18463 6307
rect 18685 6273 18719 6307
rect 20361 6273 20395 6307
rect 21097 6273 21131 6307
rect 8217 6205 8251 6239
rect 11989 6205 12023 6239
rect 12081 6205 12115 6239
rect 13185 6205 13219 6239
rect 13369 6205 13403 6239
rect 14657 6205 14691 6239
rect 20269 6205 20303 6239
rect 7021 6137 7055 6171
rect 18153 6137 18187 6171
rect 19809 6137 19843 6171
rect 6009 6069 6043 6103
rect 6561 6069 6595 6103
rect 10057 6069 10091 6103
rect 11161 6069 11195 6103
rect 12725 6069 12759 6103
rect 14289 6069 14323 6103
rect 16037 6069 16071 6103
rect 20821 6069 20855 6103
rect 5181 5865 5215 5899
rect 5641 5865 5675 5899
rect 6009 5865 6043 5899
rect 8585 5865 8619 5899
rect 8953 5865 8987 5899
rect 13093 5865 13127 5899
rect 14105 5865 14139 5899
rect 17693 5865 17727 5899
rect 20637 5865 20671 5899
rect 10149 5797 10183 5831
rect 9505 5729 9539 5763
rect 14749 5729 14783 5763
rect 18245 5729 18279 5763
rect 6929 5661 6963 5695
rect 7205 5661 7239 5695
rect 9965 5661 9999 5695
rect 12173 5661 12207 5695
rect 12449 5661 12483 5695
rect 13461 5661 13495 5695
rect 15117 5661 15151 5695
rect 15669 5661 15703 5695
rect 18889 5661 18923 5695
rect 19257 5661 19291 5695
rect 20913 5661 20947 5695
rect 6285 5593 6319 5627
rect 7450 5593 7484 5627
rect 17417 5593 17451 5627
rect 19524 5593 19558 5627
rect 4813 5525 4847 5559
rect 9321 5525 9355 5559
rect 9413 5525 9447 5559
rect 10885 5525 10919 5559
rect 13645 5525 13679 5559
rect 14473 5525 14507 5559
rect 14565 5525 14599 5559
rect 15301 5525 15335 5559
rect 18061 5525 18095 5559
rect 18153 5525 18187 5559
rect 18705 5525 18739 5559
rect 21097 5525 21131 5559
rect 6009 5321 6043 5355
rect 6929 5321 6963 5355
rect 9781 5321 9815 5355
rect 12265 5321 12299 5355
rect 13921 5321 13955 5355
rect 18337 5321 18371 5355
rect 20361 5321 20395 5355
rect 20729 5321 20763 5355
rect 6469 5253 6503 5287
rect 14381 5253 14415 5287
rect 16046 5253 16080 5287
rect 18797 5253 18831 5287
rect 5365 5185 5399 5219
rect 6745 5185 6779 5219
rect 8329 5185 8363 5219
rect 8585 5185 8619 5219
rect 9505 5185 9539 5219
rect 10905 5185 10939 5219
rect 11161 5185 11195 5219
rect 11989 5185 12023 5219
rect 13389 5185 13423 5219
rect 13645 5185 13679 5219
rect 14289 5185 14323 5219
rect 16313 5185 16347 5219
rect 17049 5185 17083 5219
rect 17693 5185 17727 5219
rect 18705 5185 18739 5219
rect 19717 5185 19751 5219
rect 8861 5117 8895 5151
rect 14565 5117 14599 5151
rect 16773 5117 16807 5151
rect 16957 5117 16991 5151
rect 18889 5117 18923 5151
rect 19533 5117 19567 5151
rect 19625 5117 19659 5151
rect 20821 5117 20855 5151
rect 21005 5117 21039 5151
rect 3617 5049 3651 5083
rect 5549 5049 5583 5083
rect 11805 5049 11839 5083
rect 17417 5049 17451 5083
rect 1409 4981 1443 5015
rect 4261 4981 4295 5015
rect 4997 4981 5031 5015
rect 7205 4981 7239 5015
rect 14933 4981 14967 5015
rect 17877 4981 17911 5015
rect 20085 4981 20119 5015
rect 3985 4777 4019 4811
rect 5181 4777 5215 4811
rect 5641 4777 5675 4811
rect 8585 4777 8619 4811
rect 9045 4777 9079 4811
rect 14749 4777 14783 4811
rect 15761 4777 15795 4811
rect 18889 4777 18923 4811
rect 20545 4777 20579 4811
rect 7021 4641 7055 4675
rect 7941 4641 7975 4675
rect 12357 4641 12391 4675
rect 15209 4641 15243 4675
rect 16313 4641 16347 4675
rect 17233 4641 17267 4675
rect 18245 4641 18279 4675
rect 19625 4641 19659 4675
rect 21005 4641 21039 4675
rect 21189 4641 21223 4675
rect 4721 4573 4755 4607
rect 4997 4573 5031 4607
rect 5457 4573 5491 4607
rect 6561 4573 6595 4607
rect 7205 4573 7239 4607
rect 8217 4573 8251 4607
rect 9505 4573 9539 4607
rect 10894 4573 10928 4607
rect 11161 4573 11195 4607
rect 12081 4573 12115 4607
rect 14105 4573 14139 4607
rect 16497 4573 16531 4607
rect 2053 4505 2087 4539
rect 4353 4505 4387 4539
rect 7113 4505 7147 4539
rect 11437 4505 11471 4539
rect 12602 4505 12636 4539
rect 18429 4505 18463 4539
rect 19901 4505 19935 4539
rect 1777 4437 1811 4471
rect 2605 4437 2639 4471
rect 3065 4437 3099 4471
rect 3433 4437 3467 4471
rect 5917 4437 5951 4471
rect 7573 4437 7607 4471
rect 8125 4437 8159 4471
rect 9321 4437 9355 4471
rect 9781 4437 9815 4471
rect 13737 4437 13771 4471
rect 15301 4437 15335 4471
rect 15393 4437 15427 4471
rect 16405 4437 16439 4471
rect 16865 4437 16899 4471
rect 17417 4437 17451 4471
rect 17509 4437 17543 4471
rect 17877 4437 17911 4471
rect 18521 4437 18555 4471
rect 19809 4437 19843 4471
rect 20269 4437 20303 4471
rect 20913 4437 20947 4471
rect 6745 4233 6779 4267
rect 18337 4233 18371 4267
rect 6009 4165 6043 4199
rect 10793 4165 10827 4199
rect 11897 4165 11931 4199
rect 13277 4165 13311 4199
rect 15577 4165 15611 4199
rect 21106 4165 21140 4199
rect 4445 4097 4479 4131
rect 4905 4097 4939 4131
rect 5365 4097 5399 4131
rect 7021 4097 7055 4131
rect 7665 4097 7699 4131
rect 8197 4097 8231 4131
rect 9873 4097 9907 4131
rect 11805 4097 11839 4131
rect 13921 4097 13955 4131
rect 14933 4097 14967 4131
rect 16313 4097 16347 4131
rect 16681 4097 16715 4131
rect 16937 4097 16971 4131
rect 19450 4097 19484 4131
rect 19717 4097 19751 4131
rect 21373 4097 21407 4131
rect 2697 4029 2731 4063
rect 4169 4029 4203 4063
rect 7941 4029 7975 4063
rect 10609 4029 10643 4063
rect 10701 4029 10735 4063
rect 11713 4029 11747 4063
rect 13093 4029 13127 4063
rect 13185 4029 13219 4063
rect 15393 4029 15427 4063
rect 15485 4029 15519 4063
rect 2329 3961 2363 3995
rect 3433 3961 3467 3995
rect 5549 3961 5583 3995
rect 13645 3961 13679 3995
rect 19993 3961 20027 3995
rect 1409 3893 1443 3927
rect 1961 3893 1995 3927
rect 3065 3893 3099 3927
rect 3801 3893 3835 3927
rect 4629 3893 4663 3927
rect 5089 3893 5123 3927
rect 9321 3893 9355 3927
rect 10057 3893 10091 3927
rect 11161 3893 11195 3927
rect 12265 3893 12299 3927
rect 12633 3893 12667 3927
rect 14565 3893 14599 3927
rect 15945 3893 15979 3927
rect 18061 3893 18095 3927
rect 1593 3689 1627 3723
rect 3433 3689 3467 3723
rect 5733 3689 5767 3723
rect 8953 3689 8987 3723
rect 11437 3689 11471 3723
rect 14565 3689 14599 3723
rect 16221 3689 16255 3723
rect 6929 3621 6963 3655
rect 11989 3621 12023 3655
rect 14289 3621 14323 3655
rect 3893 3553 3927 3587
rect 7941 3553 7975 3587
rect 9505 3553 9539 3587
rect 15945 3553 15979 3587
rect 16773 3553 16807 3587
rect 17693 3553 17727 3587
rect 17877 3553 17911 3587
rect 20821 3553 20855 3587
rect 1409 3485 1443 3519
rect 3065 3485 3099 3519
rect 4169 3485 4203 3519
rect 4629 3485 4663 3519
rect 5089 3485 5123 3519
rect 5549 3485 5583 3519
rect 6469 3485 6503 3519
rect 7573 3485 7607 3519
rect 8125 3485 8159 3519
rect 9321 3485 9355 3519
rect 10057 3485 10091 3519
rect 11805 3485 11839 3519
rect 13737 3485 13771 3519
rect 14105 3485 14139 3519
rect 18245 3485 18279 3519
rect 19441 3485 19475 3519
rect 19717 3485 19751 3519
rect 20545 3485 20579 3519
rect 2697 3417 2731 3451
rect 8217 3417 8251 3451
rect 10302 3417 10336 3451
rect 13492 3417 13526 3451
rect 15700 3417 15734 3451
rect 16589 3417 16623 3451
rect 18889 3417 18923 3451
rect 1961 3349 1995 3383
rect 2329 3349 2363 3383
rect 4353 3349 4387 3383
rect 4813 3349 4847 3383
rect 5273 3349 5307 3383
rect 6193 3349 6227 3383
rect 6653 3349 6687 3383
rect 8585 3349 8619 3383
rect 9413 3349 9447 3383
rect 12357 3349 12391 3383
rect 16681 3349 16715 3383
rect 17233 3349 17267 3383
rect 17601 3349 17635 3383
rect 1593 3145 1627 3179
rect 2053 3145 2087 3179
rect 2513 3145 2547 3179
rect 2973 3145 3007 3179
rect 4629 3145 4663 3179
rect 6837 3145 6871 3179
rect 9781 3145 9815 3179
rect 13461 3145 13495 3179
rect 13737 3145 13771 3179
rect 14197 3145 14231 3179
rect 14841 3145 14875 3179
rect 16681 3145 16715 3179
rect 17049 3145 17083 3179
rect 18337 3145 18371 3179
rect 18705 3145 18739 3179
rect 6009 3077 6043 3111
rect 10916 3077 10950 3111
rect 12348 3077 12382 3111
rect 15954 3077 15988 3111
rect 18797 3077 18831 3111
rect 1409 3009 1443 3043
rect 1869 3009 1903 3043
rect 2329 3009 2363 3043
rect 2789 3009 2823 3043
rect 3525 3009 3559 3043
rect 3985 3009 4019 3043
rect 4445 3009 4479 3043
rect 4905 3009 4939 3043
rect 5365 3009 5399 3043
rect 6377 3009 6411 3043
rect 7481 3009 7515 3043
rect 8013 3009 8047 3043
rect 9505 3009 9539 3043
rect 11161 3009 11195 3043
rect 11529 3009 11563 3043
rect 14105 3009 14139 3043
rect 16221 3009 16255 3043
rect 17693 3009 17727 3043
rect 19717 3009 19751 3043
rect 20545 3009 20579 3043
rect 20821 3009 20855 3043
rect 7757 2941 7791 2975
rect 12081 2941 12115 2975
rect 14289 2941 14323 2975
rect 17141 2941 17175 2975
rect 17233 2941 17267 2975
rect 18981 2941 19015 2975
rect 19441 2941 19475 2975
rect 3709 2873 3743 2907
rect 4169 2873 4203 2907
rect 6561 2873 6595 2907
rect 5089 2805 5123 2839
rect 5549 2805 5583 2839
rect 9137 2805 9171 2839
rect 11713 2805 11747 2839
rect 17877 2805 17911 2839
rect 3433 2601 3467 2635
rect 6469 2601 6503 2635
rect 6929 2601 6963 2635
rect 7205 2601 7239 2635
rect 8953 2601 8987 2635
rect 11161 2601 11195 2635
rect 13185 2601 13219 2635
rect 15669 2601 15703 2635
rect 16681 2601 16715 2635
rect 5365 2533 5399 2567
rect 10149 2533 10183 2567
rect 13553 2533 13587 2567
rect 17049 2533 17083 2567
rect 9505 2465 9539 2499
rect 10517 2465 10551 2499
rect 10701 2465 10735 2499
rect 12541 2465 12575 2499
rect 15117 2465 15151 2499
rect 17509 2465 17543 2499
rect 17693 2465 17727 2499
rect 18613 2465 18647 2499
rect 19717 2465 19751 2499
rect 2329 2397 2363 2431
rect 2789 2397 2823 2431
rect 3249 2397 3283 2431
rect 3985 2397 4019 2431
rect 4445 2397 4479 2431
rect 4905 2397 4939 2431
rect 6009 2397 6043 2431
rect 6745 2397 6779 2431
rect 8585 2397 8619 2431
rect 9413 2397 9447 2431
rect 9965 2397 9999 2431
rect 11529 2397 11563 2431
rect 13737 2397 13771 2431
rect 14381 2397 14415 2431
rect 15945 2397 15979 2431
rect 18889 2397 18923 2431
rect 19441 2397 19475 2431
rect 20545 2397 20579 2431
rect 20821 2397 20855 2431
rect 1685 2329 1719 2363
rect 8340 2329 8374 2363
rect 12173 2329 12207 2363
rect 15209 2329 15243 2363
rect 1777 2261 1811 2295
rect 2513 2261 2547 2295
rect 2973 2261 3007 2295
rect 4169 2261 4203 2295
rect 4629 2261 4663 2295
rect 5089 2261 5123 2295
rect 9321 2261 9355 2295
rect 10793 2261 10827 2295
rect 12725 2261 12759 2295
rect 12817 2261 12851 2295
rect 14197 2261 14231 2295
rect 15301 2261 15335 2295
rect 16129 2261 16163 2295
rect 17417 2261 17451 2295
<< metal1 >>
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 19613 20587 19671 20593
rect 19613 20553 19625 20587
rect 19659 20584 19671 20587
rect 19702 20584 19708 20596
rect 19659 20556 19708 20584
rect 19659 20553 19671 20556
rect 19613 20547 19671 20553
rect 19702 20544 19708 20556
rect 19760 20544 19766 20596
rect 18785 20519 18843 20525
rect 18785 20485 18797 20519
rect 18831 20516 18843 20519
rect 19242 20516 19248 20528
rect 18831 20488 19248 20516
rect 18831 20485 18843 20488
rect 18785 20479 18843 20485
rect 19242 20476 19248 20488
rect 19300 20516 19306 20528
rect 20165 20519 20223 20525
rect 20165 20516 20177 20519
rect 19300 20488 20177 20516
rect 19300 20476 19306 20488
rect 20165 20485 20177 20488
rect 20211 20485 20223 20519
rect 20165 20479 20223 20485
rect 5718 20408 5724 20460
rect 5776 20448 5782 20460
rect 5813 20451 5871 20457
rect 5813 20448 5825 20451
rect 5776 20420 5825 20448
rect 5776 20408 5782 20420
rect 5813 20417 5825 20420
rect 5859 20448 5871 20451
rect 6365 20451 6423 20457
rect 6365 20448 6377 20451
rect 5859 20420 6377 20448
rect 5859 20417 5871 20420
rect 5813 20411 5871 20417
rect 6365 20417 6377 20420
rect 6411 20417 6423 20451
rect 6365 20411 6423 20417
rect 17218 20408 17224 20460
rect 17276 20448 17282 20460
rect 17497 20451 17555 20457
rect 17497 20448 17509 20451
rect 17276 20420 17509 20448
rect 17276 20408 17282 20420
rect 17497 20417 17509 20420
rect 17543 20448 17555 20451
rect 17773 20451 17831 20457
rect 17773 20448 17785 20451
rect 17543 20420 17785 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 17773 20417 17785 20420
rect 17819 20417 17831 20451
rect 17773 20411 17831 20417
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19429 20451 19487 20457
rect 19429 20448 19441 20451
rect 18932 20420 19441 20448
rect 18932 20408 18938 20420
rect 19429 20417 19441 20420
rect 19475 20417 19487 20451
rect 20530 20448 20536 20460
rect 20491 20420 20536 20448
rect 19429 20411 19487 20417
rect 20530 20408 20536 20420
rect 20588 20408 20594 20460
rect 21082 20448 21088 20460
rect 21043 20420 21088 20448
rect 21082 20408 21088 20420
rect 21140 20408 21146 20460
rect 5994 20244 6000 20256
rect 5955 20216 6000 20244
rect 5994 20204 6000 20216
rect 6052 20204 6058 20256
rect 17310 20244 17316 20256
rect 17271 20216 17316 20244
rect 17310 20204 17316 20216
rect 17368 20204 17374 20256
rect 20073 20247 20131 20253
rect 20073 20213 20085 20247
rect 20119 20244 20131 20247
rect 20162 20244 20168 20256
rect 20119 20216 20168 20244
rect 20119 20213 20131 20216
rect 20073 20207 20131 20213
rect 20162 20204 20168 20216
rect 20220 20204 20226 20256
rect 20714 20244 20720 20256
rect 20675 20216 20720 20244
rect 20714 20204 20720 20216
rect 20772 20204 20778 20256
rect 21269 20247 21327 20253
rect 21269 20213 21281 20247
rect 21315 20244 21327 20247
rect 21358 20244 21364 20256
rect 21315 20216 21364 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 18874 20040 18880 20052
rect 18835 20012 18880 20040
rect 18874 20000 18880 20012
rect 18932 20000 18938 20052
rect 20165 20043 20223 20049
rect 20165 20009 20177 20043
rect 20211 20040 20223 20043
rect 20346 20040 20352 20052
rect 20211 20012 20352 20040
rect 20211 20009 20223 20012
rect 20165 20003 20223 20009
rect 20346 20000 20352 20012
rect 20404 20000 20410 20052
rect 20717 20043 20775 20049
rect 20717 20009 20729 20043
rect 20763 20040 20775 20043
rect 20806 20040 20812 20052
rect 20763 20012 20812 20040
rect 20763 20009 20775 20012
rect 20717 20003 20775 20009
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 13081 19975 13139 19981
rect 13081 19941 13093 19975
rect 13127 19972 13139 19975
rect 13127 19944 16574 19972
rect 13127 19941 13139 19944
rect 13081 19935 13139 19941
rect 16546 19904 16574 19944
rect 16546 19876 20576 19904
rect 5994 19796 6000 19848
rect 6052 19836 6058 19848
rect 6365 19839 6423 19845
rect 6365 19836 6377 19839
rect 6052 19808 6377 19836
rect 6052 19796 6058 19808
rect 6365 19805 6377 19808
rect 6411 19805 6423 19839
rect 12894 19836 12900 19848
rect 12855 19808 12900 19836
rect 6365 19799 6423 19805
rect 12894 19796 12900 19808
rect 12952 19796 12958 19848
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19805 18751 19839
rect 19518 19836 19524 19848
rect 19479 19808 19524 19836
rect 18693 19799 18751 19805
rect 6546 19768 6552 19780
rect 6507 19740 6552 19768
rect 6546 19728 6552 19740
rect 6604 19728 6610 19780
rect 18708 19768 18736 19799
rect 19518 19796 19524 19808
rect 19576 19796 19582 19848
rect 20548 19845 20576 19876
rect 19981 19839 20039 19845
rect 19981 19805 19993 19839
rect 20027 19805 20039 19839
rect 19981 19799 20039 19805
rect 20533 19839 20591 19845
rect 20533 19805 20545 19839
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 19886 19768 19892 19780
rect 18708 19740 19892 19768
rect 19886 19728 19892 19740
rect 19944 19728 19950 19780
rect 19705 19703 19763 19709
rect 19705 19669 19717 19703
rect 19751 19700 19763 19703
rect 19996 19700 20024 19799
rect 20806 19796 20812 19848
rect 20864 19836 20870 19848
rect 21085 19839 21143 19845
rect 21085 19836 21097 19839
rect 20864 19808 21097 19836
rect 20864 19796 20870 19808
rect 21085 19805 21097 19808
rect 21131 19805 21143 19839
rect 21085 19799 21143 19805
rect 21266 19700 21272 19712
rect 19751 19672 20024 19700
rect 21227 19672 21272 19700
rect 19751 19669 19763 19672
rect 19705 19663 19763 19669
rect 21266 19660 21272 19672
rect 21324 19660 21330 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 19518 19456 19524 19508
rect 19576 19496 19582 19508
rect 19705 19499 19763 19505
rect 19705 19496 19717 19499
rect 19576 19468 19717 19496
rect 19576 19456 19582 19468
rect 19705 19465 19717 19468
rect 19751 19465 19763 19499
rect 19705 19459 19763 19465
rect 19886 19456 19892 19508
rect 19944 19496 19950 19508
rect 19981 19499 20039 19505
rect 19981 19496 19993 19499
rect 19944 19468 19993 19496
rect 19944 19456 19950 19468
rect 19981 19465 19993 19468
rect 20027 19465 20039 19499
rect 19981 19459 20039 19465
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 21269 19499 21327 19505
rect 21269 19496 21281 19499
rect 20680 19468 21281 19496
rect 20680 19456 20686 19468
rect 21269 19465 21281 19468
rect 21315 19465 21327 19499
rect 21269 19459 21327 19465
rect 16206 19388 16212 19440
rect 16264 19428 16270 19440
rect 16264 19400 20208 19428
rect 16264 19388 16270 19400
rect 18414 19360 18420 19372
rect 18375 19332 18420 19360
rect 18414 19320 18420 19332
rect 18472 19320 18478 19372
rect 19061 19363 19119 19369
rect 19061 19360 19073 19363
rect 18616 19332 19073 19360
rect 18616 19233 18644 19332
rect 19061 19329 19073 19332
rect 19107 19329 19119 19363
rect 19518 19360 19524 19372
rect 19479 19332 19524 19360
rect 19061 19323 19119 19329
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 20180 19369 20208 19400
rect 20438 19388 20444 19440
rect 20496 19428 20502 19440
rect 20496 19400 20668 19428
rect 20496 19388 20502 19400
rect 20165 19363 20223 19369
rect 20165 19329 20177 19363
rect 20211 19329 20223 19363
rect 20533 19363 20591 19369
rect 20533 19360 20545 19363
rect 20165 19323 20223 19329
rect 20272 19332 20545 19360
rect 20272 19292 20300 19332
rect 20533 19329 20545 19332
rect 20579 19329 20591 19363
rect 20533 19323 20591 19329
rect 19260 19264 20300 19292
rect 19260 19233 19288 19264
rect 18601 19227 18659 19233
rect 18601 19193 18613 19227
rect 18647 19193 18659 19227
rect 18601 19187 18659 19193
rect 19245 19227 19303 19233
rect 19245 19193 19257 19227
rect 19291 19193 19303 19227
rect 20640 19224 20668 19400
rect 20714 19320 20720 19372
rect 20772 19360 20778 19372
rect 21085 19363 21143 19369
rect 21085 19360 21097 19363
rect 20772 19332 21097 19360
rect 20772 19320 20778 19332
rect 21085 19329 21097 19332
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 20717 19227 20775 19233
rect 20717 19224 20729 19227
rect 20640 19196 20729 19224
rect 19245 19187 19303 19193
rect 20717 19193 20729 19196
rect 20763 19193 20775 19227
rect 20717 19187 20775 19193
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 12161 18955 12219 18961
rect 12161 18921 12173 18955
rect 12207 18952 12219 18955
rect 12894 18952 12900 18964
rect 12207 18924 12900 18952
rect 12207 18921 12219 18924
rect 12161 18915 12219 18921
rect 12894 18912 12900 18924
rect 12952 18912 12958 18964
rect 20349 18955 20407 18961
rect 20349 18921 20361 18955
rect 20395 18952 20407 18955
rect 20530 18952 20536 18964
rect 20395 18924 20536 18952
rect 20395 18921 20407 18924
rect 20349 18915 20407 18921
rect 20530 18912 20536 18924
rect 20588 18912 20594 18964
rect 20809 18955 20867 18961
rect 20809 18921 20821 18955
rect 20855 18952 20867 18955
rect 21082 18952 21088 18964
rect 20855 18924 21088 18952
rect 20855 18921 20867 18924
rect 20809 18915 20867 18921
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 9493 18751 9551 18757
rect 9493 18717 9505 18751
rect 9539 18748 9551 18751
rect 9766 18748 9772 18760
rect 9539 18720 9772 18748
rect 9539 18717 9551 18720
rect 9493 18711 9551 18717
rect 9766 18708 9772 18720
rect 9824 18708 9830 18760
rect 11238 18708 11244 18760
rect 11296 18748 11302 18760
rect 11977 18751 12035 18757
rect 11977 18748 11989 18751
rect 11296 18720 11989 18748
rect 11296 18708 11302 18720
rect 11977 18717 11989 18720
rect 12023 18717 12035 18751
rect 20165 18751 20223 18757
rect 20165 18748 20177 18751
rect 11977 18711 12035 18717
rect 16546 18720 20177 18748
rect 9677 18615 9735 18621
rect 9677 18581 9689 18615
rect 9723 18612 9735 18615
rect 16546 18612 16574 18720
rect 20165 18717 20177 18720
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 20254 18708 20260 18760
rect 20312 18748 20318 18760
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 20312 18720 20637 18748
rect 20312 18708 20318 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 20990 18708 20996 18760
rect 21048 18748 21054 18760
rect 21085 18751 21143 18757
rect 21085 18748 21097 18751
rect 21048 18720 21097 18748
rect 21048 18708 21054 18720
rect 21085 18717 21097 18720
rect 21131 18717 21143 18751
rect 21085 18711 21143 18717
rect 21266 18612 21272 18624
rect 9723 18584 16574 18612
rect 21227 18584 21272 18612
rect 9723 18581 9735 18584
rect 9677 18575 9735 18581
rect 21266 18572 21272 18584
rect 21324 18572 21330 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 12437 18411 12495 18417
rect 12437 18377 12449 18411
rect 12483 18408 12495 18411
rect 20806 18408 20812 18420
rect 12483 18380 20812 18408
rect 12483 18377 12495 18380
rect 12437 18371 12495 18377
rect 20806 18368 20812 18380
rect 20864 18368 20870 18420
rect 8389 18275 8447 18281
rect 8389 18241 8401 18275
rect 8435 18272 8447 18275
rect 8570 18272 8576 18284
rect 8435 18244 8576 18272
rect 8435 18241 8447 18244
rect 8389 18235 8447 18241
rect 8570 18232 8576 18244
rect 8628 18232 8634 18284
rect 12250 18272 12256 18284
rect 12211 18244 12256 18272
rect 12250 18232 12256 18244
rect 12308 18232 12314 18284
rect 20806 18272 20812 18284
rect 20767 18244 20812 18272
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 20898 18232 20904 18284
rect 20956 18272 20962 18284
rect 21085 18275 21143 18281
rect 21085 18272 21097 18275
rect 20956 18244 21097 18272
rect 20956 18232 20962 18244
rect 21085 18241 21097 18244
rect 21131 18241 21143 18275
rect 21085 18235 21143 18241
rect 8573 18139 8631 18145
rect 8573 18105 8585 18139
rect 8619 18136 8631 18139
rect 8619 18108 16574 18136
rect 8619 18105 8631 18108
rect 8573 18099 8631 18105
rect 16546 18068 16574 18108
rect 20254 18068 20260 18080
rect 16546 18040 20260 18068
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20530 18028 20536 18080
rect 20588 18068 20594 18080
rect 20625 18071 20683 18077
rect 20625 18068 20637 18071
rect 20588 18040 20637 18068
rect 20588 18028 20594 18040
rect 20625 18037 20637 18040
rect 20671 18037 20683 18071
rect 20625 18031 20683 18037
rect 21269 18071 21327 18077
rect 21269 18037 21281 18071
rect 21315 18068 21327 18071
rect 21358 18068 21364 18080
rect 21315 18040 21364 18068
rect 21315 18037 21327 18040
rect 21269 18031 21327 18037
rect 21358 18028 21364 18040
rect 21416 18028 21422 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 11609 17867 11667 17873
rect 11609 17833 11621 17867
rect 11655 17864 11667 17867
rect 12250 17864 12256 17876
rect 11655 17836 12256 17864
rect 11655 17833 11667 17836
rect 11609 17827 11667 17833
rect 12250 17824 12256 17836
rect 12308 17824 12314 17876
rect 20257 17867 20315 17873
rect 20257 17833 20269 17867
rect 20303 17864 20315 17867
rect 20714 17864 20720 17876
rect 20303 17836 20720 17864
rect 20303 17833 20315 17836
rect 20257 17827 20315 17833
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17660 11483 17663
rect 12250 17660 12256 17672
rect 11471 17632 12256 17660
rect 11471 17629 11483 17632
rect 11425 17623 11483 17629
rect 12250 17620 12256 17632
rect 12308 17620 12314 17672
rect 20070 17660 20076 17672
rect 20031 17632 20076 17660
rect 20070 17620 20076 17632
rect 20128 17620 20134 17672
rect 20530 17660 20536 17672
rect 20491 17632 20536 17660
rect 20530 17620 20536 17632
rect 20588 17620 20594 17672
rect 21082 17660 21088 17672
rect 21043 17632 21088 17660
rect 21082 17620 21088 17632
rect 21140 17620 21146 17672
rect 20714 17524 20720 17536
rect 20675 17496 20720 17524
rect 20714 17484 20720 17496
rect 20772 17484 20778 17536
rect 21266 17524 21272 17536
rect 21227 17496 21272 17524
rect 21266 17484 21272 17496
rect 21324 17484 21330 17536
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 20070 17320 20076 17332
rect 20031 17292 20076 17320
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 20809 17323 20867 17329
rect 20809 17289 20821 17323
rect 20855 17320 20867 17323
rect 20898 17320 20904 17332
rect 20855 17292 20904 17320
rect 20855 17289 20867 17292
rect 20809 17283 20867 17289
rect 20898 17280 20904 17292
rect 20956 17280 20962 17332
rect 15102 17212 15108 17264
rect 15160 17252 15166 17264
rect 19518 17252 19524 17264
rect 15160 17224 19524 17252
rect 15160 17212 15166 17224
rect 19518 17212 19524 17224
rect 19576 17212 19582 17264
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 19889 17187 19947 17193
rect 19889 17184 19901 17187
rect 14332 17156 19901 17184
rect 14332 17144 14338 17156
rect 19889 17153 19901 17156
rect 19935 17153 19947 17187
rect 19889 17147 19947 17153
rect 20625 17187 20683 17193
rect 20625 17153 20637 17187
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 20640 17116 20668 17147
rect 20806 17144 20812 17196
rect 20864 17184 20870 17196
rect 21085 17187 21143 17193
rect 21085 17184 21097 17187
rect 20864 17156 21097 17184
rect 20864 17144 20870 17156
rect 21085 17153 21097 17156
rect 21131 17153 21143 17187
rect 21085 17147 21143 17153
rect 18012 17088 20668 17116
rect 18012 17076 18018 17088
rect 21269 16983 21327 16989
rect 21269 16949 21281 16983
rect 21315 16980 21327 16983
rect 21358 16980 21364 16992
rect 21315 16952 21364 16980
rect 21315 16949 21327 16952
rect 21269 16943 21327 16949
rect 21358 16940 21364 16952
rect 21416 16940 21422 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 20809 16779 20867 16785
rect 20809 16745 20821 16779
rect 20855 16776 20867 16779
rect 21082 16776 21088 16788
rect 20855 16748 21088 16776
rect 20855 16745 20867 16748
rect 20809 16739 20867 16745
rect 21082 16736 21088 16748
rect 21140 16736 21146 16788
rect 20088 16612 20300 16640
rect 18230 16572 18236 16584
rect 18191 16544 18236 16572
rect 18230 16532 18236 16544
rect 18288 16532 18294 16584
rect 15194 16464 15200 16516
rect 15252 16504 15258 16516
rect 20088 16504 20116 16612
rect 20165 16575 20223 16581
rect 20165 16541 20177 16575
rect 20211 16541 20223 16575
rect 20272 16572 20300 16612
rect 20625 16575 20683 16581
rect 20625 16572 20637 16575
rect 20272 16544 20637 16572
rect 20165 16535 20223 16541
rect 20625 16541 20637 16544
rect 20671 16541 20683 16575
rect 20625 16535 20683 16541
rect 15252 16476 20116 16504
rect 15252 16464 15258 16476
rect 18417 16439 18475 16445
rect 18417 16405 18429 16439
rect 18463 16436 18475 16439
rect 20180 16436 20208 16535
rect 20898 16532 20904 16584
rect 20956 16572 20962 16584
rect 21085 16575 21143 16581
rect 21085 16572 21097 16575
rect 20956 16544 21097 16572
rect 20956 16532 20962 16544
rect 21085 16541 21097 16544
rect 21131 16541 21143 16575
rect 21085 16535 21143 16541
rect 18463 16408 20208 16436
rect 20349 16439 20407 16445
rect 18463 16405 18475 16408
rect 18417 16399 18475 16405
rect 20349 16405 20361 16439
rect 20395 16436 20407 16439
rect 20990 16436 20996 16448
rect 20395 16408 20996 16436
rect 20395 16405 20407 16408
rect 20349 16399 20407 16405
rect 20990 16396 20996 16408
rect 21048 16396 21054 16448
rect 21266 16436 21272 16448
rect 21227 16408 21272 16436
rect 21266 16396 21272 16408
rect 21324 16396 21330 16448
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 14737 16235 14795 16241
rect 14737 16201 14749 16235
rect 14783 16232 14795 16235
rect 17954 16232 17960 16244
rect 14783 16204 17960 16232
rect 14783 16201 14795 16204
rect 14737 16195 14795 16201
rect 17954 16192 17960 16204
rect 18012 16192 18018 16244
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16232 20223 16235
rect 20622 16232 20628 16244
rect 20211 16204 20628 16232
rect 20211 16201 20223 16204
rect 20165 16195 20223 16201
rect 20622 16192 20628 16204
rect 20680 16192 20686 16244
rect 20806 16232 20812 16244
rect 20767 16204 20812 16232
rect 20806 16192 20812 16204
rect 20864 16192 20870 16244
rect 14458 16056 14464 16108
rect 14516 16096 14522 16108
rect 14553 16099 14611 16105
rect 14553 16096 14565 16099
rect 14516 16068 14565 16096
rect 14516 16056 14522 16068
rect 14553 16065 14565 16068
rect 14599 16065 14611 16099
rect 14553 16059 14611 16065
rect 17862 16056 17868 16108
rect 17920 16096 17926 16108
rect 19981 16099 20039 16105
rect 19981 16096 19993 16099
rect 17920 16068 19993 16096
rect 17920 16056 17926 16068
rect 19981 16065 19993 16068
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20625 16099 20683 16105
rect 20625 16065 20637 16099
rect 20671 16065 20683 16099
rect 21082 16096 21088 16108
rect 21043 16068 21088 16096
rect 20625 16059 20683 16065
rect 12986 15988 12992 16040
rect 13044 16028 13050 16040
rect 20640 16028 20668 16059
rect 21082 16056 21088 16068
rect 21140 16056 21146 16108
rect 13044 16000 20668 16028
rect 13044 15988 13050 16000
rect 19610 15852 19616 15904
rect 19668 15892 19674 15904
rect 19705 15895 19763 15901
rect 19705 15892 19717 15895
rect 19668 15864 19717 15892
rect 19668 15852 19674 15864
rect 19705 15861 19717 15864
rect 19751 15892 19763 15895
rect 20070 15892 20076 15904
rect 19751 15864 20076 15892
rect 19751 15861 19763 15864
rect 19705 15855 19763 15861
rect 20070 15852 20076 15864
rect 20128 15852 20134 15904
rect 21269 15895 21327 15901
rect 21269 15861 21281 15895
rect 21315 15892 21327 15895
rect 21358 15892 21364 15904
rect 21315 15864 21364 15892
rect 21315 15861 21327 15864
rect 21269 15855 21327 15861
rect 21358 15852 21364 15864
rect 21416 15852 21422 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 20349 15691 20407 15697
rect 20349 15657 20361 15691
rect 20395 15688 20407 15691
rect 21082 15688 21088 15700
rect 20395 15660 21088 15688
rect 20395 15657 20407 15660
rect 20349 15651 20407 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 15286 15512 15292 15564
rect 15344 15552 15350 15564
rect 15344 15524 20208 15552
rect 15344 15512 15350 15524
rect 18877 15487 18935 15493
rect 18877 15453 18889 15487
rect 18923 15484 18935 15487
rect 18966 15484 18972 15496
rect 18923 15456 18972 15484
rect 18923 15453 18935 15456
rect 18877 15447 18935 15453
rect 18966 15444 18972 15456
rect 19024 15484 19030 15496
rect 20180 15493 20208 15524
rect 19705 15487 19763 15493
rect 19705 15484 19717 15487
rect 19024 15456 19717 15484
rect 19024 15444 19030 15456
rect 19705 15453 19717 15456
rect 19751 15453 19763 15487
rect 19705 15447 19763 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20346 15444 20352 15496
rect 20404 15484 20410 15496
rect 20625 15487 20683 15493
rect 20625 15484 20637 15487
rect 20404 15456 20637 15484
rect 20404 15444 20410 15456
rect 20625 15453 20637 15456
rect 20671 15453 20683 15487
rect 20625 15447 20683 15453
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 21085 15487 21143 15493
rect 21085 15484 21097 15487
rect 20772 15456 21097 15484
rect 20772 15444 20778 15456
rect 21085 15453 21097 15456
rect 21131 15453 21143 15487
rect 21085 15447 21143 15453
rect 19429 15351 19487 15357
rect 19429 15317 19441 15351
rect 19475 15348 19487 15351
rect 19702 15348 19708 15360
rect 19475 15320 19708 15348
rect 19475 15317 19487 15320
rect 19429 15311 19487 15317
rect 19702 15308 19708 15320
rect 19760 15308 19766 15360
rect 19889 15351 19947 15357
rect 19889 15317 19901 15351
rect 19935 15348 19947 15351
rect 20254 15348 20260 15360
rect 19935 15320 20260 15348
rect 19935 15317 19947 15320
rect 19889 15311 19947 15317
rect 20254 15308 20260 15320
rect 20312 15308 20318 15360
rect 20809 15351 20867 15357
rect 20809 15317 20821 15351
rect 20855 15348 20867 15351
rect 21082 15348 21088 15360
rect 20855 15320 21088 15348
rect 20855 15317 20867 15320
rect 20809 15311 20867 15317
rect 21082 15308 21088 15320
rect 21140 15308 21146 15360
rect 21266 15348 21272 15360
rect 21227 15320 21272 15348
rect 21266 15308 21272 15320
rect 21324 15308 21330 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 9493 15147 9551 15153
rect 9493 15113 9505 15147
rect 9539 15144 9551 15147
rect 12986 15144 12992 15156
rect 9539 15116 12992 15144
rect 9539 15113 9551 15116
rect 9493 15107 9551 15113
rect 12986 15104 12992 15116
rect 13044 15104 13050 15156
rect 20349 15147 20407 15153
rect 20349 15113 20361 15147
rect 20395 15144 20407 15147
rect 20714 15144 20720 15156
rect 20395 15116 20720 15144
rect 20395 15113 20407 15116
rect 20349 15107 20407 15113
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 20809 15147 20867 15153
rect 20809 15113 20821 15147
rect 20855 15113 20867 15147
rect 20809 15107 20867 15113
rect 9309 15011 9367 15017
rect 9309 14977 9321 15011
rect 9355 15008 9367 15011
rect 9490 15008 9496 15020
rect 9355 14980 9496 15008
rect 9355 14977 9367 14980
rect 9309 14971 9367 14977
rect 9490 14968 9496 14980
rect 9548 14968 9554 15020
rect 11609 15011 11667 15017
rect 11609 14977 11621 15011
rect 11655 15008 11667 15011
rect 11698 15008 11704 15020
rect 11655 14980 11704 15008
rect 11655 14977 11667 14980
rect 11609 14971 11667 14977
rect 11698 14968 11704 14980
rect 11756 14968 11762 15020
rect 19245 15011 19303 15017
rect 19245 14977 19257 15011
rect 19291 15008 19303 15011
rect 19610 15008 19616 15020
rect 19291 14980 19616 15008
rect 19291 14977 19303 14980
rect 19245 14971 19303 14977
rect 19610 14968 19616 14980
rect 19668 14968 19674 15020
rect 19705 15011 19763 15017
rect 19705 14977 19717 15011
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 18877 14943 18935 14949
rect 18877 14909 18889 14943
rect 18923 14940 18935 14943
rect 19058 14940 19064 14952
rect 18923 14912 19064 14940
rect 18923 14909 18935 14912
rect 18877 14903 18935 14909
rect 19058 14900 19064 14912
rect 19116 14900 19122 14952
rect 11793 14875 11851 14881
rect 11793 14841 11805 14875
rect 11839 14872 11851 14875
rect 15194 14872 15200 14884
rect 11839 14844 15200 14872
rect 11839 14841 11851 14844
rect 11793 14835 11851 14841
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 17126 14832 17132 14884
rect 17184 14872 17190 14884
rect 19720 14872 19748 14971
rect 19978 14968 19984 15020
rect 20036 15008 20042 15020
rect 20165 15011 20223 15017
rect 20165 15008 20177 15011
rect 20036 14980 20177 15008
rect 20036 14968 20042 14980
rect 20165 14977 20177 14980
rect 20211 14977 20223 15011
rect 20622 15008 20628 15020
rect 20583 14980 20628 15008
rect 20165 14971 20223 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 20824 15008 20852 15107
rect 21085 15011 21143 15017
rect 21085 15008 21097 15011
rect 20824 14980 21097 15008
rect 21085 14977 21097 14980
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 17184 14844 19748 14872
rect 19889 14875 19947 14881
rect 17184 14832 17190 14844
rect 19889 14841 19901 14875
rect 19935 14872 19947 14875
rect 20898 14872 20904 14884
rect 19935 14844 20904 14872
rect 19935 14841 19947 14844
rect 19889 14835 19947 14841
rect 20898 14832 20904 14844
rect 20956 14832 20962 14884
rect 17954 14764 17960 14816
rect 18012 14804 18018 14816
rect 18233 14807 18291 14813
rect 18233 14804 18245 14807
rect 18012 14776 18245 14804
rect 18012 14764 18018 14776
rect 18233 14773 18245 14776
rect 18279 14773 18291 14807
rect 18233 14767 18291 14773
rect 19429 14807 19487 14813
rect 19429 14773 19441 14807
rect 19475 14804 19487 14807
rect 19794 14804 19800 14816
rect 19475 14776 19800 14804
rect 19475 14773 19487 14776
rect 19429 14767 19487 14773
rect 19794 14764 19800 14776
rect 19852 14764 19858 14816
rect 21266 14804 21272 14816
rect 21227 14776 21272 14804
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 15470 14560 15476 14612
rect 15528 14600 15534 14612
rect 20073 14603 20131 14609
rect 15528 14572 18736 14600
rect 15528 14560 15534 14572
rect 17957 14535 18015 14541
rect 17957 14501 17969 14535
rect 18003 14501 18015 14535
rect 17957 14495 18015 14501
rect 17972 14464 18000 14495
rect 18046 14492 18052 14544
rect 18104 14532 18110 14544
rect 18598 14532 18604 14544
rect 18104 14504 18604 14532
rect 18104 14492 18110 14504
rect 18598 14492 18604 14504
rect 18656 14492 18662 14544
rect 17972 14436 18644 14464
rect 8662 14356 8668 14408
rect 8720 14396 8726 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 8720 14368 8953 14396
rect 8720 14356 8726 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 17497 14399 17555 14405
rect 17497 14365 17509 14399
rect 17543 14396 17555 14399
rect 17773 14399 17831 14405
rect 17773 14396 17785 14399
rect 17543 14368 17785 14396
rect 17543 14365 17555 14368
rect 17497 14359 17555 14365
rect 17773 14365 17785 14368
rect 17819 14396 17831 14399
rect 18046 14396 18052 14408
rect 17819 14368 18052 14396
rect 17819 14365 17831 14368
rect 17773 14359 17831 14365
rect 18046 14356 18052 14368
rect 18104 14356 18110 14408
rect 18138 14356 18144 14408
rect 18196 14396 18202 14408
rect 18417 14399 18475 14405
rect 18417 14396 18429 14399
rect 18196 14368 18429 14396
rect 18196 14356 18202 14368
rect 18417 14365 18429 14368
rect 18463 14365 18475 14399
rect 18417 14359 18475 14365
rect 17126 14328 17132 14340
rect 9140 14300 17132 14328
rect 9140 14269 9168 14300
rect 17126 14288 17132 14300
rect 17184 14288 17190 14340
rect 18616 14328 18644 14436
rect 18708 14405 18736 14572
rect 20073 14569 20085 14603
rect 20119 14600 20131 14603
rect 20622 14600 20628 14612
rect 20119 14572 20628 14600
rect 20119 14569 20131 14572
rect 20073 14563 20131 14569
rect 20622 14560 20628 14572
rect 20680 14560 20686 14612
rect 19610 14492 19616 14544
rect 19668 14532 19674 14544
rect 20349 14535 20407 14541
rect 20349 14532 20361 14535
rect 19668 14504 20361 14532
rect 19668 14492 19674 14504
rect 20349 14501 20361 14504
rect 20395 14501 20407 14535
rect 20349 14495 20407 14501
rect 20530 14492 20536 14544
rect 20588 14492 20594 14544
rect 19702 14464 19708 14476
rect 19615 14436 19708 14464
rect 18693 14399 18751 14405
rect 18693 14365 18705 14399
rect 18739 14365 18751 14399
rect 19518 14396 19524 14408
rect 18693 14359 18751 14365
rect 18800 14368 19524 14396
rect 18800 14328 18828 14368
rect 19518 14356 19524 14368
rect 19576 14356 19582 14408
rect 19628 14405 19656 14436
rect 19702 14424 19708 14436
rect 19760 14464 19766 14476
rect 20548 14464 20576 14492
rect 19760 14436 20576 14464
rect 19760 14424 19766 14436
rect 19613 14399 19671 14405
rect 19613 14365 19625 14399
rect 19659 14365 19671 14399
rect 19886 14396 19892 14408
rect 19847 14368 19892 14396
rect 19613 14359 19671 14365
rect 19886 14356 19892 14368
rect 19944 14356 19950 14408
rect 20438 14356 20444 14408
rect 20496 14396 20502 14408
rect 20533 14399 20591 14405
rect 20533 14396 20545 14399
rect 20496 14368 20545 14396
rect 20496 14356 20502 14368
rect 20533 14365 20545 14368
rect 20579 14365 20591 14399
rect 21082 14396 21088 14408
rect 21043 14368 21088 14396
rect 20533 14359 20591 14365
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 20990 14328 20996 14340
rect 17328 14300 18276 14328
rect 18616 14300 18828 14328
rect 18892 14300 20996 14328
rect 9125 14263 9183 14269
rect 9125 14229 9137 14263
rect 9171 14229 9183 14263
rect 9125 14223 9183 14229
rect 12802 14220 12808 14272
rect 12860 14260 12866 14272
rect 17328 14260 17356 14300
rect 18248 14269 18276 14300
rect 18892 14269 18920 14300
rect 20990 14288 20996 14300
rect 21048 14288 21054 14340
rect 12860 14232 17356 14260
rect 18233 14263 18291 14269
rect 12860 14220 12866 14232
rect 18233 14229 18245 14263
rect 18279 14229 18291 14263
rect 18233 14223 18291 14229
rect 18877 14263 18935 14269
rect 18877 14229 18889 14263
rect 18923 14229 18935 14263
rect 18877 14223 18935 14229
rect 19429 14263 19487 14269
rect 19429 14229 19441 14263
rect 19475 14260 19487 14263
rect 19518 14260 19524 14272
rect 19475 14232 19524 14260
rect 19475 14229 19487 14232
rect 19429 14223 19487 14229
rect 19518 14220 19524 14232
rect 19576 14220 19582 14272
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20622 14260 20628 14272
rect 20128 14232 20628 14260
rect 20128 14220 20134 14232
rect 20622 14220 20628 14232
rect 20680 14220 20686 14272
rect 21266 14260 21272 14272
rect 21227 14232 21272 14260
rect 21266 14220 21272 14232
rect 21324 14220 21330 14272
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 11701 14059 11759 14065
rect 11701 14025 11713 14059
rect 11747 14056 11759 14059
rect 15286 14056 15292 14068
rect 11747 14028 15292 14056
rect 11747 14025 11759 14028
rect 11701 14019 11759 14025
rect 15286 14016 15292 14028
rect 15344 14016 15350 14068
rect 18138 14056 18144 14068
rect 18099 14028 18144 14056
rect 18138 14016 18144 14028
rect 18196 14016 18202 14068
rect 19061 14059 19119 14065
rect 19061 14025 19073 14059
rect 19107 14056 19119 14059
rect 20346 14056 20352 14068
rect 19107 14028 20352 14056
rect 19107 14025 19119 14028
rect 19061 14019 19119 14025
rect 20346 14016 20352 14028
rect 20404 14016 20410 14068
rect 16114 13948 16120 14000
rect 16172 13988 16178 14000
rect 20441 13991 20499 13997
rect 20441 13988 20453 13991
rect 16172 13960 20453 13988
rect 16172 13948 16178 13960
rect 20441 13957 20453 13960
rect 20487 13957 20499 13991
rect 20441 13951 20499 13957
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13920 11575 13923
rect 12066 13920 12072 13932
rect 11563 13892 12072 13920
rect 11563 13889 11575 13892
rect 11517 13883 11575 13889
rect 12066 13880 12072 13892
rect 12124 13880 12130 13932
rect 17129 13923 17187 13929
rect 17129 13889 17141 13923
rect 17175 13920 17187 13923
rect 17954 13920 17960 13932
rect 17175 13892 17816 13920
rect 17915 13892 17960 13920
rect 17175 13889 17187 13892
rect 17129 13883 17187 13889
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 15436 13824 16681 13852
rect 15436 13812 15442 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 17402 13852 17408 13864
rect 17363 13824 17408 13852
rect 16669 13815 16727 13821
rect 17402 13812 17408 13824
rect 17460 13812 17466 13864
rect 17788 13852 17816 13892
rect 17954 13880 17960 13892
rect 18012 13880 18018 13932
rect 18506 13880 18512 13932
rect 18564 13920 18570 13932
rect 18877 13923 18935 13929
rect 18877 13920 18889 13923
rect 18564 13892 18889 13920
rect 18564 13880 18570 13892
rect 18877 13889 18889 13892
rect 18923 13889 18935 13923
rect 18877 13883 18935 13889
rect 19337 13923 19395 13929
rect 19337 13889 19349 13923
rect 19383 13920 19395 13923
rect 19981 13923 20039 13929
rect 19383 13892 19932 13920
rect 19383 13889 19395 13892
rect 19337 13883 19395 13889
rect 18046 13852 18052 13864
rect 17788 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 18601 13855 18659 13861
rect 18601 13821 18613 13855
rect 18647 13852 18659 13855
rect 19702 13852 19708 13864
rect 18647 13824 19708 13852
rect 18647 13821 18659 13824
rect 18601 13815 18659 13821
rect 19702 13812 19708 13824
rect 19760 13812 19766 13864
rect 19904 13852 19932 13892
rect 19981 13889 19993 13923
rect 20027 13920 20039 13923
rect 20027 13892 20208 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 20070 13852 20076 13864
rect 19904 13824 20076 13852
rect 20070 13812 20076 13824
rect 20128 13812 20134 13864
rect 20180 13852 20208 13892
rect 20622 13880 20628 13932
rect 20680 13920 20686 13932
rect 21085 13923 21143 13929
rect 21085 13920 21097 13923
rect 20680 13892 21097 13920
rect 20680 13880 20686 13892
rect 21085 13889 21097 13892
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21634 13852 21640 13864
rect 20180 13824 21640 13852
rect 21634 13812 21640 13824
rect 21692 13812 21698 13864
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 19978 13512 19984 13524
rect 13771 13484 19984 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 19978 13472 19984 13484
rect 20036 13472 20042 13524
rect 20346 13512 20352 13524
rect 20307 13484 20352 13512
rect 20346 13472 20352 13484
rect 20404 13472 20410 13524
rect 14918 13404 14924 13456
rect 14976 13444 14982 13456
rect 16117 13447 16175 13453
rect 16117 13444 16129 13447
rect 14976 13416 16129 13444
rect 14976 13404 14982 13416
rect 16117 13413 16129 13416
rect 16163 13413 16175 13447
rect 16117 13407 16175 13413
rect 19518 13376 19524 13388
rect 18432 13348 19524 13376
rect 13538 13308 13544 13320
rect 13499 13280 13544 13308
rect 13538 13268 13544 13280
rect 13596 13268 13602 13320
rect 17218 13308 17224 13320
rect 17276 13317 17282 13320
rect 17188 13280 17224 13308
rect 17218 13268 17224 13280
rect 17276 13271 17288 13317
rect 17494 13308 17500 13320
rect 17455 13280 17500 13308
rect 17276 13268 17282 13271
rect 17494 13268 17500 13280
rect 17552 13268 17558 13320
rect 17957 13311 18015 13317
rect 17957 13277 17969 13311
rect 18003 13308 18015 13311
rect 18046 13308 18052 13320
rect 18003 13280 18052 13308
rect 18003 13277 18015 13280
rect 17957 13271 18015 13277
rect 18046 13268 18052 13280
rect 18104 13268 18110 13320
rect 18432 13317 18460 13348
rect 19518 13336 19524 13348
rect 19576 13336 19582 13388
rect 18417 13311 18475 13317
rect 18417 13277 18429 13311
rect 18463 13277 18475 13311
rect 18417 13271 18475 13277
rect 18874 13268 18880 13320
rect 18932 13308 18938 13320
rect 19245 13311 19303 13317
rect 19245 13308 19257 13311
rect 18932 13280 19257 13308
rect 18932 13268 18938 13280
rect 19245 13277 19257 13280
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19794 13268 19800 13320
rect 19852 13308 19858 13320
rect 20165 13311 20223 13317
rect 20165 13308 20177 13311
rect 19852 13280 20177 13308
rect 19852 13268 19858 13280
rect 20165 13277 20177 13280
rect 20211 13277 20223 13311
rect 20714 13308 20720 13320
rect 20675 13280 20720 13308
rect 20165 13271 20223 13277
rect 20714 13268 20720 13280
rect 20772 13268 20778 13320
rect 17310 13200 17316 13252
rect 17368 13240 17374 13252
rect 17368 13212 18276 13240
rect 17368 13200 17374 13212
rect 15378 13132 15384 13184
rect 15436 13172 15442 13184
rect 15749 13175 15807 13181
rect 15749 13172 15761 13175
rect 15436 13144 15761 13172
rect 15436 13132 15442 13144
rect 15749 13141 15761 13144
rect 15795 13141 15807 13175
rect 15749 13135 15807 13141
rect 17218 13132 17224 13184
rect 17276 13172 17282 13184
rect 18248 13181 18276 13212
rect 17773 13175 17831 13181
rect 17773 13172 17785 13175
rect 17276 13144 17785 13172
rect 17276 13132 17282 13144
rect 17773 13141 17785 13144
rect 17819 13141 17831 13175
rect 17773 13135 17831 13141
rect 18233 13175 18291 13181
rect 18233 13141 18245 13175
rect 18279 13141 18291 13175
rect 18690 13172 18696 13184
rect 18651 13144 18696 13172
rect 18233 13135 18291 13141
rect 18690 13132 18696 13144
rect 18748 13132 18754 13184
rect 19886 13172 19892 13184
rect 19847 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 21082 13132 21088 13184
rect 21140 13172 21146 13184
rect 21361 13175 21419 13181
rect 21361 13172 21373 13175
rect 21140 13144 21373 13172
rect 21140 13132 21146 13144
rect 21361 13141 21373 13144
rect 21407 13141 21419 13175
rect 21361 13135 21419 13141
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 18049 12971 18107 12977
rect 18049 12937 18061 12971
rect 18095 12968 18107 12971
rect 18690 12968 18696 12980
rect 18095 12940 18696 12968
rect 18095 12937 18107 12940
rect 18049 12931 18107 12937
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 15841 12903 15899 12909
rect 15841 12869 15853 12903
rect 15887 12900 15899 12903
rect 16942 12900 16948 12912
rect 15887 12872 16948 12900
rect 15887 12869 15899 12872
rect 15841 12863 15899 12869
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 17034 12792 17040 12844
rect 17092 12832 17098 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 17092 12804 17417 12832
rect 17092 12792 17098 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 17678 12792 17684 12844
rect 17736 12832 17742 12844
rect 17957 12835 18015 12841
rect 17957 12832 17969 12835
rect 17736 12804 17969 12832
rect 17736 12792 17742 12804
rect 17957 12801 17969 12804
rect 18003 12801 18015 12835
rect 18782 12832 18788 12844
rect 17957 12795 18015 12801
rect 18432 12804 18788 12832
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 16301 12767 16359 12773
rect 16301 12764 16313 12767
rect 15896 12736 16313 12764
rect 15896 12724 15902 12736
rect 16301 12733 16313 12736
rect 16347 12733 16359 12767
rect 16301 12727 16359 12733
rect 17865 12767 17923 12773
rect 17865 12733 17877 12767
rect 17911 12764 17923 12767
rect 18432 12764 18460 12804
rect 18782 12792 18788 12804
rect 18840 12792 18846 12844
rect 20346 12832 20352 12844
rect 20307 12804 20352 12832
rect 20346 12792 20352 12804
rect 20404 12792 20410 12844
rect 20622 12832 20628 12844
rect 20583 12804 20628 12832
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 17911 12736 18460 12764
rect 17911 12733 17923 12736
rect 17865 12727 17923 12733
rect 18414 12696 18420 12708
rect 18375 12668 18420 12696
rect 18414 12656 18420 12668
rect 18472 12656 18478 12708
rect 15010 12588 15016 12640
rect 15068 12628 15074 12640
rect 15197 12631 15255 12637
rect 15197 12628 15209 12631
rect 15068 12600 15209 12628
rect 15068 12588 15074 12600
rect 15197 12597 15209 12600
rect 15243 12597 15255 12631
rect 15197 12591 15255 12597
rect 16761 12631 16819 12637
rect 16761 12597 16773 12631
rect 16807 12628 16819 12631
rect 17586 12628 17592 12640
rect 16807 12600 17592 12628
rect 16807 12597 16819 12600
rect 16761 12591 16819 12597
rect 17586 12588 17592 12600
rect 17644 12588 17650 12640
rect 17862 12588 17868 12640
rect 17920 12628 17926 12640
rect 18138 12628 18144 12640
rect 17920 12600 18144 12628
rect 17920 12588 17926 12600
rect 18138 12588 18144 12600
rect 18196 12588 18202 12640
rect 18322 12588 18328 12640
rect 18380 12628 18386 12640
rect 19429 12631 19487 12637
rect 19429 12628 19441 12631
rect 18380 12600 19441 12628
rect 18380 12588 18386 12600
rect 19429 12597 19441 12600
rect 19475 12597 19487 12631
rect 19429 12591 19487 12597
rect 19518 12588 19524 12640
rect 19576 12628 19582 12640
rect 19705 12631 19763 12637
rect 19705 12628 19717 12631
rect 19576 12600 19717 12628
rect 19576 12588 19582 12600
rect 19705 12597 19717 12600
rect 19751 12597 19763 12631
rect 19705 12591 19763 12597
rect 20898 12588 20904 12640
rect 20956 12628 20962 12640
rect 21269 12631 21327 12637
rect 21269 12628 21281 12631
rect 20956 12600 21281 12628
rect 20956 12588 20962 12600
rect 21269 12597 21281 12600
rect 21315 12597 21327 12631
rect 21269 12591 21327 12597
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 15470 12424 15476 12436
rect 15431 12396 15476 12424
rect 15470 12384 15476 12396
rect 15528 12384 15534 12436
rect 18782 12424 18788 12436
rect 15764 12396 18644 12424
rect 18743 12396 18788 12424
rect 12434 12316 12440 12368
rect 12492 12356 12498 12368
rect 15764 12356 15792 12396
rect 12492 12328 15792 12356
rect 12492 12316 12498 12328
rect 18616 12288 18644 12396
rect 18782 12384 18788 12396
rect 18840 12384 18846 12436
rect 21266 12424 21272 12436
rect 21227 12396 21272 12424
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 18616 12260 19380 12288
rect 15010 12220 15016 12232
rect 14971 12192 15016 12220
rect 15010 12180 15016 12192
rect 15068 12180 15074 12232
rect 15289 12223 15347 12229
rect 15289 12189 15301 12223
rect 15335 12189 15347 12223
rect 15289 12183 15347 12189
rect 15749 12223 15807 12229
rect 15749 12189 15761 12223
rect 15795 12220 15807 12223
rect 17405 12223 17463 12229
rect 17405 12220 17417 12223
rect 15795 12192 17417 12220
rect 15795 12189 15807 12192
rect 15749 12183 15807 12189
rect 17405 12189 17417 12192
rect 17451 12220 17463 12223
rect 17494 12220 17500 12232
rect 17451 12192 17500 12220
rect 17451 12189 17463 12192
rect 17405 12183 17463 12189
rect 7190 12112 7196 12164
rect 7248 12152 7254 12164
rect 15194 12152 15200 12164
rect 7248 12124 15200 12152
rect 7248 12112 7254 12124
rect 15194 12112 15200 12124
rect 15252 12112 15258 12164
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 14366 12044 14372 12096
rect 14424 12084 14430 12096
rect 14461 12087 14519 12093
rect 14461 12084 14473 12087
rect 14424 12056 14473 12084
rect 14424 12044 14430 12056
rect 14461 12053 14473 12056
rect 14507 12053 14519 12087
rect 14826 12084 14832 12096
rect 14787 12056 14832 12084
rect 14461 12047 14519 12053
rect 14826 12044 14832 12056
rect 14884 12044 14890 12096
rect 15304 12084 15332 12183
rect 17494 12180 17500 12192
rect 17552 12220 17558 12232
rect 19245 12223 19303 12229
rect 17552 12192 17908 12220
rect 17552 12180 17558 12192
rect 17880 12164 17908 12192
rect 19245 12189 19257 12223
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 16016 12155 16074 12161
rect 16016 12121 16028 12155
rect 16062 12152 16074 12155
rect 17672 12155 17730 12161
rect 16062 12124 17632 12152
rect 16062 12121 16074 12124
rect 16016 12115 16074 12121
rect 16298 12084 16304 12096
rect 15304 12056 16304 12084
rect 16298 12044 16304 12056
rect 16356 12044 16362 12096
rect 17126 12084 17132 12096
rect 17087 12056 17132 12084
rect 17126 12044 17132 12056
rect 17184 12044 17190 12096
rect 17604 12084 17632 12124
rect 17672 12121 17684 12155
rect 17718 12152 17730 12155
rect 17770 12152 17776 12164
rect 17718 12124 17776 12152
rect 17718 12121 17730 12124
rect 17672 12115 17730 12121
rect 17770 12112 17776 12124
rect 17828 12112 17834 12164
rect 17862 12112 17868 12164
rect 17920 12152 17926 12164
rect 19260 12152 19288 12183
rect 17920 12124 19288 12152
rect 19352 12152 19380 12260
rect 19518 12229 19524 12232
rect 19512 12183 19524 12229
rect 19576 12220 19582 12232
rect 19576 12192 19612 12220
rect 19518 12180 19524 12183
rect 19576 12180 19582 12192
rect 20990 12180 20996 12232
rect 21048 12220 21054 12232
rect 21085 12223 21143 12229
rect 21085 12220 21097 12223
rect 21048 12192 21097 12220
rect 21048 12180 21054 12192
rect 21085 12189 21097 12192
rect 21131 12189 21143 12223
rect 21085 12183 21143 12189
rect 19794 12152 19800 12164
rect 19352 12124 19800 12152
rect 17920 12112 17926 12124
rect 19794 12112 19800 12124
rect 19852 12112 19858 12164
rect 18598 12084 18604 12096
rect 17604 12056 18604 12084
rect 18598 12044 18604 12056
rect 18656 12044 18662 12096
rect 20622 12084 20628 12096
rect 20583 12056 20628 12084
rect 20622 12044 20628 12056
rect 20680 12044 20686 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 12158 11840 12164 11892
rect 12216 11880 12222 11892
rect 15013 11883 15071 11889
rect 15013 11880 15025 11883
rect 12216 11852 15025 11880
rect 12216 11840 12222 11852
rect 15013 11849 15025 11852
rect 15059 11849 15071 11883
rect 16206 11880 16212 11892
rect 16167 11852 16212 11880
rect 15013 11843 15071 11849
rect 16206 11840 16212 11852
rect 16264 11840 16270 11892
rect 17770 11880 17776 11892
rect 17731 11852 17776 11880
rect 17770 11840 17776 11852
rect 17828 11840 17834 11892
rect 17880 11852 18460 11880
rect 16574 11772 16580 11824
rect 16632 11812 16638 11824
rect 17218 11812 17224 11824
rect 16632 11784 17224 11812
rect 16632 11772 16638 11784
rect 17218 11772 17224 11784
rect 17276 11772 17282 11824
rect 17494 11772 17500 11824
rect 17552 11812 17558 11824
rect 17880 11812 17908 11852
rect 18322 11821 18328 11824
rect 18316 11812 18328 11821
rect 17552 11784 17908 11812
rect 18283 11784 18328 11812
rect 17552 11772 17558 11784
rect 18316 11775 18328 11784
rect 18322 11772 18328 11775
rect 18380 11772 18386 11824
rect 18432 11812 18460 11852
rect 20254 11840 20260 11892
rect 20312 11880 20318 11892
rect 20441 11883 20499 11889
rect 20441 11880 20453 11883
rect 20312 11852 20453 11880
rect 20312 11840 20318 11852
rect 20441 11849 20453 11852
rect 20487 11849 20499 11883
rect 20441 11843 20499 11849
rect 18432 11784 21128 11812
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11744 1731 11747
rect 1719 11716 2084 11744
rect 1719 11713 1731 11716
rect 1673 11707 1731 11713
rect 2056 11617 2084 11716
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 13909 11747 13967 11753
rect 13909 11744 13921 11747
rect 13872 11716 13921 11744
rect 13872 11704 13878 11716
rect 13909 11713 13921 11716
rect 13955 11713 13967 11747
rect 13909 11707 13967 11713
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 15194 11744 15200 11756
rect 14332 11716 15056 11744
rect 15155 11716 15200 11744
rect 14332 11704 14338 11716
rect 5258 11636 5264 11688
rect 5316 11676 5322 11688
rect 14826 11676 14832 11688
rect 5316 11648 14832 11676
rect 5316 11636 5322 11648
rect 14826 11636 14832 11648
rect 14884 11636 14890 11688
rect 15028 11676 15056 11716
rect 15194 11704 15200 11716
rect 15252 11704 15258 11756
rect 15841 11747 15899 11753
rect 15841 11713 15853 11747
rect 15887 11744 15899 11747
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15887 11716 16681 11744
rect 15887 11713 15899 11716
rect 15841 11707 15899 11713
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 17126 11744 17132 11756
rect 17087 11716 17132 11744
rect 16669 11707 16727 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 17770 11704 17776 11756
rect 17828 11744 17834 11756
rect 18138 11744 18144 11756
rect 17828 11716 18144 11744
rect 17828 11704 17834 11716
rect 18138 11704 18144 11716
rect 18196 11704 18202 11756
rect 19518 11704 19524 11756
rect 19576 11744 19582 11756
rect 21100 11753 21128 11784
rect 20349 11747 20407 11753
rect 20349 11744 20361 11747
rect 19576 11716 20361 11744
rect 19576 11704 19582 11716
rect 20349 11713 20361 11716
rect 20395 11713 20407 11747
rect 20349 11707 20407 11713
rect 21085 11747 21143 11753
rect 21085 11713 21097 11747
rect 21131 11713 21143 11747
rect 21085 11707 21143 11713
rect 15470 11676 15476 11688
rect 15028 11648 15476 11676
rect 15470 11636 15476 11648
rect 15528 11636 15534 11688
rect 15565 11679 15623 11685
rect 15565 11645 15577 11679
rect 15611 11645 15623 11679
rect 15746 11676 15752 11688
rect 15707 11648 15752 11676
rect 15565 11639 15623 11645
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 12434 11608 12440 11620
rect 2087 11580 12440 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 12434 11568 12440 11580
rect 12492 11568 12498 11620
rect 13633 11611 13691 11617
rect 13633 11577 13645 11611
rect 13679 11608 13691 11611
rect 15194 11608 15200 11620
rect 13679 11580 15200 11608
rect 13679 11577 13691 11580
rect 13633 11571 13691 11577
rect 15194 11568 15200 11580
rect 15252 11568 15258 11620
rect 15580 11608 15608 11639
rect 15746 11636 15752 11648
rect 15804 11636 15810 11688
rect 17862 11636 17868 11688
rect 17920 11676 17926 11688
rect 18049 11679 18107 11685
rect 18049 11676 18061 11679
rect 17920 11648 18061 11676
rect 17920 11636 17926 11648
rect 18049 11645 18061 11648
rect 18095 11645 18107 11679
rect 18049 11639 18107 11645
rect 20533 11679 20591 11685
rect 20533 11645 20545 11679
rect 20579 11645 20591 11679
rect 20533 11639 20591 11645
rect 15838 11608 15844 11620
rect 15580 11580 15844 11608
rect 15838 11568 15844 11580
rect 15896 11568 15902 11620
rect 19429 11611 19487 11617
rect 16868 11580 18000 11608
rect 1486 11540 1492 11552
rect 1447 11512 1492 11540
rect 1486 11500 1492 11512
rect 1544 11500 1550 11552
rect 13262 11540 13268 11552
rect 13223 11512 13268 11540
rect 13262 11500 13268 11512
rect 13320 11500 13326 11552
rect 14550 11540 14556 11552
rect 14511 11512 14556 11540
rect 14550 11500 14556 11512
rect 14608 11500 14614 11552
rect 14642 11500 14648 11552
rect 14700 11540 14706 11552
rect 16868 11540 16896 11580
rect 17972 11552 18000 11580
rect 19429 11577 19441 11611
rect 19475 11608 19487 11611
rect 20346 11608 20352 11620
rect 19475 11580 20352 11608
rect 19475 11577 19487 11580
rect 19429 11571 19487 11577
rect 20346 11568 20352 11580
rect 20404 11608 20410 11620
rect 20548 11608 20576 11639
rect 20404 11580 20576 11608
rect 20404 11568 20410 11580
rect 14700 11512 16896 11540
rect 14700 11500 14706 11512
rect 16942 11500 16948 11552
rect 17000 11540 17006 11552
rect 17218 11540 17224 11552
rect 17000 11512 17224 11540
rect 17000 11500 17006 11512
rect 17218 11500 17224 11512
rect 17276 11500 17282 11552
rect 17954 11500 17960 11552
rect 18012 11500 18018 11552
rect 19978 11540 19984 11552
rect 19939 11512 19984 11540
rect 19978 11500 19984 11512
rect 20036 11500 20042 11552
rect 21269 11543 21327 11549
rect 21269 11509 21281 11543
rect 21315 11540 21327 11543
rect 21450 11540 21456 11552
rect 21315 11512 21456 11540
rect 21315 11509 21327 11512
rect 21269 11503 21327 11509
rect 21450 11500 21456 11512
rect 21508 11500 21514 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 16574 11336 16580 11348
rect 12492 11308 12537 11336
rect 13096 11308 16580 11336
rect 12492 11296 12498 11308
rect 13096 11141 13124 11308
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 16666 11296 16672 11348
rect 16724 11336 16730 11348
rect 16724 11308 16769 11336
rect 16724 11296 16730 11308
rect 18322 11296 18328 11348
rect 18380 11336 18386 11348
rect 19797 11339 19855 11345
rect 18380 11308 19748 11336
rect 18380 11296 18386 11308
rect 13265 11271 13323 11277
rect 13265 11237 13277 11271
rect 13311 11268 13323 11271
rect 14274 11268 14280 11280
rect 13311 11240 14280 11268
rect 13311 11237 13323 11240
rect 13265 11231 13323 11237
rect 14274 11228 14280 11240
rect 14332 11228 14338 11280
rect 15838 11228 15844 11280
rect 15896 11268 15902 11280
rect 16117 11271 16175 11277
rect 16117 11268 16129 11271
rect 15896 11240 16129 11268
rect 15896 11228 15902 11240
rect 16117 11237 16129 11240
rect 16163 11268 16175 11271
rect 18598 11268 18604 11280
rect 16163 11240 17264 11268
rect 18559 11240 18604 11268
rect 16163 11237 16175 11240
rect 16117 11231 16175 11237
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11200 13783 11203
rect 14642 11200 14648 11212
rect 13771 11172 14648 11200
rect 13771 11169 13783 11172
rect 13725 11163 13783 11169
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 17126 11200 17132 11212
rect 17087 11172 17132 11200
rect 17126 11160 17132 11172
rect 17184 11160 17190 11212
rect 13081 11135 13139 11141
rect 13081 11101 13093 11135
rect 13127 11101 13139 11135
rect 14737 11135 14795 11141
rect 13081 11095 13139 11101
rect 14108 11104 14688 11132
rect 12805 11067 12863 11073
rect 12805 11033 12817 11067
rect 12851 11064 12863 11067
rect 14108 11064 14136 11104
rect 12851 11036 14136 11064
rect 12851 11033 12863 11036
rect 12805 11027 12863 11033
rect 14274 10956 14280 11008
rect 14332 10996 14338 11008
rect 14660 10996 14688 11104
rect 14737 11101 14749 11135
rect 14783 11132 14795 11135
rect 14826 11132 14832 11144
rect 14783 11104 14832 11132
rect 14783 11101 14795 11104
rect 14737 11095 14795 11101
rect 14826 11092 14832 11104
rect 14884 11132 14890 11144
rect 16485 11135 16543 11141
rect 14884 11104 16436 11132
rect 14884 11092 14890 11104
rect 15004 11067 15062 11073
rect 15004 11033 15016 11067
rect 15050 11064 15062 11067
rect 16408 11064 16436 11104
rect 16485 11101 16497 11135
rect 16531 11132 16543 11135
rect 16942 11132 16948 11144
rect 16531 11104 16948 11132
rect 16531 11101 16543 11104
rect 16485 11095 16543 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 17236 11132 17264 11240
rect 18598 11228 18604 11240
rect 18656 11228 18662 11280
rect 18782 11228 18788 11280
rect 18840 11268 18846 11280
rect 19245 11271 19303 11277
rect 19245 11268 19257 11271
rect 18840 11240 19257 11268
rect 18840 11228 18846 11240
rect 19245 11237 19257 11240
rect 19291 11237 19303 11271
rect 19245 11231 19303 11237
rect 17494 11160 17500 11212
rect 17552 11200 17558 11212
rect 17678 11200 17684 11212
rect 17552 11172 17684 11200
rect 17552 11160 17558 11172
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 18966 11160 18972 11212
rect 19024 11200 19030 11212
rect 19024 11172 19472 11200
rect 19024 11160 19030 11172
rect 19444 11141 19472 11172
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17236 11104 17969 11132
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 17862 11064 17868 11076
rect 15050 11036 16344 11064
rect 16408 11036 17868 11064
rect 15050 11033 15062 11036
rect 15004 11027 15062 11033
rect 15378 10996 15384 11008
rect 14332 10968 14377 10996
rect 14660 10968 15384 10996
rect 14332 10956 14338 10968
rect 15378 10956 15384 10968
rect 15436 10956 15442 11008
rect 16316 10996 16344 11036
rect 17862 11024 17868 11036
rect 17920 11024 17926 11076
rect 19720 11064 19748 11308
rect 19797 11305 19809 11339
rect 19843 11336 19855 11339
rect 20990 11336 20996 11348
rect 19843 11308 20996 11336
rect 19843 11305 19855 11308
rect 19797 11299 19855 11305
rect 20990 11296 20996 11308
rect 21048 11296 21054 11348
rect 20070 11092 20076 11144
rect 20128 11132 20134 11144
rect 21177 11135 21235 11141
rect 21177 11132 21189 11135
rect 20128 11104 21189 11132
rect 20128 11092 20134 11104
rect 21177 11101 21189 11104
rect 21223 11101 21235 11135
rect 21177 11095 21235 11101
rect 20714 11064 20720 11076
rect 19720 11036 20720 11064
rect 20714 11024 20720 11036
rect 20772 11024 20778 11076
rect 20898 11064 20904 11076
rect 20956 11073 20962 11076
rect 20868 11036 20904 11064
rect 20898 11024 20904 11036
rect 20956 11027 20968 11073
rect 20956 11024 20962 11027
rect 16390 10996 16396 11008
rect 16316 10968 16396 10996
rect 16390 10956 16396 10968
rect 16448 10956 16454 11008
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 17221 10999 17279 11005
rect 17221 10996 17233 10999
rect 17184 10968 17233 10996
rect 17184 10956 17190 10968
rect 17221 10965 17233 10968
rect 17267 10965 17279 10999
rect 17221 10959 17279 10965
rect 17313 10999 17371 11005
rect 17313 10965 17325 10999
rect 17359 10996 17371 10999
rect 17494 10996 17500 11008
rect 17359 10968 17500 10996
rect 17359 10965 17371 10968
rect 17313 10959 17371 10965
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 17681 10999 17739 11005
rect 17681 10965 17693 10999
rect 17727 10996 17739 10999
rect 18138 10996 18144 11008
rect 17727 10968 18144 10996
rect 17727 10965 17739 10968
rect 17681 10959 17739 10965
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 13909 10795 13967 10801
rect 13909 10792 13921 10795
rect 13872 10764 13921 10792
rect 13872 10752 13878 10764
rect 13909 10761 13921 10764
rect 13955 10761 13967 10795
rect 19429 10795 19487 10801
rect 19429 10792 19441 10795
rect 13909 10755 13967 10761
rect 14384 10764 19441 10792
rect 14384 10724 14412 10764
rect 19429 10761 19441 10764
rect 19475 10761 19487 10795
rect 19429 10755 19487 10761
rect 19702 10752 19708 10804
rect 19760 10792 19766 10804
rect 19797 10795 19855 10801
rect 19797 10792 19809 10795
rect 19760 10764 19809 10792
rect 19760 10752 19766 10764
rect 19797 10761 19809 10764
rect 19843 10761 19855 10795
rect 19797 10755 19855 10761
rect 19889 10795 19947 10801
rect 19889 10761 19901 10795
rect 19935 10792 19947 10795
rect 19978 10792 19984 10804
rect 19935 10764 19984 10792
rect 19935 10761 19947 10764
rect 19889 10755 19947 10761
rect 19978 10752 19984 10764
rect 20036 10752 20042 10804
rect 20714 10752 20720 10804
rect 20772 10792 20778 10804
rect 20901 10795 20959 10801
rect 20901 10792 20913 10795
rect 20772 10764 20913 10792
rect 20772 10752 20778 10764
rect 20901 10761 20913 10764
rect 20947 10761 20959 10795
rect 20901 10755 20959 10761
rect 12406 10696 14412 10724
rect 14452 10727 14510 10733
rect 12253 10659 12311 10665
rect 12253 10625 12265 10659
rect 12299 10656 12311 10659
rect 12406 10656 12434 10696
rect 14452 10693 14464 10727
rect 14498 10724 14510 10727
rect 14550 10724 14556 10736
rect 14498 10696 14556 10724
rect 14498 10693 14510 10696
rect 14452 10687 14510 10693
rect 14550 10684 14556 10696
rect 14608 10684 14614 10736
rect 15378 10684 15384 10736
rect 15436 10724 15442 10736
rect 18322 10724 18328 10736
rect 15436 10696 18328 10724
rect 15436 10684 15442 10696
rect 12299 10628 12434 10656
rect 12796 10659 12854 10665
rect 12299 10625 12311 10628
rect 12253 10619 12311 10625
rect 12796 10625 12808 10659
rect 12842 10656 12854 10659
rect 13078 10656 13084 10668
rect 12842 10628 13084 10656
rect 12842 10625 12854 10628
rect 12796 10619 12854 10625
rect 13078 10616 13084 10628
rect 13136 10616 13142 10668
rect 14185 10659 14243 10665
rect 14185 10625 14197 10659
rect 14231 10656 14243 10659
rect 14826 10656 14832 10668
rect 14231 10628 14832 10656
rect 14231 10625 14243 10628
rect 14185 10619 14243 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 16316 10665 16344 10696
rect 18322 10684 18328 10696
rect 18380 10684 18386 10736
rect 18782 10684 18788 10736
rect 18840 10724 18846 10736
rect 19061 10727 19119 10733
rect 19061 10724 19073 10727
rect 18840 10696 19073 10724
rect 18840 10684 18846 10696
rect 19061 10693 19073 10696
rect 19107 10724 19119 10727
rect 19150 10724 19156 10736
rect 19107 10696 19156 10724
rect 19107 10693 19119 10696
rect 19061 10687 19119 10693
rect 19150 10684 19156 10696
rect 19208 10684 19214 10736
rect 19518 10684 19524 10736
rect 19576 10724 19582 10736
rect 20809 10727 20867 10733
rect 20809 10724 20821 10727
rect 19576 10696 20821 10724
rect 19576 10684 19582 10696
rect 20809 10693 20821 10696
rect 20855 10693 20867 10727
rect 20809 10687 20867 10693
rect 16301 10659 16359 10665
rect 16301 10625 16313 10659
rect 16347 10625 16359 10659
rect 16301 10619 16359 10625
rect 18069 10659 18127 10665
rect 18069 10625 18081 10659
rect 18115 10656 18127 10659
rect 20346 10656 20352 10668
rect 18115 10628 20352 10656
rect 18115 10625 18127 10628
rect 18069 10619 18127 10625
rect 20346 10616 20352 10628
rect 20404 10616 20410 10668
rect 20824 10656 20852 10687
rect 20898 10656 20904 10668
rect 20824 10628 20904 10656
rect 20898 10616 20904 10628
rect 20956 10616 20962 10668
rect 6546 10548 6552 10600
rect 6604 10588 6610 10600
rect 6604 10560 12204 10588
rect 6604 10548 6610 10560
rect 6730 10480 6736 10532
rect 6788 10520 6794 10532
rect 12069 10523 12127 10529
rect 12069 10520 12081 10523
rect 6788 10492 12081 10520
rect 6788 10480 6794 10492
rect 12069 10489 12081 10492
rect 12115 10489 12127 10523
rect 12069 10483 12127 10489
rect 11793 10455 11851 10461
rect 11793 10421 11805 10455
rect 11839 10452 11851 10455
rect 11974 10452 11980 10464
rect 11839 10424 11980 10452
rect 11839 10421 11851 10424
rect 11793 10415 11851 10421
rect 11974 10412 11980 10424
rect 12032 10412 12038 10464
rect 12176 10452 12204 10560
rect 12342 10548 12348 10600
rect 12400 10588 12406 10600
rect 12529 10591 12587 10597
rect 12529 10588 12541 10591
rect 12400 10560 12541 10588
rect 12400 10548 12406 10560
rect 12529 10557 12541 10560
rect 12575 10557 12587 10591
rect 12529 10551 12587 10557
rect 15838 10548 15844 10600
rect 15896 10588 15902 10600
rect 18325 10591 18383 10597
rect 15896 10560 17172 10588
rect 15896 10548 15902 10560
rect 17034 10520 17040 10532
rect 15396 10492 17040 10520
rect 15396 10452 15424 10492
rect 17034 10480 17040 10492
rect 17092 10480 17098 10532
rect 15562 10452 15568 10464
rect 12176 10424 15424 10452
rect 15523 10424 15568 10452
rect 15562 10412 15568 10424
rect 15620 10412 15626 10464
rect 15654 10412 15660 10464
rect 15712 10452 15718 10464
rect 16117 10455 16175 10461
rect 16117 10452 16129 10455
rect 15712 10424 16129 10452
rect 15712 10412 15718 10424
rect 16117 10421 16129 10424
rect 16163 10421 16175 10455
rect 16942 10452 16948 10464
rect 16903 10424 16948 10452
rect 16117 10415 16175 10421
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 17144 10452 17172 10560
rect 18325 10557 18337 10591
rect 18371 10557 18383 10591
rect 18598 10588 18604 10600
rect 18559 10560 18604 10588
rect 18325 10551 18383 10557
rect 18340 10520 18368 10551
rect 18598 10548 18604 10560
rect 18656 10548 18662 10600
rect 19981 10591 20039 10597
rect 19981 10557 19993 10591
rect 20027 10588 20039 10591
rect 20622 10588 20628 10600
rect 20027 10560 20628 10588
rect 20027 10557 20039 10560
rect 19981 10551 20039 10557
rect 20622 10548 20628 10560
rect 20680 10548 20686 10600
rect 20990 10548 20996 10600
rect 21048 10588 21054 10600
rect 21048 10560 21093 10588
rect 21048 10548 21054 10560
rect 20070 10520 20076 10532
rect 18340 10492 20076 10520
rect 20070 10480 20076 10492
rect 20128 10480 20134 10532
rect 19518 10452 19524 10464
rect 17144 10424 19524 10452
rect 19518 10412 19524 10424
rect 19576 10412 19582 10464
rect 19702 10412 19708 10464
rect 19760 10452 19766 10464
rect 20441 10455 20499 10461
rect 20441 10452 20453 10455
rect 19760 10424 20453 10452
rect 19760 10412 19766 10424
rect 20441 10421 20453 10424
rect 20487 10421 20499 10455
rect 20441 10415 20499 10421
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 7374 10208 7380 10260
rect 7432 10248 7438 10260
rect 14366 10248 14372 10260
rect 7432 10220 14372 10248
rect 7432 10208 7438 10220
rect 14366 10208 14372 10220
rect 14424 10208 14430 10260
rect 14829 10251 14887 10257
rect 14829 10217 14841 10251
rect 14875 10248 14887 10251
rect 15102 10248 15108 10260
rect 14875 10220 15108 10248
rect 14875 10217 14887 10220
rect 14829 10211 14887 10217
rect 15102 10208 15108 10220
rect 15160 10208 15166 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 15841 10251 15899 10257
rect 15841 10248 15853 10251
rect 15804 10220 15853 10248
rect 15804 10208 15810 10220
rect 15841 10217 15853 10220
rect 15887 10217 15899 10251
rect 15841 10211 15899 10217
rect 16574 10208 16580 10260
rect 16632 10248 16638 10260
rect 16761 10251 16819 10257
rect 16761 10248 16773 10251
rect 16632 10220 16773 10248
rect 16632 10208 16638 10220
rect 16761 10217 16773 10220
rect 16807 10217 16819 10251
rect 17034 10248 17040 10260
rect 16995 10220 17040 10248
rect 16761 10211 16819 10217
rect 17034 10208 17040 10220
rect 17092 10208 17098 10260
rect 20346 10248 20352 10260
rect 20307 10220 20352 10248
rect 20346 10208 20352 10220
rect 20404 10208 20410 10260
rect 5442 10140 5448 10192
rect 5500 10180 5506 10192
rect 15654 10180 15660 10192
rect 5500 10152 15660 10180
rect 5500 10140 5506 10152
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 17126 10140 17132 10192
rect 17184 10180 17190 10192
rect 17494 10180 17500 10192
rect 17184 10152 17500 10180
rect 17184 10140 17190 10152
rect 17494 10140 17500 10152
rect 17552 10140 17558 10192
rect 18877 10183 18935 10189
rect 18877 10149 18889 10183
rect 18923 10180 18935 10183
rect 18923 10152 19932 10180
rect 18923 10149 18935 10152
rect 18877 10143 18935 10149
rect 13814 10072 13820 10124
rect 13872 10112 13878 10124
rect 14185 10115 14243 10121
rect 14185 10112 14197 10115
rect 13872 10084 14197 10112
rect 13872 10072 13878 10084
rect 14185 10081 14197 10084
rect 14231 10081 14243 10115
rect 14185 10075 14243 10081
rect 15289 10115 15347 10121
rect 15289 10081 15301 10115
rect 15335 10081 15347 10115
rect 15289 10075 15347 10081
rect 11146 10044 11152 10056
rect 11107 10016 11152 10044
rect 11146 10004 11152 10016
rect 11204 10004 11210 10056
rect 13538 10044 13544 10056
rect 13499 10016 13544 10044
rect 13538 10004 13544 10016
rect 13596 10004 13602 10056
rect 14274 10004 14280 10056
rect 14332 10044 14338 10056
rect 14461 10047 14519 10053
rect 14461 10044 14473 10047
rect 14332 10016 14473 10044
rect 14332 10004 14338 10016
rect 14461 10013 14473 10016
rect 14507 10013 14519 10047
rect 15304 10044 15332 10075
rect 19610 10072 19616 10124
rect 19668 10112 19674 10124
rect 19904 10121 19932 10152
rect 19797 10115 19855 10121
rect 19797 10112 19809 10115
rect 19668 10084 19809 10112
rect 19668 10072 19674 10084
rect 19797 10081 19809 10084
rect 19843 10081 19855 10115
rect 19797 10075 19855 10081
rect 19889 10115 19947 10121
rect 19889 10081 19901 10115
rect 19935 10112 19947 10115
rect 20346 10112 20352 10124
rect 19935 10084 20352 10112
rect 19935 10081 19947 10084
rect 19889 10075 19947 10081
rect 20346 10072 20352 10084
rect 20404 10072 20410 10124
rect 15562 10044 15568 10056
rect 15304 10016 15568 10044
rect 14461 10007 14519 10013
rect 15562 10004 15568 10016
rect 15620 10044 15626 10056
rect 16117 10047 16175 10053
rect 16117 10044 16129 10047
rect 15620 10016 16129 10044
rect 15620 10004 15626 10016
rect 16117 10013 16129 10016
rect 16163 10013 16175 10047
rect 16117 10007 16175 10013
rect 17221 10047 17279 10053
rect 17221 10013 17233 10047
rect 17267 10013 17279 10047
rect 17221 10007 17279 10013
rect 17497 10047 17555 10053
rect 17497 10013 17509 10047
rect 17543 10044 17555 10047
rect 17543 10016 17908 10044
rect 17543 10013 17555 10016
rect 17497 10007 17555 10013
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 15473 9979 15531 9985
rect 15473 9976 15485 9979
rect 15344 9948 15485 9976
rect 15344 9936 15350 9948
rect 15473 9945 15485 9948
rect 15519 9945 15531 9979
rect 15473 9939 15531 9945
rect 11790 9908 11796 9920
rect 11751 9880 11796 9908
rect 11790 9868 11796 9880
rect 11848 9868 11854 9920
rect 12066 9908 12072 9920
rect 12027 9880 12072 9908
rect 12066 9868 12072 9880
rect 12124 9868 12130 9920
rect 12434 9868 12440 9920
rect 12492 9908 12498 9920
rect 12529 9911 12587 9917
rect 12529 9908 12541 9911
rect 12492 9880 12541 9908
rect 12492 9868 12498 9880
rect 12529 9877 12541 9880
rect 12575 9877 12587 9911
rect 12894 9908 12900 9920
rect 12855 9880 12900 9908
rect 12529 9871 12587 9877
rect 12894 9868 12900 9880
rect 12952 9868 12958 9920
rect 14366 9908 14372 9920
rect 14327 9880 14372 9908
rect 14366 9868 14372 9880
rect 14424 9868 14430 9920
rect 15381 9911 15439 9917
rect 15381 9877 15393 9911
rect 15427 9908 15439 9911
rect 17126 9908 17132 9920
rect 15427 9880 17132 9908
rect 15427 9877 15439 9880
rect 15381 9871 15439 9877
rect 17126 9868 17132 9880
rect 17184 9868 17190 9920
rect 17236 9908 17264 10007
rect 17880 9988 17908 10016
rect 19518 10004 19524 10056
rect 19576 10044 19582 10056
rect 19705 10047 19763 10053
rect 19705 10044 19717 10047
rect 19576 10016 19717 10044
rect 19576 10004 19582 10016
rect 19705 10013 19717 10016
rect 19751 10013 19763 10047
rect 20990 10044 20996 10056
rect 20951 10016 20996 10044
rect 19705 10007 19763 10013
rect 20990 10004 20996 10016
rect 21048 10004 21054 10056
rect 17586 9936 17592 9988
rect 17644 9976 17650 9988
rect 17742 9979 17800 9985
rect 17742 9976 17754 9979
rect 17644 9948 17754 9976
rect 17644 9936 17650 9948
rect 17742 9945 17754 9948
rect 17788 9945 17800 9979
rect 17742 9939 17800 9945
rect 17862 9936 17868 9988
rect 17920 9936 17926 9988
rect 17972 9948 21404 9976
rect 17972 9908 18000 9948
rect 21376 9920 21404 9948
rect 17236 9880 18000 9908
rect 19337 9911 19395 9917
rect 19337 9877 19349 9911
rect 19383 9908 19395 9911
rect 19518 9908 19524 9920
rect 19383 9880 19524 9908
rect 19383 9877 19395 9880
rect 19337 9871 19395 9877
rect 19518 9868 19524 9880
rect 19576 9868 19582 9920
rect 21358 9908 21364 9920
rect 21319 9880 21364 9908
rect 21358 9868 21364 9880
rect 21416 9868 21422 9920
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 11146 9704 11152 9716
rect 11107 9676 11152 9704
rect 11146 9664 11152 9676
rect 11204 9664 11210 9716
rect 12897 9707 12955 9713
rect 12897 9673 12909 9707
rect 12943 9704 12955 9707
rect 12986 9704 12992 9716
rect 12943 9676 12992 9704
rect 12943 9673 12955 9676
rect 12897 9667 12955 9673
rect 12986 9664 12992 9676
rect 13044 9704 13050 9716
rect 13538 9704 13544 9716
rect 13044 9676 13544 9704
rect 13044 9664 13050 9676
rect 13538 9664 13544 9676
rect 13596 9664 13602 9716
rect 15470 9664 15476 9716
rect 15528 9704 15534 9716
rect 17678 9704 17684 9716
rect 15528 9676 17684 9704
rect 15528 9664 15534 9676
rect 17678 9664 17684 9676
rect 17736 9664 17742 9716
rect 18049 9707 18107 9713
rect 18049 9673 18061 9707
rect 18095 9704 18107 9707
rect 18598 9704 18604 9716
rect 18095 9676 18604 9704
rect 18095 9673 18107 9676
rect 18049 9667 18107 9673
rect 18598 9664 18604 9676
rect 18656 9664 18662 9716
rect 8386 9596 8392 9648
rect 8444 9636 8450 9648
rect 9033 9639 9091 9645
rect 9033 9636 9045 9639
rect 8444 9608 9045 9636
rect 8444 9596 8450 9608
rect 9033 9605 9045 9608
rect 9079 9605 9091 9639
rect 12342 9636 12348 9648
rect 9033 9599 9091 9605
rect 9784 9608 12348 9636
rect 9784 9580 9812 9608
rect 7650 9528 7656 9580
rect 7708 9568 7714 9580
rect 9125 9571 9183 9577
rect 9125 9568 9137 9571
rect 7708 9540 9137 9568
rect 7708 9528 7714 9540
rect 9125 9537 9137 9540
rect 9171 9537 9183 9571
rect 9766 9568 9772 9580
rect 9679 9540 9772 9568
rect 9125 9531 9183 9537
rect 9766 9528 9772 9540
rect 9824 9528 9830 9580
rect 10036 9571 10094 9577
rect 10036 9537 10048 9571
rect 10082 9568 10094 9571
rect 11238 9568 11244 9580
rect 10082 9540 11244 9568
rect 10082 9537 10094 9540
rect 10036 9531 10094 9537
rect 11238 9528 11244 9540
rect 11296 9528 11302 9580
rect 11532 9577 11560 9608
rect 12342 9596 12348 9608
rect 12400 9596 12406 9648
rect 14185 9639 14243 9645
rect 14185 9605 14197 9639
rect 14231 9636 14243 9639
rect 15749 9639 15807 9645
rect 15749 9636 15761 9639
rect 14231 9608 15761 9636
rect 14231 9605 14243 9608
rect 14185 9599 14243 9605
rect 15749 9605 15761 9608
rect 15795 9605 15807 9639
rect 15749 9599 15807 9605
rect 17037 9639 17095 9645
rect 17037 9605 17049 9639
rect 17083 9636 17095 9639
rect 17402 9636 17408 9648
rect 17083 9608 17408 9636
rect 17083 9605 17095 9608
rect 17037 9599 17095 9605
rect 17402 9596 17408 9608
rect 17460 9596 17466 9648
rect 18141 9639 18199 9645
rect 18141 9605 18153 9639
rect 18187 9636 18199 9639
rect 19702 9636 19708 9648
rect 18187 9608 19708 9636
rect 18187 9605 18199 9608
rect 18141 9599 18199 9605
rect 19702 9596 19708 9608
rect 19760 9596 19766 9648
rect 19828 9639 19886 9645
rect 19828 9605 19840 9639
rect 19874 9636 19886 9639
rect 20993 9639 21051 9645
rect 20993 9636 21005 9639
rect 19874 9608 21005 9636
rect 19874 9605 19886 9608
rect 19828 9599 19886 9605
rect 20993 9605 21005 9608
rect 21039 9605 21051 9639
rect 20993 9599 21051 9605
rect 11790 9577 11796 9580
rect 11517 9571 11575 9577
rect 11517 9537 11529 9571
rect 11563 9537 11575 9571
rect 11784 9568 11796 9577
rect 11751 9540 11796 9568
rect 11517 9531 11575 9537
rect 11784 9531 11796 9540
rect 11790 9528 11796 9531
rect 11848 9528 11854 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9537 13599 9571
rect 14829 9571 14887 9577
rect 14829 9568 14841 9571
rect 13541 9531 13599 9537
rect 14016 9540 14841 9568
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 8849 9503 8907 9509
rect 8849 9500 8861 9503
rect 7984 9472 8861 9500
rect 7984 9460 7990 9472
rect 8849 9469 8861 9472
rect 8895 9469 8907 9503
rect 8849 9463 8907 9469
rect 9490 9432 9496 9444
rect 9451 9404 9496 9432
rect 9490 9392 9496 9404
rect 9548 9392 9554 9444
rect 10778 9392 10784 9444
rect 10836 9432 10842 9444
rect 13357 9435 13415 9441
rect 13357 9432 13369 9435
rect 10836 9404 11008 9432
rect 10836 9392 10842 9404
rect 1578 9324 1584 9376
rect 1636 9364 1642 9376
rect 10870 9364 10876 9376
rect 1636 9336 10876 9364
rect 1636 9324 1642 9336
rect 10870 9324 10876 9336
rect 10928 9324 10934 9376
rect 10980 9364 11008 9404
rect 12820 9404 13369 9432
rect 12820 9364 12848 9404
rect 13357 9401 13369 9404
rect 13403 9401 13415 9435
rect 13357 9395 13415 9401
rect 10980 9336 12848 9364
rect 13556 9364 13584 9531
rect 13722 9460 13728 9512
rect 13780 9500 13786 9512
rect 14016 9509 14044 9540
rect 14829 9537 14841 9540
rect 14875 9537 14887 9571
rect 14829 9531 14887 9537
rect 15010 9528 15016 9580
rect 15068 9568 15074 9580
rect 18046 9568 18052 9580
rect 15068 9540 18052 9568
rect 15068 9528 15074 9540
rect 18046 9528 18052 9540
rect 18104 9528 18110 9580
rect 20346 9568 20352 9580
rect 20307 9540 20352 9568
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 14001 9503 14059 9509
rect 14001 9500 14013 9503
rect 13780 9472 14013 9500
rect 13780 9460 13786 9472
rect 14001 9469 14013 9472
rect 14047 9469 14059 9503
rect 14001 9463 14059 9469
rect 14093 9503 14151 9509
rect 14093 9469 14105 9503
rect 14139 9469 14151 9503
rect 14093 9463 14151 9469
rect 14200 9472 14688 9500
rect 13630 9392 13636 9444
rect 13688 9432 13694 9444
rect 14108 9432 14136 9463
rect 13688 9404 14136 9432
rect 13688 9392 13694 9404
rect 14200 9364 14228 9472
rect 14458 9392 14464 9444
rect 14516 9432 14522 9444
rect 14553 9435 14611 9441
rect 14553 9432 14565 9435
rect 14516 9404 14565 9432
rect 14516 9392 14522 9404
rect 14553 9401 14565 9404
rect 14599 9401 14611 9435
rect 14660 9432 14688 9472
rect 15286 9460 15292 9512
rect 15344 9500 15350 9512
rect 16209 9503 16267 9509
rect 16209 9500 16221 9503
rect 15344 9472 16221 9500
rect 15344 9460 15350 9472
rect 16209 9469 16221 9472
rect 16255 9469 16267 9503
rect 16758 9500 16764 9512
rect 16719 9472 16764 9500
rect 16209 9463 16267 9469
rect 16758 9460 16764 9472
rect 16816 9460 16822 9512
rect 16942 9500 16948 9512
rect 16903 9472 16948 9500
rect 16942 9460 16948 9472
rect 17000 9460 17006 9512
rect 17034 9460 17040 9512
rect 17092 9500 17098 9512
rect 18233 9503 18291 9509
rect 18233 9500 18245 9503
rect 17092 9472 18245 9500
rect 17092 9460 17098 9472
rect 18233 9469 18245 9472
rect 18279 9469 18291 9503
rect 20070 9500 20076 9512
rect 20031 9472 20076 9500
rect 18233 9463 18291 9469
rect 20070 9460 20076 9472
rect 20128 9460 20134 9512
rect 17681 9435 17739 9441
rect 17681 9432 17693 9435
rect 14660 9404 17693 9432
rect 14553 9395 14611 9401
rect 17681 9401 17693 9404
rect 17727 9401 17739 9435
rect 17681 9395 17739 9401
rect 18693 9435 18751 9441
rect 18693 9401 18705 9435
rect 18739 9432 18751 9435
rect 18874 9432 18880 9444
rect 18739 9404 18880 9432
rect 18739 9401 18751 9404
rect 18693 9395 18751 9401
rect 18874 9392 18880 9404
rect 18932 9392 18938 9444
rect 13556 9336 14228 9364
rect 14642 9324 14648 9376
rect 14700 9364 14706 9376
rect 15473 9367 15531 9373
rect 15473 9364 15485 9367
rect 14700 9336 15485 9364
rect 14700 9324 14706 9336
rect 15473 9333 15485 9336
rect 15519 9333 15531 9367
rect 15473 9327 15531 9333
rect 17405 9367 17463 9373
rect 17405 9333 17417 9367
rect 17451 9364 17463 9367
rect 17770 9364 17776 9376
rect 17451 9336 17776 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 17770 9324 17776 9336
rect 17828 9324 17834 9376
rect 20898 9324 20904 9376
rect 20956 9364 20962 9376
rect 21269 9367 21327 9373
rect 21269 9364 21281 9367
rect 20956 9336 21281 9364
rect 20956 9324 20962 9336
rect 21269 9333 21281 9336
rect 21315 9333 21327 9367
rect 21269 9327 21327 9333
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 7098 9120 7104 9172
rect 7156 9160 7162 9172
rect 10778 9160 10784 9172
rect 7156 9132 10784 9160
rect 7156 9120 7162 9132
rect 10778 9120 10784 9132
rect 10836 9120 10842 9172
rect 10870 9120 10876 9172
rect 10928 9160 10934 9172
rect 13538 9160 13544 9172
rect 10928 9132 13544 9160
rect 10928 9120 10934 9132
rect 13538 9120 13544 9132
rect 13596 9120 13602 9172
rect 13722 9160 13728 9172
rect 13683 9132 13728 9160
rect 13722 9120 13728 9132
rect 13780 9120 13786 9172
rect 18141 9163 18199 9169
rect 18141 9160 18153 9163
rect 13924 9132 18153 9160
rect 10689 9095 10747 9101
rect 10689 9061 10701 9095
rect 10735 9092 10747 9095
rect 11974 9092 11980 9104
rect 10735 9064 11980 9092
rect 10735 9061 10747 9064
rect 10689 9055 10747 9061
rect 11974 9052 11980 9064
rect 12032 9052 12038 9104
rect 7650 9024 7656 9036
rect 7611 8996 7656 9024
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 11146 9024 11152 9036
rect 11107 8996 11152 9024
rect 11146 8984 11152 8996
rect 11204 8984 11210 9036
rect 11256 8996 12480 9024
rect 7926 8956 7932 8968
rect 7887 8928 7932 8956
rect 7926 8916 7932 8928
rect 7984 8916 7990 8968
rect 8941 8959 8999 8965
rect 8941 8925 8953 8959
rect 8987 8956 8999 8959
rect 9490 8956 9496 8968
rect 8987 8928 9496 8956
rect 8987 8925 8999 8928
rect 8941 8919 8999 8925
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 11256 8956 11284 8996
rect 12452 8968 12480 8996
rect 9600 8928 11284 8956
rect 11333 8959 11391 8965
rect 8573 8891 8631 8897
rect 8573 8857 8585 8891
rect 8619 8888 8631 8891
rect 9186 8891 9244 8897
rect 9186 8888 9198 8891
rect 8619 8860 9198 8888
rect 8619 8857 8631 8860
rect 8573 8851 8631 8857
rect 9186 8857 9198 8860
rect 9232 8857 9244 8891
rect 9186 8851 9244 8857
rect 4614 8780 4620 8832
rect 4672 8820 4678 8832
rect 9600 8820 9628 8928
rect 11333 8925 11345 8959
rect 11379 8956 11391 8959
rect 12066 8956 12072 8968
rect 11379 8928 12072 8956
rect 11379 8925 11391 8928
rect 11333 8919 11391 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 12434 8916 12440 8968
rect 12492 8916 12498 8968
rect 12612 8959 12670 8965
rect 12612 8925 12624 8959
rect 12658 8956 12670 8959
rect 12894 8956 12900 8968
rect 12658 8928 12900 8956
rect 12658 8925 12670 8928
rect 12612 8919 12670 8925
rect 12894 8916 12900 8928
rect 12952 8916 12958 8968
rect 13924 8956 13952 9132
rect 18141 9129 18153 9132
rect 18187 9129 18199 9163
rect 19794 9160 19800 9172
rect 18141 9123 18199 9129
rect 18524 9132 19800 9160
rect 17773 9095 17831 9101
rect 17773 9061 17785 9095
rect 17819 9092 17831 9095
rect 18524 9092 18552 9132
rect 19794 9120 19800 9132
rect 19852 9120 19858 9172
rect 20806 9120 20812 9172
rect 20864 9160 20870 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 20864 9132 20913 9160
rect 20864 9120 20870 9132
rect 20901 9129 20913 9132
rect 20947 9129 20959 9163
rect 20901 9123 20959 9129
rect 19518 9092 19524 9104
rect 17819 9064 18552 9092
rect 18616 9064 19524 9092
rect 17819 9061 17831 9064
rect 17773 9055 17831 9061
rect 16758 8984 16764 9036
rect 16816 9024 16822 9036
rect 18616 9033 18644 9064
rect 19518 9052 19524 9064
rect 19576 9052 19582 9104
rect 18601 9027 18659 9033
rect 16816 8996 17724 9024
rect 16816 8984 16822 8996
rect 13372 8928 13952 8956
rect 14093 8959 14151 8965
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 13372 8888 13400 8928
rect 14093 8925 14105 8959
rect 14139 8956 14151 8959
rect 15749 8959 15807 8965
rect 15749 8956 15761 8959
rect 14139 8928 15761 8956
rect 14139 8925 14151 8928
rect 14093 8919 14151 8925
rect 15749 8925 15761 8928
rect 15795 8956 15807 8959
rect 16390 8956 16396 8968
rect 15795 8928 16396 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 16390 8916 16396 8928
rect 16448 8916 16454 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 17052 8928 17601 8956
rect 10008 8860 13400 8888
rect 14360 8891 14418 8897
rect 10008 8848 10014 8860
rect 14360 8857 14372 8891
rect 14406 8888 14418 8891
rect 14642 8888 14648 8900
rect 14406 8860 14648 8888
rect 14406 8857 14418 8860
rect 14360 8851 14418 8857
rect 14642 8848 14648 8860
rect 14700 8848 14706 8900
rect 16016 8891 16074 8897
rect 16016 8857 16028 8891
rect 16062 8888 16074 8891
rect 16206 8888 16212 8900
rect 16062 8860 16212 8888
rect 16062 8857 16074 8860
rect 16016 8851 16074 8857
rect 16206 8848 16212 8860
rect 16264 8848 16270 8900
rect 4672 8792 9628 8820
rect 10321 8823 10379 8829
rect 4672 8780 4678 8792
rect 10321 8789 10333 8823
rect 10367 8820 10379 8823
rect 10502 8820 10508 8832
rect 10367 8792 10508 8820
rect 10367 8789 10379 8792
rect 10321 8783 10379 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 11204 8792 11253 8820
rect 11204 8780 11210 8792
rect 11241 8789 11253 8792
rect 11287 8789 11299 8823
rect 11698 8820 11704 8832
rect 11659 8792 11704 8820
rect 11241 8783 11299 8789
rect 11698 8780 11704 8792
rect 11756 8780 11762 8832
rect 12069 8823 12127 8829
rect 12069 8789 12081 8823
rect 12115 8820 12127 8823
rect 12894 8820 12900 8832
rect 12115 8792 12900 8820
rect 12115 8789 12127 8792
rect 12069 8783 12127 8789
rect 12894 8780 12900 8792
rect 12952 8780 12958 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 15286 8820 15292 8832
rect 13596 8792 15292 8820
rect 13596 8780 13602 8792
rect 15286 8780 15292 8792
rect 15344 8780 15350 8832
rect 15470 8820 15476 8832
rect 15431 8792 15476 8820
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 15654 8780 15660 8832
rect 15712 8820 15718 8832
rect 17052 8820 17080 8928
rect 17589 8925 17601 8928
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 17696 8888 17724 8996
rect 18601 8993 18613 9027
rect 18647 8993 18659 9027
rect 18601 8987 18659 8993
rect 18785 9027 18843 9033
rect 18785 8993 18797 9027
rect 18831 9024 18843 9027
rect 18874 9024 18880 9036
rect 18831 8996 18880 9024
rect 18831 8993 18843 8996
rect 18785 8987 18843 8993
rect 18874 8984 18880 8996
rect 18932 8984 18938 9036
rect 20714 8984 20720 9036
rect 20772 9024 20778 9036
rect 20772 8996 21404 9024
rect 20772 8984 20778 8996
rect 17862 8916 17868 8968
rect 17920 8956 17926 8968
rect 19518 8956 19524 8968
rect 17920 8928 19524 8956
rect 17920 8916 17926 8928
rect 19518 8916 19524 8928
rect 19576 8956 19582 8968
rect 20070 8956 20076 8968
rect 19576 8928 20076 8956
rect 19576 8916 19582 8928
rect 20070 8916 20076 8928
rect 20128 8916 20134 8968
rect 21376 8965 21404 8996
rect 21361 8959 21419 8965
rect 21361 8925 21373 8959
rect 21407 8956 21419 8959
rect 21726 8956 21732 8968
rect 21407 8928 21732 8956
rect 21407 8925 21419 8928
rect 21361 8919 21419 8925
rect 21726 8916 21732 8928
rect 21784 8916 21790 8968
rect 18598 8888 18604 8900
rect 17144 8860 18604 8888
rect 17144 8829 17172 8860
rect 18598 8848 18604 8860
rect 18656 8848 18662 8900
rect 19788 8891 19846 8897
rect 19788 8857 19800 8891
rect 19834 8888 19846 8891
rect 19886 8888 19892 8900
rect 19834 8860 19892 8888
rect 19834 8857 19846 8860
rect 19788 8851 19846 8857
rect 19886 8848 19892 8860
rect 19944 8848 19950 8900
rect 15712 8792 17080 8820
rect 17129 8823 17187 8829
rect 15712 8780 15718 8792
rect 17129 8789 17141 8823
rect 17175 8789 17187 8823
rect 17129 8783 17187 8789
rect 17218 8780 17224 8832
rect 17276 8820 17282 8832
rect 18509 8823 18567 8829
rect 18509 8820 18521 8823
rect 17276 8792 18521 8820
rect 17276 8780 17282 8792
rect 18509 8789 18521 8792
rect 18555 8789 18567 8823
rect 18509 8783 18567 8789
rect 20070 8780 20076 8832
rect 20128 8820 20134 8832
rect 20254 8820 20260 8832
rect 20128 8792 20260 8820
rect 20128 8780 20134 8792
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 21174 8820 21180 8832
rect 21135 8792 21180 8820
rect 21174 8780 21180 8792
rect 21232 8780 21238 8832
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 7926 8576 7932 8628
rect 7984 8616 7990 8628
rect 8113 8619 8171 8625
rect 8113 8616 8125 8619
rect 7984 8588 8125 8616
rect 7984 8576 7990 8588
rect 8113 8585 8125 8588
rect 8159 8585 8171 8619
rect 11146 8616 11152 8628
rect 8113 8579 8171 8585
rect 8312 8588 10916 8616
rect 11107 8588 11152 8616
rect 4154 8508 4160 8560
rect 4212 8548 4218 8560
rect 8312 8548 8340 8588
rect 4212 8520 8340 8548
rect 4212 8508 4218 8520
rect 10686 8508 10692 8560
rect 10744 8548 10750 8560
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 10744 8520 10793 8548
rect 10744 8508 10750 8520
rect 10781 8517 10793 8520
rect 10827 8517 10839 8551
rect 10888 8548 10916 8588
rect 11146 8576 11152 8588
rect 11204 8576 11210 8628
rect 11238 8576 11244 8628
rect 11296 8616 11302 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 11296 8588 12173 8616
rect 11296 8576 11302 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12161 8579 12219 8585
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 13630 8616 13636 8628
rect 12492 8588 13400 8616
rect 13591 8588 13636 8616
rect 12492 8576 12498 8588
rect 13265 8551 13323 8557
rect 13265 8548 13277 8551
rect 10888 8520 13277 8548
rect 10781 8511 10839 8517
rect 13265 8517 13277 8520
rect 13311 8517 13323 8551
rect 13372 8548 13400 8588
rect 13630 8576 13636 8588
rect 13688 8576 13694 8628
rect 14366 8576 14372 8628
rect 14424 8616 14430 8628
rect 14829 8619 14887 8625
rect 14829 8616 14841 8619
rect 14424 8588 14841 8616
rect 14424 8576 14430 8588
rect 14829 8585 14841 8588
rect 14875 8585 14887 8619
rect 14829 8579 14887 8585
rect 16025 8619 16083 8625
rect 16025 8585 16037 8619
rect 16071 8616 16083 8619
rect 16942 8616 16948 8628
rect 16071 8588 16948 8616
rect 16071 8585 16083 8588
rect 16025 8579 16083 8585
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18325 8619 18383 8625
rect 18325 8616 18337 8619
rect 18288 8588 18337 8616
rect 18288 8576 18294 8588
rect 18325 8585 18337 8588
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 19521 8619 19579 8625
rect 19521 8585 19533 8619
rect 19567 8616 19579 8619
rect 19610 8616 19616 8628
rect 19567 8588 19616 8616
rect 19567 8585 19579 8588
rect 19521 8579 19579 8585
rect 19610 8576 19616 8588
rect 19668 8576 19674 8628
rect 19702 8576 19708 8628
rect 19760 8616 19766 8628
rect 19981 8619 20039 8625
rect 19981 8616 19993 8619
rect 19760 8588 19993 8616
rect 19760 8576 19766 8588
rect 19981 8585 19993 8588
rect 20027 8616 20039 8619
rect 20254 8616 20260 8628
rect 20027 8588 20260 8616
rect 20027 8585 20039 8588
rect 19981 8579 20039 8585
rect 20254 8576 20260 8588
rect 20312 8576 20318 8628
rect 14461 8551 14519 8557
rect 14461 8548 14473 8551
rect 13372 8520 14473 8548
rect 13265 8511 13323 8517
rect 14461 8517 14473 8520
rect 14507 8517 14519 8551
rect 15930 8548 15936 8560
rect 14461 8511 14519 8517
rect 15212 8520 15936 8548
rect 7282 8440 7288 8492
rect 7340 8480 7346 8492
rect 9226 8483 9284 8489
rect 9226 8480 9238 8483
rect 7340 8452 9238 8480
rect 7340 8440 7346 8452
rect 9226 8449 9238 8452
rect 9272 8449 9284 8483
rect 9490 8480 9496 8492
rect 9451 8452 9496 8480
rect 9226 8443 9284 8449
rect 9490 8440 9496 8452
rect 9548 8480 9554 8492
rect 9766 8480 9772 8492
rect 9548 8452 9772 8480
rect 9548 8440 9554 8452
rect 9766 8440 9772 8452
rect 9824 8440 9830 8492
rect 9950 8480 9956 8492
rect 9911 8452 9956 8480
rect 9950 8440 9956 8452
rect 10008 8440 10014 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 10520 8452 11529 8480
rect 10520 8424 10548 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8480 13231 8483
rect 14369 8483 14427 8489
rect 14369 8480 14381 8483
rect 13219 8452 14381 8480
rect 13219 8449 13231 8452
rect 13173 8443 13231 8449
rect 14369 8449 14381 8452
rect 14415 8480 14427 8483
rect 15212 8480 15240 8520
rect 15930 8508 15936 8520
rect 15988 8508 15994 8560
rect 16390 8508 16396 8560
rect 16448 8548 16454 8560
rect 17862 8548 17868 8560
rect 16448 8520 17868 8548
rect 16448 8508 16454 8520
rect 14415 8452 15240 8480
rect 14415 8449 14427 8452
rect 14369 8443 14427 8449
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 16684 8489 16712 8520
rect 17862 8508 17868 8520
rect 17920 8508 17926 8560
rect 17954 8508 17960 8560
rect 18012 8548 18018 8560
rect 18693 8551 18751 8557
rect 18693 8548 18705 8551
rect 18012 8520 18705 8548
rect 18012 8508 18018 8520
rect 18693 8517 18705 8520
rect 18739 8517 18751 8551
rect 18693 8511 18751 8517
rect 21082 8508 21088 8560
rect 21140 8557 21146 8560
rect 21140 8548 21152 8557
rect 21140 8520 21185 8548
rect 21140 8511 21152 8520
rect 21140 8508 21146 8511
rect 15657 8483 15715 8489
rect 15657 8480 15669 8483
rect 15344 8452 15669 8480
rect 15344 8440 15350 8452
rect 15657 8449 15669 8452
rect 15703 8449 15715 8483
rect 15657 8443 15715 8449
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16936 8483 16994 8489
rect 16936 8449 16948 8483
rect 16982 8480 16994 8483
rect 18506 8480 18512 8492
rect 16982 8452 18512 8480
rect 16982 8449 16994 8452
rect 16936 8443 16994 8449
rect 18506 8440 18512 8452
rect 18564 8440 18570 8492
rect 18966 8440 18972 8492
rect 19024 8480 19030 8492
rect 19337 8483 19395 8489
rect 19337 8480 19349 8483
rect 19024 8452 19349 8480
rect 19024 8440 19030 8452
rect 19337 8449 19349 8452
rect 19383 8449 19395 8483
rect 19337 8443 19395 8449
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 21361 8483 21419 8489
rect 21361 8480 21373 8483
rect 19576 8452 21373 8480
rect 19576 8440 19582 8452
rect 21361 8449 21373 8452
rect 21407 8449 21419 8483
rect 21361 8443 21419 8449
rect 10502 8412 10508 8424
rect 10463 8384 10508 8412
rect 10502 8372 10508 8384
rect 10560 8372 10566 8424
rect 10689 8415 10747 8421
rect 10689 8381 10701 8415
rect 10735 8412 10747 8415
rect 10778 8412 10784 8424
rect 10735 8384 10784 8412
rect 10735 8381 10747 8384
rect 10689 8375 10747 8381
rect 10778 8372 10784 8384
rect 10836 8372 10842 8424
rect 12526 8372 12532 8424
rect 12584 8412 12590 8424
rect 12621 8415 12679 8421
rect 12621 8412 12633 8415
rect 12584 8384 12633 8412
rect 12584 8372 12590 8384
rect 12621 8381 12633 8384
rect 12667 8381 12679 8415
rect 12986 8412 12992 8424
rect 12947 8384 12992 8412
rect 12621 8375 12679 8381
rect 12986 8372 12992 8384
rect 13044 8372 13050 8424
rect 13722 8372 13728 8424
rect 13780 8412 13786 8424
rect 14185 8415 14243 8421
rect 14185 8412 14197 8415
rect 13780 8384 14197 8412
rect 13780 8372 13786 8384
rect 14185 8381 14197 8384
rect 14231 8381 14243 8415
rect 15470 8412 15476 8424
rect 15431 8384 15476 8412
rect 14185 8375 14243 8381
rect 15470 8372 15476 8384
rect 15528 8372 15534 8424
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8412 15623 8415
rect 15611 8384 16712 8412
rect 15611 8381 15623 8384
rect 15565 8375 15623 8381
rect 11146 8304 11152 8356
rect 11204 8344 11210 8356
rect 15654 8344 15660 8356
rect 11204 8316 15660 8344
rect 11204 8304 11210 8316
rect 15654 8304 15660 8316
rect 15712 8304 15718 8356
rect 10134 8276 10140 8288
rect 10095 8248 10140 8276
rect 10134 8236 10140 8248
rect 10192 8236 10198 8288
rect 16684 8276 16712 8384
rect 17954 8372 17960 8424
rect 18012 8412 18018 8424
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18012 8384 18797 8412
rect 18012 8372 18018 8384
rect 18785 8381 18797 8384
rect 18831 8381 18843 8415
rect 18785 8375 18843 8381
rect 18874 8372 18880 8424
rect 18932 8412 18938 8424
rect 18932 8384 18977 8412
rect 18932 8372 18938 8384
rect 17678 8304 17684 8356
rect 17736 8344 17742 8356
rect 18049 8347 18107 8353
rect 18049 8344 18061 8347
rect 17736 8316 18061 8344
rect 17736 8304 17742 8316
rect 18049 8313 18061 8316
rect 18095 8344 18107 8347
rect 18095 8316 20484 8344
rect 18095 8313 18107 8316
rect 18049 8307 18107 8313
rect 17034 8276 17040 8288
rect 16684 8248 17040 8276
rect 17034 8236 17040 8248
rect 17092 8236 17098 8288
rect 20456 8276 20484 8316
rect 20714 8276 20720 8288
rect 20456 8248 20720 8276
rect 20714 8236 20720 8248
rect 20772 8236 20778 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 10873 8075 10931 8081
rect 10873 8072 10885 8075
rect 10560 8044 10885 8072
rect 10560 8032 10566 8044
rect 10873 8041 10885 8044
rect 10919 8072 10931 8075
rect 12342 8072 12348 8084
rect 10919 8044 12348 8072
rect 10919 8041 10931 8044
rect 10873 8035 10931 8041
rect 12342 8032 12348 8044
rect 12400 8032 12406 8084
rect 13078 8072 13084 8084
rect 13039 8044 13084 8072
rect 13078 8032 13084 8044
rect 13136 8032 13142 8084
rect 17862 8072 17868 8084
rect 17823 8044 17868 8072
rect 17862 8032 17868 8044
rect 17920 8032 17926 8084
rect 18138 8072 18144 8084
rect 17972 8044 18144 8072
rect 8294 7964 8300 8016
rect 8352 8004 8358 8016
rect 13630 8004 13636 8016
rect 8352 7976 13636 8004
rect 8352 7964 8358 7976
rect 13630 7964 13636 7976
rect 13688 7964 13694 8016
rect 17972 8004 18000 8044
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 15488 7976 18000 8004
rect 9585 7939 9643 7945
rect 9585 7936 9597 7939
rect 8588 7908 9597 7936
rect 7466 7868 7472 7880
rect 7427 7840 7472 7868
rect 7466 7828 7472 7840
rect 7524 7828 7530 7880
rect 8588 7877 8616 7908
rect 9585 7905 9597 7908
rect 9631 7936 9643 7939
rect 10594 7936 10600 7948
rect 9631 7908 10600 7936
rect 9631 7905 9643 7908
rect 9585 7899 9643 7905
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 15488 7936 15516 7976
rect 18046 7964 18052 8016
rect 18104 8004 18110 8016
rect 19705 8007 19763 8013
rect 19705 8004 19717 8007
rect 18104 7976 19717 8004
rect 18104 7964 18110 7976
rect 19705 7973 19717 7976
rect 19751 7973 19763 8007
rect 19705 7967 19763 7973
rect 10888 7908 15516 7936
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7837 8631 7871
rect 8573 7831 8631 7837
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9677 7871 9735 7877
rect 8812 7840 9628 7868
rect 8812 7828 8818 7840
rect 6914 7800 6920 7812
rect 6875 7772 6920 7800
rect 6914 7760 6920 7772
rect 6972 7760 6978 7812
rect 8938 7760 8944 7812
rect 8996 7800 9002 7812
rect 9490 7800 9496 7812
rect 8996 7772 9496 7800
rect 8996 7760 9002 7772
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 7653 7735 7711 7741
rect 7653 7701 7665 7735
rect 7699 7732 7711 7735
rect 7834 7732 7840 7744
rect 7699 7704 7840 7732
rect 7699 7701 7711 7704
rect 7653 7695 7711 7701
rect 7834 7692 7840 7704
rect 7892 7692 7898 7744
rect 7929 7735 7987 7741
rect 7929 7701 7941 7735
rect 7975 7732 7987 7735
rect 8478 7732 8484 7744
rect 7975 7704 8484 7732
rect 7975 7701 7987 7704
rect 7929 7695 7987 7701
rect 8478 7692 8484 7704
rect 8536 7692 8542 7744
rect 9122 7732 9128 7744
rect 9083 7704 9128 7732
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 9600 7732 9628 7840
rect 9677 7837 9689 7871
rect 9723 7868 9735 7871
rect 10778 7868 10784 7880
rect 9723 7840 10784 7868
rect 9723 7837 9735 7840
rect 9677 7831 9735 7837
rect 10778 7828 10784 7840
rect 10836 7828 10842 7880
rect 10888 7800 10916 7908
rect 15562 7896 15568 7948
rect 15620 7936 15626 7948
rect 19245 7939 19303 7945
rect 19245 7936 19257 7939
rect 15620 7908 19257 7936
rect 15620 7896 15626 7908
rect 19245 7905 19257 7908
rect 19291 7905 19303 7939
rect 20254 7936 20260 7948
rect 20215 7908 20260 7936
rect 19245 7899 19303 7905
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 12805 7871 12863 7877
rect 12805 7837 12817 7871
rect 12851 7868 12863 7871
rect 12894 7868 12900 7880
rect 12851 7840 12900 7868
rect 12851 7837 12863 7840
rect 12805 7831 12863 7837
rect 12894 7828 12900 7840
rect 12952 7828 12958 7880
rect 13722 7868 13728 7880
rect 13683 7840 13728 7868
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 16114 7868 16120 7880
rect 16075 7840 16120 7868
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 18046 7828 18052 7880
rect 18104 7868 18110 7880
rect 18601 7871 18659 7877
rect 18601 7868 18613 7871
rect 18104 7840 18613 7868
rect 18104 7828 18110 7840
rect 18601 7837 18613 7840
rect 18647 7837 18659 7871
rect 18601 7831 18659 7837
rect 19058 7828 19064 7880
rect 19116 7868 19122 7880
rect 20073 7871 20131 7877
rect 20073 7868 20085 7871
rect 19116 7840 20085 7868
rect 19116 7828 19122 7840
rect 20073 7837 20085 7840
rect 20119 7837 20131 7871
rect 20714 7868 20720 7880
rect 20675 7840 20720 7868
rect 20073 7831 20131 7837
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 9692 7772 10916 7800
rect 9692 7732 9720 7772
rect 10962 7760 10968 7812
rect 11020 7800 11026 7812
rect 12158 7800 12164 7812
rect 11020 7772 11376 7800
rect 12119 7772 12164 7800
rect 11020 7760 11026 7772
rect 9600 7704 9720 7732
rect 9766 7692 9772 7744
rect 9824 7732 9830 7744
rect 10137 7735 10195 7741
rect 9824 7704 9869 7732
rect 9824 7692 9830 7704
rect 10137 7701 10149 7735
rect 10183 7732 10195 7735
rect 11238 7732 11244 7744
rect 10183 7704 11244 7732
rect 10183 7701 10195 7704
rect 10137 7695 10195 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 11348 7732 11376 7772
rect 12158 7760 12164 7772
rect 12216 7800 12222 7812
rect 14369 7803 14427 7809
rect 14369 7800 14381 7803
rect 12216 7772 14381 7800
rect 12216 7760 12222 7772
rect 14369 7769 14381 7772
rect 14415 7800 14427 7803
rect 15654 7800 15660 7812
rect 14415 7772 15660 7800
rect 14415 7769 14427 7772
rect 14369 7763 14427 7769
rect 15654 7760 15660 7772
rect 15712 7800 15718 7812
rect 16393 7803 16451 7809
rect 16393 7800 16405 7803
rect 15712 7772 16405 7800
rect 15712 7760 15718 7772
rect 16393 7769 16405 7772
rect 16439 7769 16451 7803
rect 21542 7800 21548 7812
rect 16393 7763 16451 7769
rect 18800 7772 21548 7800
rect 12621 7735 12679 7741
rect 12621 7732 12633 7735
rect 11348 7704 12633 7732
rect 12621 7701 12633 7704
rect 12667 7701 12679 7735
rect 12621 7695 12679 7701
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 15838 7732 15844 7744
rect 13044 7704 15844 7732
rect 13044 7692 13050 7704
rect 15838 7692 15844 7704
rect 15896 7692 15902 7744
rect 18800 7741 18828 7772
rect 21542 7760 21548 7772
rect 21600 7760 21606 7812
rect 18785 7735 18843 7741
rect 18785 7701 18797 7735
rect 18831 7701 18843 7735
rect 18785 7695 18843 7701
rect 20165 7735 20223 7741
rect 20165 7701 20177 7735
rect 20211 7732 20223 7735
rect 20530 7732 20536 7744
rect 20211 7704 20536 7732
rect 20211 7701 20223 7704
rect 20165 7695 20223 7701
rect 20530 7692 20536 7704
rect 20588 7692 20594 7744
rect 21358 7732 21364 7744
rect 21319 7704 21364 7732
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 7984 7500 8892 7528
rect 7984 7488 7990 7500
rect 6641 7463 6699 7469
rect 6641 7429 6653 7463
rect 6687 7460 6699 7463
rect 8294 7460 8300 7472
rect 6687 7432 7880 7460
rect 8255 7432 8300 7460
rect 6687 7429 6699 7432
rect 6641 7423 6699 7429
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 7852 7401 7880 7432
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 8864 7460 8892 7500
rect 9214 7488 9220 7540
rect 9272 7528 9278 7540
rect 9766 7528 9772 7540
rect 9272 7500 9772 7528
rect 9272 7488 9278 7500
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 10594 7528 10600 7540
rect 10555 7500 10600 7528
rect 10594 7488 10600 7500
rect 10652 7488 10658 7540
rect 11146 7528 11152 7540
rect 11107 7500 11152 7528
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 13633 7531 13691 7537
rect 13633 7497 13645 7531
rect 13679 7528 13691 7531
rect 13722 7528 13728 7540
rect 13679 7500 13728 7528
rect 13679 7497 13691 7500
rect 13633 7491 13691 7497
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 16206 7528 16212 7540
rect 16167 7500 16212 7528
rect 16206 7488 16212 7500
rect 16264 7488 16270 7540
rect 18325 7531 18383 7537
rect 18325 7497 18337 7531
rect 18371 7528 18383 7531
rect 18874 7528 18880 7540
rect 18371 7500 18880 7528
rect 18371 7497 18383 7500
rect 18325 7491 18383 7497
rect 18874 7488 18880 7500
rect 18932 7488 18938 7540
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 19981 7531 20039 7537
rect 19981 7528 19993 7531
rect 19944 7500 19993 7528
rect 19944 7488 19950 7500
rect 19981 7497 19993 7500
rect 20027 7528 20039 7531
rect 20070 7528 20076 7540
rect 20027 7500 20076 7528
rect 20027 7497 20039 7500
rect 19981 7491 20039 7497
rect 20070 7488 20076 7500
rect 20128 7488 20134 7540
rect 20530 7528 20536 7540
rect 20491 7500 20536 7528
rect 20530 7488 20536 7500
rect 20588 7488 20594 7540
rect 20898 7528 20904 7540
rect 20859 7500 20904 7528
rect 20898 7488 20904 7500
rect 20956 7488 20962 7540
rect 9473 7463 9531 7469
rect 9473 7460 9485 7463
rect 8864 7432 9485 7460
rect 9473 7429 9485 7432
rect 9519 7429 9531 7463
rect 12342 7460 12348 7472
rect 12255 7432 12348 7460
rect 9473 7423 9531 7429
rect 7377 7395 7435 7401
rect 7377 7392 7389 7395
rect 5592 7364 7389 7392
rect 5592 7352 5598 7364
rect 7377 7361 7389 7364
rect 7423 7361 7435 7395
rect 7377 7355 7435 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8754 7392 8760 7404
rect 7883 7364 8760 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 8941 7395 8999 7401
rect 8941 7361 8953 7395
rect 8987 7392 8999 7395
rect 10042 7392 10048 7404
rect 8987 7364 10048 7392
rect 8987 7361 8999 7364
rect 8941 7355 8999 7361
rect 10042 7352 10048 7364
rect 10100 7352 10106 7404
rect 10962 7392 10968 7404
rect 10923 7364 10968 7392
rect 10962 7352 10968 7364
rect 11020 7352 11026 7404
rect 11974 7392 11980 7404
rect 11935 7364 11980 7392
rect 11974 7352 11980 7364
rect 12032 7352 12038 7404
rect 12268 7401 12296 7432
rect 12342 7420 12348 7432
rect 12400 7460 12406 7472
rect 14176 7463 14234 7469
rect 12400 7432 13952 7460
rect 12400 7420 12406 7432
rect 12253 7395 12311 7401
rect 12253 7361 12265 7395
rect 12299 7361 12311 7395
rect 12253 7355 12311 7361
rect 12520 7395 12578 7401
rect 12520 7361 12532 7395
rect 12566 7392 12578 7395
rect 13078 7392 13084 7404
rect 12566 7364 13084 7392
rect 12566 7361 12578 7364
rect 12520 7355 12578 7361
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 13924 7401 13952 7432
rect 14176 7429 14188 7463
rect 14222 7460 14234 7463
rect 17212 7463 17270 7469
rect 14222 7432 17172 7460
rect 14222 7429 14234 7432
rect 14176 7423 14234 7429
rect 13909 7395 13967 7401
rect 13909 7361 13921 7395
rect 13955 7361 13967 7395
rect 13909 7355 13967 7361
rect 15470 7352 15476 7404
rect 15528 7392 15534 7404
rect 15565 7395 15623 7401
rect 15565 7392 15577 7395
rect 15528 7364 15577 7392
rect 15528 7352 15534 7364
rect 15565 7361 15577 7364
rect 15611 7361 15623 7395
rect 17144 7392 17172 7432
rect 17212 7429 17224 7463
rect 17258 7460 17270 7463
rect 21358 7460 21364 7472
rect 17258 7432 21364 7460
rect 17258 7429 17270 7432
rect 17212 7423 17270 7429
rect 21358 7420 21364 7432
rect 21416 7420 21422 7472
rect 18230 7392 18236 7404
rect 17144 7364 18236 7392
rect 15565 7355 15623 7361
rect 18230 7352 18236 7364
rect 18288 7352 18294 7404
rect 18598 7392 18604 7404
rect 18559 7364 18604 7392
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 19889 7395 19947 7401
rect 19889 7361 19901 7395
rect 19935 7392 19947 7395
rect 20070 7392 20076 7404
rect 19935 7364 20076 7392
rect 19935 7361 19947 7364
rect 19889 7355 19947 7361
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20990 7352 20996 7404
rect 21048 7392 21054 7404
rect 21048 7364 21093 7392
rect 21048 7352 21054 7364
rect 7101 7327 7159 7333
rect 7101 7293 7113 7327
rect 7147 7324 7159 7327
rect 7650 7324 7656 7336
rect 7147 7296 7656 7324
rect 7147 7293 7159 7296
rect 7101 7287 7159 7293
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 9030 7284 9036 7336
rect 9088 7324 9094 7336
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 9088 7296 9229 7324
rect 9088 7284 9094 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 16942 7324 16948 7336
rect 16903 7296 16948 7324
rect 9217 7287 9275 7293
rect 16942 7284 16948 7296
rect 17000 7284 17006 7336
rect 18506 7284 18512 7336
rect 18564 7324 18570 7336
rect 19245 7327 19303 7333
rect 19245 7324 19257 7327
rect 18564 7296 19257 7324
rect 18564 7284 18570 7296
rect 19245 7293 19257 7296
rect 19291 7293 19303 7327
rect 19245 7287 19303 7293
rect 20165 7327 20223 7333
rect 20165 7293 20177 7327
rect 20211 7293 20223 7327
rect 20165 7287 20223 7293
rect 8018 7256 8024 7268
rect 7979 7228 8024 7256
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 20180 7256 20208 7287
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21085 7327 21143 7333
rect 21085 7324 21097 7327
rect 20864 7296 21097 7324
rect 20864 7284 20870 7296
rect 21085 7293 21097 7296
rect 21131 7293 21143 7327
rect 21085 7287 21143 7293
rect 21266 7256 21272 7268
rect 15120 7228 15424 7256
rect 20180 7228 21272 7256
rect 7561 7191 7619 7197
rect 7561 7157 7573 7191
rect 7607 7188 7619 7191
rect 9490 7188 9496 7200
rect 7607 7160 9496 7188
rect 7607 7157 7619 7160
rect 7561 7151 7619 7157
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 10778 7148 10784 7200
rect 10836 7188 10842 7200
rect 11606 7188 11612 7200
rect 10836 7160 11612 7188
rect 10836 7148 10842 7160
rect 11606 7148 11612 7160
rect 11664 7148 11670 7200
rect 11790 7188 11796 7200
rect 11751 7160 11796 7188
rect 11790 7148 11796 7160
rect 11848 7148 11854 7200
rect 11974 7148 11980 7200
rect 12032 7188 12038 7200
rect 15120 7188 15148 7228
rect 12032 7160 15148 7188
rect 12032 7148 12038 7160
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15289 7191 15347 7197
rect 15289 7188 15301 7191
rect 15252 7160 15301 7188
rect 15252 7148 15258 7160
rect 15289 7157 15301 7160
rect 15335 7157 15347 7191
rect 15396 7188 15424 7228
rect 21266 7216 21272 7228
rect 21324 7216 21330 7268
rect 18506 7188 18512 7200
rect 15396 7160 18512 7188
rect 15289 7151 15347 7157
rect 18506 7148 18512 7160
rect 18564 7148 18570 7200
rect 19521 7191 19579 7197
rect 19521 7157 19533 7191
rect 19567 7188 19579 7191
rect 19794 7188 19800 7200
rect 19567 7160 19800 7188
rect 19567 7157 19579 7160
rect 19521 7151 19579 7157
rect 19794 7148 19800 7160
rect 19852 7148 19858 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 5166 6944 5172 6996
rect 5224 6984 5230 6996
rect 10870 6984 10876 6996
rect 5224 6956 10876 6984
rect 5224 6944 5230 6956
rect 10870 6944 10876 6956
rect 10928 6944 10934 6996
rect 11606 6944 11612 6996
rect 11664 6984 11670 6996
rect 11664 6956 12848 6984
rect 11664 6944 11670 6956
rect 3142 6876 3148 6928
rect 3200 6916 3206 6928
rect 7006 6916 7012 6928
rect 3200 6888 7012 6916
rect 3200 6876 3206 6888
rect 7006 6876 7012 6888
rect 7064 6876 7070 6928
rect 7926 6916 7932 6928
rect 7887 6888 7932 6916
rect 7926 6876 7932 6888
rect 7984 6876 7990 6928
rect 9677 6919 9735 6925
rect 8496 6888 9168 6916
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5859 6820 7052 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 6549 6783 6607 6789
rect 6549 6749 6561 6783
rect 6595 6780 6607 6783
rect 6914 6780 6920 6792
rect 6595 6752 6920 6780
rect 6595 6749 6607 6752
rect 6549 6743 6607 6749
rect 6914 6740 6920 6752
rect 6972 6740 6978 6792
rect 7024 6789 7052 6820
rect 7009 6783 7067 6789
rect 7009 6749 7021 6783
rect 7055 6780 7067 6783
rect 8496 6780 8524 6888
rect 9030 6848 9036 6860
rect 8588 6820 9036 6848
rect 8588 6789 8616 6820
rect 9030 6808 9036 6820
rect 9088 6808 9094 6860
rect 9140 6848 9168 6888
rect 9677 6885 9689 6919
rect 9723 6916 9735 6919
rect 9858 6916 9864 6928
rect 9723 6888 9864 6916
rect 9723 6885 9735 6888
rect 9677 6879 9735 6885
rect 9858 6876 9864 6888
rect 9916 6876 9922 6928
rect 11885 6919 11943 6925
rect 11885 6885 11897 6919
rect 11931 6885 11943 6919
rect 12820 6916 12848 6956
rect 12894 6944 12900 6996
rect 12952 6984 12958 6996
rect 18782 6984 18788 6996
rect 12952 6956 18788 6984
rect 12952 6944 12958 6956
rect 18782 6944 18788 6956
rect 18840 6944 18846 6996
rect 16390 6916 16396 6928
rect 12820 6888 16396 6916
rect 11885 6879 11943 6885
rect 9766 6848 9772 6860
rect 9140 6820 9772 6848
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 10502 6848 10508 6860
rect 10463 6820 10508 6848
rect 10502 6808 10508 6820
rect 10560 6808 10566 6860
rect 11900 6848 11928 6879
rect 16390 6876 16396 6888
rect 16448 6876 16454 6928
rect 12434 6848 12440 6860
rect 11900 6820 12440 6848
rect 12434 6808 12440 6820
rect 12492 6848 12498 6860
rect 12713 6851 12771 6857
rect 12713 6848 12725 6851
rect 12492 6820 12725 6848
rect 12492 6808 12498 6820
rect 12713 6817 12725 6820
rect 12759 6817 12771 6851
rect 12713 6811 12771 6817
rect 15381 6851 15439 6857
rect 15381 6817 15393 6851
rect 15427 6848 15439 6851
rect 16022 6848 16028 6860
rect 15427 6820 16028 6848
rect 15427 6817 15439 6820
rect 15381 6811 15439 6817
rect 16022 6808 16028 6820
rect 16080 6808 16086 6860
rect 16761 6851 16819 6857
rect 16761 6817 16773 6851
rect 16807 6817 16819 6851
rect 16761 6811 16819 6817
rect 17405 6851 17463 6857
rect 17405 6817 17417 6851
rect 17451 6848 17463 6851
rect 17678 6848 17684 6860
rect 17451 6820 17684 6848
rect 17451 6817 17463 6820
rect 17405 6811 17463 6817
rect 7055 6752 8524 6780
rect 8573 6783 8631 6789
rect 7055 6749 7067 6752
rect 7009 6743 7067 6749
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9309 6783 9367 6789
rect 9309 6780 9321 6783
rect 9180 6752 9321 6780
rect 9180 6740 9186 6752
rect 9309 6749 9321 6752
rect 9355 6749 9367 6783
rect 9309 6743 9367 6749
rect 10045 6783 10103 6789
rect 10045 6749 10057 6783
rect 10091 6780 10103 6783
rect 11790 6780 11796 6792
rect 10091 6752 11796 6780
rect 10091 6749 10103 6752
rect 10045 6743 10103 6749
rect 11790 6740 11796 6752
rect 11848 6740 11854 6792
rect 12526 6780 12532 6792
rect 12487 6752 12532 6780
rect 12526 6740 12532 6752
rect 12584 6740 12590 6792
rect 13446 6780 13452 6792
rect 13407 6752 13452 6780
rect 13446 6740 13452 6752
rect 13504 6740 13510 6792
rect 14921 6783 14979 6789
rect 14921 6749 14933 6783
rect 14967 6780 14979 6783
rect 15194 6780 15200 6792
rect 14967 6752 15200 6780
rect 14967 6749 14979 6752
rect 14921 6743 14979 6749
rect 15194 6740 15200 6752
rect 15252 6740 15258 6792
rect 15562 6780 15568 6792
rect 15523 6752 15568 6780
rect 15562 6740 15568 6752
rect 15620 6740 15626 6792
rect 15746 6740 15752 6792
rect 15804 6780 15810 6792
rect 16776 6780 16804 6811
rect 17678 6808 17684 6820
rect 17736 6808 17742 6860
rect 18230 6848 18236 6860
rect 18191 6820 18236 6848
rect 18230 6808 18236 6820
rect 18288 6808 18294 6860
rect 15804 6752 16804 6780
rect 15804 6740 15810 6752
rect 17494 6740 17500 6792
rect 17552 6780 17558 6792
rect 17589 6783 17647 6789
rect 17589 6780 17601 6783
rect 17552 6752 17601 6780
rect 17552 6740 17558 6752
rect 17589 6749 17601 6752
rect 17635 6749 17647 6783
rect 18874 6780 18880 6792
rect 18835 6752 18880 6780
rect 17589 6743 17647 6749
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19245 6783 19303 6789
rect 19245 6749 19257 6783
rect 19291 6749 19303 6783
rect 19245 6743 19303 6749
rect 6270 6712 6276 6724
rect 6231 6684 6276 6712
rect 6270 6672 6276 6684
rect 6328 6672 6334 6724
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 10750 6715 10808 6721
rect 10750 6712 10762 6715
rect 8536 6684 10762 6712
rect 8536 6672 8542 6684
rect 10750 6681 10762 6684
rect 10796 6681 10808 6715
rect 10750 6675 10808 6681
rect 11238 6672 11244 6724
rect 11296 6712 11302 6724
rect 12621 6715 12679 6721
rect 12621 6712 12633 6715
rect 11296 6684 12633 6712
rect 11296 6672 11302 6684
rect 12621 6681 12633 6684
rect 12667 6681 12679 6715
rect 15838 6712 15844 6724
rect 12621 6675 12679 6681
rect 13648 6684 15844 6712
rect 6733 6647 6791 6653
rect 6733 6613 6745 6647
rect 6779 6644 6791 6647
rect 6822 6644 6828 6656
rect 6779 6616 6828 6644
rect 6779 6613 6791 6616
rect 6733 6607 6791 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7190 6644 7196 6656
rect 7151 6616 7196 6644
rect 7190 6604 7196 6616
rect 7248 6604 7254 6656
rect 7466 6604 7472 6656
rect 7524 6644 7530 6656
rect 7653 6647 7711 6653
rect 7653 6644 7665 6647
rect 7524 6616 7665 6644
rect 7524 6604 7530 6616
rect 7653 6613 7665 6616
rect 7699 6613 7711 6647
rect 9214 6644 9220 6656
rect 9175 6616 9220 6644
rect 7653 6607 7711 6613
rect 9214 6604 9220 6616
rect 9272 6604 9278 6656
rect 10226 6644 10232 6656
rect 10187 6616 10232 6644
rect 10226 6604 10232 6616
rect 10284 6604 10290 6656
rect 11054 6604 11060 6656
rect 11112 6644 11118 6656
rect 13648 6653 13676 6684
rect 15838 6672 15844 6684
rect 15896 6672 15902 6724
rect 16577 6715 16635 6721
rect 16577 6712 16589 6715
rect 15948 6684 16589 6712
rect 12161 6647 12219 6653
rect 12161 6644 12173 6647
rect 11112 6616 12173 6644
rect 11112 6604 11118 6616
rect 12161 6613 12173 6616
rect 12207 6613 12219 6647
rect 12161 6607 12219 6613
rect 13633 6647 13691 6653
rect 13633 6613 13645 6647
rect 13679 6613 13691 6647
rect 13633 6607 13691 6613
rect 13814 6604 13820 6656
rect 13872 6644 13878 6656
rect 14277 6647 14335 6653
rect 14277 6644 14289 6647
rect 13872 6616 14289 6644
rect 13872 6604 13878 6616
rect 14277 6613 14289 6616
rect 14323 6613 14335 6647
rect 15470 6644 15476 6656
rect 15431 6616 15476 6644
rect 14277 6607 14335 6613
rect 15470 6604 15476 6616
rect 15528 6604 15534 6656
rect 15562 6604 15568 6656
rect 15620 6644 15626 6656
rect 15746 6644 15752 6656
rect 15620 6616 15752 6644
rect 15620 6604 15626 6616
rect 15746 6604 15752 6616
rect 15804 6604 15810 6656
rect 15948 6653 15976 6684
rect 16577 6681 16589 6684
rect 16623 6681 16635 6715
rect 16577 6675 16635 6681
rect 17034 6672 17040 6724
rect 17092 6712 17098 6724
rect 19260 6712 19288 6743
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 19392 6752 19809 6780
rect 19392 6740 19398 6752
rect 19797 6749 19809 6752
rect 19843 6780 19855 6783
rect 20530 6780 20536 6792
rect 19843 6752 20536 6780
rect 19843 6749 19855 6752
rect 19797 6743 19855 6749
rect 20530 6740 20536 6752
rect 20588 6740 20594 6792
rect 17092 6684 19288 6712
rect 20064 6715 20122 6721
rect 17092 6672 17098 6684
rect 20064 6681 20076 6715
rect 20110 6712 20122 6715
rect 20162 6712 20168 6724
rect 20110 6684 20168 6712
rect 20110 6681 20122 6684
rect 20064 6675 20122 6681
rect 20162 6672 20168 6684
rect 20220 6672 20226 6724
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6613 15991 6647
rect 15933 6607 15991 6613
rect 16209 6647 16267 6653
rect 16209 6613 16221 6647
rect 16255 6644 16267 6647
rect 16298 6644 16304 6656
rect 16255 6616 16304 6644
rect 16255 6613 16267 6616
rect 16209 6607 16267 6613
rect 16298 6604 16304 6616
rect 16356 6604 16362 6656
rect 16669 6647 16727 6653
rect 16669 6613 16681 6647
rect 16715 6644 16727 6647
rect 17402 6644 17408 6656
rect 16715 6616 17408 6644
rect 16715 6613 16727 6616
rect 16669 6607 16727 6613
rect 17402 6604 17408 6616
rect 17460 6604 17466 6656
rect 17497 6647 17555 6653
rect 17497 6613 17509 6647
rect 17543 6644 17555 6647
rect 17586 6644 17592 6656
rect 17543 6616 17592 6644
rect 17543 6613 17555 6616
rect 17497 6607 17555 6613
rect 17586 6604 17592 6616
rect 17644 6604 17650 6656
rect 17954 6644 17960 6656
rect 17915 6616 17960 6644
rect 17954 6604 17960 6616
rect 18012 6604 18018 6656
rect 18322 6604 18328 6656
rect 18380 6644 18386 6656
rect 19429 6647 19487 6653
rect 19429 6644 19441 6647
rect 18380 6616 19441 6644
rect 18380 6604 18386 6616
rect 19429 6613 19441 6616
rect 19475 6613 19487 6647
rect 19429 6607 19487 6613
rect 21177 6647 21235 6653
rect 21177 6613 21189 6647
rect 21223 6644 21235 6647
rect 21266 6644 21272 6656
rect 21223 6616 21272 6644
rect 21223 6613 21235 6616
rect 21177 6607 21235 6613
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6696 6412 8616 6440
rect 6696 6400 6702 6412
rect 7285 6375 7343 6381
rect 7285 6341 7297 6375
rect 7331 6372 7343 6375
rect 8450 6375 8508 6381
rect 8450 6372 8462 6375
rect 7331 6344 8462 6372
rect 7331 6341 7343 6344
rect 7285 6335 7343 6341
rect 8450 6341 8462 6344
rect 8496 6341 8508 6375
rect 8588 6372 8616 6412
rect 9030 6400 9036 6452
rect 9088 6440 9094 6452
rect 9585 6443 9643 6449
rect 9585 6440 9597 6443
rect 9088 6412 9597 6440
rect 9088 6400 9094 6412
rect 9585 6409 9597 6412
rect 9631 6409 9643 6443
rect 9585 6403 9643 6409
rect 11517 6443 11575 6449
rect 11517 6409 11529 6443
rect 11563 6440 11575 6443
rect 12250 6440 12256 6452
rect 11563 6412 12256 6440
rect 11563 6409 11575 6412
rect 11517 6403 11575 6409
rect 12250 6400 12256 6412
rect 12308 6400 12314 6452
rect 13446 6440 13452 6452
rect 12406 6412 13452 6440
rect 11885 6375 11943 6381
rect 11885 6372 11897 6375
rect 8588 6344 11897 6372
rect 8450 6335 8508 6341
rect 11885 6341 11897 6344
rect 11931 6341 11943 6375
rect 12406 6372 12434 6412
rect 13446 6400 13452 6412
rect 13504 6400 13510 6452
rect 13817 6443 13875 6449
rect 13817 6409 13829 6443
rect 13863 6440 13875 6443
rect 14734 6440 14740 6452
rect 13863 6412 14740 6440
rect 13863 6409 13875 6412
rect 13817 6403 13875 6409
rect 14734 6400 14740 6412
rect 14792 6400 14798 6452
rect 14826 6400 14832 6452
rect 14884 6440 14890 6452
rect 14884 6412 20300 6440
rect 14884 6400 14890 6412
rect 11885 6335 11943 6341
rect 11992 6344 12434 6372
rect 6365 6307 6423 6313
rect 6365 6273 6377 6307
rect 6411 6304 6423 6307
rect 6546 6304 6552 6316
rect 6411 6276 6552 6304
rect 6411 6273 6423 6276
rect 6365 6267 6423 6273
rect 6546 6264 6552 6276
rect 6604 6264 6610 6316
rect 6822 6304 6828 6316
rect 6783 6276 6828 6304
rect 6822 6264 6828 6276
rect 6880 6264 6886 6316
rect 7926 6304 7932 6316
rect 7887 6276 7932 6304
rect 7926 6264 7932 6276
rect 7984 6264 7990 6316
rect 8036 6276 9260 6304
rect 5074 6196 5080 6248
rect 5132 6236 5138 6248
rect 8036 6236 8064 6276
rect 5132 6208 8064 6236
rect 5132 6196 5138 6208
rect 8110 6196 8116 6248
rect 8168 6236 8174 6248
rect 8205 6239 8263 6245
rect 8205 6236 8217 6239
rect 8168 6208 8217 6236
rect 8168 6196 8174 6208
rect 8205 6205 8217 6208
rect 8251 6205 8263 6239
rect 9232 6236 9260 6276
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 10229 6307 10287 6313
rect 10229 6304 10241 6307
rect 9456 6276 10241 6304
rect 9456 6264 9462 6276
rect 10229 6273 10241 6276
rect 10275 6273 10287 6307
rect 10502 6304 10508 6316
rect 10463 6276 10508 6304
rect 10229 6267 10287 6273
rect 10502 6264 10508 6276
rect 10560 6264 10566 6316
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11992 6304 12020 6344
rect 13630 6332 13636 6384
rect 13688 6372 13694 6384
rect 16850 6372 16856 6384
rect 13688 6344 15700 6372
rect 13688 6332 13694 6344
rect 11204 6276 12020 6304
rect 12529 6307 12587 6313
rect 11204 6264 11210 6276
rect 12529 6273 12541 6307
rect 12575 6273 12587 6307
rect 13446 6304 13452 6316
rect 13407 6276 13452 6304
rect 12529 6267 12587 6273
rect 11974 6236 11980 6248
rect 9232 6208 11376 6236
rect 11935 6208 11980 6236
rect 8205 6199 8263 6205
rect 4890 6128 4896 6180
rect 4948 6168 4954 6180
rect 7006 6168 7012 6180
rect 4948 6140 6684 6168
rect 6967 6140 7012 6168
rect 4948 6128 4954 6140
rect 5994 6100 6000 6112
rect 5955 6072 6000 6100
rect 5994 6060 6000 6072
rect 6052 6060 6058 6112
rect 6546 6100 6552 6112
rect 6507 6072 6552 6100
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 6656 6100 6684 6140
rect 7006 6128 7012 6140
rect 7064 6128 7070 6180
rect 10045 6103 10103 6109
rect 10045 6100 10057 6103
rect 6656 6072 10057 6100
rect 10045 6069 10057 6072
rect 10091 6069 10103 6103
rect 10045 6063 10103 6069
rect 10870 6060 10876 6112
rect 10928 6100 10934 6112
rect 11149 6103 11207 6109
rect 11149 6100 11161 6103
rect 10928 6072 11161 6100
rect 10928 6060 10934 6072
rect 11149 6069 11161 6072
rect 11195 6069 11207 6103
rect 11348 6100 11376 6208
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 12069 6239 12127 6245
rect 12069 6205 12081 6239
rect 12115 6205 12127 6239
rect 12544 6236 12572 6267
rect 13446 6264 13452 6276
rect 13504 6264 13510 6316
rect 14918 6313 14924 6316
rect 14093 6307 14151 6313
rect 14093 6304 14105 6307
rect 13556 6276 14105 6304
rect 13170 6236 13176 6248
rect 12069 6199 12127 6205
rect 12176 6208 12572 6236
rect 13131 6208 13176 6236
rect 11606 6128 11612 6180
rect 11664 6168 11670 6180
rect 12084 6168 12112 6199
rect 11664 6140 12112 6168
rect 11664 6128 11670 6140
rect 12176 6100 12204 6208
rect 13170 6196 13176 6208
rect 13228 6196 13234 6248
rect 13354 6236 13360 6248
rect 13315 6208 13360 6236
rect 13354 6196 13360 6208
rect 13412 6196 13418 6248
rect 12250 6128 12256 6180
rect 12308 6168 12314 6180
rect 13556 6168 13584 6276
rect 14093 6273 14105 6276
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 14912 6267 14924 6313
rect 14976 6304 14982 6316
rect 14976 6276 15012 6304
rect 14918 6264 14924 6267
rect 14976 6264 14982 6276
rect 13630 6196 13636 6248
rect 13688 6236 13694 6248
rect 14645 6239 14703 6245
rect 14645 6236 14657 6239
rect 13688 6208 14657 6236
rect 13688 6196 13694 6208
rect 14645 6205 14657 6208
rect 14691 6205 14703 6239
rect 15672 6236 15700 6344
rect 16776 6344 16856 6372
rect 16776 6313 16804 6344
rect 16850 6332 16856 6344
rect 16908 6372 16914 6384
rect 19334 6372 19340 6384
rect 16908 6344 19340 6372
rect 16908 6332 16914 6344
rect 18432 6313 18460 6344
rect 19334 6332 19340 6344
rect 19392 6332 19398 6384
rect 20272 6372 20300 6412
rect 20346 6400 20352 6452
rect 20404 6440 20410 6452
rect 20441 6443 20499 6449
rect 20441 6440 20453 6443
rect 20404 6412 20453 6440
rect 20404 6400 20410 6412
rect 20441 6409 20453 6412
rect 20487 6409 20499 6443
rect 20441 6403 20499 6409
rect 20622 6400 20628 6452
rect 20680 6440 20686 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 20680 6412 21281 6440
rect 20680 6400 20686 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21269 6403 21327 6409
rect 20714 6372 20720 6384
rect 20272 6344 20720 6372
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 16761 6307 16819 6313
rect 16761 6273 16773 6307
rect 16807 6273 16819 6307
rect 17017 6307 17075 6313
rect 17017 6304 17029 6307
rect 16761 6267 16819 6273
rect 16868 6276 17029 6304
rect 16868 6236 16896 6276
rect 17017 6273 17029 6276
rect 17063 6273 17075 6307
rect 17017 6267 17075 6273
rect 18417 6307 18475 6313
rect 18417 6273 18429 6307
rect 18463 6273 18475 6307
rect 18673 6307 18731 6313
rect 18673 6304 18685 6307
rect 18417 6267 18475 6273
rect 18524 6276 18685 6304
rect 18524 6236 18552 6276
rect 18673 6273 18685 6276
rect 18719 6304 18731 6307
rect 19518 6304 19524 6316
rect 18719 6276 19524 6304
rect 18719 6273 18731 6276
rect 18673 6267 18731 6273
rect 19518 6264 19524 6276
rect 19576 6264 19582 6316
rect 20349 6307 20407 6313
rect 20349 6304 20361 6307
rect 19628 6276 20361 6304
rect 15672 6208 16896 6236
rect 18156 6208 18552 6236
rect 14645 6199 14703 6205
rect 18156 6177 18184 6208
rect 18141 6171 18199 6177
rect 12308 6140 13584 6168
rect 14200 6140 14688 6168
rect 12308 6128 12314 6140
rect 11348 6072 12204 6100
rect 12713 6103 12771 6109
rect 11149 6063 11207 6069
rect 12713 6069 12725 6103
rect 12759 6100 12771 6103
rect 14200 6100 14228 6140
rect 12759 6072 14228 6100
rect 14277 6103 14335 6109
rect 12759 6069 12771 6072
rect 12713 6063 12771 6069
rect 14277 6069 14289 6103
rect 14323 6100 14335 6103
rect 14550 6100 14556 6112
rect 14323 6072 14556 6100
rect 14323 6069 14335 6072
rect 14277 6063 14335 6069
rect 14550 6060 14556 6072
rect 14608 6060 14614 6112
rect 14660 6100 14688 6140
rect 18141 6137 18153 6171
rect 18187 6137 18199 6171
rect 18141 6131 18199 6137
rect 15746 6100 15752 6112
rect 14660 6072 15752 6100
rect 15746 6060 15752 6072
rect 15804 6060 15810 6112
rect 16022 6100 16028 6112
rect 15983 6072 16028 6100
rect 16022 6060 16028 6072
rect 16080 6060 16086 6112
rect 16114 6060 16120 6112
rect 16172 6100 16178 6112
rect 19628 6100 19656 6276
rect 20349 6273 20361 6276
rect 20395 6273 20407 6307
rect 21082 6304 21088 6316
rect 21043 6276 21088 6304
rect 20349 6267 20407 6273
rect 21082 6264 21088 6276
rect 21140 6264 21146 6316
rect 20257 6239 20315 6245
rect 20257 6205 20269 6239
rect 20303 6205 20315 6239
rect 20257 6199 20315 6205
rect 19797 6171 19855 6177
rect 19797 6137 19809 6171
rect 19843 6168 19855 6171
rect 20272 6168 20300 6199
rect 21174 6168 21180 6180
rect 19843 6140 21180 6168
rect 19843 6137 19855 6140
rect 19797 6131 19855 6137
rect 21174 6128 21180 6140
rect 21232 6128 21238 6180
rect 20806 6100 20812 6112
rect 16172 6072 19656 6100
rect 20767 6072 20812 6100
rect 16172 6060 16178 6072
rect 20806 6060 20812 6072
rect 20864 6060 20870 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 4522 5856 4528 5908
rect 4580 5896 4586 5908
rect 4982 5896 4988 5908
rect 4580 5868 4988 5896
rect 4580 5856 4586 5868
rect 4982 5856 4988 5868
rect 5040 5896 5046 5908
rect 5169 5899 5227 5905
rect 5169 5896 5181 5899
rect 5040 5868 5181 5896
rect 5040 5856 5046 5868
rect 5169 5865 5181 5868
rect 5215 5865 5227 5899
rect 5626 5896 5632 5908
rect 5587 5868 5632 5896
rect 5169 5859 5227 5865
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 5997 5899 6055 5905
rect 5997 5865 6009 5899
rect 6043 5896 6055 5899
rect 7834 5896 7840 5908
rect 6043 5868 7840 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 7834 5856 7840 5868
rect 7892 5856 7898 5908
rect 7926 5856 7932 5908
rect 7984 5896 7990 5908
rect 8573 5899 8631 5905
rect 8573 5896 8585 5899
rect 7984 5868 8585 5896
rect 7984 5856 7990 5868
rect 8573 5865 8585 5868
rect 8619 5865 8631 5899
rect 8573 5859 8631 5865
rect 8941 5899 8999 5905
rect 8941 5865 8953 5899
rect 8987 5896 8999 5899
rect 9214 5896 9220 5908
rect 8987 5868 9220 5896
rect 8987 5865 8999 5868
rect 8941 5859 8999 5865
rect 2498 5788 2504 5840
rect 2556 5828 2562 5840
rect 2556 5800 2774 5828
rect 2556 5788 2562 5800
rect 2746 5624 2774 5800
rect 5902 5720 5908 5772
rect 5960 5760 5966 5772
rect 8588 5760 8616 5859
rect 9214 5856 9220 5868
rect 9272 5856 9278 5908
rect 12250 5896 12256 5908
rect 9324 5868 12256 5896
rect 8754 5788 8760 5840
rect 8812 5828 8818 5840
rect 9324 5828 9352 5868
rect 12250 5856 12256 5868
rect 12308 5856 12314 5908
rect 13078 5896 13084 5908
rect 13039 5868 13084 5896
rect 13078 5856 13084 5868
rect 13136 5856 13142 5908
rect 13446 5856 13452 5908
rect 13504 5896 13510 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13504 5868 14105 5896
rect 13504 5856 13510 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 17034 5896 17040 5908
rect 14093 5859 14151 5865
rect 14384 5868 17040 5896
rect 8812 5800 9352 5828
rect 10137 5831 10195 5837
rect 8812 5788 8818 5800
rect 10137 5797 10149 5831
rect 10183 5828 10195 5831
rect 14384 5828 14412 5868
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17402 5856 17408 5908
rect 17460 5896 17466 5908
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 17460 5868 17693 5896
rect 17460 5856 17466 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 17770 5856 17776 5908
rect 17828 5896 17834 5908
rect 20625 5899 20683 5905
rect 17828 5868 20576 5896
rect 17828 5856 17834 5868
rect 18874 5828 18880 5840
rect 10183 5800 14412 5828
rect 14476 5800 18880 5828
rect 10183 5797 10195 5800
rect 10137 5791 10195 5797
rect 9493 5763 9551 5769
rect 9493 5760 9505 5763
rect 5960 5732 7328 5760
rect 8588 5732 9505 5760
rect 5960 5720 5966 5732
rect 6914 5692 6920 5704
rect 6875 5664 6920 5692
rect 6914 5652 6920 5664
rect 6972 5652 6978 5704
rect 7190 5692 7196 5704
rect 7151 5664 7196 5692
rect 7190 5652 7196 5664
rect 7248 5652 7254 5704
rect 7300 5692 7328 5732
rect 9493 5729 9505 5732
rect 9539 5729 9551 5763
rect 14476 5760 14504 5800
rect 18874 5788 18880 5800
rect 18932 5788 18938 5840
rect 20548 5828 20576 5868
rect 20625 5865 20637 5899
rect 20671 5896 20683 5899
rect 20990 5896 20996 5908
rect 20671 5868 20996 5896
rect 20671 5865 20683 5868
rect 20625 5859 20683 5865
rect 20990 5856 20996 5868
rect 21048 5896 21054 5908
rect 21634 5896 21640 5908
rect 21048 5868 21640 5896
rect 21048 5856 21054 5868
rect 21634 5856 21640 5868
rect 21692 5856 21698 5908
rect 22646 5828 22652 5840
rect 20548 5800 22652 5828
rect 22646 5788 22652 5800
rect 22704 5788 22710 5840
rect 9493 5723 9551 5729
rect 9600 5732 14504 5760
rect 7300 5664 7604 5692
rect 6273 5627 6331 5633
rect 2746 5596 6040 5624
rect 1854 5516 1860 5568
rect 1912 5556 1918 5568
rect 4614 5556 4620 5568
rect 1912 5528 4620 5556
rect 1912 5516 1918 5528
rect 4614 5516 4620 5528
rect 4672 5516 4678 5568
rect 4798 5556 4804 5568
rect 4759 5528 4804 5556
rect 4798 5516 4804 5528
rect 4856 5516 4862 5568
rect 6012 5556 6040 5596
rect 6273 5593 6285 5627
rect 6319 5624 6331 5627
rect 7438 5627 7496 5633
rect 7438 5624 7450 5627
rect 6319 5596 7450 5624
rect 6319 5593 6331 5596
rect 6273 5587 6331 5593
rect 7438 5593 7450 5596
rect 7484 5593 7496 5627
rect 7576 5624 7604 5664
rect 7834 5652 7840 5704
rect 7892 5692 7898 5704
rect 9600 5692 9628 5732
rect 14550 5720 14556 5772
rect 14608 5760 14614 5772
rect 14737 5763 14795 5769
rect 14737 5760 14749 5763
rect 14608 5732 14749 5760
rect 14608 5720 14614 5732
rect 14737 5729 14749 5732
rect 14783 5760 14795 5763
rect 15194 5760 15200 5772
rect 14783 5732 15200 5760
rect 14783 5729 14795 5732
rect 14737 5723 14795 5729
rect 15194 5720 15200 5732
rect 15252 5720 15258 5772
rect 16022 5720 16028 5772
rect 16080 5760 16086 5772
rect 18233 5763 18291 5769
rect 18233 5760 18245 5763
rect 16080 5732 18245 5760
rect 16080 5720 16086 5732
rect 18233 5729 18245 5732
rect 18279 5729 18291 5763
rect 18233 5723 18291 5729
rect 7892 5664 9628 5692
rect 7892 5652 7898 5664
rect 9674 5652 9680 5704
rect 9732 5692 9738 5704
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9732 5664 9965 5692
rect 9732 5652 9738 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10502 5652 10508 5704
rect 10560 5692 10566 5704
rect 11606 5692 11612 5704
rect 10560 5664 11612 5692
rect 10560 5652 10566 5664
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 12158 5692 12164 5704
rect 12119 5664 12164 5692
rect 12158 5652 12164 5664
rect 12216 5652 12222 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 12492 5664 12537 5692
rect 12492 5652 12498 5664
rect 12618 5652 12624 5704
rect 12676 5692 12682 5704
rect 13449 5695 13507 5701
rect 13449 5692 13461 5695
rect 12676 5664 13461 5692
rect 12676 5652 12682 5664
rect 13449 5661 13461 5664
rect 13495 5661 13507 5695
rect 15102 5692 15108 5704
rect 15063 5664 15108 5692
rect 13449 5655 13507 5661
rect 15102 5652 15108 5664
rect 15160 5652 15166 5704
rect 15654 5692 15660 5704
rect 15615 5664 15660 5692
rect 15654 5652 15660 5664
rect 15712 5652 15718 5704
rect 18138 5692 18144 5704
rect 17328 5664 18144 5692
rect 8754 5624 8760 5636
rect 7576 5596 8760 5624
rect 7438 5587 7496 5593
rect 8754 5584 8760 5596
rect 8812 5584 8818 5636
rect 9490 5584 9496 5636
rect 9548 5624 9554 5636
rect 17328 5624 17356 5664
rect 18138 5652 18144 5664
rect 18196 5652 18202 5704
rect 18874 5692 18880 5704
rect 18835 5664 18880 5692
rect 18874 5652 18880 5664
rect 18932 5652 18938 5704
rect 19245 5695 19303 5701
rect 19245 5661 19257 5695
rect 19291 5692 19303 5695
rect 20530 5692 20536 5704
rect 19291 5664 20536 5692
rect 19291 5661 19303 5664
rect 19245 5655 19303 5661
rect 9548 5596 17356 5624
rect 9548 5584 9554 5596
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 19260 5624 19288 5655
rect 20530 5652 20536 5664
rect 20588 5652 20594 5704
rect 20898 5692 20904 5704
rect 20859 5664 20904 5692
rect 20898 5652 20904 5664
rect 20956 5652 20962 5704
rect 17460 5596 19288 5624
rect 19512 5627 19570 5633
rect 17460 5584 17466 5596
rect 19512 5593 19524 5627
rect 19558 5624 19570 5627
rect 21174 5624 21180 5636
rect 19558 5596 19656 5624
rect 19558 5593 19570 5596
rect 19512 5587 19570 5593
rect 9309 5559 9367 5565
rect 9309 5556 9321 5559
rect 6012 5528 9321 5556
rect 9309 5525 9321 5528
rect 9355 5525 9367 5559
rect 9309 5519 9367 5525
rect 9401 5559 9459 5565
rect 9401 5525 9413 5559
rect 9447 5556 9459 5559
rect 9582 5556 9588 5568
rect 9447 5528 9588 5556
rect 9447 5525 9459 5528
rect 9401 5519 9459 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10873 5559 10931 5565
rect 10873 5525 10885 5559
rect 10919 5556 10931 5559
rect 11054 5556 11060 5568
rect 10919 5528 11060 5556
rect 10919 5525 10931 5528
rect 10873 5519 10931 5525
rect 11054 5516 11060 5528
rect 11112 5516 11118 5568
rect 13633 5559 13691 5565
rect 13633 5525 13645 5559
rect 13679 5556 13691 5559
rect 13722 5556 13728 5568
rect 13679 5528 13728 5556
rect 13679 5525 13691 5528
rect 13633 5519 13691 5525
rect 13722 5516 13728 5528
rect 13780 5516 13786 5568
rect 14458 5556 14464 5568
rect 14419 5528 14464 5556
rect 14458 5516 14464 5528
rect 14516 5516 14522 5568
rect 14553 5559 14611 5565
rect 14553 5525 14565 5559
rect 14599 5556 14611 5559
rect 14642 5556 14648 5568
rect 14599 5528 14648 5556
rect 14599 5525 14611 5528
rect 14553 5519 14611 5525
rect 14642 5516 14648 5528
rect 14700 5516 14706 5568
rect 15289 5559 15347 5565
rect 15289 5525 15301 5559
rect 15335 5556 15347 5559
rect 17586 5556 17592 5568
rect 15335 5528 17592 5556
rect 15335 5525 15347 5528
rect 15289 5519 15347 5525
rect 17586 5516 17592 5528
rect 17644 5516 17650 5568
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18049 5559 18107 5565
rect 18049 5556 18061 5559
rect 17828 5528 18061 5556
rect 17828 5516 17834 5528
rect 18049 5525 18061 5528
rect 18095 5525 18107 5559
rect 18049 5519 18107 5525
rect 18138 5516 18144 5568
rect 18196 5556 18202 5568
rect 18690 5556 18696 5568
rect 18196 5528 18241 5556
rect 18651 5528 18696 5556
rect 18196 5516 18202 5528
rect 18690 5516 18696 5528
rect 18748 5516 18754 5568
rect 19628 5556 19656 5596
rect 19812 5596 21180 5624
rect 19812 5556 19840 5596
rect 21174 5584 21180 5596
rect 21232 5584 21238 5636
rect 21082 5556 21088 5568
rect 19628 5528 19840 5556
rect 21043 5528 21088 5556
rect 21082 5516 21088 5528
rect 21140 5516 21146 5568
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 5997 5355 6055 5361
rect 5997 5321 6009 5355
rect 6043 5352 6055 5355
rect 6638 5352 6644 5364
rect 6043 5324 6644 5352
rect 6043 5321 6055 5324
rect 5997 5315 6055 5321
rect 6638 5312 6644 5324
rect 6696 5312 6702 5364
rect 6917 5355 6975 5361
rect 6917 5321 6929 5355
rect 6963 5352 6975 5355
rect 8202 5352 8208 5364
rect 6963 5324 8208 5352
rect 6963 5321 6975 5324
rect 6917 5315 6975 5321
rect 8202 5312 8208 5324
rect 8260 5312 8266 5364
rect 9769 5355 9827 5361
rect 9769 5321 9781 5355
rect 9815 5352 9827 5355
rect 10502 5352 10508 5364
rect 9815 5324 10508 5352
rect 9815 5321 9827 5324
rect 9769 5315 9827 5321
rect 10502 5312 10508 5324
rect 10560 5312 10566 5364
rect 12066 5312 12072 5364
rect 12124 5352 12130 5364
rect 12253 5355 12311 5361
rect 12253 5352 12265 5355
rect 12124 5324 12265 5352
rect 12124 5312 12130 5324
rect 12253 5321 12265 5324
rect 12299 5352 12311 5355
rect 13170 5352 13176 5364
rect 12299 5324 13176 5352
rect 12299 5321 12311 5324
rect 12253 5315 12311 5321
rect 13170 5312 13176 5324
rect 13228 5312 13234 5364
rect 13354 5312 13360 5364
rect 13412 5352 13418 5364
rect 13909 5355 13967 5361
rect 13909 5352 13921 5355
rect 13412 5324 13921 5352
rect 13412 5312 13418 5324
rect 13909 5321 13921 5324
rect 13955 5321 13967 5355
rect 13909 5315 13967 5321
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18325 5355 18383 5361
rect 18325 5352 18337 5355
rect 18196 5324 18337 5352
rect 18196 5312 18202 5324
rect 18325 5321 18337 5324
rect 18371 5321 18383 5355
rect 19886 5352 19892 5364
rect 18325 5315 18383 5321
rect 18800 5324 19892 5352
rect 6454 5284 6460 5296
rect 6415 5256 6460 5284
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 7190 5244 7196 5296
rect 7248 5284 7254 5296
rect 7742 5284 7748 5296
rect 7248 5256 7748 5284
rect 7248 5244 7254 5256
rect 7742 5244 7748 5256
rect 7800 5284 7806 5296
rect 8110 5284 8116 5296
rect 7800 5256 8116 5284
rect 7800 5244 7806 5256
rect 8110 5244 8116 5256
rect 8168 5284 8174 5296
rect 11054 5284 11060 5296
rect 8168 5256 11060 5284
rect 8168 5244 8174 5256
rect 5353 5219 5411 5225
rect 5353 5185 5365 5219
rect 5399 5216 5411 5219
rect 5442 5216 5448 5228
rect 5399 5188 5448 5216
rect 5399 5185 5411 5188
rect 5353 5179 5411 5185
rect 5442 5176 5448 5188
rect 5500 5176 5506 5228
rect 6730 5216 6736 5228
rect 6691 5188 6736 5216
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 8588 5225 8616 5256
rect 11054 5244 11060 5256
rect 11112 5284 11118 5296
rect 13814 5284 13820 5296
rect 11112 5256 11192 5284
rect 11112 5244 11118 5256
rect 8317 5219 8375 5225
rect 8317 5185 8329 5219
rect 8363 5216 8375 5219
rect 8573 5219 8631 5225
rect 8363 5188 8524 5216
rect 8363 5185 8375 5188
rect 8317 5179 8375 5185
rect 8496 5148 8524 5188
rect 8573 5185 8585 5219
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 9582 5216 9588 5228
rect 9539 5188 9588 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 11164 5225 11192 5256
rect 13464 5256 13820 5284
rect 10893 5219 10951 5225
rect 10893 5185 10905 5219
rect 10939 5216 10951 5219
rect 11149 5219 11207 5225
rect 10939 5188 11100 5216
rect 10939 5185 10951 5188
rect 10893 5179 10951 5185
rect 8849 5151 8907 5157
rect 8849 5148 8861 5151
rect 8496 5120 8861 5148
rect 8849 5117 8861 5120
rect 8895 5117 8907 5151
rect 11072 5148 11100 5188
rect 11149 5185 11161 5219
rect 11195 5185 11207 5219
rect 11149 5179 11207 5185
rect 11977 5219 12035 5225
rect 11977 5185 11989 5219
rect 12023 5216 12035 5219
rect 12158 5216 12164 5228
rect 12023 5188 12164 5216
rect 12023 5185 12035 5188
rect 11977 5179 12035 5185
rect 12158 5176 12164 5188
rect 12216 5176 12222 5228
rect 13377 5219 13435 5225
rect 13377 5185 13389 5219
rect 13423 5216 13435 5219
rect 13464 5216 13492 5256
rect 13814 5244 13820 5256
rect 13872 5244 13878 5296
rect 14182 5244 14188 5296
rect 14240 5284 14246 5296
rect 14369 5287 14427 5293
rect 14369 5284 14381 5287
rect 14240 5256 14381 5284
rect 14240 5244 14246 5256
rect 14369 5253 14381 5256
rect 14415 5284 14427 5287
rect 14826 5284 14832 5296
rect 14415 5256 14832 5284
rect 14415 5253 14427 5256
rect 14369 5247 14427 5253
rect 14826 5244 14832 5256
rect 14884 5244 14890 5296
rect 16022 5244 16028 5296
rect 16080 5293 16086 5296
rect 16080 5284 16092 5293
rect 17402 5284 17408 5296
rect 16080 5256 16125 5284
rect 16316 5256 17408 5284
rect 16080 5247 16092 5256
rect 16080 5244 16086 5247
rect 13630 5216 13636 5228
rect 13423 5188 13492 5216
rect 13591 5188 13636 5216
rect 13423 5185 13435 5188
rect 13377 5179 13435 5185
rect 13630 5176 13636 5188
rect 13688 5176 13694 5228
rect 14274 5216 14280 5228
rect 14235 5188 14280 5216
rect 14274 5176 14280 5188
rect 14332 5176 14338 5228
rect 15010 5176 15016 5228
rect 15068 5216 15074 5228
rect 16316 5225 16344 5256
rect 17402 5244 17408 5256
rect 17460 5244 17466 5296
rect 18230 5244 18236 5296
rect 18288 5284 18294 5296
rect 18800 5293 18828 5324
rect 19886 5312 19892 5324
rect 19944 5312 19950 5364
rect 20349 5355 20407 5361
rect 20349 5321 20361 5355
rect 20395 5352 20407 5355
rect 20438 5352 20444 5364
rect 20395 5324 20444 5352
rect 20395 5321 20407 5324
rect 20349 5315 20407 5321
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 20717 5355 20775 5361
rect 20717 5321 20729 5355
rect 20763 5352 20775 5355
rect 20806 5352 20812 5364
rect 20763 5324 20812 5352
rect 20763 5321 20775 5324
rect 20717 5315 20775 5321
rect 20806 5312 20812 5324
rect 20864 5312 20870 5364
rect 18785 5287 18843 5293
rect 18785 5284 18797 5287
rect 18288 5256 18797 5284
rect 18288 5244 18294 5256
rect 18785 5253 18797 5256
rect 18831 5253 18843 5287
rect 18785 5247 18843 5253
rect 16301 5219 16359 5225
rect 15068 5188 16252 5216
rect 15068 5176 15074 5188
rect 11606 5148 11612 5160
rect 11072 5120 11612 5148
rect 8849 5111 8907 5117
rect 11606 5108 11612 5120
rect 11664 5108 11670 5160
rect 14550 5148 14556 5160
rect 14511 5120 14556 5148
rect 14550 5108 14556 5120
rect 14608 5108 14614 5160
rect 16224 5148 16252 5188
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16390 5176 16396 5228
rect 16448 5216 16454 5228
rect 17034 5216 17040 5228
rect 16448 5188 16896 5216
rect 16995 5188 17040 5216
rect 16448 5176 16454 5188
rect 16868 5160 16896 5188
rect 17034 5176 17040 5188
rect 17092 5176 17098 5228
rect 17678 5216 17684 5228
rect 17639 5188 17684 5216
rect 17678 5176 17684 5188
rect 17736 5176 17742 5228
rect 18598 5176 18604 5228
rect 18656 5216 18662 5228
rect 18693 5219 18751 5225
rect 18693 5216 18705 5219
rect 18656 5188 18705 5216
rect 18656 5176 18662 5188
rect 18693 5185 18705 5188
rect 18739 5185 18751 5219
rect 19702 5216 19708 5228
rect 19663 5188 19708 5216
rect 18693 5179 18751 5185
rect 19702 5176 19708 5188
rect 19760 5176 19766 5228
rect 16761 5151 16819 5157
rect 16761 5148 16773 5151
rect 16224 5120 16773 5148
rect 16761 5117 16773 5120
rect 16807 5117 16819 5151
rect 16761 5111 16819 5117
rect 3605 5083 3663 5089
rect 3605 5049 3617 5083
rect 3651 5080 3663 5083
rect 4338 5080 4344 5092
rect 3651 5052 4344 5080
rect 3651 5049 3663 5052
rect 3605 5043 3663 5049
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 5537 5083 5595 5089
rect 5537 5049 5549 5083
rect 5583 5080 5595 5083
rect 11793 5083 11851 5089
rect 5583 5052 7696 5080
rect 5583 5049 5595 5052
rect 5537 5043 5595 5049
rect 1394 5012 1400 5024
rect 1355 4984 1400 5012
rect 1394 4972 1400 4984
rect 1452 4972 1458 5024
rect 4246 5012 4252 5024
rect 4207 4984 4252 5012
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 4982 5012 4988 5024
rect 4943 4984 4988 5012
rect 4982 4972 4988 4984
rect 5040 4972 5046 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6972 4984 7205 5012
rect 6972 4972 6978 4984
rect 7193 4981 7205 4984
rect 7239 5012 7251 5015
rect 7558 5012 7564 5024
rect 7239 4984 7564 5012
rect 7239 4981 7251 4984
rect 7193 4975 7251 4981
rect 7558 4972 7564 4984
rect 7616 4972 7622 5024
rect 7668 5012 7696 5052
rect 11793 5049 11805 5083
rect 11839 5080 11851 5083
rect 12434 5080 12440 5092
rect 11839 5052 12440 5080
rect 11839 5049 11851 5052
rect 11793 5043 11851 5049
rect 12434 5040 12440 5052
rect 12492 5040 12498 5092
rect 16776 5080 16804 5111
rect 16850 5108 16856 5160
rect 16908 5148 16914 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16908 5120 16957 5148
rect 16908 5108 16914 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 18877 5151 18935 5157
rect 16945 5111 17003 5117
rect 17052 5120 18736 5148
rect 17052 5080 17080 5120
rect 16776 5052 17080 5080
rect 17405 5083 17463 5089
rect 17405 5049 17417 5083
rect 17451 5080 17463 5083
rect 17770 5080 17776 5092
rect 17451 5052 17776 5080
rect 17451 5049 17463 5052
rect 17405 5043 17463 5049
rect 17770 5040 17776 5052
rect 17828 5040 17834 5092
rect 18708 5080 18736 5120
rect 18877 5117 18889 5151
rect 18923 5117 18935 5151
rect 19518 5148 19524 5160
rect 19479 5120 19524 5148
rect 18877 5111 18935 5117
rect 18892 5080 18920 5111
rect 19518 5108 19524 5120
rect 19576 5108 19582 5160
rect 19613 5151 19671 5157
rect 19613 5117 19625 5151
rect 19659 5148 19671 5151
rect 20254 5148 20260 5160
rect 19659 5120 20260 5148
rect 19659 5117 19671 5120
rect 19613 5111 19671 5117
rect 20254 5108 20260 5120
rect 20312 5108 20318 5160
rect 20530 5108 20536 5160
rect 20588 5148 20594 5160
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20588 5120 20821 5148
rect 20588 5108 20594 5120
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20990 5148 20996 5160
rect 20951 5120 20996 5148
rect 20809 5111 20867 5117
rect 20990 5108 20996 5120
rect 21048 5108 21054 5160
rect 18708 5052 18920 5080
rect 9858 5012 9864 5024
rect 7668 4984 9864 5012
rect 9858 4972 9864 4984
rect 9916 4972 9922 5024
rect 10042 4972 10048 5024
rect 10100 5012 10106 5024
rect 14921 5015 14979 5021
rect 14921 5012 14933 5015
rect 10100 4984 14933 5012
rect 10100 4972 10106 4984
rect 14921 4981 14933 4984
rect 14967 5012 14979 5015
rect 15562 5012 15568 5024
rect 14967 4984 15568 5012
rect 14967 4981 14979 4984
rect 14921 4975 14979 4981
rect 15562 4972 15568 4984
rect 15620 4972 15626 5024
rect 16942 4972 16948 5024
rect 17000 5012 17006 5024
rect 17865 5015 17923 5021
rect 17865 5012 17877 5015
rect 17000 4984 17877 5012
rect 17000 4972 17006 4984
rect 17865 4981 17877 4984
rect 17911 4981 17923 5015
rect 20070 5012 20076 5024
rect 20031 4984 20076 5012
rect 17865 4975 17923 4981
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 3970 4808 3976 4820
rect 3931 4780 3976 4808
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 5169 4811 5227 4817
rect 5169 4777 5181 4811
rect 5215 4808 5227 4811
rect 5534 4808 5540 4820
rect 5215 4780 5540 4808
rect 5215 4777 5227 4780
rect 5169 4771 5227 4777
rect 5534 4768 5540 4780
rect 5592 4768 5598 4820
rect 5629 4811 5687 4817
rect 5629 4777 5641 4811
rect 5675 4808 5687 4811
rect 8570 4808 8576 4820
rect 5675 4780 8493 4808
rect 8531 4780 8576 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 4430 4700 4436 4752
rect 4488 4740 4494 4752
rect 8294 4740 8300 4752
rect 4488 4712 8300 4740
rect 4488 4700 4494 4712
rect 8294 4700 8300 4712
rect 8352 4700 8358 4752
rect 8465 4740 8493 4780
rect 8570 4768 8576 4780
rect 8628 4768 8634 4820
rect 9033 4811 9091 4817
rect 9033 4777 9045 4811
rect 9079 4808 9091 4811
rect 9398 4808 9404 4820
rect 9079 4780 9404 4808
rect 9079 4777 9091 4780
rect 9033 4771 9091 4777
rect 9398 4768 9404 4780
rect 9456 4768 9462 4820
rect 11146 4808 11152 4820
rect 9646 4780 11152 4808
rect 9646 4740 9674 4780
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 11606 4768 11612 4820
rect 11664 4808 11670 4820
rect 14737 4811 14795 4817
rect 14737 4808 14749 4811
rect 11664 4780 14749 4808
rect 11664 4768 11670 4780
rect 14737 4777 14749 4780
rect 14783 4777 14795 4811
rect 14737 4771 14795 4777
rect 15470 4768 15476 4820
rect 15528 4808 15534 4820
rect 15749 4811 15807 4817
rect 15749 4808 15761 4811
rect 15528 4780 15761 4808
rect 15528 4768 15534 4780
rect 15749 4777 15761 4780
rect 15795 4777 15807 4811
rect 15749 4771 15807 4777
rect 16316 4780 18276 4808
rect 8465 4712 9674 4740
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 7009 4675 7067 4681
rect 3016 4644 6684 4672
rect 3016 4632 3022 4644
rect 4709 4607 4767 4613
rect 4709 4573 4721 4607
rect 4755 4604 4767 4607
rect 4985 4607 5043 4613
rect 4985 4604 4997 4607
rect 4755 4576 4997 4604
rect 4755 4573 4767 4576
rect 4709 4567 4767 4573
rect 4985 4573 4997 4576
rect 5031 4604 5043 4607
rect 5350 4604 5356 4616
rect 5031 4576 5356 4604
rect 5031 4573 5043 4576
rect 4985 4567 5043 4573
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5442 4564 5448 4616
rect 5500 4604 5506 4616
rect 6546 4604 6552 4616
rect 5500 4576 5545 4604
rect 6507 4576 6552 4604
rect 5500 4564 5506 4576
rect 6546 4564 6552 4576
rect 6604 4564 6610 4616
rect 6656 4604 6684 4644
rect 7009 4641 7021 4675
rect 7055 4672 7067 4675
rect 7055 4644 7512 4672
rect 7055 4641 7067 4644
rect 7009 4635 7067 4641
rect 7193 4607 7251 4613
rect 7193 4604 7205 4607
rect 6656 4576 7205 4604
rect 7193 4573 7205 4576
rect 7239 4573 7251 4607
rect 7193 4567 7251 4573
rect 1670 4496 1676 4548
rect 1728 4536 1734 4548
rect 2041 4539 2099 4545
rect 2041 4536 2053 4539
rect 1728 4508 2053 4536
rect 1728 4496 1734 4508
rect 2041 4505 2053 4508
rect 2087 4505 2099 4539
rect 2041 4499 2099 4505
rect 4341 4539 4399 4545
rect 4341 4505 4353 4539
rect 4387 4536 4399 4539
rect 5810 4536 5816 4548
rect 4387 4508 5816 4536
rect 4387 4505 4399 4508
rect 4341 4499 4399 4505
rect 5810 4496 5816 4508
rect 5868 4496 5874 4548
rect 7098 4536 7104 4548
rect 7059 4508 7104 4536
rect 7098 4496 7104 4508
rect 7156 4496 7162 4548
rect 7484 4536 7512 4644
rect 7558 4632 7564 4684
rect 7616 4672 7622 4684
rect 7929 4675 7987 4681
rect 7929 4672 7941 4675
rect 7616 4644 7941 4672
rect 7616 4632 7622 4644
rect 7929 4641 7941 4644
rect 7975 4641 7987 4675
rect 12345 4675 12403 4681
rect 12345 4672 12357 4675
rect 7929 4635 7987 4641
rect 11164 4644 12357 4672
rect 7650 4564 7656 4616
rect 7708 4604 7714 4616
rect 8205 4607 8263 4613
rect 8205 4604 8217 4607
rect 7708 4576 8217 4604
rect 7708 4564 7714 4576
rect 8205 4573 8217 4576
rect 8251 4573 8263 4607
rect 8205 4567 8263 4573
rect 8386 4564 8392 4616
rect 8444 4604 8450 4616
rect 9122 4604 9128 4616
rect 8444 4576 9128 4604
rect 8444 4564 8450 4576
rect 9122 4564 9128 4576
rect 9180 4564 9186 4616
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9456 4576 9505 4604
rect 9456 4564 9462 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 10870 4564 10876 4616
rect 10928 4613 10934 4616
rect 10928 4604 10940 4613
rect 10928 4576 10973 4604
rect 10928 4567 10940 4576
rect 10928 4564 10934 4567
rect 11054 4564 11060 4616
rect 11112 4604 11118 4616
rect 11164 4613 11192 4644
rect 12345 4641 12357 4644
rect 12391 4641 12403 4675
rect 12345 4635 12403 4641
rect 11149 4607 11207 4613
rect 11149 4604 11161 4607
rect 11112 4576 11161 4604
rect 11112 4564 11118 4576
rect 11149 4573 11161 4576
rect 11195 4573 11207 4607
rect 12066 4604 12072 4616
rect 12027 4576 12072 4604
rect 11149 4567 11207 4573
rect 12066 4564 12072 4576
rect 12124 4564 12130 4616
rect 12360 4604 12388 4635
rect 14918 4632 14924 4684
rect 14976 4672 14982 4684
rect 16316 4681 16344 4780
rect 17126 4740 17132 4752
rect 16592 4712 17132 4740
rect 15197 4675 15255 4681
rect 15197 4672 15209 4675
rect 14976 4644 15209 4672
rect 14976 4632 14982 4644
rect 15197 4641 15209 4644
rect 15243 4641 15255 4675
rect 15197 4635 15255 4641
rect 16301 4675 16359 4681
rect 16301 4641 16313 4675
rect 16347 4641 16359 4675
rect 16301 4635 16359 4641
rect 13630 4604 13636 4616
rect 12360 4576 13636 4604
rect 13630 4564 13636 4576
rect 13688 4564 13694 4616
rect 14093 4607 14151 4613
rect 14093 4604 14105 4607
rect 13740 4576 14105 4604
rect 9582 4536 9588 4548
rect 7484 4508 9588 4536
rect 9582 4496 9588 4508
rect 9640 4536 9646 4548
rect 11425 4539 11483 4545
rect 9640 4508 9812 4536
rect 9640 4496 9646 4508
rect 1762 4468 1768 4480
rect 1723 4440 1768 4468
rect 1762 4428 1768 4440
rect 1820 4428 1826 4480
rect 2314 4428 2320 4480
rect 2372 4468 2378 4480
rect 2593 4471 2651 4477
rect 2593 4468 2605 4471
rect 2372 4440 2605 4468
rect 2372 4428 2378 4440
rect 2593 4437 2605 4440
rect 2639 4437 2651 4471
rect 3050 4468 3056 4480
rect 3011 4440 3056 4468
rect 2593 4431 2651 4437
rect 3050 4428 3056 4440
rect 3108 4428 3114 4480
rect 3418 4468 3424 4480
rect 3379 4440 3424 4468
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 5905 4471 5963 4477
rect 5905 4437 5917 4471
rect 5951 4468 5963 4471
rect 7006 4468 7012 4480
rect 5951 4440 7012 4468
rect 5951 4437 5963 4440
rect 5905 4431 5963 4437
rect 7006 4428 7012 4440
rect 7064 4428 7070 4480
rect 7561 4471 7619 4477
rect 7561 4437 7573 4471
rect 7607 4468 7619 4471
rect 8113 4471 8171 4477
rect 8113 4468 8125 4471
rect 7607 4440 8125 4468
rect 7607 4437 7619 4440
rect 7561 4431 7619 4437
rect 8113 4437 8125 4440
rect 8159 4437 8171 4471
rect 8113 4431 8171 4437
rect 8294 4428 8300 4480
rect 8352 4468 8358 4480
rect 9784 4477 9812 4508
rect 11425 4505 11437 4539
rect 11471 4536 11483 4539
rect 12590 4539 12648 4545
rect 12590 4536 12602 4539
rect 11471 4508 12602 4536
rect 11471 4505 11483 4508
rect 11425 4499 11483 4505
rect 12590 4505 12602 4508
rect 12636 4505 12648 4539
rect 13354 4536 13360 4548
rect 12590 4499 12648 4505
rect 12728 4508 13360 4536
rect 9309 4471 9367 4477
rect 9309 4468 9321 4471
rect 8352 4440 9321 4468
rect 8352 4428 8358 4440
rect 9309 4437 9321 4440
rect 9355 4437 9367 4471
rect 9309 4431 9367 4437
rect 9769 4471 9827 4477
rect 9769 4437 9781 4471
rect 9815 4437 9827 4471
rect 9769 4431 9827 4437
rect 12434 4428 12440 4480
rect 12492 4468 12498 4480
rect 12728 4468 12756 4508
rect 13354 4496 13360 4508
rect 13412 4496 13418 4548
rect 12492 4440 12756 4468
rect 12492 4428 12498 4440
rect 12986 4428 12992 4480
rect 13044 4468 13050 4480
rect 13740 4477 13768 4576
rect 14093 4573 14105 4576
rect 14139 4573 14151 4607
rect 14093 4567 14151 4573
rect 16390 4564 16396 4616
rect 16448 4604 16454 4616
rect 16485 4607 16543 4613
rect 16485 4604 16497 4607
rect 16448 4576 16497 4604
rect 16448 4564 16454 4576
rect 16485 4573 16497 4576
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 16592 4536 16620 4712
rect 17126 4700 17132 4712
rect 17184 4700 17190 4752
rect 18248 4740 18276 4780
rect 18414 4768 18420 4820
rect 18472 4808 18478 4820
rect 18877 4811 18935 4817
rect 18877 4808 18889 4811
rect 18472 4780 18889 4808
rect 18472 4768 18478 4780
rect 18877 4777 18889 4780
rect 18923 4777 18935 4811
rect 20530 4808 20536 4820
rect 20491 4780 20536 4808
rect 18877 4771 18935 4777
rect 20530 4768 20536 4780
rect 20588 4768 20594 4820
rect 18966 4740 18972 4752
rect 18248 4712 18972 4740
rect 18966 4700 18972 4712
rect 19024 4700 19030 4752
rect 17218 4672 17224 4684
rect 17179 4644 17224 4672
rect 17218 4632 17224 4644
rect 17276 4632 17282 4684
rect 18230 4672 18236 4684
rect 17420 4644 17908 4672
rect 18191 4644 18236 4672
rect 17420 4604 17448 4644
rect 15304 4508 16620 4536
rect 16776 4576 17448 4604
rect 17880 4604 17908 4644
rect 18230 4632 18236 4644
rect 18288 4632 18294 4684
rect 19518 4632 19524 4684
rect 19576 4672 19582 4684
rect 19613 4675 19671 4681
rect 19613 4672 19625 4675
rect 19576 4644 19625 4672
rect 19576 4632 19582 4644
rect 19613 4641 19625 4644
rect 19659 4641 19671 4675
rect 19613 4635 19671 4641
rect 20070 4632 20076 4684
rect 20128 4672 20134 4684
rect 20993 4675 21051 4681
rect 20993 4672 21005 4675
rect 20128 4644 21005 4672
rect 20128 4632 20134 4644
rect 20993 4641 21005 4644
rect 21039 4641 21051 4675
rect 21174 4672 21180 4684
rect 21135 4644 21180 4672
rect 20993 4635 21051 4641
rect 21174 4632 21180 4644
rect 21232 4632 21238 4684
rect 19794 4604 19800 4616
rect 17880 4576 19800 4604
rect 13725 4471 13783 4477
rect 13725 4468 13737 4471
rect 13044 4440 13737 4468
rect 13044 4428 13050 4440
rect 13725 4437 13737 4440
rect 13771 4437 13783 4471
rect 13725 4431 13783 4437
rect 14274 4428 14280 4480
rect 14332 4468 14338 4480
rect 15304 4477 15332 4508
rect 15289 4471 15347 4477
rect 15289 4468 15301 4471
rect 14332 4440 15301 4468
rect 14332 4428 14338 4440
rect 15289 4437 15301 4440
rect 15335 4437 15347 4471
rect 15289 4431 15347 4437
rect 15378 4428 15384 4480
rect 15436 4468 15442 4480
rect 16393 4471 16451 4477
rect 15436 4440 15481 4468
rect 15436 4428 15442 4440
rect 16393 4437 16405 4471
rect 16439 4468 16451 4471
rect 16776 4468 16804 4576
rect 19794 4564 19800 4576
rect 19852 4564 19858 4616
rect 18417 4539 18475 4545
rect 18417 4536 18429 4539
rect 16868 4508 18429 4536
rect 16868 4477 16896 4508
rect 18417 4505 18429 4508
rect 18463 4505 18475 4539
rect 18417 4499 18475 4505
rect 18874 4496 18880 4548
rect 18932 4536 18938 4548
rect 19889 4539 19947 4545
rect 19889 4536 19901 4539
rect 18932 4508 19901 4536
rect 18932 4496 18938 4508
rect 19889 4505 19901 4508
rect 19935 4505 19947 4539
rect 19889 4499 19947 4505
rect 16439 4440 16804 4468
rect 16853 4471 16911 4477
rect 16439 4437 16451 4440
rect 16393 4431 16451 4437
rect 16853 4437 16865 4471
rect 16899 4437 16911 4471
rect 16853 4431 16911 4437
rect 17126 4428 17132 4480
rect 17184 4468 17190 4480
rect 17405 4471 17463 4477
rect 17405 4468 17417 4471
rect 17184 4440 17417 4468
rect 17184 4428 17190 4440
rect 17405 4437 17417 4440
rect 17451 4437 17463 4471
rect 17405 4431 17463 4437
rect 17494 4428 17500 4480
rect 17552 4468 17558 4480
rect 17865 4471 17923 4477
rect 17552 4440 17597 4468
rect 17552 4428 17558 4440
rect 17865 4437 17877 4471
rect 17911 4468 17923 4471
rect 18230 4468 18236 4480
rect 17911 4440 18236 4468
rect 17911 4437 17923 4440
rect 17865 4431 17923 4437
rect 18230 4428 18236 4440
rect 18288 4428 18294 4480
rect 18506 4428 18512 4480
rect 18564 4468 18570 4480
rect 18564 4440 18609 4468
rect 18564 4428 18570 4440
rect 19610 4428 19616 4480
rect 19668 4468 19674 4480
rect 19797 4471 19855 4477
rect 19797 4468 19809 4471
rect 19668 4440 19809 4468
rect 19668 4428 19674 4440
rect 19797 4437 19809 4440
rect 19843 4437 19855 4471
rect 19797 4431 19855 4437
rect 20257 4471 20315 4477
rect 20257 4437 20269 4471
rect 20303 4468 20315 4471
rect 20901 4471 20959 4477
rect 20901 4468 20913 4471
rect 20303 4440 20913 4468
rect 20303 4437 20315 4440
rect 20257 4431 20315 4437
rect 20901 4437 20913 4440
rect 20947 4437 20959 4471
rect 20901 4431 20959 4437
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 6733 4267 6791 4273
rect 6733 4233 6745 4267
rect 6779 4264 6791 4267
rect 14458 4264 14464 4276
rect 6779 4236 14464 4264
rect 6779 4233 6791 4236
rect 6733 4227 6791 4233
rect 14458 4224 14464 4236
rect 14516 4224 14522 4276
rect 17678 4264 17684 4276
rect 14568 4236 17684 4264
rect 5997 4199 6055 4205
rect 5997 4165 6009 4199
rect 6043 4196 6055 4199
rect 10781 4199 10839 4205
rect 10781 4196 10793 4199
rect 6043 4168 10793 4196
rect 6043 4165 6055 4168
rect 5997 4159 6055 4165
rect 10781 4165 10793 4168
rect 10827 4165 10839 4199
rect 10781 4159 10839 4165
rect 11885 4199 11943 4205
rect 11885 4165 11897 4199
rect 11931 4196 11943 4199
rect 12066 4196 12072 4208
rect 11931 4168 12072 4196
rect 11931 4165 11943 4168
rect 11885 4159 11943 4165
rect 12066 4156 12072 4168
rect 12124 4156 12130 4208
rect 13262 4196 13268 4208
rect 13223 4168 13268 4196
rect 13262 4156 13268 4168
rect 13320 4156 13326 4208
rect 13354 4156 13360 4208
rect 13412 4196 13418 4208
rect 14568 4196 14596 4236
rect 17678 4224 17684 4236
rect 17736 4224 17742 4276
rect 18138 4224 18144 4276
rect 18196 4264 18202 4276
rect 18325 4267 18383 4273
rect 18325 4264 18337 4267
rect 18196 4236 18337 4264
rect 18196 4224 18202 4236
rect 18325 4233 18337 4236
rect 18371 4233 18383 4267
rect 18325 4227 18383 4233
rect 18598 4224 18604 4276
rect 18656 4264 18662 4276
rect 20162 4264 20168 4276
rect 18656 4236 20168 4264
rect 18656 4224 18662 4236
rect 20162 4224 20168 4236
rect 20220 4264 20226 4276
rect 20438 4264 20444 4276
rect 20220 4236 20444 4264
rect 20220 4224 20226 4236
rect 20438 4224 20444 4236
rect 20496 4224 20502 4276
rect 15562 4196 15568 4208
rect 13412 4168 14596 4196
rect 15523 4168 15568 4196
rect 13412 4156 13418 4168
rect 15562 4156 15568 4168
rect 15620 4156 15626 4208
rect 16206 4156 16212 4208
rect 16264 4196 16270 4208
rect 16482 4196 16488 4208
rect 16264 4168 16488 4196
rect 16264 4156 16270 4168
rect 16482 4156 16488 4168
rect 16540 4156 16546 4208
rect 17402 4196 17408 4208
rect 16684 4168 17408 4196
rect 16684 4140 16712 4168
rect 17402 4156 17408 4168
rect 17460 4156 17466 4208
rect 18414 4196 18420 4208
rect 17512 4168 18420 4196
rect 4430 4128 4436 4140
rect 4391 4100 4436 4128
rect 4430 4088 4436 4100
rect 4488 4088 4494 4140
rect 4890 4128 4896 4140
rect 4851 4100 4896 4128
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 7009 4131 7067 4137
rect 7009 4097 7021 4131
rect 7055 4128 7067 4131
rect 7282 4128 7288 4140
rect 7055 4100 7288 4128
rect 7055 4097 7067 4100
rect 7009 4091 7067 4097
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 4062 4060 4068 4072
rect 2731 4032 4068 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 4062 4020 4068 4032
rect 4120 4020 4126 4072
rect 4157 4063 4215 4069
rect 4157 4029 4169 4063
rect 4203 4060 4215 4063
rect 5368 4060 5396 4091
rect 7282 4088 7288 4100
rect 7340 4088 7346 4140
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7558 4060 7564 4072
rect 4203 4032 7564 4060
rect 4203 4029 4215 4032
rect 4157 4023 4215 4029
rect 7558 4020 7564 4032
rect 7616 4020 7622 4072
rect 2317 3995 2375 4001
rect 2317 3961 2329 3995
rect 2363 3992 2375 3995
rect 2866 3992 2872 4004
rect 2363 3964 2872 3992
rect 2363 3961 2375 3964
rect 2317 3955 2375 3961
rect 2866 3952 2872 3964
rect 2924 3952 2930 4004
rect 3421 3995 3479 4001
rect 3421 3961 3433 3995
rect 3467 3992 3479 3995
rect 4890 3992 4896 4004
rect 3467 3964 4896 3992
rect 3467 3961 3479 3964
rect 3421 3955 3479 3961
rect 4890 3952 4896 3964
rect 4948 3952 4954 4004
rect 4982 3952 4988 4004
rect 5040 3992 5046 4004
rect 5534 3992 5540 4004
rect 5040 3964 5212 3992
rect 5495 3964 5540 3992
rect 5040 3952 5046 3964
rect 1302 3884 1308 3936
rect 1360 3924 1366 3936
rect 1397 3927 1455 3933
rect 1397 3924 1409 3927
rect 1360 3896 1409 3924
rect 1360 3884 1366 3896
rect 1397 3893 1409 3896
rect 1443 3893 1455 3927
rect 1946 3924 1952 3936
rect 1907 3896 1952 3924
rect 1397 3887 1455 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 3053 3927 3111 3933
rect 3053 3893 3065 3927
rect 3099 3924 3111 3927
rect 3234 3924 3240 3936
rect 3099 3896 3240 3924
rect 3099 3893 3111 3896
rect 3053 3887 3111 3893
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3789 3927 3847 3933
rect 3789 3893 3801 3927
rect 3835 3924 3847 3927
rect 3970 3924 3976 3936
rect 3835 3896 3976 3924
rect 3835 3893 3847 3896
rect 3789 3887 3847 3893
rect 3970 3884 3976 3896
rect 4028 3884 4034 3936
rect 4614 3924 4620 3936
rect 4575 3896 4620 3924
rect 4614 3884 4620 3896
rect 4672 3884 4678 3936
rect 5074 3924 5080 3936
rect 5035 3896 5080 3924
rect 5074 3884 5080 3896
rect 5132 3884 5138 3936
rect 5184 3924 5212 3964
rect 5534 3952 5540 3964
rect 5592 3952 5598 4004
rect 7282 3924 7288 3936
rect 5184 3896 7288 3924
rect 7282 3884 7288 3896
rect 7340 3884 7346 3936
rect 7668 3924 7696 4091
rect 7834 4088 7840 4140
rect 7892 4128 7898 4140
rect 8185 4131 8243 4137
rect 8185 4128 8197 4131
rect 7892 4100 8197 4128
rect 7892 4088 7898 4100
rect 8185 4097 8197 4100
rect 8231 4097 8243 4131
rect 9858 4128 9864 4140
rect 9819 4100 9864 4128
rect 8185 4091 8243 4097
rect 9858 4088 9864 4100
rect 9916 4088 9922 4140
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11793 4131 11851 4137
rect 11793 4128 11805 4131
rect 10928 4100 11805 4128
rect 10928 4088 10934 4100
rect 11793 4097 11805 4100
rect 11839 4128 11851 4131
rect 12526 4128 12532 4140
rect 11839 4100 12532 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 13446 4128 13452 4140
rect 13096 4100 13452 4128
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 7929 4063 7987 4069
rect 7929 4060 7941 4063
rect 7800 4032 7941 4060
rect 7800 4020 7806 4032
rect 7929 4029 7941 4032
rect 7975 4029 7987 4063
rect 7929 4023 7987 4029
rect 10597 4063 10655 4069
rect 10597 4029 10609 4063
rect 10643 4029 10655 4063
rect 10597 4023 10655 4029
rect 10689 4063 10747 4069
rect 10689 4029 10701 4063
rect 10735 4060 10747 4063
rect 11054 4060 11060 4072
rect 10735 4032 11060 4060
rect 10735 4029 10747 4032
rect 10689 4023 10747 4029
rect 10612 3992 10640 4023
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11701 4063 11759 4069
rect 11701 4029 11713 4063
rect 11747 4029 11759 4063
rect 12986 4060 12992 4072
rect 11701 4023 11759 4029
rect 12406 4032 12992 4060
rect 11422 3992 11428 4004
rect 10612 3964 11428 3992
rect 11422 3952 11428 3964
rect 11480 3952 11486 4004
rect 11716 3992 11744 4023
rect 12406 3992 12434 4032
rect 12986 4020 12992 4032
rect 13044 4020 13050 4072
rect 13096 4069 13124 4100
rect 13446 4088 13452 4100
rect 13504 4128 13510 4140
rect 13909 4131 13967 4137
rect 13909 4128 13921 4131
rect 13504 4100 13921 4128
rect 13504 4088 13510 4100
rect 13909 4097 13921 4100
rect 13955 4097 13967 4131
rect 13909 4091 13967 4097
rect 14921 4131 14979 4137
rect 14921 4097 14933 4131
rect 14967 4128 14979 4131
rect 15102 4128 15108 4140
rect 14967 4100 15108 4128
rect 14967 4097 14979 4100
rect 14921 4091 14979 4097
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 15746 4128 15752 4140
rect 15212 4100 15752 4128
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 13081 4023 13139 4029
rect 13173 4063 13231 4069
rect 13173 4029 13185 4063
rect 13219 4060 13231 4063
rect 13722 4060 13728 4072
rect 13219 4032 13728 4060
rect 13219 4029 13231 4032
rect 13173 4023 13231 4029
rect 13722 4020 13728 4032
rect 13780 4020 13786 4072
rect 14826 4020 14832 4072
rect 14884 4060 14890 4072
rect 15212 4060 15240 4100
rect 15746 4088 15752 4100
rect 15804 4128 15810 4140
rect 16301 4131 16359 4137
rect 16301 4128 16313 4131
rect 15804 4100 16313 4128
rect 15804 4088 15810 4100
rect 16301 4097 16313 4100
rect 16347 4097 16359 4131
rect 16666 4128 16672 4140
rect 16579 4100 16672 4128
rect 16301 4091 16359 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16758 4088 16764 4140
rect 16816 4128 16822 4140
rect 16925 4131 16983 4137
rect 16925 4128 16937 4131
rect 16816 4100 16937 4128
rect 16816 4088 16822 4100
rect 16925 4097 16937 4100
rect 16971 4097 16983 4131
rect 16925 4091 16983 4097
rect 17218 4088 17224 4140
rect 17276 4128 17282 4140
rect 17512 4128 17540 4168
rect 18414 4156 18420 4168
rect 18472 4196 18478 4208
rect 21094 4199 21152 4205
rect 21094 4196 21106 4199
rect 18472 4168 21106 4196
rect 18472 4156 18478 4168
rect 21094 4165 21106 4168
rect 21140 4196 21152 4199
rect 21266 4196 21272 4208
rect 21140 4168 21272 4196
rect 21140 4165 21152 4168
rect 21094 4159 21152 4165
rect 21266 4156 21272 4168
rect 21324 4156 21330 4208
rect 17276 4100 17540 4128
rect 17276 4088 17282 4100
rect 18966 4088 18972 4140
rect 19024 4128 19030 4140
rect 19438 4131 19496 4137
rect 19438 4128 19450 4131
rect 19024 4100 19450 4128
rect 19024 4088 19030 4100
rect 19438 4097 19450 4100
rect 19484 4128 19496 4131
rect 19705 4131 19763 4137
rect 19484 4100 19656 4128
rect 19484 4097 19496 4100
rect 19438 4091 19496 4097
rect 14884 4032 15240 4060
rect 15381 4063 15439 4069
rect 14884 4020 14890 4032
rect 15381 4029 15393 4063
rect 15427 4029 15439 4063
rect 15381 4023 15439 4029
rect 15473 4063 15531 4069
rect 15473 4029 15485 4063
rect 15519 4060 15531 4063
rect 16206 4060 16212 4072
rect 15519 4032 16212 4060
rect 15519 4029 15531 4032
rect 15473 4023 15531 4029
rect 11716 3964 12434 3992
rect 13538 3952 13544 4004
rect 13596 3992 13602 4004
rect 13633 3995 13691 4001
rect 13633 3992 13645 3995
rect 13596 3964 13645 3992
rect 13596 3952 13602 3964
rect 13633 3961 13645 3964
rect 13679 3961 13691 3995
rect 13633 3955 13691 3961
rect 14734 3952 14740 4004
rect 14792 3992 14798 4004
rect 15396 3992 15424 4023
rect 16206 4020 16212 4032
rect 16264 4020 16270 4072
rect 19628 4060 19656 4100
rect 19705 4097 19717 4131
rect 19751 4128 19763 4131
rect 20530 4128 20536 4140
rect 19751 4100 20536 4128
rect 19751 4097 19763 4100
rect 19705 4091 19763 4097
rect 20530 4088 20536 4100
rect 20588 4128 20594 4140
rect 21361 4131 21419 4137
rect 21361 4128 21373 4131
rect 20588 4100 21373 4128
rect 20588 4088 20594 4100
rect 21361 4097 21373 4100
rect 21407 4097 21419 4131
rect 21361 4091 21419 4097
rect 19628 4032 20024 4060
rect 19996 4001 20024 4032
rect 19981 3995 20039 4001
rect 14792 3964 16344 3992
rect 14792 3952 14798 3964
rect 9309 3927 9367 3933
rect 9309 3924 9321 3927
rect 7668 3896 9321 3924
rect 9309 3893 9321 3896
rect 9355 3924 9367 3927
rect 9490 3924 9496 3936
rect 9355 3896 9496 3924
rect 9355 3893 9367 3896
rect 9309 3887 9367 3893
rect 9490 3884 9496 3896
rect 9548 3884 9554 3936
rect 10045 3927 10103 3933
rect 10045 3893 10057 3927
rect 10091 3924 10103 3927
rect 10962 3924 10968 3936
rect 10091 3896 10968 3924
rect 10091 3893 10103 3896
rect 10045 3887 10103 3893
rect 10962 3884 10968 3896
rect 11020 3884 11026 3936
rect 11149 3927 11207 3933
rect 11149 3893 11161 3927
rect 11195 3924 11207 3927
rect 11882 3924 11888 3936
rect 11195 3896 11888 3924
rect 11195 3893 11207 3896
rect 11149 3887 11207 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12253 3927 12311 3933
rect 12253 3924 12265 3927
rect 12032 3896 12265 3924
rect 12032 3884 12038 3896
rect 12253 3893 12265 3896
rect 12299 3893 12311 3927
rect 12253 3887 12311 3893
rect 12621 3927 12679 3933
rect 12621 3893 12633 3927
rect 12667 3924 12679 3927
rect 12894 3924 12900 3936
rect 12667 3896 12900 3924
rect 12667 3893 12679 3896
rect 12621 3887 12679 3893
rect 12894 3884 12900 3896
rect 12952 3884 12958 3936
rect 13170 3884 13176 3936
rect 13228 3924 13234 3936
rect 14553 3927 14611 3933
rect 14553 3924 14565 3927
rect 13228 3896 14565 3924
rect 13228 3884 13234 3896
rect 14553 3893 14565 3896
rect 14599 3893 14611 3927
rect 14553 3887 14611 3893
rect 15470 3884 15476 3936
rect 15528 3924 15534 3936
rect 15933 3927 15991 3933
rect 15933 3924 15945 3927
rect 15528 3896 15945 3924
rect 15528 3884 15534 3896
rect 15933 3893 15945 3896
rect 15979 3893 15991 3927
rect 16316 3924 16344 3964
rect 19981 3961 19993 3995
rect 20027 3961 20039 3995
rect 19981 3955 20039 3961
rect 17402 3924 17408 3936
rect 16316 3896 17408 3924
rect 15933 3887 15991 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 17862 3884 17868 3936
rect 17920 3924 17926 3936
rect 18049 3927 18107 3933
rect 18049 3924 18061 3927
rect 17920 3896 18061 3924
rect 17920 3884 17926 3896
rect 18049 3893 18061 3896
rect 18095 3893 18107 3927
rect 18049 3887 18107 3893
rect 18782 3884 18788 3936
rect 18840 3924 18846 3936
rect 19518 3924 19524 3936
rect 18840 3896 19524 3924
rect 18840 3884 18846 3896
rect 19518 3884 19524 3896
rect 19576 3884 19582 3936
rect 19886 3884 19892 3936
rect 19944 3924 19950 3936
rect 21450 3924 21456 3936
rect 19944 3896 21456 3924
rect 19944 3884 19950 3896
rect 21450 3884 21456 3896
rect 21508 3884 21514 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 1578 3720 1584 3732
rect 1539 3692 1584 3720
rect 1578 3680 1584 3692
rect 1636 3680 1642 3732
rect 3421 3723 3479 3729
rect 3421 3689 3433 3723
rect 3467 3720 3479 3723
rect 5534 3720 5540 3732
rect 3467 3692 5540 3720
rect 3467 3689 3479 3692
rect 3421 3683 3479 3689
rect 5534 3680 5540 3692
rect 5592 3680 5598 3732
rect 5718 3720 5724 3732
rect 5679 3692 5724 3720
rect 5718 3680 5724 3692
rect 5776 3680 5782 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 8941 3723 8999 3729
rect 6880 3692 8708 3720
rect 6880 3680 6886 3692
rect 3970 3612 3976 3664
rect 4028 3652 4034 3664
rect 5074 3652 5080 3664
rect 4028 3624 5080 3652
rect 4028 3612 4034 3624
rect 5074 3612 5080 3624
rect 5132 3612 5138 3664
rect 6917 3655 6975 3661
rect 6917 3621 6929 3655
rect 6963 3652 6975 3655
rect 8386 3652 8392 3664
rect 6963 3624 8392 3652
rect 6963 3621 6975 3624
rect 6917 3615 6975 3621
rect 8386 3612 8392 3624
rect 8444 3612 8450 3664
rect 8680 3652 8708 3692
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 9122 3720 9128 3732
rect 8987 3692 9128 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 9582 3680 9588 3732
rect 9640 3720 9646 3732
rect 11422 3720 11428 3732
rect 9640 3692 11284 3720
rect 11383 3692 11428 3720
rect 9640 3680 9646 3692
rect 10042 3652 10048 3664
rect 8680 3624 10048 3652
rect 10042 3612 10048 3624
rect 10100 3612 10106 3664
rect 11256 3652 11284 3692
rect 11422 3680 11428 3692
rect 11480 3680 11486 3732
rect 14458 3720 14464 3732
rect 11900 3692 14464 3720
rect 11900 3652 11928 3692
rect 14458 3680 14464 3692
rect 14516 3680 14522 3732
rect 14553 3723 14611 3729
rect 14553 3689 14565 3723
rect 14599 3720 14611 3723
rect 14734 3720 14740 3732
rect 14599 3692 14740 3720
rect 14599 3689 14611 3692
rect 14553 3683 14611 3689
rect 14734 3680 14740 3692
rect 14792 3680 14798 3732
rect 16206 3720 16212 3732
rect 16167 3692 16212 3720
rect 16206 3680 16212 3692
rect 16264 3680 16270 3732
rect 16298 3680 16304 3732
rect 16356 3720 16362 3732
rect 16942 3720 16948 3732
rect 16356 3692 16948 3720
rect 16356 3680 16362 3692
rect 16942 3680 16948 3692
rect 17000 3680 17006 3732
rect 17126 3680 17132 3732
rect 17184 3720 17190 3732
rect 20622 3720 20628 3732
rect 17184 3692 20628 3720
rect 17184 3680 17190 3692
rect 20622 3680 20628 3692
rect 20680 3680 20686 3732
rect 11256 3624 11928 3652
rect 11977 3655 12035 3661
rect 11977 3621 11989 3655
rect 12023 3652 12035 3655
rect 12710 3652 12716 3664
rect 12023 3624 12716 3652
rect 12023 3621 12035 3624
rect 11977 3615 12035 3621
rect 12710 3612 12716 3624
rect 12768 3612 12774 3664
rect 14277 3655 14335 3661
rect 14277 3621 14289 3655
rect 14323 3652 14335 3655
rect 14366 3652 14372 3664
rect 14323 3624 14372 3652
rect 14323 3621 14335 3624
rect 14277 3615 14335 3621
rect 14366 3612 14372 3624
rect 14424 3612 14430 3664
rect 16022 3612 16028 3664
rect 16080 3652 16086 3664
rect 16080 3624 16804 3652
rect 16080 3612 16086 3624
rect 3881 3587 3939 3593
rect 3881 3553 3893 3587
rect 3927 3584 3939 3587
rect 5350 3584 5356 3596
rect 3927 3556 5356 3584
rect 3927 3553 3939 3556
rect 3881 3547 3939 3553
rect 5350 3544 5356 3556
rect 5408 3544 5414 3596
rect 7926 3584 7932 3596
rect 7887 3556 7932 3584
rect 7926 3544 7932 3556
rect 7984 3544 7990 3596
rect 9490 3584 9496 3596
rect 8312 3556 9352 3584
rect 9451 3556 9496 3584
rect 658 3476 664 3528
rect 716 3516 722 3528
rect 1302 3516 1308 3528
rect 716 3488 1308 3516
rect 716 3476 722 3488
rect 1302 3476 1308 3488
rect 1360 3516 1366 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 1360 3488 1409 3516
rect 1360 3476 1366 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 3053 3519 3111 3525
rect 3053 3485 3065 3519
rect 3099 3516 3111 3519
rect 3326 3516 3332 3528
rect 3099 3488 3332 3516
rect 3099 3485 3111 3488
rect 3053 3479 3111 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3485 4215 3519
rect 4157 3479 4215 3485
rect 2685 3451 2743 3457
rect 2685 3417 2697 3451
rect 2731 3448 2743 3451
rect 4172 3448 4200 3479
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4430 3516 4436 3528
rect 4304 3488 4436 3516
rect 4304 3476 4310 3488
rect 4430 3476 4436 3488
rect 4488 3476 4494 3528
rect 4617 3519 4675 3525
rect 4617 3485 4629 3519
rect 4663 3516 4675 3519
rect 4982 3516 4988 3528
rect 4663 3488 4988 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 4982 3476 4988 3488
rect 5040 3476 5046 3528
rect 5074 3476 5080 3528
rect 5132 3516 5138 3528
rect 5132 3488 5177 3516
rect 5132 3476 5138 3488
rect 5534 3476 5540 3528
rect 5592 3516 5598 3528
rect 5718 3516 5724 3528
rect 5592 3488 5724 3516
rect 5592 3476 5598 3488
rect 5718 3476 5724 3488
rect 5776 3476 5782 3528
rect 6457 3519 6515 3525
rect 6457 3485 6469 3519
rect 6503 3512 6515 3519
rect 6914 3516 6920 3528
rect 6564 3512 6920 3516
rect 6503 3488 6920 3512
rect 6503 3485 6592 3488
rect 6457 3484 6592 3485
rect 6457 3479 6515 3484
rect 6914 3476 6920 3488
rect 6972 3476 6978 3528
rect 7561 3519 7619 3525
rect 7561 3485 7573 3519
rect 7607 3516 7619 3519
rect 7650 3516 7656 3528
rect 7607 3488 7656 3516
rect 7607 3485 7619 3488
rect 7561 3479 7619 3485
rect 7650 3476 7656 3488
rect 7708 3476 7714 3528
rect 8110 3516 8116 3528
rect 8071 3488 8116 3516
rect 8110 3476 8116 3488
rect 8168 3476 8174 3528
rect 4706 3448 4712 3460
rect 2731 3420 4712 3448
rect 2731 3417 2743 3420
rect 2685 3411 2743 3417
rect 4706 3408 4712 3420
rect 4764 3408 4770 3460
rect 8205 3451 8263 3457
rect 8205 3448 8217 3451
rect 4816 3420 8217 3448
rect 1949 3383 2007 3389
rect 1949 3349 1961 3383
rect 1995 3380 2007 3383
rect 2130 3380 2136 3392
rect 1995 3352 2136 3380
rect 1995 3349 2007 3352
rect 1949 3343 2007 3349
rect 2130 3340 2136 3352
rect 2188 3340 2194 3392
rect 2317 3383 2375 3389
rect 2317 3349 2329 3383
rect 2363 3380 2375 3383
rect 2590 3380 2596 3392
rect 2363 3352 2596 3380
rect 2363 3349 2375 3352
rect 2317 3343 2375 3349
rect 2590 3340 2596 3352
rect 2648 3340 2654 3392
rect 4341 3383 4399 3389
rect 4341 3349 4353 3383
rect 4387 3380 4399 3383
rect 4614 3380 4620 3392
rect 4387 3352 4620 3380
rect 4387 3349 4399 3352
rect 4341 3343 4399 3349
rect 4614 3340 4620 3352
rect 4672 3340 4678 3392
rect 4816 3389 4844 3420
rect 8205 3417 8217 3420
rect 8251 3417 8263 3451
rect 8205 3411 8263 3417
rect 4801 3383 4859 3389
rect 4801 3349 4813 3383
rect 4847 3349 4859 3383
rect 5258 3380 5264 3392
rect 5219 3352 5264 3380
rect 4801 3343 4859 3349
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6181 3383 6239 3389
rect 6181 3380 6193 3383
rect 6052 3352 6193 3380
rect 6052 3340 6058 3352
rect 6181 3349 6193 3352
rect 6227 3349 6239 3383
rect 6638 3380 6644 3392
rect 6599 3352 6644 3380
rect 6181 3343 6239 3349
rect 6638 3340 6644 3352
rect 6696 3340 6702 3392
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 8312 3380 8340 3556
rect 9324 3525 9352 3556
rect 9490 3544 9496 3556
rect 9548 3544 9554 3596
rect 15933 3587 15991 3593
rect 15933 3553 15945 3587
rect 15979 3584 15991 3587
rect 16666 3584 16672 3596
rect 15979 3556 16672 3584
rect 15979 3553 15991 3556
rect 15933 3547 15991 3553
rect 16666 3544 16672 3556
rect 16724 3544 16730 3596
rect 16776 3593 16804 3624
rect 16761 3587 16819 3593
rect 16761 3553 16773 3587
rect 16807 3553 16819 3587
rect 16761 3547 16819 3553
rect 17218 3544 17224 3596
rect 17276 3584 17282 3596
rect 17681 3587 17739 3593
rect 17681 3584 17693 3587
rect 17276 3556 17693 3584
rect 17276 3544 17282 3556
rect 17681 3553 17693 3556
rect 17727 3553 17739 3587
rect 17862 3584 17868 3596
rect 17823 3556 17868 3584
rect 17681 3547 17739 3553
rect 17862 3544 17868 3556
rect 17920 3544 17926 3596
rect 20438 3544 20444 3596
rect 20496 3584 20502 3596
rect 20809 3587 20867 3593
rect 20809 3584 20821 3587
rect 20496 3556 20821 3584
rect 20496 3544 20502 3556
rect 20809 3553 20821 3556
rect 20855 3553 20867 3587
rect 20809 3547 20867 3553
rect 9309 3519 9367 3525
rect 9309 3485 9321 3519
rect 9355 3485 9367 3519
rect 9309 3479 9367 3485
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 11146 3516 11152 3528
rect 10091 3488 11152 3516
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 11146 3476 11152 3488
rect 11204 3476 11210 3528
rect 11790 3516 11796 3528
rect 11751 3488 11796 3516
rect 11790 3476 11796 3488
rect 11848 3476 11854 3528
rect 13630 3476 13636 3528
rect 13688 3516 13694 3528
rect 13725 3519 13783 3525
rect 13725 3516 13737 3519
rect 13688 3488 13737 3516
rect 13688 3476 13694 3488
rect 13725 3485 13737 3488
rect 13771 3485 13783 3519
rect 13725 3479 13783 3485
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3516 14151 3519
rect 15194 3516 15200 3528
rect 14139 3488 15200 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 15194 3476 15200 3488
rect 15252 3476 15258 3528
rect 15580 3488 17356 3516
rect 8386 3408 8392 3460
rect 8444 3448 8450 3460
rect 10290 3451 10348 3457
rect 10290 3448 10302 3451
rect 8444 3420 10302 3448
rect 8444 3408 8450 3420
rect 10290 3417 10302 3420
rect 10336 3417 10348 3451
rect 10290 3411 10348 3417
rect 10962 3408 10968 3460
rect 11020 3448 11026 3460
rect 13480 3451 13538 3457
rect 11020 3420 13400 3448
rect 11020 3408 11026 3420
rect 6788 3352 8340 3380
rect 6788 3340 6794 3352
rect 8570 3340 8576 3392
rect 8628 3380 8634 3392
rect 9401 3383 9459 3389
rect 8628 3352 8673 3380
rect 8628 3340 8634 3352
rect 9401 3349 9413 3383
rect 9447 3380 9459 3383
rect 9582 3380 9588 3392
rect 9447 3352 9588 3380
rect 9447 3349 9459 3352
rect 9401 3343 9459 3349
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 12345 3383 12403 3389
rect 12345 3349 12357 3383
rect 12391 3380 12403 3383
rect 12434 3380 12440 3392
rect 12391 3352 12440 3380
rect 12391 3349 12403 3352
rect 12345 3343 12403 3349
rect 12434 3340 12440 3352
rect 12492 3340 12498 3392
rect 13372 3380 13400 3420
rect 13480 3417 13492 3451
rect 13526 3448 13538 3451
rect 15580 3448 15608 3488
rect 13526 3420 15608 3448
rect 13526 3417 13538 3420
rect 13480 3411 13538 3417
rect 15654 3408 15660 3460
rect 15712 3457 15718 3460
rect 15712 3451 15746 3457
rect 15734 3448 15746 3451
rect 16022 3448 16028 3460
rect 15734 3420 16028 3448
rect 15734 3417 15746 3420
rect 15712 3411 15746 3417
rect 15712 3408 15718 3411
rect 16022 3408 16028 3420
rect 16080 3408 16086 3460
rect 16114 3408 16120 3460
rect 16172 3448 16178 3460
rect 16577 3451 16635 3457
rect 16172 3420 16436 3448
rect 16172 3408 16178 3420
rect 13906 3380 13912 3392
rect 13372 3352 13912 3380
rect 13906 3340 13912 3352
rect 13964 3340 13970 3392
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 16298 3380 16304 3392
rect 15528 3352 16304 3380
rect 15528 3340 15534 3352
rect 16298 3340 16304 3352
rect 16356 3340 16362 3392
rect 16408 3380 16436 3420
rect 16577 3417 16589 3451
rect 16623 3448 16635 3451
rect 17328 3448 17356 3488
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 18233 3519 18291 3525
rect 18233 3516 18245 3519
rect 17460 3488 18245 3516
rect 17460 3476 17466 3488
rect 18233 3485 18245 3488
rect 18279 3485 18291 3519
rect 18233 3479 18291 3485
rect 19429 3519 19487 3525
rect 19429 3485 19441 3519
rect 19475 3516 19487 3519
rect 19518 3516 19524 3528
rect 19475 3488 19524 3516
rect 19475 3485 19487 3488
rect 19429 3479 19487 3485
rect 19518 3476 19524 3488
rect 19576 3476 19582 3528
rect 19702 3516 19708 3528
rect 19663 3488 19708 3516
rect 19702 3476 19708 3488
rect 19760 3476 19766 3528
rect 20346 3476 20352 3528
rect 20404 3516 20410 3528
rect 20533 3519 20591 3525
rect 20533 3516 20545 3519
rect 20404 3488 20545 3516
rect 20404 3476 20410 3488
rect 20533 3485 20545 3488
rect 20579 3516 20591 3519
rect 20622 3516 20628 3528
rect 20579 3488 20628 3516
rect 20579 3485 20591 3488
rect 20533 3479 20591 3485
rect 20622 3476 20628 3488
rect 20680 3476 20686 3528
rect 18877 3451 18935 3457
rect 18877 3448 18889 3451
rect 16623 3420 17264 3448
rect 17328 3420 18889 3448
rect 16623 3417 16635 3420
rect 16577 3411 16635 3417
rect 17236 3389 17264 3420
rect 18877 3417 18889 3420
rect 18923 3417 18935 3451
rect 18877 3411 18935 3417
rect 16669 3383 16727 3389
rect 16669 3380 16681 3383
rect 16408 3352 16681 3380
rect 16669 3349 16681 3352
rect 16715 3349 16727 3383
rect 16669 3343 16727 3349
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3349 17279 3383
rect 17221 3343 17279 3349
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 17589 3383 17647 3389
rect 17589 3380 17601 3383
rect 17552 3352 17601 3380
rect 17552 3340 17558 3352
rect 17589 3349 17601 3352
rect 17635 3349 17647 3383
rect 17589 3343 17647 3349
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 20530 3380 20536 3392
rect 18104 3352 20536 3380
rect 18104 3340 18110 3352
rect 20530 3340 20536 3352
rect 20588 3340 20594 3392
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 1581 3179 1639 3185
rect 1581 3145 1593 3179
rect 1627 3176 1639 3179
rect 1854 3176 1860 3188
rect 1627 3148 1860 3176
rect 1627 3145 1639 3148
rect 1581 3139 1639 3145
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 2038 3176 2044 3188
rect 1999 3148 2044 3176
rect 2038 3136 2044 3148
rect 2096 3136 2102 3188
rect 2498 3176 2504 3188
rect 2459 3148 2504 3176
rect 2498 3136 2504 3148
rect 2556 3136 2562 3188
rect 2958 3176 2964 3188
rect 2919 3148 2964 3176
rect 2958 3136 2964 3148
rect 3016 3136 3022 3188
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 3292 3148 4384 3176
rect 3292 3136 3298 3148
rect 4356 3108 4384 3148
rect 4430 3136 4436 3188
rect 4488 3176 4494 3188
rect 4617 3179 4675 3185
rect 4488 3148 4568 3176
rect 4488 3136 4494 3148
rect 4540 3108 4568 3148
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 6730 3176 6736 3188
rect 4663 3148 6736 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 6825 3179 6883 3185
rect 6825 3145 6837 3179
rect 6871 3176 6883 3179
rect 7834 3176 7840 3188
rect 6871 3148 7840 3176
rect 6871 3145 6883 3148
rect 6825 3139 6883 3145
rect 7834 3136 7840 3148
rect 7892 3136 7898 3188
rect 8018 3136 8024 3188
rect 8076 3176 8082 3188
rect 9769 3179 9827 3185
rect 9769 3176 9781 3179
rect 8076 3148 9781 3176
rect 8076 3136 8082 3148
rect 9769 3145 9781 3148
rect 9815 3176 9827 3179
rect 10502 3176 10508 3188
rect 9815 3148 10508 3176
rect 9815 3145 9827 3148
rect 9769 3139 9827 3145
rect 10502 3136 10508 3148
rect 10560 3136 10566 3188
rect 13170 3176 13176 3188
rect 11164 3148 13176 3176
rect 5626 3108 5632 3120
rect 4356 3080 4476 3108
rect 4540 3080 5632 3108
rect 1210 3000 1216 3052
rect 1268 3040 1274 3052
rect 1397 3043 1455 3049
rect 1397 3040 1409 3043
rect 1268 3012 1409 3040
rect 1268 3000 1274 3012
rect 1397 3009 1409 3012
rect 1443 3040 1455 3043
rect 1670 3040 1676 3052
rect 1443 3012 1676 3040
rect 1443 3009 1455 3012
rect 1397 3003 1455 3009
rect 1670 3000 1676 3012
rect 1728 3000 1734 3052
rect 1762 3000 1768 3052
rect 1820 3040 1826 3052
rect 1857 3043 1915 3049
rect 1857 3040 1869 3043
rect 1820 3012 1869 3040
rect 1820 3000 1826 3012
rect 1857 3009 1869 3012
rect 1903 3009 1915 3043
rect 2314 3040 2320 3052
rect 2275 3012 2320 3040
rect 1857 3003 1915 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2777 3043 2835 3049
rect 2777 3009 2789 3043
rect 2823 3040 2835 3043
rect 2866 3040 2872 3052
rect 2823 3012 2872 3040
rect 2823 3009 2835 3012
rect 2777 3003 2835 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 3418 3000 3424 3052
rect 3476 3040 3482 3052
rect 3513 3043 3571 3049
rect 3513 3040 3525 3043
rect 3476 3012 3525 3040
rect 3476 3000 3482 3012
rect 3513 3009 3525 3012
rect 3559 3009 3571 3043
rect 3513 3003 3571 3009
rect 3973 3043 4031 3049
rect 3973 3009 3985 3043
rect 4019 3040 4031 3043
rect 4246 3040 4252 3052
rect 4019 3012 4252 3040
rect 4019 3009 4031 3012
rect 3973 3003 4031 3009
rect 3528 2972 3556 3003
rect 4246 3000 4252 3012
rect 4304 3000 4310 3052
rect 4448 3049 4476 3080
rect 5626 3068 5632 3080
rect 5684 3068 5690 3120
rect 5997 3111 6055 3117
rect 5997 3077 6009 3111
rect 6043 3108 6055 3111
rect 7650 3108 7656 3120
rect 6043 3080 7656 3108
rect 6043 3077 6055 3080
rect 5997 3071 6055 3077
rect 7650 3068 7656 3080
rect 7708 3068 7714 3120
rect 8202 3068 8208 3120
rect 8260 3108 8266 3120
rect 10904 3111 10962 3117
rect 8260 3080 9628 3108
rect 8260 3068 8266 3080
rect 4433 3043 4491 3049
rect 4433 3009 4445 3043
rect 4479 3040 4491 3043
rect 4890 3040 4896 3052
rect 4479 3012 4752 3040
rect 4851 3012 4896 3040
rect 4479 3009 4491 3012
rect 4433 3003 4491 3009
rect 4522 2972 4528 2984
rect 3528 2944 4528 2972
rect 4522 2932 4528 2944
rect 4580 2932 4586 2984
rect 3694 2904 3700 2916
rect 3655 2876 3700 2904
rect 3694 2864 3700 2876
rect 3752 2864 3758 2916
rect 4154 2904 4160 2916
rect 4115 2876 4160 2904
rect 4154 2864 4160 2876
rect 4212 2864 4218 2916
rect 4430 2864 4436 2916
rect 4488 2864 4494 2916
rect 4724 2904 4752 3012
rect 4890 3000 4896 3012
rect 4948 3000 4954 3052
rect 5166 3000 5172 3052
rect 5224 3040 5230 3052
rect 5353 3043 5411 3049
rect 5353 3040 5365 3043
rect 5224 3012 5365 3040
rect 5224 3000 5230 3012
rect 5353 3009 5365 3012
rect 5399 3009 5411 3043
rect 5353 3003 5411 3009
rect 6365 3043 6423 3049
rect 6365 3009 6377 3043
rect 6411 3040 6423 3043
rect 6822 3040 6828 3052
rect 6411 3012 6828 3040
rect 6411 3009 6423 3012
rect 6365 3003 6423 3009
rect 6822 3000 6828 3012
rect 6880 3000 6886 3052
rect 7469 3043 7527 3049
rect 7469 3009 7481 3043
rect 7515 3009 7527 3043
rect 7469 3003 7527 3009
rect 4908 2972 4936 3000
rect 6638 2972 6644 2984
rect 4908 2944 6644 2972
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 6546 2904 6552 2916
rect 4724 2876 6408 2904
rect 6507 2876 6552 2904
rect 4448 2836 4476 2864
rect 4890 2836 4896 2848
rect 4448 2808 4896 2836
rect 4890 2796 4896 2808
rect 4948 2796 4954 2848
rect 5077 2839 5135 2845
rect 5077 2805 5089 2839
rect 5123 2836 5135 2839
rect 5442 2836 5448 2848
rect 5123 2808 5448 2836
rect 5123 2805 5135 2808
rect 5077 2799 5135 2805
rect 5442 2796 5448 2808
rect 5500 2796 5506 2848
rect 5537 2839 5595 2845
rect 5537 2805 5549 2839
rect 5583 2836 5595 2839
rect 5902 2836 5908 2848
rect 5583 2808 5908 2836
rect 5583 2805 5595 2808
rect 5537 2799 5595 2805
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6380 2836 6408 2876
rect 6546 2864 6552 2876
rect 6604 2864 6610 2916
rect 6454 2836 6460 2848
rect 6380 2808 6460 2836
rect 6454 2796 6460 2808
rect 6512 2796 6518 2848
rect 7484 2836 7512 3003
rect 7558 3000 7564 3052
rect 7616 3040 7622 3052
rect 8001 3043 8059 3049
rect 8001 3040 8013 3043
rect 7616 3012 8013 3040
rect 7616 3000 7622 3012
rect 8001 3009 8013 3012
rect 8047 3009 8059 3043
rect 9490 3040 9496 3052
rect 9451 3012 9496 3040
rect 8001 3003 8059 3009
rect 9490 3000 9496 3012
rect 9548 3000 9554 3052
rect 9600 3040 9628 3080
rect 10904 3077 10916 3111
rect 10950 3108 10962 3111
rect 11164 3108 11192 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 13446 3176 13452 3188
rect 13407 3148 13452 3176
rect 13446 3136 13452 3148
rect 13504 3136 13510 3188
rect 13722 3176 13728 3188
rect 13683 3148 13728 3176
rect 13722 3136 13728 3148
rect 13780 3136 13786 3188
rect 14185 3179 14243 3185
rect 14185 3145 14197 3179
rect 14231 3176 14243 3179
rect 14734 3176 14740 3188
rect 14231 3148 14740 3176
rect 14231 3145 14243 3148
rect 14185 3139 14243 3145
rect 14734 3136 14740 3148
rect 14792 3136 14798 3188
rect 14829 3179 14887 3185
rect 14829 3145 14841 3179
rect 14875 3176 14887 3179
rect 15194 3176 15200 3188
rect 14875 3148 15200 3176
rect 14875 3145 14887 3148
rect 14829 3139 14887 3145
rect 15194 3136 15200 3148
rect 15252 3176 15258 3188
rect 15654 3176 15660 3188
rect 15252 3148 15660 3176
rect 15252 3136 15258 3148
rect 15654 3136 15660 3148
rect 15712 3136 15718 3188
rect 16114 3136 16120 3188
rect 16172 3176 16178 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 16172 3148 16681 3176
rect 16172 3136 16178 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 17037 3179 17095 3185
rect 17037 3176 17049 3179
rect 16669 3139 16727 3145
rect 16776 3148 17049 3176
rect 10950 3080 11192 3108
rect 12336 3111 12394 3117
rect 10950 3077 10962 3080
rect 10904 3071 10962 3077
rect 12336 3077 12348 3111
rect 12382 3108 12394 3111
rect 12434 3108 12440 3120
rect 12382 3080 12440 3108
rect 12382 3077 12394 3080
rect 12336 3071 12394 3077
rect 12434 3068 12440 3080
rect 12492 3108 12498 3120
rect 13354 3108 13360 3120
rect 12492 3080 13360 3108
rect 12492 3068 12498 3080
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 14274 3108 14280 3120
rect 14108 3080 14280 3108
rect 11146 3040 11152 3052
rect 9600 3012 9674 3040
rect 11107 3012 11152 3040
rect 7742 2972 7748 2984
rect 7703 2944 7748 2972
rect 7742 2932 7748 2944
rect 7800 2932 7806 2984
rect 9490 2904 9496 2916
rect 9140 2876 9496 2904
rect 9140 2845 9168 2876
rect 9490 2864 9496 2876
rect 9548 2864 9554 2916
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 7484 2808 9137 2836
rect 9125 2805 9137 2808
rect 9171 2805 9183 2839
rect 9646 2836 9674 3012
rect 11146 3000 11152 3012
rect 11204 3000 11210 3052
rect 11514 3040 11520 3052
rect 11475 3012 11520 3040
rect 11514 3000 11520 3012
rect 11572 3000 11578 3052
rect 13722 3000 13728 3052
rect 13780 3040 13786 3052
rect 14108 3049 14136 3080
rect 14274 3068 14280 3080
rect 14332 3068 14338 3120
rect 15942 3111 16000 3117
rect 15942 3077 15954 3111
rect 15988 3108 16000 3111
rect 15988 3080 16059 3108
rect 15988 3077 16000 3080
rect 15942 3071 16000 3077
rect 14093 3043 14151 3049
rect 14093 3040 14105 3043
rect 13780 3012 14105 3040
rect 13780 3000 13786 3012
rect 14093 3009 14105 3012
rect 14139 3009 14151 3043
rect 16031 3040 16059 3080
rect 16298 3068 16304 3120
rect 16356 3108 16362 3120
rect 16776 3108 16804 3148
rect 17037 3145 17049 3148
rect 17083 3176 17095 3179
rect 18325 3179 18383 3185
rect 17083 3148 18092 3176
rect 17083 3145 17095 3148
rect 17037 3139 17095 3145
rect 17862 3108 17868 3120
rect 16356 3080 16804 3108
rect 17032 3080 17868 3108
rect 16356 3068 16362 3080
rect 16209 3043 16267 3049
rect 16031 3012 16160 3040
rect 14093 3003 14151 3009
rect 11164 2972 11192 3000
rect 12069 2975 12127 2981
rect 12069 2972 12081 2975
rect 11164 2944 12081 2972
rect 12069 2941 12081 2944
rect 12115 2941 12127 2975
rect 12069 2935 12127 2941
rect 13354 2932 13360 2984
rect 13412 2972 13418 2984
rect 14277 2975 14335 2981
rect 14277 2972 14289 2975
rect 13412 2944 14289 2972
rect 13412 2932 13418 2944
rect 14277 2941 14289 2944
rect 14323 2941 14335 2975
rect 16132 2972 16160 3012
rect 16209 3009 16221 3043
rect 16255 3040 16267 3043
rect 16850 3040 16856 3052
rect 16255 3012 16856 3040
rect 16255 3009 16267 3012
rect 16209 3003 16267 3009
rect 16850 3000 16856 3012
rect 16908 3000 16914 3052
rect 17032 2972 17060 3080
rect 17236 2981 17264 3080
rect 17862 3068 17868 3080
rect 17920 3068 17926 3120
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3040 17739 3043
rect 17954 3040 17960 3052
rect 17727 3012 17960 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 17954 3000 17960 3012
rect 18012 3000 18018 3052
rect 18064 3040 18092 3148
rect 18325 3145 18337 3179
rect 18371 3176 18383 3179
rect 18506 3176 18512 3188
rect 18371 3148 18512 3176
rect 18371 3145 18383 3148
rect 18325 3139 18383 3145
rect 18506 3136 18512 3148
rect 18564 3136 18570 3188
rect 18598 3136 18604 3188
rect 18656 3176 18662 3188
rect 18693 3179 18751 3185
rect 18693 3176 18705 3179
rect 18656 3148 18705 3176
rect 18656 3136 18662 3148
rect 18693 3145 18705 3148
rect 18739 3145 18751 3179
rect 18693 3139 18751 3145
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 20070 3176 20076 3188
rect 19392 3148 20076 3176
rect 19392 3136 19398 3148
rect 20070 3136 20076 3148
rect 20128 3136 20134 3188
rect 18230 3068 18236 3120
rect 18288 3108 18294 3120
rect 18785 3111 18843 3117
rect 18785 3108 18797 3111
rect 18288 3080 18797 3108
rect 18288 3068 18294 3080
rect 18785 3077 18797 3080
rect 18831 3077 18843 3111
rect 18785 3071 18843 3077
rect 18874 3068 18880 3120
rect 18932 3108 18938 3120
rect 18932 3080 20852 3108
rect 18932 3068 18938 3080
rect 19705 3043 19763 3049
rect 19705 3040 19717 3043
rect 18064 3012 19717 3040
rect 19705 3009 19717 3012
rect 19751 3040 19763 3043
rect 19794 3040 19800 3052
rect 19751 3012 19800 3040
rect 19751 3009 19763 3012
rect 19705 3003 19763 3009
rect 19794 3000 19800 3012
rect 19852 3000 19858 3052
rect 20530 3040 20536 3052
rect 20491 3012 20536 3040
rect 20530 3000 20536 3012
rect 20588 3000 20594 3052
rect 20824 3049 20852 3080
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3009 20867 3043
rect 20809 3003 20867 3009
rect 16132 2944 17060 2972
rect 17129 2975 17187 2981
rect 14277 2935 14335 2941
rect 17129 2941 17141 2975
rect 17175 2941 17187 2975
rect 17129 2935 17187 2941
rect 17221 2975 17279 2981
rect 17221 2941 17233 2975
rect 17267 2941 17279 2975
rect 17221 2935 17279 2941
rect 13906 2864 13912 2916
rect 13964 2904 13970 2916
rect 14918 2904 14924 2916
rect 13964 2876 14924 2904
rect 13964 2864 13970 2876
rect 14918 2864 14924 2876
rect 14976 2864 14982 2916
rect 16206 2864 16212 2916
rect 16264 2904 16270 2916
rect 17144 2904 17172 2935
rect 17494 2932 17500 2984
rect 17552 2972 17558 2984
rect 17770 2972 17776 2984
rect 17552 2944 17776 2972
rect 17552 2932 17558 2944
rect 17770 2932 17776 2944
rect 17828 2932 17834 2984
rect 18966 2972 18972 2984
rect 18927 2944 18972 2972
rect 18966 2932 18972 2944
rect 19024 2932 19030 2984
rect 19426 2972 19432 2984
rect 19387 2944 19432 2972
rect 19426 2932 19432 2944
rect 19484 2932 19490 2984
rect 16264 2876 18000 2904
rect 16264 2864 16270 2876
rect 11514 2836 11520 2848
rect 9646 2808 11520 2836
rect 9125 2799 9183 2805
rect 11514 2796 11520 2808
rect 11572 2796 11578 2848
rect 11698 2836 11704 2848
rect 11659 2808 11704 2836
rect 11698 2796 11704 2808
rect 11756 2796 11762 2848
rect 13354 2796 13360 2848
rect 13412 2836 13418 2848
rect 17865 2839 17923 2845
rect 17865 2836 17877 2839
rect 13412 2808 17877 2836
rect 13412 2796 13418 2808
rect 17865 2805 17877 2808
rect 17911 2805 17923 2839
rect 17972 2836 18000 2876
rect 18138 2864 18144 2916
rect 18196 2904 18202 2916
rect 21082 2904 21088 2916
rect 18196 2876 21088 2904
rect 18196 2864 18202 2876
rect 21082 2864 21088 2876
rect 21140 2864 21146 2916
rect 20254 2836 20260 2848
rect 17972 2808 20260 2836
rect 17865 2799 17923 2805
rect 20254 2796 20260 2808
rect 20312 2796 20318 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 3234 2592 3240 2644
rect 3292 2632 3298 2644
rect 3421 2635 3479 2641
rect 3421 2632 3433 2635
rect 3292 2604 3433 2632
rect 3292 2592 3298 2604
rect 3421 2601 3433 2604
rect 3467 2601 3479 2635
rect 3421 2595 3479 2601
rect 6457 2635 6515 2641
rect 6457 2601 6469 2635
rect 6503 2632 6515 2635
rect 6730 2632 6736 2644
rect 6503 2604 6736 2632
rect 6503 2601 6515 2604
rect 6457 2595 6515 2601
rect 6730 2592 6736 2604
rect 6788 2592 6794 2644
rect 6917 2635 6975 2641
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7098 2632 7104 2644
rect 6963 2604 7104 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7098 2592 7104 2604
rect 7156 2592 7162 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7926 2632 7932 2644
rect 7248 2604 7932 2632
rect 7248 2592 7254 2604
rect 7926 2592 7932 2604
rect 7984 2592 7990 2644
rect 8662 2592 8668 2644
rect 8720 2632 8726 2644
rect 8941 2635 8999 2641
rect 8941 2632 8953 2635
rect 8720 2604 8953 2632
rect 8720 2592 8726 2604
rect 8941 2601 8953 2604
rect 8987 2601 8999 2635
rect 8941 2595 8999 2601
rect 11054 2592 11060 2644
rect 11112 2632 11118 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 11112 2604 11161 2632
rect 11112 2592 11118 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 12526 2632 12532 2644
rect 11149 2595 11207 2601
rect 11808 2604 12532 2632
rect 3326 2564 3332 2576
rect 2516 2536 3332 2564
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2317 2431 2375 2437
rect 2317 2428 2329 2431
rect 2004 2400 2329 2428
rect 2004 2388 2010 2400
rect 2317 2397 2329 2400
rect 2363 2428 2375 2431
rect 2516 2428 2544 2536
rect 3326 2524 3332 2536
rect 3384 2524 3390 2576
rect 5353 2567 5411 2573
rect 5353 2533 5365 2567
rect 5399 2564 5411 2567
rect 7558 2564 7564 2576
rect 5399 2536 7564 2564
rect 5399 2533 5411 2536
rect 5353 2527 5411 2533
rect 7558 2524 7564 2536
rect 7616 2524 7622 2576
rect 10137 2567 10195 2573
rect 10137 2533 10149 2567
rect 10183 2564 10195 2567
rect 11808 2564 11836 2604
rect 12526 2592 12532 2604
rect 12584 2592 12590 2644
rect 13173 2635 13231 2641
rect 13173 2601 13185 2635
rect 13219 2632 13231 2635
rect 13262 2632 13268 2644
rect 13219 2604 13268 2632
rect 13219 2601 13231 2604
rect 13173 2595 13231 2601
rect 13262 2592 13268 2604
rect 13320 2592 13326 2644
rect 15562 2592 15568 2644
rect 15620 2632 15626 2644
rect 15657 2635 15715 2641
rect 15657 2632 15669 2635
rect 15620 2604 15669 2632
rect 15620 2592 15626 2604
rect 15657 2601 15669 2604
rect 15703 2601 15715 2635
rect 15657 2595 15715 2601
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 16669 2635 16727 2641
rect 16669 2632 16681 2635
rect 15804 2604 16681 2632
rect 15804 2592 15810 2604
rect 16669 2601 16681 2604
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 17494 2592 17500 2644
rect 17552 2632 17558 2644
rect 19702 2632 19708 2644
rect 17552 2604 19708 2632
rect 17552 2592 17558 2604
rect 19702 2592 19708 2604
rect 19760 2592 19766 2644
rect 10183 2536 11836 2564
rect 10183 2533 10195 2536
rect 10137 2527 10195 2533
rect 12158 2524 12164 2576
rect 12216 2564 12222 2576
rect 13541 2567 13599 2573
rect 13541 2564 13553 2567
rect 12216 2536 13553 2564
rect 12216 2524 12222 2536
rect 13541 2533 13553 2536
rect 13587 2533 13599 2567
rect 13541 2527 13599 2533
rect 14384 2536 16344 2564
rect 3050 2496 3056 2508
rect 2792 2468 3056 2496
rect 2792 2437 2820 2468
rect 3050 2456 3056 2468
rect 3108 2496 3114 2508
rect 3878 2496 3884 2508
rect 3108 2468 3884 2496
rect 3108 2456 3114 2468
rect 3878 2456 3884 2468
rect 3936 2456 3942 2508
rect 7190 2496 7196 2508
rect 6012 2468 7196 2496
rect 2363 2400 2544 2428
rect 2777 2431 2835 2437
rect 2363 2397 2375 2400
rect 2317 2391 2375 2397
rect 2777 2397 2789 2431
rect 2823 2397 2835 2431
rect 3234 2428 3240 2440
rect 3195 2400 3240 2428
rect 2777 2391 2835 2397
rect 3234 2388 3240 2400
rect 3292 2388 3298 2440
rect 3973 2431 4031 2437
rect 3973 2397 3985 2431
rect 4019 2428 4031 2431
rect 4062 2428 4068 2440
rect 4019 2400 4068 2428
rect 4019 2397 4031 2400
rect 3973 2391 4031 2397
rect 4062 2388 4068 2400
rect 4120 2388 4126 2440
rect 4433 2431 4491 2437
rect 4433 2397 4445 2431
rect 4479 2428 4491 2431
rect 4614 2428 4620 2440
rect 4479 2400 4620 2428
rect 4479 2397 4491 2400
rect 4433 2391 4491 2397
rect 4614 2388 4620 2400
rect 4672 2388 4678 2440
rect 4890 2428 4896 2440
rect 4851 2400 4896 2428
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 5074 2388 5080 2440
rect 5132 2428 5138 2440
rect 6012 2437 6040 2468
rect 7190 2456 7196 2468
rect 7248 2456 7254 2508
rect 9490 2496 9496 2508
rect 9451 2468 9496 2496
rect 9490 2456 9496 2468
rect 9548 2456 9554 2508
rect 10502 2496 10508 2508
rect 10463 2468 10508 2496
rect 10502 2456 10508 2468
rect 10560 2456 10566 2508
rect 10689 2499 10747 2505
rect 10689 2465 10701 2499
rect 10735 2496 10747 2499
rect 10778 2496 10784 2508
rect 10735 2468 10784 2496
rect 10735 2465 10747 2468
rect 10689 2459 10747 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 10870 2456 10876 2508
rect 10928 2496 10934 2508
rect 10928 2468 12296 2496
rect 10928 2456 10934 2468
rect 5997 2431 6055 2437
rect 5132 2400 5672 2428
rect 5132 2388 5138 2400
rect 198 2320 204 2372
rect 256 2360 262 2372
rect 1394 2360 1400 2372
rect 256 2332 1400 2360
rect 256 2320 262 2332
rect 1394 2320 1400 2332
rect 1452 2360 1458 2372
rect 1673 2363 1731 2369
rect 1673 2360 1685 2363
rect 1452 2332 1685 2360
rect 1452 2320 1458 2332
rect 1673 2329 1685 2332
rect 1719 2329 1731 2363
rect 5534 2360 5540 2372
rect 1673 2323 1731 2329
rect 2516 2332 5540 2360
rect 1765 2295 1823 2301
rect 1765 2261 1777 2295
rect 1811 2292 1823 2295
rect 2406 2292 2412 2304
rect 1811 2264 2412 2292
rect 1811 2261 1823 2264
rect 1765 2255 1823 2261
rect 2406 2252 2412 2264
rect 2464 2252 2470 2304
rect 2516 2301 2544 2332
rect 5534 2320 5540 2332
rect 5592 2320 5598 2372
rect 5644 2360 5672 2400
rect 5997 2397 6009 2431
rect 6043 2397 6055 2431
rect 6730 2428 6736 2440
rect 6691 2400 6736 2428
rect 5997 2391 6055 2397
rect 6730 2388 6736 2400
rect 6788 2388 6794 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8573 2431 8631 2437
rect 8573 2428 8585 2431
rect 7800 2400 8585 2428
rect 7800 2388 7806 2400
rect 8573 2397 8585 2400
rect 8619 2397 8631 2431
rect 8573 2391 8631 2397
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 9401 2431 9459 2437
rect 9401 2428 9413 2431
rect 8720 2400 9413 2428
rect 8720 2388 8726 2400
rect 9401 2397 9413 2400
rect 9447 2397 9459 2431
rect 9401 2391 9459 2397
rect 9953 2431 10011 2437
rect 9953 2397 9965 2431
rect 9999 2428 10011 2431
rect 10134 2428 10140 2440
rect 9999 2400 10140 2428
rect 9999 2397 10011 2400
rect 9953 2391 10011 2397
rect 10134 2388 10140 2400
rect 10192 2388 10198 2440
rect 11238 2388 11244 2440
rect 11296 2428 11302 2440
rect 11517 2431 11575 2437
rect 11517 2428 11529 2431
rect 11296 2400 11529 2428
rect 11296 2388 11302 2400
rect 11517 2397 11529 2400
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 7834 2360 7840 2372
rect 5644 2332 7840 2360
rect 7834 2320 7840 2332
rect 7892 2320 7898 2372
rect 8328 2363 8386 2369
rect 8328 2329 8340 2363
rect 8374 2360 8386 2363
rect 12161 2363 12219 2369
rect 12161 2360 12173 2363
rect 8374 2332 12173 2360
rect 8374 2329 8386 2332
rect 8328 2323 8386 2329
rect 12161 2329 12173 2332
rect 12207 2329 12219 2363
rect 12268 2360 12296 2468
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12529 2499 12587 2505
rect 12529 2496 12541 2499
rect 12492 2468 12541 2496
rect 12492 2456 12498 2468
rect 12529 2465 12541 2468
rect 12575 2465 12587 2499
rect 12529 2459 12587 2465
rect 12802 2388 12808 2440
rect 12860 2428 12866 2440
rect 14384 2437 14412 2536
rect 15105 2499 15163 2505
rect 15105 2465 15117 2499
rect 15151 2496 15163 2499
rect 15194 2496 15200 2508
rect 15151 2468 15200 2496
rect 15151 2465 15163 2468
rect 15105 2459 15163 2465
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 16316 2496 16344 2536
rect 16390 2524 16396 2576
rect 16448 2564 16454 2576
rect 17037 2567 17095 2573
rect 17037 2564 17049 2567
rect 16448 2536 17049 2564
rect 16448 2524 16454 2536
rect 17037 2533 17049 2536
rect 17083 2533 17095 2567
rect 17037 2527 17095 2533
rect 17770 2524 17776 2576
rect 17828 2564 17834 2576
rect 17828 2536 18644 2564
rect 17828 2524 17834 2536
rect 17310 2496 17316 2508
rect 16316 2468 17316 2496
rect 17310 2456 17316 2468
rect 17368 2456 17374 2508
rect 17494 2496 17500 2508
rect 17455 2468 17500 2496
rect 17494 2456 17500 2468
rect 17552 2456 17558 2508
rect 17681 2499 17739 2505
rect 17681 2465 17693 2499
rect 17727 2496 17739 2499
rect 18414 2496 18420 2508
rect 17727 2468 18420 2496
rect 17727 2465 17739 2468
rect 17681 2459 17739 2465
rect 18414 2456 18420 2468
rect 18472 2456 18478 2508
rect 18616 2505 18644 2536
rect 18601 2499 18659 2505
rect 18601 2465 18613 2499
rect 18647 2496 18659 2499
rect 19610 2496 19616 2508
rect 18647 2468 19616 2496
rect 18647 2465 18659 2468
rect 18601 2459 18659 2465
rect 19610 2456 19616 2468
rect 19668 2456 19674 2508
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 20254 2496 20260 2508
rect 19751 2468 20260 2496
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 20254 2456 20260 2468
rect 20312 2456 20318 2508
rect 13725 2431 13783 2437
rect 13725 2428 13737 2431
rect 12860 2400 13737 2428
rect 12860 2388 12866 2400
rect 13725 2397 13737 2400
rect 13771 2397 13783 2431
rect 13725 2391 13783 2397
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2397 14427 2431
rect 14369 2391 14427 2397
rect 14458 2388 14464 2440
rect 14516 2428 14522 2440
rect 15930 2428 15936 2440
rect 14516 2400 15332 2428
rect 15891 2400 15936 2428
rect 14516 2388 14522 2400
rect 15197 2363 15255 2369
rect 15197 2360 15209 2363
rect 12268 2332 15209 2360
rect 12161 2323 12219 2329
rect 15197 2329 15209 2332
rect 15243 2329 15255 2363
rect 15304 2360 15332 2400
rect 15930 2388 15936 2400
rect 15988 2388 15994 2440
rect 18874 2428 18880 2440
rect 18835 2400 18880 2428
rect 18874 2388 18880 2400
rect 18932 2388 18938 2440
rect 19426 2428 19432 2440
rect 19387 2400 19432 2428
rect 19426 2388 19432 2400
rect 19484 2388 19490 2440
rect 20530 2428 20536 2440
rect 20443 2400 20536 2428
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 20809 2431 20867 2437
rect 20809 2397 20821 2431
rect 20855 2397 20867 2431
rect 20809 2391 20867 2397
rect 15304 2332 16160 2360
rect 15197 2323 15255 2329
rect 2501 2295 2559 2301
rect 2501 2261 2513 2295
rect 2547 2261 2559 2295
rect 2958 2292 2964 2304
rect 2919 2264 2964 2292
rect 2501 2255 2559 2261
rect 2958 2252 2964 2264
rect 3016 2252 3022 2304
rect 4154 2292 4160 2304
rect 4115 2264 4160 2292
rect 4154 2252 4160 2264
rect 4212 2252 4218 2304
rect 4614 2292 4620 2304
rect 4575 2264 4620 2292
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 5074 2292 5080 2304
rect 5035 2264 5080 2292
rect 5074 2252 5080 2264
rect 5132 2252 5138 2304
rect 7650 2252 7656 2304
rect 7708 2292 7714 2304
rect 9309 2295 9367 2301
rect 9309 2292 9321 2295
rect 7708 2264 9321 2292
rect 7708 2252 7714 2264
rect 9309 2261 9321 2264
rect 9355 2261 9367 2295
rect 9309 2255 9367 2261
rect 10778 2252 10784 2304
rect 10836 2292 10842 2304
rect 10836 2264 10881 2292
rect 10836 2252 10842 2264
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 12713 2295 12771 2301
rect 12713 2292 12725 2295
rect 11020 2264 12725 2292
rect 11020 2252 11026 2264
rect 12713 2261 12725 2264
rect 12759 2261 12771 2295
rect 12713 2255 12771 2261
rect 12802 2252 12808 2304
rect 12860 2292 12866 2304
rect 14182 2292 14188 2304
rect 12860 2264 12905 2292
rect 14143 2264 14188 2292
rect 12860 2252 12866 2264
rect 14182 2252 14188 2264
rect 14240 2252 14246 2304
rect 15286 2292 15292 2304
rect 15247 2264 15292 2292
rect 15286 2252 15292 2264
rect 15344 2252 15350 2304
rect 16132 2301 16160 2332
rect 18414 2320 18420 2372
rect 18472 2360 18478 2372
rect 20548 2360 20576 2388
rect 18472 2332 20576 2360
rect 18472 2320 18478 2332
rect 16117 2295 16175 2301
rect 16117 2261 16129 2295
rect 16163 2261 16175 2295
rect 16117 2255 16175 2261
rect 17034 2252 17040 2304
rect 17092 2292 17098 2304
rect 17405 2295 17463 2301
rect 17405 2292 17417 2295
rect 17092 2264 17417 2292
rect 17092 2252 17098 2264
rect 17405 2261 17417 2264
rect 17451 2292 17463 2295
rect 20824 2292 20852 2391
rect 17451 2264 20852 2292
rect 17451 2261 17463 2264
rect 17405 2255 17463 2261
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
rect 3234 2048 3240 2100
rect 3292 2088 3298 2100
rect 4430 2088 4436 2100
rect 3292 2060 4436 2088
rect 3292 2048 3298 2060
rect 4430 2048 4436 2060
rect 4488 2088 4494 2100
rect 4982 2088 4988 2100
rect 4488 2060 4988 2088
rect 4488 2048 4494 2060
rect 4982 2048 4988 2060
rect 5040 2048 5046 2100
rect 5350 2048 5356 2100
rect 5408 2088 5414 2100
rect 6730 2088 6736 2100
rect 5408 2060 6736 2088
rect 5408 2048 5414 2060
rect 6730 2048 6736 2060
rect 6788 2088 6794 2100
rect 11146 2088 11152 2100
rect 6788 2060 11152 2088
rect 6788 2048 6794 2060
rect 11146 2048 11152 2060
rect 11204 2048 11210 2100
rect 14182 2048 14188 2100
rect 14240 2088 14246 2100
rect 22094 2088 22100 2100
rect 14240 2060 22100 2088
rect 14240 2048 14246 2060
rect 22094 2048 22100 2060
rect 22152 2048 22158 2100
rect 5074 1980 5080 2032
rect 5132 2020 5138 2032
rect 15930 2020 15936 2032
rect 5132 1992 15936 2020
rect 5132 1980 5138 1992
rect 15930 1980 15936 1992
rect 15988 1980 15994 2032
rect 2406 1912 2412 1964
rect 2464 1952 2470 1964
rect 7190 1952 7196 1964
rect 2464 1924 7196 1952
rect 2464 1912 2470 1924
rect 7190 1912 7196 1924
rect 7248 1912 7254 1964
rect 7466 1912 7472 1964
rect 7524 1952 7530 1964
rect 15286 1952 15292 1964
rect 7524 1924 15292 1952
rect 7524 1912 7530 1924
rect 15286 1912 15292 1924
rect 15344 1912 15350 1964
rect 4614 1844 4620 1896
rect 4672 1884 4678 1896
rect 10962 1884 10968 1896
rect 4672 1856 10968 1884
rect 4672 1844 4678 1856
rect 10962 1844 10968 1856
rect 11020 1844 11026 1896
rect 5994 1776 6000 1828
rect 6052 1816 6058 1828
rect 12802 1816 12808 1828
rect 6052 1788 12808 1816
rect 6052 1776 6058 1788
rect 12802 1776 12808 1788
rect 12860 1776 12866 1828
rect 19334 1776 19340 1828
rect 19392 1816 19398 1828
rect 20070 1816 20076 1828
rect 19392 1788 20076 1816
rect 19392 1776 19398 1788
rect 20070 1776 20076 1788
rect 20128 1776 20134 1828
rect 5258 1708 5264 1760
rect 5316 1748 5322 1760
rect 10778 1748 10784 1760
rect 5316 1720 10784 1748
rect 5316 1708 5322 1720
rect 10778 1708 10784 1720
rect 10836 1708 10842 1760
rect 4154 1640 4160 1692
rect 4212 1680 4218 1692
rect 10686 1680 10692 1692
rect 4212 1652 10692 1680
rect 4212 1640 4218 1652
rect 10686 1640 10692 1652
rect 10744 1640 10750 1692
rect 4062 1572 4068 1624
rect 4120 1612 4126 1624
rect 6178 1612 6184 1624
rect 4120 1584 6184 1612
rect 4120 1572 4126 1584
rect 6178 1572 6184 1584
rect 6236 1572 6242 1624
rect 7190 1572 7196 1624
rect 7248 1612 7254 1624
rect 12894 1612 12900 1624
rect 7248 1584 12900 1612
rect 7248 1572 7254 1584
rect 12894 1572 12900 1584
rect 12952 1572 12958 1624
rect 5718 1504 5724 1556
rect 5776 1544 5782 1556
rect 9490 1544 9496 1556
rect 5776 1516 9496 1544
rect 5776 1504 5782 1516
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 19518 1368 19524 1420
rect 19576 1368 19582 1420
rect 2590 1300 2596 1352
rect 2648 1340 2654 1352
rect 19426 1340 19432 1352
rect 2648 1312 19432 1340
rect 2648 1300 2654 1312
rect 19426 1300 19432 1312
rect 19484 1300 19490 1352
rect 3510 1232 3516 1284
rect 3568 1272 3574 1284
rect 19536 1272 19564 1368
rect 3568 1244 19564 1272
rect 3568 1232 3574 1244
rect 16574 1096 16580 1148
rect 16632 1136 16638 1148
rect 18138 1136 18144 1148
rect 16632 1108 18144 1136
rect 16632 1096 16638 1108
rect 18138 1096 18144 1108
rect 18196 1096 18202 1148
<< via1 >>
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 19708 20544 19760 20596
rect 19248 20476 19300 20528
rect 5724 20408 5776 20460
rect 17224 20408 17276 20460
rect 18880 20408 18932 20460
rect 20536 20451 20588 20460
rect 20536 20417 20545 20451
rect 20545 20417 20579 20451
rect 20579 20417 20588 20451
rect 20536 20408 20588 20417
rect 21088 20451 21140 20460
rect 21088 20417 21097 20451
rect 21097 20417 21131 20451
rect 21131 20417 21140 20451
rect 21088 20408 21140 20417
rect 6000 20247 6052 20256
rect 6000 20213 6009 20247
rect 6009 20213 6043 20247
rect 6043 20213 6052 20247
rect 6000 20204 6052 20213
rect 17316 20247 17368 20256
rect 17316 20213 17325 20247
rect 17325 20213 17359 20247
rect 17359 20213 17368 20247
rect 17316 20204 17368 20213
rect 20168 20204 20220 20256
rect 20720 20247 20772 20256
rect 20720 20213 20729 20247
rect 20729 20213 20763 20247
rect 20763 20213 20772 20247
rect 20720 20204 20772 20213
rect 21364 20204 21416 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 20352 20000 20404 20052
rect 20812 20000 20864 20052
rect 6000 19796 6052 19848
rect 12900 19839 12952 19848
rect 12900 19805 12909 19839
rect 12909 19805 12943 19839
rect 12943 19805 12952 19839
rect 12900 19796 12952 19805
rect 19524 19839 19576 19848
rect 6552 19771 6604 19780
rect 6552 19737 6561 19771
rect 6561 19737 6595 19771
rect 6595 19737 6604 19771
rect 6552 19728 6604 19737
rect 19524 19805 19533 19839
rect 19533 19805 19567 19839
rect 19567 19805 19576 19839
rect 19524 19796 19576 19805
rect 19892 19728 19944 19780
rect 20812 19796 20864 19848
rect 21272 19703 21324 19712
rect 21272 19669 21281 19703
rect 21281 19669 21315 19703
rect 21315 19669 21324 19703
rect 21272 19660 21324 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 19524 19456 19576 19508
rect 19892 19456 19944 19508
rect 20628 19456 20680 19508
rect 16212 19388 16264 19440
rect 18420 19363 18472 19372
rect 18420 19329 18429 19363
rect 18429 19329 18463 19363
rect 18463 19329 18472 19363
rect 18420 19320 18472 19329
rect 19524 19363 19576 19372
rect 19524 19329 19533 19363
rect 19533 19329 19567 19363
rect 19567 19329 19576 19363
rect 19524 19320 19576 19329
rect 20444 19388 20496 19440
rect 20720 19320 20772 19372
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 12900 18912 12952 18964
rect 20536 18912 20588 18964
rect 21088 18912 21140 18964
rect 9772 18708 9824 18760
rect 11244 18708 11296 18760
rect 20260 18708 20312 18760
rect 20996 18708 21048 18760
rect 21272 18615 21324 18624
rect 21272 18581 21281 18615
rect 21281 18581 21315 18615
rect 21315 18581 21324 18615
rect 21272 18572 21324 18581
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 20812 18368 20864 18420
rect 8576 18232 8628 18284
rect 12256 18275 12308 18284
rect 12256 18241 12265 18275
rect 12265 18241 12299 18275
rect 12299 18241 12308 18275
rect 12256 18232 12308 18241
rect 20812 18275 20864 18284
rect 20812 18241 20821 18275
rect 20821 18241 20855 18275
rect 20855 18241 20864 18275
rect 20812 18232 20864 18241
rect 20904 18232 20956 18284
rect 20260 18028 20312 18080
rect 20536 18028 20588 18080
rect 21364 18028 21416 18080
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 12256 17824 12308 17876
rect 20720 17824 20772 17876
rect 12256 17620 12308 17672
rect 20076 17663 20128 17672
rect 20076 17629 20085 17663
rect 20085 17629 20119 17663
rect 20119 17629 20128 17663
rect 20076 17620 20128 17629
rect 20536 17663 20588 17672
rect 20536 17629 20545 17663
rect 20545 17629 20579 17663
rect 20579 17629 20588 17663
rect 20536 17620 20588 17629
rect 21088 17663 21140 17672
rect 21088 17629 21097 17663
rect 21097 17629 21131 17663
rect 21131 17629 21140 17663
rect 21088 17620 21140 17629
rect 20720 17527 20772 17536
rect 20720 17493 20729 17527
rect 20729 17493 20763 17527
rect 20763 17493 20772 17527
rect 20720 17484 20772 17493
rect 21272 17527 21324 17536
rect 21272 17493 21281 17527
rect 21281 17493 21315 17527
rect 21315 17493 21324 17527
rect 21272 17484 21324 17493
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 20076 17323 20128 17332
rect 20076 17289 20085 17323
rect 20085 17289 20119 17323
rect 20119 17289 20128 17323
rect 20076 17280 20128 17289
rect 20904 17280 20956 17332
rect 15108 17212 15160 17264
rect 19524 17212 19576 17264
rect 14280 17144 14332 17196
rect 17960 17076 18012 17128
rect 20812 17144 20864 17196
rect 21364 16940 21416 16992
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 21088 16736 21140 16788
rect 18236 16575 18288 16584
rect 18236 16541 18245 16575
rect 18245 16541 18279 16575
rect 18279 16541 18288 16575
rect 18236 16532 18288 16541
rect 15200 16464 15252 16516
rect 20904 16532 20956 16584
rect 20996 16396 21048 16448
rect 21272 16439 21324 16448
rect 21272 16405 21281 16439
rect 21281 16405 21315 16439
rect 21315 16405 21324 16439
rect 21272 16396 21324 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 17960 16192 18012 16244
rect 20628 16192 20680 16244
rect 20812 16235 20864 16244
rect 20812 16201 20821 16235
rect 20821 16201 20855 16235
rect 20855 16201 20864 16235
rect 20812 16192 20864 16201
rect 14464 16056 14516 16108
rect 17868 16056 17920 16108
rect 21088 16099 21140 16108
rect 12992 15988 13044 16040
rect 21088 16065 21097 16099
rect 21097 16065 21131 16099
rect 21131 16065 21140 16099
rect 21088 16056 21140 16065
rect 19616 15852 19668 15904
rect 20076 15852 20128 15904
rect 21364 15852 21416 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 21088 15648 21140 15700
rect 15292 15512 15344 15564
rect 18972 15444 19024 15496
rect 20352 15444 20404 15496
rect 20720 15444 20772 15496
rect 19708 15308 19760 15360
rect 20260 15308 20312 15360
rect 21088 15308 21140 15360
rect 21272 15351 21324 15360
rect 21272 15317 21281 15351
rect 21281 15317 21315 15351
rect 21315 15317 21324 15351
rect 21272 15308 21324 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 12992 15104 13044 15156
rect 20720 15104 20772 15156
rect 9496 14968 9548 15020
rect 11704 14968 11756 15020
rect 19616 14968 19668 15020
rect 19064 14900 19116 14952
rect 15200 14832 15252 14884
rect 17132 14832 17184 14884
rect 19984 14968 20036 15020
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 20904 14832 20956 14884
rect 17960 14764 18012 14816
rect 19800 14764 19852 14816
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 15476 14560 15528 14612
rect 18052 14492 18104 14544
rect 18604 14492 18656 14544
rect 8668 14356 8720 14408
rect 18052 14356 18104 14408
rect 18144 14356 18196 14408
rect 17132 14288 17184 14340
rect 20628 14560 20680 14612
rect 19616 14492 19668 14544
rect 20536 14492 20588 14544
rect 19524 14356 19576 14408
rect 19708 14424 19760 14476
rect 19892 14399 19944 14408
rect 19892 14365 19901 14399
rect 19901 14365 19935 14399
rect 19935 14365 19944 14399
rect 19892 14356 19944 14365
rect 20444 14356 20496 14408
rect 21088 14399 21140 14408
rect 21088 14365 21097 14399
rect 21097 14365 21131 14399
rect 21131 14365 21140 14399
rect 21088 14356 21140 14365
rect 12808 14220 12860 14272
rect 20996 14288 21048 14340
rect 19524 14220 19576 14272
rect 20076 14220 20128 14272
rect 20628 14220 20680 14272
rect 21272 14263 21324 14272
rect 21272 14229 21281 14263
rect 21281 14229 21315 14263
rect 21315 14229 21324 14263
rect 21272 14220 21324 14229
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 15292 14016 15344 14068
rect 18144 14059 18196 14068
rect 18144 14025 18153 14059
rect 18153 14025 18187 14059
rect 18187 14025 18196 14059
rect 18144 14016 18196 14025
rect 20352 14016 20404 14068
rect 16120 13948 16172 14000
rect 12072 13880 12124 13932
rect 17960 13923 18012 13932
rect 15384 13812 15436 13864
rect 17408 13855 17460 13864
rect 17408 13821 17417 13855
rect 17417 13821 17451 13855
rect 17451 13821 17460 13855
rect 17408 13812 17460 13821
rect 17960 13889 17969 13923
rect 17969 13889 18003 13923
rect 18003 13889 18012 13923
rect 17960 13880 18012 13889
rect 18512 13880 18564 13932
rect 18052 13812 18104 13864
rect 19708 13812 19760 13864
rect 20076 13812 20128 13864
rect 20628 13880 20680 13932
rect 21640 13812 21692 13864
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 19984 13472 20036 13524
rect 20352 13515 20404 13524
rect 20352 13481 20361 13515
rect 20361 13481 20395 13515
rect 20395 13481 20404 13515
rect 20352 13472 20404 13481
rect 14924 13404 14976 13456
rect 13544 13311 13596 13320
rect 13544 13277 13553 13311
rect 13553 13277 13587 13311
rect 13587 13277 13596 13311
rect 13544 13268 13596 13277
rect 17224 13311 17276 13320
rect 17224 13277 17242 13311
rect 17242 13277 17276 13311
rect 17224 13268 17276 13277
rect 17500 13311 17552 13320
rect 17500 13277 17509 13311
rect 17509 13277 17543 13311
rect 17543 13277 17552 13311
rect 17500 13268 17552 13277
rect 18052 13268 18104 13320
rect 19524 13336 19576 13388
rect 18880 13268 18932 13320
rect 19800 13268 19852 13320
rect 20720 13311 20772 13320
rect 20720 13277 20729 13311
rect 20729 13277 20763 13311
rect 20763 13277 20772 13311
rect 20720 13268 20772 13277
rect 17316 13200 17368 13252
rect 15384 13132 15436 13184
rect 17224 13132 17276 13184
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 18696 13132 18748 13141
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 21088 13132 21140 13184
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 18696 12928 18748 12980
rect 16948 12860 17000 12912
rect 17040 12792 17092 12844
rect 17684 12792 17736 12844
rect 18788 12835 18840 12844
rect 15844 12724 15896 12776
rect 18788 12801 18797 12835
rect 18797 12801 18831 12835
rect 18831 12801 18840 12835
rect 18788 12792 18840 12801
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 20628 12835 20680 12844
rect 20628 12801 20637 12835
rect 20637 12801 20671 12835
rect 20671 12801 20680 12835
rect 20628 12792 20680 12801
rect 18420 12699 18472 12708
rect 18420 12665 18429 12699
rect 18429 12665 18463 12699
rect 18463 12665 18472 12699
rect 18420 12656 18472 12665
rect 15016 12588 15068 12640
rect 17592 12588 17644 12640
rect 17868 12588 17920 12640
rect 18144 12588 18196 12640
rect 18328 12588 18380 12640
rect 19524 12588 19576 12640
rect 20904 12588 20956 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 15476 12427 15528 12436
rect 15476 12393 15485 12427
rect 15485 12393 15519 12427
rect 15519 12393 15528 12427
rect 15476 12384 15528 12393
rect 18788 12427 18840 12436
rect 12440 12316 12492 12368
rect 18788 12393 18797 12427
rect 18797 12393 18831 12427
rect 18831 12393 18840 12427
rect 18788 12384 18840 12393
rect 21272 12427 21324 12436
rect 21272 12393 21281 12427
rect 21281 12393 21315 12427
rect 21315 12393 21324 12427
rect 21272 12384 21324 12393
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 7196 12112 7248 12164
rect 15200 12112 15252 12164
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 14372 12044 14424 12096
rect 14832 12087 14884 12096
rect 14832 12053 14841 12087
rect 14841 12053 14875 12087
rect 14875 12053 14884 12087
rect 14832 12044 14884 12053
rect 17500 12180 17552 12232
rect 16304 12044 16356 12096
rect 17132 12087 17184 12096
rect 17132 12053 17141 12087
rect 17141 12053 17175 12087
rect 17175 12053 17184 12087
rect 17132 12044 17184 12053
rect 17776 12112 17828 12164
rect 17868 12112 17920 12164
rect 19524 12223 19576 12232
rect 19524 12189 19558 12223
rect 19558 12189 19576 12223
rect 19524 12180 19576 12189
rect 20996 12180 21048 12232
rect 19800 12112 19852 12164
rect 18604 12044 18656 12096
rect 20628 12087 20680 12096
rect 20628 12053 20637 12087
rect 20637 12053 20671 12087
rect 20671 12053 20680 12087
rect 20628 12044 20680 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 12164 11840 12216 11892
rect 16212 11883 16264 11892
rect 16212 11849 16221 11883
rect 16221 11849 16255 11883
rect 16255 11849 16264 11883
rect 16212 11840 16264 11849
rect 17776 11883 17828 11892
rect 17776 11849 17785 11883
rect 17785 11849 17819 11883
rect 17819 11849 17828 11883
rect 17776 11840 17828 11849
rect 16580 11772 16632 11824
rect 17224 11772 17276 11824
rect 17500 11772 17552 11824
rect 18328 11815 18380 11824
rect 18328 11781 18362 11815
rect 18362 11781 18380 11815
rect 18328 11772 18380 11781
rect 20260 11840 20312 11892
rect 13820 11704 13872 11756
rect 14280 11704 14332 11756
rect 15200 11747 15252 11756
rect 5264 11636 5316 11688
rect 14832 11636 14884 11688
rect 15200 11713 15209 11747
rect 15209 11713 15243 11747
rect 15243 11713 15252 11747
rect 15200 11704 15252 11713
rect 17132 11747 17184 11756
rect 17132 11713 17141 11747
rect 17141 11713 17175 11747
rect 17175 11713 17184 11747
rect 17132 11704 17184 11713
rect 17776 11704 17828 11756
rect 18144 11704 18196 11756
rect 19524 11704 19576 11756
rect 15476 11636 15528 11688
rect 15752 11679 15804 11688
rect 12440 11568 12492 11620
rect 15200 11568 15252 11620
rect 15752 11645 15761 11679
rect 15761 11645 15795 11679
rect 15795 11645 15804 11679
rect 15752 11636 15804 11645
rect 17868 11636 17920 11688
rect 15844 11568 15896 11620
rect 1492 11543 1544 11552
rect 1492 11509 1501 11543
rect 1501 11509 1535 11543
rect 1535 11509 1544 11543
rect 1492 11500 1544 11509
rect 13268 11543 13320 11552
rect 13268 11509 13277 11543
rect 13277 11509 13311 11543
rect 13311 11509 13320 11543
rect 13268 11500 13320 11509
rect 14556 11543 14608 11552
rect 14556 11509 14565 11543
rect 14565 11509 14599 11543
rect 14599 11509 14608 11543
rect 14556 11500 14608 11509
rect 14648 11500 14700 11552
rect 20352 11568 20404 11620
rect 16948 11500 17000 11552
rect 17224 11500 17276 11552
rect 17960 11500 18012 11552
rect 19984 11543 20036 11552
rect 19984 11509 19993 11543
rect 19993 11509 20027 11543
rect 20027 11509 20036 11543
rect 19984 11500 20036 11509
rect 21456 11500 21508 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 16580 11296 16632 11348
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 18328 11296 18380 11348
rect 14280 11228 14332 11280
rect 15844 11228 15896 11280
rect 18604 11271 18656 11280
rect 14648 11160 14700 11212
rect 17132 11203 17184 11212
rect 17132 11169 17141 11203
rect 17141 11169 17175 11203
rect 17175 11169 17184 11203
rect 17132 11160 17184 11169
rect 14280 10999 14332 11008
rect 14280 10965 14289 10999
rect 14289 10965 14323 10999
rect 14323 10965 14332 10999
rect 14832 11092 14884 11144
rect 16948 11092 17000 11144
rect 18604 11237 18613 11271
rect 18613 11237 18647 11271
rect 18647 11237 18656 11271
rect 18604 11228 18656 11237
rect 18788 11228 18840 11280
rect 17500 11160 17552 11212
rect 17684 11160 17736 11212
rect 18972 11160 19024 11212
rect 14280 10956 14332 10965
rect 15384 10956 15436 11008
rect 17868 11024 17920 11076
rect 20996 11296 21048 11348
rect 20076 11092 20128 11144
rect 20720 11024 20772 11076
rect 20904 11067 20956 11076
rect 20904 11033 20922 11067
rect 20922 11033 20956 11067
rect 20904 11024 20956 11033
rect 16396 10956 16448 11008
rect 17132 10956 17184 11008
rect 17500 10956 17552 11008
rect 18144 10956 18196 11008
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 13820 10752 13872 10804
rect 19708 10752 19760 10804
rect 19984 10752 20036 10804
rect 20720 10752 20772 10804
rect 14556 10684 14608 10736
rect 15384 10684 15436 10736
rect 13084 10616 13136 10668
rect 14832 10616 14884 10668
rect 18328 10684 18380 10736
rect 18788 10684 18840 10736
rect 19156 10684 19208 10736
rect 19524 10684 19576 10736
rect 20352 10616 20404 10668
rect 20904 10616 20956 10668
rect 6552 10548 6604 10600
rect 6736 10480 6788 10532
rect 11980 10412 12032 10464
rect 12348 10548 12400 10600
rect 15844 10548 15896 10600
rect 17040 10480 17092 10532
rect 15568 10455 15620 10464
rect 15568 10421 15577 10455
rect 15577 10421 15611 10455
rect 15611 10421 15620 10455
rect 15568 10412 15620 10421
rect 15660 10412 15712 10464
rect 16948 10455 17000 10464
rect 16948 10421 16957 10455
rect 16957 10421 16991 10455
rect 16991 10421 17000 10455
rect 16948 10412 17000 10421
rect 18604 10591 18656 10600
rect 18604 10557 18613 10591
rect 18613 10557 18647 10591
rect 18647 10557 18656 10591
rect 18604 10548 18656 10557
rect 20628 10548 20680 10600
rect 20996 10591 21048 10600
rect 20996 10557 21005 10591
rect 21005 10557 21039 10591
rect 21039 10557 21048 10591
rect 20996 10548 21048 10557
rect 20076 10480 20128 10532
rect 19524 10412 19576 10464
rect 19708 10412 19760 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 7380 10208 7432 10260
rect 14372 10208 14424 10260
rect 15108 10208 15160 10260
rect 15752 10208 15804 10260
rect 16580 10208 16632 10260
rect 17040 10251 17092 10260
rect 17040 10217 17049 10251
rect 17049 10217 17083 10251
rect 17083 10217 17092 10251
rect 17040 10208 17092 10217
rect 20352 10251 20404 10260
rect 20352 10217 20361 10251
rect 20361 10217 20395 10251
rect 20395 10217 20404 10251
rect 20352 10208 20404 10217
rect 5448 10140 5500 10192
rect 15660 10140 15712 10192
rect 17132 10140 17184 10192
rect 17500 10140 17552 10192
rect 13820 10072 13872 10124
rect 11152 10047 11204 10056
rect 11152 10013 11161 10047
rect 11161 10013 11195 10047
rect 11195 10013 11204 10047
rect 11152 10004 11204 10013
rect 13544 10047 13596 10056
rect 13544 10013 13553 10047
rect 13553 10013 13587 10047
rect 13587 10013 13596 10047
rect 13544 10004 13596 10013
rect 14280 10004 14332 10056
rect 19616 10072 19668 10124
rect 20352 10072 20404 10124
rect 15568 10004 15620 10056
rect 15292 9936 15344 9988
rect 11796 9911 11848 9920
rect 11796 9877 11805 9911
rect 11805 9877 11839 9911
rect 11839 9877 11848 9911
rect 11796 9868 11848 9877
rect 12072 9911 12124 9920
rect 12072 9877 12081 9911
rect 12081 9877 12115 9911
rect 12115 9877 12124 9911
rect 12072 9868 12124 9877
rect 12440 9868 12492 9920
rect 12900 9911 12952 9920
rect 12900 9877 12909 9911
rect 12909 9877 12943 9911
rect 12943 9877 12952 9911
rect 12900 9868 12952 9877
rect 14372 9911 14424 9920
rect 14372 9877 14381 9911
rect 14381 9877 14415 9911
rect 14415 9877 14424 9911
rect 14372 9868 14424 9877
rect 17132 9868 17184 9920
rect 19524 10004 19576 10056
rect 20996 10047 21048 10056
rect 20996 10013 21005 10047
rect 21005 10013 21039 10047
rect 21039 10013 21048 10047
rect 20996 10004 21048 10013
rect 17592 9936 17644 9988
rect 17868 9936 17920 9988
rect 19524 9868 19576 9920
rect 21364 9911 21416 9920
rect 21364 9877 21373 9911
rect 21373 9877 21407 9911
rect 21407 9877 21416 9911
rect 21364 9868 21416 9877
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 11152 9707 11204 9716
rect 11152 9673 11161 9707
rect 11161 9673 11195 9707
rect 11195 9673 11204 9707
rect 11152 9664 11204 9673
rect 12992 9664 13044 9716
rect 13544 9664 13596 9716
rect 15476 9664 15528 9716
rect 17684 9664 17736 9716
rect 18604 9664 18656 9716
rect 8392 9596 8444 9648
rect 7656 9528 7708 9580
rect 9772 9571 9824 9580
rect 9772 9537 9781 9571
rect 9781 9537 9815 9571
rect 9815 9537 9824 9571
rect 9772 9528 9824 9537
rect 11244 9528 11296 9580
rect 12348 9596 12400 9648
rect 17408 9596 17460 9648
rect 19708 9596 19760 9648
rect 11796 9571 11848 9580
rect 11796 9537 11830 9571
rect 11830 9537 11848 9571
rect 11796 9528 11848 9537
rect 7932 9460 7984 9512
rect 9496 9435 9548 9444
rect 9496 9401 9505 9435
rect 9505 9401 9539 9435
rect 9539 9401 9548 9435
rect 9496 9392 9548 9401
rect 10784 9392 10836 9444
rect 1584 9324 1636 9376
rect 10876 9324 10928 9376
rect 13728 9460 13780 9512
rect 15016 9528 15068 9580
rect 18052 9528 18104 9580
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 13636 9392 13688 9444
rect 14464 9392 14516 9444
rect 15292 9460 15344 9512
rect 16764 9503 16816 9512
rect 16764 9469 16773 9503
rect 16773 9469 16807 9503
rect 16807 9469 16816 9503
rect 16764 9460 16816 9469
rect 16948 9503 17000 9512
rect 16948 9469 16957 9503
rect 16957 9469 16991 9503
rect 16991 9469 17000 9503
rect 16948 9460 17000 9469
rect 17040 9460 17092 9512
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 18880 9392 18932 9444
rect 14648 9324 14700 9376
rect 17776 9324 17828 9376
rect 20904 9324 20956 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 7104 9120 7156 9172
rect 10784 9120 10836 9172
rect 10876 9120 10928 9172
rect 13544 9120 13596 9172
rect 13728 9163 13780 9172
rect 13728 9129 13737 9163
rect 13737 9129 13771 9163
rect 13771 9129 13780 9163
rect 13728 9120 13780 9129
rect 11980 9052 12032 9104
rect 7656 9027 7708 9036
rect 7656 8993 7665 9027
rect 7665 8993 7699 9027
rect 7699 8993 7708 9027
rect 7656 8984 7708 8993
rect 11152 9027 11204 9036
rect 11152 8993 11161 9027
rect 11161 8993 11195 9027
rect 11195 8993 11204 9027
rect 11152 8984 11204 8993
rect 7932 8959 7984 8968
rect 7932 8925 7941 8959
rect 7941 8925 7975 8959
rect 7975 8925 7984 8959
rect 7932 8916 7984 8925
rect 9496 8916 9548 8968
rect 4620 8780 4672 8832
rect 12072 8916 12124 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 12440 8916 12492 8968
rect 12900 8916 12952 8968
rect 19800 9120 19852 9172
rect 20812 9120 20864 9172
rect 16764 8984 16816 9036
rect 19524 9052 19576 9104
rect 9956 8848 10008 8900
rect 16396 8916 16448 8968
rect 14648 8848 14700 8900
rect 16212 8848 16264 8900
rect 10508 8780 10560 8832
rect 11152 8780 11204 8832
rect 11704 8823 11756 8832
rect 11704 8789 11713 8823
rect 11713 8789 11747 8823
rect 11747 8789 11756 8823
rect 11704 8780 11756 8789
rect 12900 8780 12952 8832
rect 13544 8780 13596 8832
rect 15292 8780 15344 8832
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 15660 8780 15712 8832
rect 18880 8984 18932 9036
rect 20720 8984 20772 9036
rect 17868 8916 17920 8968
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 20076 8916 20128 8968
rect 21732 8916 21784 8968
rect 18604 8848 18656 8900
rect 19892 8848 19944 8900
rect 17224 8780 17276 8832
rect 20076 8780 20128 8832
rect 20260 8780 20312 8832
rect 21180 8823 21232 8832
rect 21180 8789 21189 8823
rect 21189 8789 21223 8823
rect 21223 8789 21232 8823
rect 21180 8780 21232 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 7932 8576 7984 8628
rect 11152 8619 11204 8628
rect 4160 8508 4212 8560
rect 10692 8508 10744 8560
rect 11152 8585 11161 8619
rect 11161 8585 11195 8619
rect 11195 8585 11204 8619
rect 11152 8576 11204 8585
rect 11244 8576 11296 8628
rect 12440 8576 12492 8628
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 14372 8576 14424 8628
rect 16948 8576 17000 8628
rect 18236 8576 18288 8628
rect 19616 8576 19668 8628
rect 19708 8576 19760 8628
rect 20260 8576 20312 8628
rect 7288 8440 7340 8492
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 9772 8440 9824 8492
rect 9956 8483 10008 8492
rect 9956 8449 9965 8483
rect 9965 8449 9999 8483
rect 9999 8449 10008 8483
rect 9956 8440 10008 8449
rect 15936 8508 15988 8560
rect 16396 8508 16448 8560
rect 15292 8440 15344 8492
rect 17868 8508 17920 8560
rect 17960 8508 18012 8560
rect 21088 8551 21140 8560
rect 21088 8517 21106 8551
rect 21106 8517 21140 8551
rect 21088 8508 21140 8517
rect 18512 8440 18564 8492
rect 18972 8440 19024 8492
rect 19524 8440 19576 8492
rect 10508 8415 10560 8424
rect 10508 8381 10517 8415
rect 10517 8381 10551 8415
rect 10551 8381 10560 8415
rect 10508 8372 10560 8381
rect 10784 8372 10836 8424
rect 12532 8372 12584 8424
rect 12992 8415 13044 8424
rect 12992 8381 13001 8415
rect 13001 8381 13035 8415
rect 13035 8381 13044 8415
rect 12992 8372 13044 8381
rect 13728 8372 13780 8424
rect 15476 8415 15528 8424
rect 15476 8381 15485 8415
rect 15485 8381 15519 8415
rect 15519 8381 15528 8415
rect 15476 8372 15528 8381
rect 11152 8304 11204 8356
rect 15660 8304 15712 8356
rect 10140 8279 10192 8288
rect 10140 8245 10149 8279
rect 10149 8245 10183 8279
rect 10183 8245 10192 8279
rect 10140 8236 10192 8245
rect 17960 8372 18012 8424
rect 18880 8415 18932 8424
rect 18880 8381 18889 8415
rect 18889 8381 18923 8415
rect 18923 8381 18932 8415
rect 18880 8372 18932 8381
rect 17684 8304 17736 8356
rect 17040 8236 17092 8288
rect 20720 8236 20772 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 10508 8032 10560 8084
rect 12348 8032 12400 8084
rect 13084 8075 13136 8084
rect 13084 8041 13093 8075
rect 13093 8041 13127 8075
rect 13127 8041 13136 8075
rect 13084 8032 13136 8041
rect 17868 8075 17920 8084
rect 17868 8041 17877 8075
rect 17877 8041 17911 8075
rect 17911 8041 17920 8075
rect 17868 8032 17920 8041
rect 8300 7964 8352 8016
rect 13636 7964 13688 8016
rect 18144 8032 18196 8084
rect 7472 7871 7524 7880
rect 7472 7837 7481 7871
rect 7481 7837 7515 7871
rect 7515 7837 7524 7871
rect 7472 7828 7524 7837
rect 10600 7896 10652 7948
rect 18052 7964 18104 8016
rect 8760 7828 8812 7880
rect 6920 7803 6972 7812
rect 6920 7769 6929 7803
rect 6929 7769 6963 7803
rect 6963 7769 6972 7803
rect 6920 7760 6972 7769
rect 8944 7760 8996 7812
rect 9496 7760 9548 7812
rect 7840 7692 7892 7744
rect 8484 7692 8536 7744
rect 9128 7735 9180 7744
rect 9128 7701 9137 7735
rect 9137 7701 9171 7735
rect 9171 7701 9180 7735
rect 9128 7692 9180 7701
rect 10784 7828 10836 7880
rect 15568 7896 15620 7948
rect 20260 7939 20312 7948
rect 20260 7905 20269 7939
rect 20269 7905 20303 7939
rect 20303 7905 20312 7939
rect 20260 7896 20312 7905
rect 12900 7828 12952 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 18052 7828 18104 7880
rect 19064 7828 19116 7880
rect 20720 7871 20772 7880
rect 20720 7837 20729 7871
rect 20729 7837 20763 7871
rect 20763 7837 20772 7871
rect 20720 7828 20772 7837
rect 10968 7760 11020 7812
rect 12164 7803 12216 7812
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 11244 7692 11296 7744
rect 12164 7769 12173 7803
rect 12173 7769 12207 7803
rect 12207 7769 12216 7803
rect 12164 7760 12216 7769
rect 15660 7760 15712 7812
rect 12992 7692 13044 7744
rect 15844 7692 15896 7744
rect 21548 7760 21600 7812
rect 20536 7692 20588 7744
rect 21364 7735 21416 7744
rect 21364 7701 21373 7735
rect 21373 7701 21407 7735
rect 21407 7701 21416 7735
rect 21364 7692 21416 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 7932 7488 7984 7540
rect 8300 7463 8352 7472
rect 5540 7352 5592 7404
rect 8300 7429 8309 7463
rect 8309 7429 8343 7463
rect 8343 7429 8352 7463
rect 8300 7420 8352 7429
rect 9220 7488 9272 7540
rect 9772 7488 9824 7540
rect 10600 7531 10652 7540
rect 10600 7497 10609 7531
rect 10609 7497 10643 7531
rect 10643 7497 10652 7531
rect 10600 7488 10652 7497
rect 11152 7531 11204 7540
rect 11152 7497 11161 7531
rect 11161 7497 11195 7531
rect 11195 7497 11204 7531
rect 11152 7488 11204 7497
rect 13728 7488 13780 7540
rect 16212 7531 16264 7540
rect 16212 7497 16221 7531
rect 16221 7497 16255 7531
rect 16255 7497 16264 7531
rect 16212 7488 16264 7497
rect 18880 7488 18932 7540
rect 19892 7488 19944 7540
rect 20076 7488 20128 7540
rect 20536 7531 20588 7540
rect 20536 7497 20545 7531
rect 20545 7497 20579 7531
rect 20579 7497 20588 7531
rect 20536 7488 20588 7497
rect 20904 7531 20956 7540
rect 20904 7497 20913 7531
rect 20913 7497 20947 7531
rect 20947 7497 20956 7531
rect 20904 7488 20956 7497
rect 8760 7352 8812 7404
rect 10048 7352 10100 7404
rect 10968 7395 11020 7404
rect 10968 7361 10977 7395
rect 10977 7361 11011 7395
rect 11011 7361 11020 7395
rect 10968 7352 11020 7361
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12348 7420 12400 7472
rect 13084 7352 13136 7404
rect 15476 7352 15528 7404
rect 21364 7420 21416 7472
rect 18236 7352 18288 7404
rect 18604 7395 18656 7404
rect 18604 7361 18613 7395
rect 18613 7361 18647 7395
rect 18647 7361 18656 7395
rect 18604 7352 18656 7361
rect 20076 7352 20128 7404
rect 20996 7395 21048 7404
rect 20996 7361 21005 7395
rect 21005 7361 21039 7395
rect 21039 7361 21048 7395
rect 20996 7352 21048 7361
rect 7656 7284 7708 7336
rect 9036 7284 9088 7336
rect 16948 7327 17000 7336
rect 16948 7293 16957 7327
rect 16957 7293 16991 7327
rect 16991 7293 17000 7327
rect 16948 7284 17000 7293
rect 18512 7284 18564 7336
rect 8024 7259 8076 7268
rect 8024 7225 8033 7259
rect 8033 7225 8067 7259
rect 8067 7225 8076 7259
rect 8024 7216 8076 7225
rect 20812 7284 20864 7336
rect 9496 7148 9548 7200
rect 10784 7148 10836 7200
rect 11612 7148 11664 7200
rect 11796 7191 11848 7200
rect 11796 7157 11805 7191
rect 11805 7157 11839 7191
rect 11839 7157 11848 7191
rect 11796 7148 11848 7157
rect 11980 7148 12032 7200
rect 15200 7148 15252 7200
rect 21272 7216 21324 7268
rect 18512 7148 18564 7200
rect 19800 7148 19852 7200
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 5172 6944 5224 6996
rect 10876 6944 10928 6996
rect 11612 6944 11664 6996
rect 3148 6876 3200 6928
rect 7012 6876 7064 6928
rect 7932 6919 7984 6928
rect 7932 6885 7941 6919
rect 7941 6885 7975 6919
rect 7975 6885 7984 6919
rect 7932 6876 7984 6885
rect 6920 6740 6972 6792
rect 9036 6851 9088 6860
rect 9036 6817 9045 6851
rect 9045 6817 9079 6851
rect 9079 6817 9088 6851
rect 9036 6808 9088 6817
rect 9864 6876 9916 6928
rect 12900 6944 12952 6996
rect 18788 6944 18840 6996
rect 9772 6808 9824 6860
rect 10508 6851 10560 6860
rect 10508 6817 10517 6851
rect 10517 6817 10551 6851
rect 10551 6817 10560 6851
rect 10508 6808 10560 6817
rect 16396 6876 16448 6928
rect 12440 6808 12492 6860
rect 16028 6808 16080 6860
rect 9128 6740 9180 6792
rect 11796 6740 11848 6792
rect 12532 6783 12584 6792
rect 12532 6749 12541 6783
rect 12541 6749 12575 6783
rect 12575 6749 12584 6783
rect 12532 6740 12584 6749
rect 13452 6783 13504 6792
rect 13452 6749 13461 6783
rect 13461 6749 13495 6783
rect 13495 6749 13504 6783
rect 13452 6740 13504 6749
rect 15200 6740 15252 6792
rect 15568 6783 15620 6792
rect 15568 6749 15577 6783
rect 15577 6749 15611 6783
rect 15611 6749 15620 6783
rect 15568 6740 15620 6749
rect 15752 6740 15804 6792
rect 17684 6808 17736 6860
rect 18236 6851 18288 6860
rect 18236 6817 18245 6851
rect 18245 6817 18279 6851
rect 18279 6817 18288 6851
rect 18236 6808 18288 6817
rect 17500 6740 17552 6792
rect 18880 6783 18932 6792
rect 18880 6749 18889 6783
rect 18889 6749 18923 6783
rect 18923 6749 18932 6783
rect 18880 6740 18932 6749
rect 6276 6715 6328 6724
rect 6276 6681 6285 6715
rect 6285 6681 6319 6715
rect 6319 6681 6328 6715
rect 6276 6672 6328 6681
rect 8484 6672 8536 6724
rect 11244 6672 11296 6724
rect 6828 6604 6880 6656
rect 7196 6647 7248 6656
rect 7196 6613 7205 6647
rect 7205 6613 7239 6647
rect 7239 6613 7248 6647
rect 7196 6604 7248 6613
rect 7472 6604 7524 6656
rect 9220 6647 9272 6656
rect 9220 6613 9229 6647
rect 9229 6613 9263 6647
rect 9263 6613 9272 6647
rect 9220 6604 9272 6613
rect 10232 6647 10284 6656
rect 10232 6613 10241 6647
rect 10241 6613 10275 6647
rect 10275 6613 10284 6647
rect 10232 6604 10284 6613
rect 11060 6604 11112 6656
rect 15844 6672 15896 6724
rect 13820 6604 13872 6656
rect 15476 6647 15528 6656
rect 15476 6613 15485 6647
rect 15485 6613 15519 6647
rect 15519 6613 15528 6647
rect 15476 6604 15528 6613
rect 15568 6604 15620 6656
rect 15752 6604 15804 6656
rect 17040 6672 17092 6724
rect 19340 6740 19392 6792
rect 20536 6740 20588 6792
rect 20168 6672 20220 6724
rect 16304 6604 16356 6656
rect 17408 6604 17460 6656
rect 17592 6604 17644 6656
rect 17960 6647 18012 6656
rect 17960 6613 17969 6647
rect 17969 6613 18003 6647
rect 18003 6613 18012 6647
rect 17960 6604 18012 6613
rect 18328 6604 18380 6656
rect 21272 6604 21324 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 6644 6400 6696 6452
rect 9036 6400 9088 6452
rect 12256 6400 12308 6452
rect 13452 6400 13504 6452
rect 14740 6400 14792 6452
rect 14832 6400 14884 6452
rect 6552 6264 6604 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7932 6307 7984 6316
rect 7932 6273 7941 6307
rect 7941 6273 7975 6307
rect 7975 6273 7984 6307
rect 7932 6264 7984 6273
rect 5080 6196 5132 6248
rect 8116 6196 8168 6248
rect 9404 6264 9456 6316
rect 10508 6307 10560 6316
rect 10508 6273 10517 6307
rect 10517 6273 10551 6307
rect 10551 6273 10560 6307
rect 10508 6264 10560 6273
rect 11152 6264 11204 6316
rect 13636 6332 13688 6384
rect 13452 6307 13504 6316
rect 11980 6239 12032 6248
rect 4896 6128 4948 6180
rect 7012 6171 7064 6180
rect 6000 6103 6052 6112
rect 6000 6069 6009 6103
rect 6009 6069 6043 6103
rect 6043 6069 6052 6103
rect 6000 6060 6052 6069
rect 6552 6103 6604 6112
rect 6552 6069 6561 6103
rect 6561 6069 6595 6103
rect 6595 6069 6604 6103
rect 6552 6060 6604 6069
rect 7012 6137 7021 6171
rect 7021 6137 7055 6171
rect 7055 6137 7064 6171
rect 7012 6128 7064 6137
rect 10876 6060 10928 6112
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 11980 6196 12032 6205
rect 13452 6273 13461 6307
rect 13461 6273 13495 6307
rect 13495 6273 13504 6307
rect 13452 6264 13504 6273
rect 13176 6239 13228 6248
rect 11612 6128 11664 6180
rect 13176 6205 13185 6239
rect 13185 6205 13219 6239
rect 13219 6205 13228 6239
rect 13176 6196 13228 6205
rect 13360 6239 13412 6248
rect 13360 6205 13369 6239
rect 13369 6205 13403 6239
rect 13403 6205 13412 6239
rect 13360 6196 13412 6205
rect 12256 6128 12308 6180
rect 14924 6307 14976 6316
rect 14924 6273 14958 6307
rect 14958 6273 14976 6307
rect 14924 6264 14976 6273
rect 13636 6196 13688 6248
rect 16856 6332 16908 6384
rect 19340 6332 19392 6384
rect 20352 6400 20404 6452
rect 20628 6400 20680 6452
rect 20720 6332 20772 6384
rect 19524 6264 19576 6316
rect 14556 6060 14608 6112
rect 15752 6060 15804 6112
rect 16028 6103 16080 6112
rect 16028 6069 16037 6103
rect 16037 6069 16071 6103
rect 16071 6069 16080 6103
rect 16028 6060 16080 6069
rect 16120 6060 16172 6112
rect 21088 6307 21140 6316
rect 21088 6273 21097 6307
rect 21097 6273 21131 6307
rect 21131 6273 21140 6307
rect 21088 6264 21140 6273
rect 21180 6128 21232 6180
rect 20812 6103 20864 6112
rect 20812 6069 20821 6103
rect 20821 6069 20855 6103
rect 20855 6069 20864 6103
rect 20812 6060 20864 6069
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 4528 5856 4580 5908
rect 4988 5856 5040 5908
rect 5632 5899 5684 5908
rect 5632 5865 5641 5899
rect 5641 5865 5675 5899
rect 5675 5865 5684 5899
rect 5632 5856 5684 5865
rect 7840 5856 7892 5908
rect 7932 5856 7984 5908
rect 2504 5788 2556 5840
rect 5908 5720 5960 5772
rect 9220 5856 9272 5908
rect 8760 5788 8812 5840
rect 12256 5856 12308 5908
rect 13084 5899 13136 5908
rect 13084 5865 13093 5899
rect 13093 5865 13127 5899
rect 13127 5865 13136 5899
rect 13084 5856 13136 5865
rect 13452 5856 13504 5908
rect 17040 5856 17092 5908
rect 17408 5856 17460 5908
rect 17776 5856 17828 5908
rect 6920 5695 6972 5704
rect 6920 5661 6929 5695
rect 6929 5661 6963 5695
rect 6963 5661 6972 5695
rect 6920 5652 6972 5661
rect 7196 5695 7248 5704
rect 7196 5661 7205 5695
rect 7205 5661 7239 5695
rect 7239 5661 7248 5695
rect 7196 5652 7248 5661
rect 18880 5788 18932 5840
rect 20996 5856 21048 5908
rect 21640 5856 21692 5908
rect 22652 5788 22704 5840
rect 1860 5516 1912 5568
rect 4620 5516 4672 5568
rect 4804 5559 4856 5568
rect 4804 5525 4813 5559
rect 4813 5525 4847 5559
rect 4847 5525 4856 5559
rect 4804 5516 4856 5525
rect 7840 5652 7892 5704
rect 14556 5720 14608 5772
rect 15200 5720 15252 5772
rect 16028 5720 16080 5772
rect 9680 5652 9732 5704
rect 10508 5652 10560 5704
rect 11612 5652 11664 5704
rect 12164 5695 12216 5704
rect 12164 5661 12173 5695
rect 12173 5661 12207 5695
rect 12207 5661 12216 5695
rect 12164 5652 12216 5661
rect 12440 5695 12492 5704
rect 12440 5661 12449 5695
rect 12449 5661 12483 5695
rect 12483 5661 12492 5695
rect 12440 5652 12492 5661
rect 12624 5652 12676 5704
rect 15108 5695 15160 5704
rect 15108 5661 15117 5695
rect 15117 5661 15151 5695
rect 15151 5661 15160 5695
rect 15108 5652 15160 5661
rect 15660 5695 15712 5704
rect 15660 5661 15669 5695
rect 15669 5661 15703 5695
rect 15703 5661 15712 5695
rect 15660 5652 15712 5661
rect 8760 5584 8812 5636
rect 9496 5584 9548 5636
rect 18144 5652 18196 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 17408 5627 17460 5636
rect 17408 5593 17417 5627
rect 17417 5593 17451 5627
rect 17451 5593 17460 5627
rect 20536 5652 20588 5704
rect 20904 5695 20956 5704
rect 20904 5661 20913 5695
rect 20913 5661 20947 5695
rect 20947 5661 20956 5695
rect 20904 5652 20956 5661
rect 17408 5584 17460 5593
rect 9588 5516 9640 5568
rect 11060 5516 11112 5568
rect 13728 5516 13780 5568
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 14464 5516 14516 5525
rect 14648 5516 14700 5568
rect 17592 5516 17644 5568
rect 17776 5516 17828 5568
rect 18144 5559 18196 5568
rect 18144 5525 18153 5559
rect 18153 5525 18187 5559
rect 18187 5525 18196 5559
rect 18696 5559 18748 5568
rect 18144 5516 18196 5525
rect 18696 5525 18705 5559
rect 18705 5525 18739 5559
rect 18739 5525 18748 5559
rect 18696 5516 18748 5525
rect 21180 5584 21232 5636
rect 21088 5559 21140 5568
rect 21088 5525 21097 5559
rect 21097 5525 21131 5559
rect 21131 5525 21140 5559
rect 21088 5516 21140 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 6644 5312 6696 5364
rect 8208 5312 8260 5364
rect 10508 5312 10560 5364
rect 12072 5312 12124 5364
rect 13176 5312 13228 5364
rect 13360 5312 13412 5364
rect 18144 5312 18196 5364
rect 6460 5287 6512 5296
rect 6460 5253 6469 5287
rect 6469 5253 6503 5287
rect 6503 5253 6512 5287
rect 6460 5244 6512 5253
rect 7196 5244 7248 5296
rect 7748 5244 7800 5296
rect 8116 5244 8168 5296
rect 5448 5176 5500 5228
rect 6736 5219 6788 5228
rect 6736 5185 6745 5219
rect 6745 5185 6779 5219
rect 6779 5185 6788 5219
rect 6736 5176 6788 5185
rect 11060 5244 11112 5296
rect 9588 5176 9640 5228
rect 12164 5176 12216 5228
rect 13820 5244 13872 5296
rect 14188 5244 14240 5296
rect 14832 5244 14884 5296
rect 16028 5287 16080 5296
rect 16028 5253 16046 5287
rect 16046 5253 16080 5287
rect 16028 5244 16080 5253
rect 13636 5219 13688 5228
rect 13636 5185 13645 5219
rect 13645 5185 13679 5219
rect 13679 5185 13688 5219
rect 13636 5176 13688 5185
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 15016 5176 15068 5228
rect 17408 5244 17460 5296
rect 18236 5244 18288 5296
rect 19892 5312 19944 5364
rect 20444 5312 20496 5364
rect 20812 5312 20864 5364
rect 11612 5108 11664 5160
rect 14556 5151 14608 5160
rect 14556 5117 14565 5151
rect 14565 5117 14599 5151
rect 14599 5117 14608 5151
rect 14556 5108 14608 5117
rect 16396 5176 16448 5228
rect 17040 5219 17092 5228
rect 17040 5185 17049 5219
rect 17049 5185 17083 5219
rect 17083 5185 17092 5219
rect 17040 5176 17092 5185
rect 17684 5219 17736 5228
rect 17684 5185 17693 5219
rect 17693 5185 17727 5219
rect 17727 5185 17736 5219
rect 17684 5176 17736 5185
rect 18604 5176 18656 5228
rect 19708 5219 19760 5228
rect 19708 5185 19717 5219
rect 19717 5185 19751 5219
rect 19751 5185 19760 5219
rect 19708 5176 19760 5185
rect 4344 5040 4396 5092
rect 1400 5015 1452 5024
rect 1400 4981 1409 5015
rect 1409 4981 1443 5015
rect 1443 4981 1452 5015
rect 1400 4972 1452 4981
rect 4252 5015 4304 5024
rect 4252 4981 4261 5015
rect 4261 4981 4295 5015
rect 4295 4981 4304 5015
rect 4252 4972 4304 4981
rect 4988 5015 5040 5024
rect 4988 4981 4997 5015
rect 4997 4981 5031 5015
rect 5031 4981 5040 5015
rect 4988 4972 5040 4981
rect 6920 4972 6972 5024
rect 7564 4972 7616 5024
rect 12440 5040 12492 5092
rect 16856 5108 16908 5160
rect 17776 5040 17828 5092
rect 19524 5151 19576 5160
rect 19524 5117 19533 5151
rect 19533 5117 19567 5151
rect 19567 5117 19576 5151
rect 19524 5108 19576 5117
rect 20260 5108 20312 5160
rect 20536 5108 20588 5160
rect 20996 5151 21048 5160
rect 20996 5117 21005 5151
rect 21005 5117 21039 5151
rect 21039 5117 21048 5151
rect 20996 5108 21048 5117
rect 9864 4972 9916 5024
rect 10048 4972 10100 5024
rect 15568 4972 15620 5024
rect 16948 4972 17000 5024
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 5540 4768 5592 4820
rect 8576 4811 8628 4820
rect 4436 4700 4488 4752
rect 8300 4700 8352 4752
rect 8576 4777 8585 4811
rect 8585 4777 8619 4811
rect 8619 4777 8628 4811
rect 8576 4768 8628 4777
rect 9404 4768 9456 4820
rect 11152 4768 11204 4820
rect 11612 4768 11664 4820
rect 15476 4768 15528 4820
rect 2964 4632 3016 4684
rect 5356 4564 5408 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 6552 4607 6604 4616
rect 5448 4564 5500 4573
rect 6552 4573 6561 4607
rect 6561 4573 6595 4607
rect 6595 4573 6604 4607
rect 6552 4564 6604 4573
rect 1676 4496 1728 4548
rect 5816 4496 5868 4548
rect 7104 4539 7156 4548
rect 7104 4505 7113 4539
rect 7113 4505 7147 4539
rect 7147 4505 7156 4539
rect 7104 4496 7156 4505
rect 7564 4632 7616 4684
rect 7656 4564 7708 4616
rect 8392 4564 8444 4616
rect 9128 4564 9180 4616
rect 9404 4564 9456 4616
rect 10876 4607 10928 4616
rect 10876 4573 10894 4607
rect 10894 4573 10928 4607
rect 10876 4564 10928 4573
rect 11060 4564 11112 4616
rect 12072 4607 12124 4616
rect 12072 4573 12081 4607
rect 12081 4573 12115 4607
rect 12115 4573 12124 4607
rect 12072 4564 12124 4573
rect 14924 4632 14976 4684
rect 13636 4564 13688 4616
rect 9588 4496 9640 4548
rect 1768 4471 1820 4480
rect 1768 4437 1777 4471
rect 1777 4437 1811 4471
rect 1811 4437 1820 4471
rect 1768 4428 1820 4437
rect 2320 4428 2372 4480
rect 3056 4471 3108 4480
rect 3056 4437 3065 4471
rect 3065 4437 3099 4471
rect 3099 4437 3108 4471
rect 3056 4428 3108 4437
rect 3424 4471 3476 4480
rect 3424 4437 3433 4471
rect 3433 4437 3467 4471
rect 3467 4437 3476 4471
rect 3424 4428 3476 4437
rect 7012 4428 7064 4480
rect 8300 4428 8352 4480
rect 12440 4428 12492 4480
rect 13360 4496 13412 4548
rect 12992 4428 13044 4480
rect 16396 4564 16448 4616
rect 17132 4700 17184 4752
rect 18420 4768 18472 4820
rect 20536 4811 20588 4820
rect 20536 4777 20545 4811
rect 20545 4777 20579 4811
rect 20579 4777 20588 4811
rect 20536 4768 20588 4777
rect 18972 4700 19024 4752
rect 17224 4675 17276 4684
rect 17224 4641 17233 4675
rect 17233 4641 17267 4675
rect 17267 4641 17276 4675
rect 17224 4632 17276 4641
rect 18236 4675 18288 4684
rect 18236 4641 18245 4675
rect 18245 4641 18279 4675
rect 18279 4641 18288 4675
rect 18236 4632 18288 4641
rect 19524 4632 19576 4684
rect 20076 4632 20128 4684
rect 21180 4675 21232 4684
rect 21180 4641 21189 4675
rect 21189 4641 21223 4675
rect 21223 4641 21232 4675
rect 21180 4632 21232 4641
rect 14280 4428 14332 4480
rect 15384 4471 15436 4480
rect 15384 4437 15393 4471
rect 15393 4437 15427 4471
rect 15427 4437 15436 4471
rect 15384 4428 15436 4437
rect 19800 4564 19852 4616
rect 18880 4496 18932 4548
rect 17132 4428 17184 4480
rect 17500 4471 17552 4480
rect 17500 4437 17509 4471
rect 17509 4437 17543 4471
rect 17543 4437 17552 4471
rect 17500 4428 17552 4437
rect 18236 4428 18288 4480
rect 18512 4471 18564 4480
rect 18512 4437 18521 4471
rect 18521 4437 18555 4471
rect 18555 4437 18564 4471
rect 18512 4428 18564 4437
rect 19616 4428 19668 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 14464 4224 14516 4276
rect 12072 4156 12124 4208
rect 13268 4199 13320 4208
rect 13268 4165 13277 4199
rect 13277 4165 13311 4199
rect 13311 4165 13320 4199
rect 13268 4156 13320 4165
rect 13360 4156 13412 4208
rect 17684 4224 17736 4276
rect 18144 4224 18196 4276
rect 18604 4224 18656 4276
rect 20168 4224 20220 4276
rect 20444 4224 20496 4276
rect 15568 4199 15620 4208
rect 15568 4165 15577 4199
rect 15577 4165 15611 4199
rect 15611 4165 15620 4199
rect 15568 4156 15620 4165
rect 16212 4156 16264 4208
rect 16488 4156 16540 4208
rect 17408 4156 17460 4208
rect 4436 4131 4488 4140
rect 4436 4097 4445 4131
rect 4445 4097 4479 4131
rect 4479 4097 4488 4131
rect 4436 4088 4488 4097
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 4068 4020 4120 4072
rect 7288 4088 7340 4140
rect 7564 4020 7616 4072
rect 2872 3952 2924 4004
rect 4896 3952 4948 4004
rect 4988 3952 5040 4004
rect 5540 3995 5592 4004
rect 1308 3884 1360 3936
rect 1952 3927 2004 3936
rect 1952 3893 1961 3927
rect 1961 3893 1995 3927
rect 1995 3893 2004 3927
rect 1952 3884 2004 3893
rect 3240 3884 3292 3936
rect 3976 3884 4028 3936
rect 4620 3927 4672 3936
rect 4620 3893 4629 3927
rect 4629 3893 4663 3927
rect 4663 3893 4672 3927
rect 4620 3884 4672 3893
rect 5080 3927 5132 3936
rect 5080 3893 5089 3927
rect 5089 3893 5123 3927
rect 5123 3893 5132 3927
rect 5080 3884 5132 3893
rect 5540 3961 5549 3995
rect 5549 3961 5583 3995
rect 5583 3961 5592 3995
rect 5540 3952 5592 3961
rect 7288 3884 7340 3936
rect 7840 4088 7892 4140
rect 9864 4131 9916 4140
rect 9864 4097 9873 4131
rect 9873 4097 9907 4131
rect 9907 4097 9916 4131
rect 9864 4088 9916 4097
rect 10876 4088 10928 4140
rect 12532 4088 12584 4140
rect 7748 4020 7800 4072
rect 11060 4020 11112 4072
rect 11428 3952 11480 4004
rect 12992 4020 13044 4072
rect 13452 4088 13504 4140
rect 15108 4088 15160 4140
rect 13728 4020 13780 4072
rect 14832 4020 14884 4072
rect 15752 4088 15804 4140
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 16764 4088 16816 4140
rect 17224 4088 17276 4140
rect 18420 4156 18472 4208
rect 21272 4156 21324 4208
rect 18972 4088 19024 4140
rect 13544 3952 13596 4004
rect 14740 3952 14792 4004
rect 16212 4020 16264 4072
rect 20536 4088 20588 4140
rect 9496 3884 9548 3936
rect 10968 3884 11020 3936
rect 11888 3884 11940 3936
rect 11980 3884 12032 3936
rect 12900 3884 12952 3936
rect 13176 3884 13228 3936
rect 15476 3884 15528 3936
rect 17408 3884 17460 3936
rect 17868 3884 17920 3936
rect 18788 3884 18840 3936
rect 19524 3884 19576 3936
rect 19892 3884 19944 3936
rect 21456 3884 21508 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 5540 3680 5592 3732
rect 5724 3723 5776 3732
rect 5724 3689 5733 3723
rect 5733 3689 5767 3723
rect 5767 3689 5776 3723
rect 5724 3680 5776 3689
rect 6828 3680 6880 3732
rect 3976 3612 4028 3664
rect 5080 3612 5132 3664
rect 8392 3612 8444 3664
rect 9128 3680 9180 3732
rect 9588 3680 9640 3732
rect 11428 3723 11480 3732
rect 10048 3612 10100 3664
rect 11428 3689 11437 3723
rect 11437 3689 11471 3723
rect 11471 3689 11480 3723
rect 11428 3680 11480 3689
rect 14464 3680 14516 3732
rect 14740 3680 14792 3732
rect 16212 3723 16264 3732
rect 16212 3689 16221 3723
rect 16221 3689 16255 3723
rect 16255 3689 16264 3723
rect 16212 3680 16264 3689
rect 16304 3680 16356 3732
rect 16948 3680 17000 3732
rect 17132 3680 17184 3732
rect 20628 3680 20680 3732
rect 12716 3612 12768 3664
rect 14372 3612 14424 3664
rect 16028 3612 16080 3664
rect 5356 3544 5408 3596
rect 7932 3587 7984 3596
rect 7932 3553 7941 3587
rect 7941 3553 7975 3587
rect 7975 3553 7984 3587
rect 7932 3544 7984 3553
rect 9496 3587 9548 3596
rect 664 3476 716 3528
rect 1308 3476 1360 3528
rect 3332 3476 3384 3528
rect 4252 3476 4304 3528
rect 4436 3476 4488 3528
rect 4988 3476 5040 3528
rect 5080 3519 5132 3528
rect 5080 3485 5089 3519
rect 5089 3485 5123 3519
rect 5123 3485 5132 3519
rect 5080 3476 5132 3485
rect 5540 3519 5592 3528
rect 5540 3485 5549 3519
rect 5549 3485 5583 3519
rect 5583 3485 5592 3519
rect 5540 3476 5592 3485
rect 5724 3476 5776 3528
rect 6920 3476 6972 3528
rect 7656 3476 7708 3528
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 4712 3408 4764 3460
rect 2136 3340 2188 3392
rect 2596 3340 2648 3392
rect 4620 3340 4672 3392
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 6000 3340 6052 3392
rect 6644 3383 6696 3392
rect 6644 3349 6653 3383
rect 6653 3349 6687 3383
rect 6687 3349 6696 3383
rect 6644 3340 6696 3349
rect 6736 3340 6788 3392
rect 9496 3553 9505 3587
rect 9505 3553 9539 3587
rect 9539 3553 9548 3587
rect 9496 3544 9548 3553
rect 16672 3544 16724 3596
rect 17224 3544 17276 3596
rect 17868 3587 17920 3596
rect 17868 3553 17877 3587
rect 17877 3553 17911 3587
rect 17911 3553 17920 3587
rect 17868 3544 17920 3553
rect 20444 3544 20496 3596
rect 11152 3476 11204 3528
rect 11796 3519 11848 3528
rect 11796 3485 11805 3519
rect 11805 3485 11839 3519
rect 11839 3485 11848 3519
rect 11796 3476 11848 3485
rect 13636 3476 13688 3528
rect 15200 3476 15252 3528
rect 8392 3408 8444 3460
rect 10968 3408 11020 3460
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9588 3340 9640 3392
rect 12440 3340 12492 3392
rect 15660 3451 15712 3460
rect 15660 3417 15700 3451
rect 15700 3417 15712 3451
rect 15660 3408 15712 3417
rect 16028 3408 16080 3460
rect 16120 3408 16172 3460
rect 13912 3340 13964 3392
rect 15476 3340 15528 3392
rect 16304 3340 16356 3392
rect 17408 3476 17460 3528
rect 19524 3476 19576 3528
rect 19708 3519 19760 3528
rect 19708 3485 19717 3519
rect 19717 3485 19751 3519
rect 19751 3485 19760 3519
rect 19708 3476 19760 3485
rect 20352 3476 20404 3528
rect 20628 3476 20680 3528
rect 17500 3340 17552 3392
rect 18052 3340 18104 3392
rect 20536 3340 20588 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 1860 3136 1912 3188
rect 2044 3179 2096 3188
rect 2044 3145 2053 3179
rect 2053 3145 2087 3179
rect 2087 3145 2096 3179
rect 2044 3136 2096 3145
rect 2504 3179 2556 3188
rect 2504 3145 2513 3179
rect 2513 3145 2547 3179
rect 2547 3145 2556 3179
rect 2504 3136 2556 3145
rect 2964 3179 3016 3188
rect 2964 3145 2973 3179
rect 2973 3145 3007 3179
rect 3007 3145 3016 3179
rect 2964 3136 3016 3145
rect 3240 3136 3292 3188
rect 4436 3136 4488 3188
rect 6736 3136 6788 3188
rect 7840 3136 7892 3188
rect 8024 3136 8076 3188
rect 10508 3136 10560 3188
rect 1216 3000 1268 3052
rect 1676 3000 1728 3052
rect 1768 3000 1820 3052
rect 2320 3043 2372 3052
rect 2320 3009 2329 3043
rect 2329 3009 2363 3043
rect 2363 3009 2372 3043
rect 2320 3000 2372 3009
rect 2872 3000 2924 3052
rect 3424 3000 3476 3052
rect 4252 3000 4304 3052
rect 5632 3068 5684 3120
rect 7656 3068 7708 3120
rect 8208 3068 8260 3120
rect 4896 3043 4948 3052
rect 4528 2932 4580 2984
rect 3700 2907 3752 2916
rect 3700 2873 3709 2907
rect 3709 2873 3743 2907
rect 3743 2873 3752 2907
rect 3700 2864 3752 2873
rect 4160 2907 4212 2916
rect 4160 2873 4169 2907
rect 4169 2873 4203 2907
rect 4203 2873 4212 2907
rect 4160 2864 4212 2873
rect 4436 2864 4488 2916
rect 4896 3009 4905 3043
rect 4905 3009 4939 3043
rect 4939 3009 4948 3043
rect 4896 3000 4948 3009
rect 5172 3000 5224 3052
rect 6828 3000 6880 3052
rect 6644 2932 6696 2984
rect 6552 2907 6604 2916
rect 4896 2796 4948 2848
rect 5448 2796 5500 2848
rect 5908 2796 5960 2848
rect 6552 2873 6561 2907
rect 6561 2873 6595 2907
rect 6595 2873 6604 2907
rect 6552 2864 6604 2873
rect 6460 2796 6512 2848
rect 7564 3000 7616 3052
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 13176 3136 13228 3188
rect 13452 3179 13504 3188
rect 13452 3145 13461 3179
rect 13461 3145 13495 3179
rect 13495 3145 13504 3179
rect 13452 3136 13504 3145
rect 13728 3179 13780 3188
rect 13728 3145 13737 3179
rect 13737 3145 13771 3179
rect 13771 3145 13780 3179
rect 13728 3136 13780 3145
rect 14740 3136 14792 3188
rect 15200 3136 15252 3188
rect 15660 3136 15712 3188
rect 16120 3136 16172 3188
rect 12440 3068 12492 3120
rect 13360 3068 13412 3120
rect 11152 3043 11204 3052
rect 7748 2975 7800 2984
rect 7748 2941 7757 2975
rect 7757 2941 7791 2975
rect 7791 2941 7800 2975
rect 7748 2932 7800 2941
rect 9496 2864 9548 2916
rect 11152 3009 11161 3043
rect 11161 3009 11195 3043
rect 11195 3009 11204 3043
rect 11152 3000 11204 3009
rect 11520 3043 11572 3052
rect 11520 3009 11529 3043
rect 11529 3009 11563 3043
rect 11563 3009 11572 3043
rect 11520 3000 11572 3009
rect 13728 3000 13780 3052
rect 14280 3068 14332 3120
rect 16304 3068 16356 3120
rect 13360 2932 13412 2984
rect 16856 3000 16908 3052
rect 17868 3068 17920 3120
rect 17960 3000 18012 3052
rect 18512 3136 18564 3188
rect 18604 3136 18656 3188
rect 19340 3136 19392 3188
rect 20076 3136 20128 3188
rect 18236 3068 18288 3120
rect 18880 3068 18932 3120
rect 19800 3000 19852 3052
rect 20536 3043 20588 3052
rect 20536 3009 20545 3043
rect 20545 3009 20579 3043
rect 20579 3009 20588 3043
rect 20536 3000 20588 3009
rect 13912 2864 13964 2916
rect 14924 2864 14976 2916
rect 16212 2864 16264 2916
rect 17500 2932 17552 2984
rect 17776 2932 17828 2984
rect 18972 2975 19024 2984
rect 18972 2941 18981 2975
rect 18981 2941 19015 2975
rect 19015 2941 19024 2975
rect 18972 2932 19024 2941
rect 19432 2975 19484 2984
rect 19432 2941 19441 2975
rect 19441 2941 19475 2975
rect 19475 2941 19484 2975
rect 19432 2932 19484 2941
rect 11520 2796 11572 2848
rect 11704 2839 11756 2848
rect 11704 2805 11713 2839
rect 11713 2805 11747 2839
rect 11747 2805 11756 2839
rect 11704 2796 11756 2805
rect 13360 2796 13412 2848
rect 18144 2864 18196 2916
rect 21088 2864 21140 2916
rect 20260 2796 20312 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 3240 2592 3292 2644
rect 6736 2592 6788 2644
rect 7104 2592 7156 2644
rect 7196 2635 7248 2644
rect 7196 2601 7205 2635
rect 7205 2601 7239 2635
rect 7239 2601 7248 2635
rect 7196 2592 7248 2601
rect 7932 2592 7984 2644
rect 8668 2592 8720 2644
rect 11060 2592 11112 2644
rect 1952 2388 2004 2440
rect 3332 2524 3384 2576
rect 7564 2524 7616 2576
rect 12532 2592 12584 2644
rect 13268 2592 13320 2644
rect 15568 2592 15620 2644
rect 15752 2592 15804 2644
rect 17500 2592 17552 2644
rect 19708 2592 19760 2644
rect 12164 2524 12216 2576
rect 3056 2456 3108 2508
rect 3884 2456 3936 2508
rect 3240 2431 3292 2440
rect 3240 2397 3249 2431
rect 3249 2397 3283 2431
rect 3283 2397 3292 2431
rect 3240 2388 3292 2397
rect 4068 2388 4120 2440
rect 4620 2388 4672 2440
rect 4896 2431 4948 2440
rect 4896 2397 4905 2431
rect 4905 2397 4939 2431
rect 4939 2397 4948 2431
rect 4896 2388 4948 2397
rect 5080 2388 5132 2440
rect 7196 2456 7248 2508
rect 9496 2499 9548 2508
rect 9496 2465 9505 2499
rect 9505 2465 9539 2499
rect 9539 2465 9548 2499
rect 9496 2456 9548 2465
rect 10508 2499 10560 2508
rect 10508 2465 10517 2499
rect 10517 2465 10551 2499
rect 10551 2465 10560 2499
rect 10508 2456 10560 2465
rect 10784 2456 10836 2508
rect 10876 2456 10928 2508
rect 204 2320 256 2372
rect 1400 2320 1452 2372
rect 2412 2252 2464 2304
rect 5540 2320 5592 2372
rect 6736 2431 6788 2440
rect 6736 2397 6745 2431
rect 6745 2397 6779 2431
rect 6779 2397 6788 2431
rect 6736 2388 6788 2397
rect 7748 2388 7800 2440
rect 8668 2388 8720 2440
rect 10140 2388 10192 2440
rect 11244 2388 11296 2440
rect 7840 2320 7892 2372
rect 12440 2456 12492 2508
rect 12808 2388 12860 2440
rect 15200 2456 15252 2508
rect 16396 2524 16448 2576
rect 17776 2524 17828 2576
rect 17316 2456 17368 2508
rect 17500 2499 17552 2508
rect 17500 2465 17509 2499
rect 17509 2465 17543 2499
rect 17543 2465 17552 2499
rect 17500 2456 17552 2465
rect 18420 2456 18472 2508
rect 19616 2456 19668 2508
rect 20260 2456 20312 2508
rect 14464 2388 14516 2440
rect 15936 2431 15988 2440
rect 15936 2397 15945 2431
rect 15945 2397 15979 2431
rect 15979 2397 15988 2431
rect 15936 2388 15988 2397
rect 18880 2431 18932 2440
rect 18880 2397 18889 2431
rect 18889 2397 18923 2431
rect 18923 2397 18932 2431
rect 18880 2388 18932 2397
rect 19432 2431 19484 2440
rect 19432 2397 19441 2431
rect 19441 2397 19475 2431
rect 19475 2397 19484 2431
rect 19432 2388 19484 2397
rect 20536 2431 20588 2440
rect 20536 2397 20545 2431
rect 20545 2397 20579 2431
rect 20579 2397 20588 2431
rect 20536 2388 20588 2397
rect 2964 2295 3016 2304
rect 2964 2261 2973 2295
rect 2973 2261 3007 2295
rect 3007 2261 3016 2295
rect 2964 2252 3016 2261
rect 4160 2295 4212 2304
rect 4160 2261 4169 2295
rect 4169 2261 4203 2295
rect 4203 2261 4212 2295
rect 4160 2252 4212 2261
rect 4620 2295 4672 2304
rect 4620 2261 4629 2295
rect 4629 2261 4663 2295
rect 4663 2261 4672 2295
rect 4620 2252 4672 2261
rect 5080 2295 5132 2304
rect 5080 2261 5089 2295
rect 5089 2261 5123 2295
rect 5123 2261 5132 2295
rect 5080 2252 5132 2261
rect 7656 2252 7708 2304
rect 10784 2295 10836 2304
rect 10784 2261 10793 2295
rect 10793 2261 10827 2295
rect 10827 2261 10836 2295
rect 10784 2252 10836 2261
rect 10968 2252 11020 2304
rect 12808 2295 12860 2304
rect 12808 2261 12817 2295
rect 12817 2261 12851 2295
rect 12851 2261 12860 2295
rect 14188 2295 14240 2304
rect 12808 2252 12860 2261
rect 14188 2261 14197 2295
rect 14197 2261 14231 2295
rect 14231 2261 14240 2295
rect 14188 2252 14240 2261
rect 15292 2295 15344 2304
rect 15292 2261 15301 2295
rect 15301 2261 15335 2295
rect 15335 2261 15344 2295
rect 15292 2252 15344 2261
rect 18420 2320 18472 2372
rect 17040 2252 17092 2304
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 3240 2048 3292 2100
rect 4436 2048 4488 2100
rect 4988 2048 5040 2100
rect 5356 2048 5408 2100
rect 6736 2048 6788 2100
rect 11152 2048 11204 2100
rect 14188 2048 14240 2100
rect 22100 2048 22152 2100
rect 5080 1980 5132 2032
rect 15936 1980 15988 2032
rect 2412 1912 2464 1964
rect 7196 1912 7248 1964
rect 7472 1912 7524 1964
rect 15292 1912 15344 1964
rect 4620 1844 4672 1896
rect 10968 1844 11020 1896
rect 6000 1776 6052 1828
rect 12808 1776 12860 1828
rect 19340 1776 19392 1828
rect 20076 1776 20128 1828
rect 5264 1708 5316 1760
rect 10784 1708 10836 1760
rect 4160 1640 4212 1692
rect 10692 1640 10744 1692
rect 4068 1572 4120 1624
rect 6184 1572 6236 1624
rect 7196 1572 7248 1624
rect 12900 1572 12952 1624
rect 5724 1504 5776 1556
rect 9496 1504 9548 1556
rect 19524 1368 19576 1420
rect 2596 1300 2648 1352
rect 19432 1300 19484 1352
rect 3516 1232 3568 1284
rect 16580 1096 16632 1148
rect 18144 1096 18196 1148
<< metal2 >>
rect 5722 22200 5778 23000
rect 17222 22200 17278 23000
rect 19246 22672 19302 22681
rect 19246 22607 19302 22616
rect 5736 20466 5764 22200
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 17236 20466 17264 22200
rect 19260 20534 19288 22607
rect 19614 22264 19670 22273
rect 19614 22199 19670 22208
rect 19248 20528 19300 20534
rect 19248 20470 19300 20476
rect 5724 20460 5776 20466
rect 5724 20402 5776 20408
rect 17224 20460 17276 20466
rect 17224 20402 17276 20408
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 6000 20256 6052 20262
rect 6000 20198 6052 20204
rect 17316 20256 17368 20262
rect 17316 20198 17368 20204
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 6012 19854 6040 20198
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 6000 19848 6052 19854
rect 6000 19790 6052 19796
rect 12900 19848 12952 19854
rect 12900 19790 12952 19796
rect 6552 19780 6604 19786
rect 6552 19722 6604 19728
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18448 6456 18468
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6564 17241 6592 19722
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 12912 18970 12940 19790
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 16212 19440 16264 19446
rect 16212 19382 16264 19388
rect 13945 19068 14253 19088
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 12900 18964 12952 18970
rect 12900 18906 12952 18912
rect 9772 18760 9824 18766
rect 9772 18702 9824 18708
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 8576 18284 8628 18290
rect 8576 18226 8628 18232
rect 6550 17232 6606 17241
rect 6550 17167 6606 17176
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 4986 12336 5042 12345
rect 4986 12271 5042 12280
rect 1492 11552 1544 11558
rect 1490 11520 1492 11529
rect 1544 11520 1546 11529
rect 1490 11455 1546 11464
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1308 3936 1360 3942
rect 1308 3878 1360 3884
rect 1320 3534 1348 3878
rect 664 3528 716 3534
rect 664 3470 716 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 204 2372 256 2378
rect 204 2314 256 2320
rect 216 800 244 2314
rect 676 800 704 3470
rect 1216 3052 1268 3058
rect 1216 2994 1268 3000
rect 1228 800 1256 2994
rect 1412 2378 1440 4966
rect 1596 3738 1624 9318
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3974 9072 4030 9081
rect 3974 9007 4030 9016
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 2042 7440 2098 7449
rect 2042 7375 2098 7384
rect 1860 5568 1912 5574
rect 1860 5510 1912 5516
rect 1676 4548 1728 4554
rect 1676 4490 1728 4496
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1688 3058 1716 4490
rect 1768 4480 1820 4486
rect 1768 4422 1820 4428
rect 1780 3058 1808 4422
rect 1872 3194 1900 5510
rect 1952 3936 2004 3942
rect 1952 3878 2004 3884
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1768 3052 1820 3058
rect 1768 2994 1820 3000
rect 1400 2372 1452 2378
rect 1400 2314 1452 2320
rect 1780 800 1808 2994
rect 1964 2446 1992 3878
rect 2056 3194 2084 7375
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3148 6928 3200 6934
rect 3148 6870 3200 6876
rect 2504 5840 2556 5846
rect 2504 5782 2556 5788
rect 2320 4480 2372 4486
rect 2320 4422 2372 4428
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2148 1873 2176 3334
rect 2332 3058 2360 4422
rect 2516 3194 2544 5782
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 2872 4004 2924 4010
rect 2872 3946 2924 3952
rect 2596 3392 2648 3398
rect 2596 3334 2648 3340
rect 2504 3188 2556 3194
rect 2504 3130 2556 3136
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2134 1864 2190 1873
rect 2134 1799 2190 1808
rect 2332 800 2360 2994
rect 2412 2304 2464 2310
rect 2412 2246 2464 2252
rect 2424 1970 2452 2246
rect 2412 1964 2464 1970
rect 2412 1906 2464 1912
rect 2608 1358 2636 3334
rect 2884 3058 2912 3946
rect 2976 3194 3004 4626
rect 3056 4480 3108 4486
rect 3056 4422 3108 4428
rect 2964 3188 3016 3194
rect 2964 3130 3016 3136
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2596 1352 2648 1358
rect 2596 1294 2648 1300
rect 2884 800 2912 2994
rect 3068 2514 3096 4422
rect 3160 2774 3188 6870
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3988 4826 4016 9007
rect 4620 8832 4672 8838
rect 4620 8774 4672 8780
rect 4160 8560 4212 8566
rect 4160 8502 4212 8508
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3194 3280 3878
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3160 2746 3280 2774
rect 3252 2650 3280 2746
rect 3344 2666 3372 3470
rect 3436 3058 3464 4422
rect 4068 4072 4120 4078
rect 4068 4014 4120 4020
rect 3976 3936 4028 3942
rect 3976 3878 4028 3884
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3988 3670 4016 3878
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3424 3052 3476 3058
rect 3424 2994 3476 3000
rect 3698 2952 3754 2961
rect 3698 2887 3700 2896
rect 3752 2887 3754 2896
rect 3700 2858 3752 2864
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 3240 2644 3292 2650
rect 3344 2638 3464 2666
rect 3436 2632 3464 2638
rect 3436 2604 3556 2632
rect 3240 2586 3292 2592
rect 3332 2576 3384 2582
rect 3384 2524 3464 2530
rect 3332 2518 3464 2524
rect 3056 2508 3108 2514
rect 3344 2502 3464 2518
rect 3056 2450 3108 2456
rect 3240 2440 3292 2446
rect 2962 2408 3018 2417
rect 3240 2382 3292 2388
rect 2962 2343 3018 2352
rect 2976 2310 3004 2343
rect 2964 2304 3016 2310
rect 2964 2246 3016 2252
rect 3252 2106 3280 2382
rect 3240 2100 3292 2106
rect 3240 2042 3292 2048
rect 3436 800 3464 2502
rect 3528 1290 3556 2604
rect 3884 2508 3936 2514
rect 3936 2468 4016 2496
rect 3884 2450 3936 2456
rect 3516 1284 3568 1290
rect 3516 1226 3568 1232
rect 3988 800 4016 2468
rect 4080 2446 4108 4014
rect 4172 2922 4200 8502
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4264 3534 4292 4966
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4264 3058 4292 3470
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4160 2916 4212 2922
rect 4160 2858 4212 2864
rect 4356 2774 4384 5034
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4448 4146 4476 4694
rect 4436 4140 4488 4146
rect 4436 4082 4488 4088
rect 4436 3528 4488 3534
rect 4436 3470 4488 3476
rect 4448 3194 4476 3470
rect 4436 3188 4488 3194
rect 4436 3130 4488 3136
rect 4540 3074 4568 5850
rect 4632 5574 4660 8774
rect 4896 6180 4948 6186
rect 4896 6122 4948 6128
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4804 5568 4856 5574
rect 4804 5510 4856 5516
rect 4618 4040 4674 4049
rect 4618 3975 4674 3984
rect 4632 3942 4660 3975
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4712 3460 4764 3466
rect 4712 3402 4764 3408
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3097 4660 3334
rect 4448 3046 4568 3074
rect 4618 3088 4674 3097
rect 4448 2922 4476 3046
rect 4618 3023 4674 3032
rect 4528 2984 4580 2990
rect 4528 2926 4580 2932
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 4356 2746 4476 2774
rect 4068 2440 4120 2446
rect 4068 2382 4120 2388
rect 4080 1630 4108 2382
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 4172 1698 4200 2246
rect 4448 2106 4476 2746
rect 4436 2100 4488 2106
rect 4436 2042 4488 2048
rect 4160 1692 4212 1698
rect 4160 1634 4212 1640
rect 4068 1624 4120 1630
rect 4068 1566 4120 1572
rect 4540 800 4568 2926
rect 4618 2816 4674 2825
rect 4618 2751 4674 2760
rect 4632 2446 4660 2751
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4632 1902 4660 2246
rect 4620 1896 4672 1902
rect 4620 1838 4672 1844
rect 4724 1737 4752 3402
rect 4816 2825 4844 5510
rect 4908 4146 4936 6122
rect 5000 5914 5028 12271
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 5264 11688 5316 11694
rect 5264 11630 5316 11636
rect 5172 6996 5224 7002
rect 5172 6938 5224 6944
rect 5080 6248 5132 6254
rect 5080 6190 5132 6196
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4988 5024 5040 5030
rect 4988 4966 5040 4972
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 5000 4010 5028 4966
rect 4896 4004 4948 4010
rect 4896 3946 4948 3952
rect 4988 4004 5040 4010
rect 4988 3946 5040 3952
rect 4908 3058 4936 3946
rect 5000 3534 5028 3946
rect 5092 3942 5120 6190
rect 5080 3936 5132 3942
rect 5080 3878 5132 3884
rect 5080 3664 5132 3670
rect 5080 3606 5132 3612
rect 5092 3534 5120 3606
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 4896 3052 4948 3058
rect 4896 2994 4948 3000
rect 4896 2848 4948 2854
rect 4802 2816 4858 2825
rect 4896 2790 4948 2796
rect 4802 2751 4858 2760
rect 4908 2446 4936 2790
rect 5092 2446 5120 3470
rect 5184 3058 5212 6938
rect 5276 4468 5304 11630
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6552 10600 6604 10606
rect 6552 10542 6604 10548
rect 5448 10192 5500 10198
rect 5448 10134 5500 10140
rect 5354 6896 5410 6905
rect 5354 6831 5410 6840
rect 5368 4622 5396 6831
rect 5460 5234 5488 10134
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 5630 8936 5686 8945
rect 5630 8871 5686 8880
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5552 4826 5580 7346
rect 5644 5914 5672 8871
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6274 6760 6330 6769
rect 6274 6695 6276 6704
rect 6328 6695 6330 6704
rect 6276 6666 6328 6672
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 6564 6322 6592 10542
rect 6736 10532 6788 10538
rect 6736 10474 6788 10480
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6000 6112 6052 6118
rect 6000 6054 6052 6060
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 6012 5817 6040 6054
rect 5998 5808 6054 5817
rect 5908 5772 5960 5778
rect 5998 5743 6054 5752
rect 5908 5714 5960 5720
rect 5540 4820 5592 4826
rect 5540 4762 5592 4768
rect 5722 4720 5778 4729
rect 5722 4655 5778 4664
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5460 4468 5488 4558
rect 5276 4440 5488 4468
rect 5538 4176 5594 4185
rect 5538 4111 5594 4120
rect 5552 4010 5580 4111
rect 5540 4004 5592 4010
rect 5540 3946 5592 3952
rect 5736 3738 5764 4655
rect 5816 4548 5868 4554
rect 5816 4490 5868 4496
rect 5540 3732 5592 3738
rect 5540 3674 5592 3680
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5356 3596 5408 3602
rect 5356 3538 5408 3544
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5172 3052 5224 3058
rect 5172 2994 5224 3000
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 5080 2304 5132 2310
rect 5080 2246 5132 2252
rect 4988 2100 5040 2106
rect 4988 2042 5040 2048
rect 5000 1850 5028 2042
rect 5092 2038 5120 2246
rect 5080 2032 5132 2038
rect 5080 1974 5132 1980
rect 5000 1822 5120 1850
rect 4710 1728 4766 1737
rect 4710 1663 4766 1672
rect 5092 800 5120 1822
rect 5276 1766 5304 3334
rect 5368 2106 5396 3538
rect 5552 3534 5580 3674
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 5724 3528 5776 3534
rect 5724 3470 5776 3476
rect 5632 3120 5684 3126
rect 5632 3062 5684 3068
rect 5448 2848 5500 2854
rect 5448 2790 5500 2796
rect 5356 2100 5408 2106
rect 5356 2042 5408 2048
rect 5264 1760 5316 1766
rect 5264 1702 5316 1708
rect 5460 1601 5488 2790
rect 5540 2372 5592 2378
rect 5540 2314 5592 2320
rect 5552 2009 5580 2314
rect 5538 2000 5594 2009
rect 5538 1935 5594 1944
rect 5446 1592 5502 1601
rect 5446 1527 5502 1536
rect 5644 800 5672 3062
rect 5736 1562 5764 3470
rect 5828 2689 5856 4490
rect 5920 2854 5948 5714
rect 6564 5681 6592 6054
rect 6550 5672 6606 5681
rect 6550 5607 6606 5616
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 6656 5370 6684 6394
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6460 5296 6512 5302
rect 6458 5264 6460 5273
rect 6512 5264 6514 5273
rect 6748 5234 6776 10474
rect 7104 9172 7156 9178
rect 7104 9114 7156 9120
rect 7010 8392 7066 8401
rect 7010 8327 7066 8336
rect 6918 7848 6974 7857
rect 6918 7783 6920 7792
rect 6972 7783 6974 7792
rect 6920 7754 6972 7760
rect 6932 6798 6960 7754
rect 7024 6934 7052 8327
rect 7012 6928 7064 6934
rect 7012 6870 7064 6876
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6840 6322 6868 6598
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 7010 6216 7066 6225
rect 7010 6151 7012 6160
rect 7064 6151 7066 6160
rect 7012 6122 7064 6128
rect 6920 5704 6972 5710
rect 6920 5646 6972 5652
rect 6458 5199 6514 5208
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6550 5128 6606 5137
rect 6550 5063 6606 5072
rect 6564 4622 6592 5063
rect 6932 5030 6960 5646
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 7116 4842 7144 9114
rect 7208 6662 7236 12106
rect 7380 10260 7432 10266
rect 7380 10202 7432 10208
rect 7288 8492 7340 8498
rect 7288 8434 7340 8440
rect 7196 6656 7248 6662
rect 7196 6598 7248 6604
rect 7196 5704 7248 5710
rect 7196 5646 7248 5652
rect 7208 5302 7236 5646
rect 7196 5296 7248 5302
rect 7196 5238 7248 5244
rect 6932 4814 7144 4842
rect 6552 4616 6604 4622
rect 6552 4558 6604 4564
rect 6148 4380 6456 4400
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6550 3632 6606 3641
rect 6550 3567 6606 3576
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5908 2848 5960 2854
rect 5908 2790 5960 2796
rect 5814 2680 5870 2689
rect 5814 2615 5870 2624
rect 6012 1834 6040 3334
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 6564 2922 6592 3567
rect 6642 3496 6698 3505
rect 6642 3431 6698 3440
rect 6656 3398 6684 3431
rect 6644 3392 6696 3398
rect 6644 3334 6696 3340
rect 6736 3392 6788 3398
rect 6736 3334 6788 3340
rect 6748 3194 6776 3334
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6840 3058 6868 3674
rect 6932 3534 6960 4814
rect 7102 4584 7158 4593
rect 7102 4519 7104 4528
rect 7156 4519 7158 4528
rect 7104 4490 7156 4496
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 7024 4049 7052 4422
rect 7300 4146 7328 8434
rect 7288 4140 7340 4146
rect 7288 4082 7340 4088
rect 7010 4040 7066 4049
rect 7392 4026 7420 10202
rect 8392 9648 8444 9654
rect 8392 9590 8444 9596
rect 7656 9580 7708 9586
rect 7656 9522 7708 9528
rect 7668 9042 7696 9522
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 7944 8974 7972 9454
rect 7932 8968 7984 8974
rect 7932 8910 7984 8916
rect 7944 8634 7972 8910
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 8300 8016 8352 8022
rect 7470 7984 7526 7993
rect 8300 7958 8352 7964
rect 7470 7919 7526 7928
rect 7484 7886 7512 7919
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7840 7744 7892 7750
rect 7840 7686 7892 7692
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7472 6656 7524 6662
rect 7472 6598 7524 6604
rect 7010 3975 7066 3984
rect 7116 3998 7420 4026
rect 6920 3528 6972 3534
rect 6920 3470 6972 3476
rect 6828 3052 6880 3058
rect 6828 2994 6880 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6552 2916 6604 2922
rect 6552 2858 6604 2864
rect 6460 2848 6512 2854
rect 6512 2796 6592 2802
rect 6460 2790 6592 2796
rect 6472 2774 6592 2790
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 6564 1986 6592 2774
rect 6656 2553 6684 2926
rect 6840 2774 6868 2994
rect 6748 2746 6868 2774
rect 6748 2650 6776 2746
rect 6826 2680 6882 2689
rect 6736 2644 6788 2650
rect 7116 2650 7144 3998
rect 7288 3936 7340 3942
rect 7288 3878 7340 3884
rect 6826 2615 6882 2624
rect 7104 2644 7156 2650
rect 6736 2586 6788 2592
rect 6642 2544 6698 2553
rect 6642 2479 6698 2488
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 6748 2106 6776 2382
rect 6840 2281 6868 2615
rect 7104 2586 7156 2592
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7208 2514 7236 2586
rect 7196 2508 7248 2514
rect 7196 2450 7248 2456
rect 6826 2272 6882 2281
rect 6826 2207 6882 2216
rect 6736 2100 6788 2106
rect 6736 2042 6788 2048
rect 6564 1958 6776 1986
rect 6000 1828 6052 1834
rect 6000 1770 6052 1776
rect 6184 1624 6236 1630
rect 6184 1566 6236 1572
rect 5724 1556 5776 1562
rect 5724 1498 5776 1504
rect 6196 800 6224 1566
rect 6748 800 6776 1958
rect 7196 1964 7248 1970
rect 7196 1906 7248 1912
rect 7208 1630 7236 1906
rect 7196 1624 7248 1630
rect 7196 1566 7248 1572
rect 7300 800 7328 3878
rect 7484 1970 7512 6598
rect 7564 5024 7616 5030
rect 7564 4966 7616 4972
rect 7576 4690 7604 4966
rect 7564 4684 7616 4690
rect 7564 4626 7616 4632
rect 7668 4622 7696 7278
rect 7852 6497 7880 7686
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7944 6934 7972 7482
rect 8312 7478 8340 7958
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8022 7304 8078 7313
rect 8022 7239 8024 7248
rect 8076 7239 8078 7248
rect 8024 7210 8076 7216
rect 7932 6928 7984 6934
rect 7932 6870 7984 6876
rect 7838 6488 7894 6497
rect 7838 6423 7894 6432
rect 7932 6316 7984 6322
rect 7932 6258 7984 6264
rect 7944 5914 7972 6258
rect 8116 6248 8168 6254
rect 8116 6190 8168 6196
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 7852 5710 7880 5850
rect 7840 5704 7892 5710
rect 7840 5646 7892 5652
rect 8128 5302 8156 6190
rect 8208 5364 8260 5370
rect 8208 5306 8260 5312
rect 7748 5296 7800 5302
rect 7748 5238 7800 5244
rect 8116 5296 8168 5302
rect 8116 5238 8168 5244
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7760 4078 7788 5238
rect 8114 4584 8170 4593
rect 8114 4519 8170 4528
rect 7840 4140 7892 4146
rect 7840 4082 7892 4088
rect 7564 4072 7616 4078
rect 7564 4014 7616 4020
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 7576 3233 7604 4014
rect 7654 3768 7710 3777
rect 7654 3703 7710 3712
rect 7668 3534 7696 3703
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7562 3224 7618 3233
rect 7562 3159 7618 3168
rect 7656 3120 7708 3126
rect 7656 3062 7708 3068
rect 7564 3052 7616 3058
rect 7564 2994 7616 3000
rect 7576 2582 7604 2994
rect 7564 2576 7616 2582
rect 7564 2518 7616 2524
rect 7668 2310 7696 3062
rect 7760 2990 7788 4014
rect 7852 3194 7880 4082
rect 8022 3768 8078 3777
rect 8022 3703 8078 3712
rect 7932 3596 7984 3602
rect 7932 3538 7984 3544
rect 7840 3188 7892 3194
rect 7840 3130 7892 3136
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7760 2446 7788 2926
rect 7944 2650 7972 3538
rect 8036 3194 8064 3703
rect 8128 3534 8156 4519
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8024 3188 8076 3194
rect 8024 3130 8076 3136
rect 8220 3126 8248 5306
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 4486 8340 4694
rect 8404 4622 8432 9590
rect 8484 7744 8536 7750
rect 8484 7686 8536 7692
rect 8496 6730 8524 7686
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8588 4826 8616 18226
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 9784 16574 9812 18702
rect 9692 16546 9812 16574
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 9496 15020 9548 15026
rect 9496 14962 9548 14968
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 8668 14408 8720 14414
rect 8668 14350 8720 14356
rect 8576 4820 8628 4826
rect 8576 4762 8628 4768
rect 8392 4616 8444 4622
rect 8392 4558 8444 4564
rect 8300 4480 8352 4486
rect 8300 4422 8352 4428
rect 8392 3664 8444 3670
rect 8392 3606 8444 3612
rect 8404 3466 8432 3606
rect 8392 3460 8444 3466
rect 8392 3402 8444 3408
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8208 3120 8260 3126
rect 8208 3062 8260 3068
rect 8390 2816 8446 2825
rect 8390 2751 8446 2760
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 7840 2372 7892 2378
rect 7840 2314 7892 2320
rect 7656 2304 7708 2310
rect 7656 2246 7708 2252
rect 7472 1964 7524 1970
rect 7472 1906 7524 1912
rect 7852 800 7880 2314
rect 8404 800 8432 2751
rect 8588 2428 8616 3334
rect 8680 2650 8708 14350
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 9508 9450 9536 14962
rect 9692 9674 9720 16546
rect 11256 12434 11284 18702
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 12256 18284 12308 18290
rect 12256 18226 12308 18232
rect 12268 17882 12296 18226
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 12256 17876 12308 17882
rect 12256 17818 12308 17824
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11704 15020 11756 15026
rect 11704 14962 11756 14968
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11072 12406 11284 12434
rect 10230 10160 10286 10169
rect 10230 10095 10286 10104
rect 9692 9646 9904 9674
rect 9772 9580 9824 9586
rect 9772 9522 9824 9528
rect 9496 9444 9548 9450
rect 9496 9386 9548 9392
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 9508 8498 9536 8910
rect 9784 8498 9812 9522
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9772 8492 9824 8498
rect 9772 8434 9824 8440
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8772 7410 8800 7822
rect 8944 7812 8996 7818
rect 8944 7754 8996 7760
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8956 7324 8984 7754
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 9036 7336 9088 7342
rect 8956 7296 9036 7324
rect 9036 7278 9088 7284
rect 8747 7100 9055 7120
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 9048 6458 9076 6802
rect 9140 6798 9168 7686
rect 9220 7540 9272 7546
rect 9508 7528 9536 7754
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9632 7542 9688 7551
rect 9784 7546 9812 7686
rect 9508 7500 9632 7528
rect 9220 7482 9272 7488
rect 9232 7449 9260 7482
rect 9632 7477 9688 7486
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9218 7440 9274 7449
rect 9218 7375 9274 7384
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9770 7168 9826 7177
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9220 6656 9272 6662
rect 9220 6598 9272 6604
rect 9036 6452 9088 6458
rect 9036 6394 9088 6400
rect 9126 6352 9182 6361
rect 9126 6287 9182 6296
rect 9140 6089 9168 6287
rect 9126 6080 9182 6089
rect 8747 6012 9055 6032
rect 9126 6015 9182 6024
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5936 9055 5956
rect 9232 5914 9260 6598
rect 9508 6361 9536 7142
rect 9770 7103 9826 7112
rect 9784 6866 9812 7103
rect 9876 6934 9904 9646
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9968 8498 9996 8842
rect 9956 8492 10008 8498
rect 9956 8434 10008 8440
rect 10140 8288 10192 8294
rect 10140 8230 10192 8236
rect 10048 7404 10100 7410
rect 10048 7346 10100 7352
rect 9864 6928 9916 6934
rect 9864 6870 9916 6876
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9586 6488 9642 6497
rect 9586 6423 9642 6432
rect 9494 6352 9550 6361
rect 9404 6316 9456 6322
rect 9494 6287 9550 6296
rect 9404 6258 9456 6264
rect 9220 5908 9272 5914
rect 9220 5850 9272 5856
rect 8760 5840 8812 5846
rect 8760 5782 8812 5788
rect 8772 5642 8800 5782
rect 9416 5658 9444 6258
rect 9600 5692 9628 6423
rect 9680 5704 9732 5710
rect 9600 5664 9680 5692
rect 9416 5642 9536 5658
rect 9680 5646 9732 5652
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 9416 5636 9548 5642
rect 9416 5630 9496 5636
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 9416 4826 9444 5630
rect 9496 5578 9548 5584
rect 9588 5568 9640 5574
rect 9508 5516 9588 5522
rect 9508 5510 9640 5516
rect 9508 5494 9628 5510
rect 9404 4820 9456 4826
rect 9404 4762 9456 4768
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 9140 3738 9168 4558
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9126 3088 9182 3097
rect 9416 3074 9444 4558
rect 9508 4434 9536 5494
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9600 4554 9628 5170
rect 10060 5030 10088 7346
rect 9864 5024 9916 5030
rect 9864 4966 9916 4972
rect 10048 5024 10100 5030
rect 10048 4966 10100 4972
rect 9588 4548 9640 4554
rect 9588 4490 9640 4496
rect 9508 4406 9628 4434
rect 9496 3936 9548 3942
rect 9496 3878 9548 3884
rect 9508 3602 9536 3878
rect 9600 3738 9628 4406
rect 9876 4146 9904 4966
rect 9864 4140 9916 4146
rect 9864 4082 9916 4088
rect 9588 3732 9640 3738
rect 9588 3674 9640 3680
rect 9496 3596 9548 3602
rect 9496 3538 9548 3544
rect 9600 3398 9628 3674
rect 10048 3664 10100 3670
rect 10048 3606 10100 3612
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9494 3088 9550 3097
rect 9416 3046 9494 3074
rect 9126 3023 9182 3032
rect 9494 3023 9496 3032
rect 9140 2825 9168 3023
rect 9548 3023 9550 3032
rect 9496 2994 9548 3000
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9126 2816 9182 2825
rect 8747 2748 9055 2768
rect 9126 2751 9182 2760
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 8668 2644 8720 2650
rect 8668 2586 8720 2592
rect 8942 2544 8998 2553
rect 9508 2514 9536 2858
rect 8942 2479 8998 2488
rect 9496 2508 9548 2514
rect 8668 2440 8720 2446
rect 8588 2400 8668 2428
rect 8668 2382 8720 2388
rect 8956 800 8984 2479
rect 9496 2450 9548 2456
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9508 800 9536 1498
rect 10060 800 10088 3606
rect 10152 2446 10180 8230
rect 10244 6662 10272 10095
rect 10784 9444 10836 9450
rect 10784 9386 10836 9392
rect 10414 9208 10470 9217
rect 10796 9178 10824 9386
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10888 9178 10916 9318
rect 10414 9143 10470 9152
rect 10784 9172 10836 9178
rect 10232 6656 10284 6662
rect 10232 6598 10284 6604
rect 10428 5273 10456 9143
rect 10784 9114 10836 9120
rect 10876 9172 10928 9178
rect 10876 9114 10928 9120
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8430 10548 8774
rect 10692 8560 10744 8566
rect 10692 8502 10744 8508
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 10520 7585 10548 8026
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10506 7576 10562 7585
rect 10612 7546 10640 7890
rect 10506 7511 10562 7520
rect 10600 7540 10652 7546
rect 10520 6866 10548 7511
rect 10600 7482 10652 7488
rect 10508 6860 10560 6866
rect 10508 6802 10560 6808
rect 10508 6316 10560 6322
rect 10508 6258 10560 6264
rect 10520 5710 10548 6258
rect 10508 5704 10560 5710
rect 10508 5646 10560 5652
rect 10520 5370 10548 5646
rect 10508 5364 10560 5370
rect 10508 5306 10560 5312
rect 10414 5264 10470 5273
rect 10414 5199 10470 5208
rect 10598 3224 10654 3233
rect 10508 3188 10560 3194
rect 10598 3159 10654 3168
rect 10508 3130 10560 3136
rect 10520 2514 10548 3130
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 10140 2440 10192 2446
rect 10140 2382 10192 2388
rect 10612 800 10640 3159
rect 10704 1698 10732 8502
rect 10784 8424 10836 8430
rect 10784 8366 10836 8372
rect 10796 7886 10824 8366
rect 10784 7880 10836 7886
rect 10784 7822 10836 7828
rect 10796 7206 10824 7822
rect 10968 7812 11020 7818
rect 10968 7754 11020 7760
rect 10980 7698 11008 7754
rect 10888 7670 11008 7698
rect 10784 7200 10836 7206
rect 10784 7142 10836 7148
rect 10888 7002 10916 7670
rect 10966 7440 11022 7449
rect 10966 7375 10968 7384
rect 11020 7375 11022 7384
rect 10968 7346 11020 7352
rect 10876 6996 10928 7002
rect 10876 6938 10928 6944
rect 11072 6662 11100 12406
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11152 10056 11204 10062
rect 11152 9998 11204 10004
rect 11164 9722 11192 9998
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11152 9716 11204 9722
rect 11152 9658 11204 9664
rect 11164 9042 11192 9658
rect 11244 9580 11296 9586
rect 11244 9522 11296 9528
rect 11152 9036 11204 9042
rect 11152 8978 11204 8984
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11164 8634 11192 8774
rect 11256 8634 11284 9522
rect 11716 8838 11744 14962
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 12084 12434 12112 13874
rect 11900 12406 12112 12434
rect 11796 9920 11848 9926
rect 11796 9862 11848 9868
rect 11808 9586 11836 9862
rect 11900 9625 11928 12406
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11980 10464 12032 10470
rect 11980 10406 12032 10412
rect 11886 9616 11942 9625
rect 11796 9580 11848 9586
rect 11886 9551 11942 9560
rect 11796 9522 11848 9528
rect 11886 9344 11942 9353
rect 11886 9279 11942 9288
rect 11704 8832 11756 8838
rect 11704 8774 11756 8780
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 11152 8628 11204 8634
rect 11152 8570 11204 8576
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11152 8356 11204 8362
rect 11152 8298 11204 8304
rect 11164 7546 11192 8298
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 11256 6730 11284 7686
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 11612 7200 11664 7206
rect 11612 7142 11664 7148
rect 11796 7200 11848 7206
rect 11796 7142 11848 7148
rect 11624 7002 11652 7142
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 11808 6798 11836 7142
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11244 6724 11296 6730
rect 11244 6666 11296 6672
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 11794 6488 11850 6497
rect 11794 6423 11850 6432
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 10876 6112 10928 6118
rect 10876 6054 10928 6060
rect 10888 4622 10916 6054
rect 11060 5568 11112 5574
rect 11060 5510 11112 5516
rect 11072 5302 11100 5510
rect 11060 5296 11112 5302
rect 11060 5238 11112 5244
rect 11072 4622 11100 5238
rect 11164 4826 11192 6258
rect 11612 6180 11664 6186
rect 11612 6122 11664 6128
rect 11624 5710 11652 6122
rect 11808 6089 11836 6423
rect 11794 6080 11850 6089
rect 11794 6015 11850 6024
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 11612 5160 11664 5166
rect 11612 5102 11664 5108
rect 11624 4826 11652 5102
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 11612 4820 11664 4826
rect 11612 4762 11664 4768
rect 10876 4616 10928 4622
rect 10876 4558 10928 4564
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4162 11100 4558
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 10876 4140 10928 4146
rect 10796 4100 10876 4128
rect 10796 2514 10824 4100
rect 11072 4134 11192 4162
rect 10876 4082 10928 4088
rect 11060 4072 11112 4078
rect 11060 4014 11112 4020
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3466 11008 3878
rect 10968 3460 11020 3466
rect 10968 3402 11020 3408
rect 11072 2650 11100 4014
rect 11164 3534 11192 4134
rect 11428 4004 11480 4010
rect 11428 3946 11480 3952
rect 11440 3738 11468 3946
rect 11900 3942 11928 9279
rect 11992 9217 12020 10406
rect 12072 9920 12124 9926
rect 12072 9862 12124 9868
rect 11978 9208 12034 9217
rect 11978 9143 12034 9152
rect 11980 9104 12032 9110
rect 11980 9046 12032 9052
rect 11992 7410 12020 9046
rect 12084 8974 12112 9862
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 12176 8786 12204 11834
rect 12084 8758 12204 8786
rect 11980 7404 12032 7410
rect 11980 7346 12032 7352
rect 11992 7206 12020 7346
rect 11980 7200 12032 7206
rect 11980 7142 12032 7148
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11992 3942 12020 6190
rect 12084 5522 12112 8758
rect 12164 7812 12216 7818
rect 12164 7754 12216 7760
rect 12176 5710 12204 7754
rect 12268 6458 12296 17614
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 14292 16574 14320 17138
rect 14292 16546 14780 16574
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 12992 16040 13044 16046
rect 12992 15982 13044 15988
rect 13004 15162 13032 15982
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 12992 15156 13044 15162
rect 12992 15098 13044 15104
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 12808 14272 12860 14278
rect 12808 14214 12860 14220
rect 12440 12368 12492 12374
rect 12440 12310 12492 12316
rect 12452 11626 12480 12310
rect 12440 11620 12492 11626
rect 12440 11562 12492 11568
rect 12452 11354 12480 11562
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12348 10600 12400 10606
rect 12348 10542 12400 10548
rect 12360 9654 12388 10542
rect 12440 9920 12492 9926
rect 12440 9862 12492 9868
rect 12348 9648 12400 9654
rect 12348 9590 12400 9596
rect 12360 8974 12388 9590
rect 12452 8974 12480 9862
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12440 8968 12492 8974
rect 12440 8910 12492 8916
rect 12360 8090 12388 8910
rect 12452 8634 12480 8910
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12532 8424 12584 8430
rect 12532 8366 12584 8372
rect 12348 8084 12400 8090
rect 12348 8026 12400 8032
rect 12360 7478 12388 8026
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12440 6860 12492 6866
rect 12440 6802 12492 6808
rect 12256 6452 12308 6458
rect 12256 6394 12308 6400
rect 12256 6180 12308 6186
rect 12256 6122 12308 6128
rect 12268 5914 12296 6122
rect 12256 5908 12308 5914
rect 12256 5850 12308 5856
rect 12452 5710 12480 6802
rect 12544 6798 12572 8366
rect 12532 6792 12584 6798
rect 12532 6734 12584 6740
rect 12164 5704 12216 5710
rect 12164 5646 12216 5652
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12084 5494 12204 5522
rect 12072 5364 12124 5370
rect 12072 5306 12124 5312
rect 12084 4622 12112 5306
rect 12176 5234 12204 5494
rect 12164 5228 12216 5234
rect 12164 5170 12216 5176
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 12072 4616 12124 4622
rect 12072 4558 12124 4564
rect 12452 4486 12480 5034
rect 12440 4480 12492 4486
rect 12440 4422 12492 4428
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11428 3732 11480 3738
rect 11428 3674 11480 3680
rect 11152 3528 11204 3534
rect 11152 3470 11204 3476
rect 11164 3058 11192 3470
rect 11440 3380 11468 3674
rect 11796 3528 11848 3534
rect 11794 3496 11796 3505
rect 11848 3496 11850 3505
rect 11794 3431 11850 3440
rect 11256 3352 11468 3380
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11060 2644 11112 2650
rect 11060 2586 11112 2592
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 10784 2304 10836 2310
rect 10784 2246 10836 2252
rect 10796 1766 10824 2246
rect 10784 1760 10836 1766
rect 10784 1702 10836 1708
rect 10692 1692 10744 1698
rect 10692 1634 10744 1640
rect 10888 1601 10916 2450
rect 11256 2446 11284 3352
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11532 2854 11560 2994
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 11704 2848 11756 2854
rect 11704 2790 11756 2796
rect 11244 2440 11296 2446
rect 11244 2382 11296 2388
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 1902 11008 2246
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 11152 2100 11204 2106
rect 11152 2042 11204 2048
rect 10968 1896 11020 1902
rect 10968 1838 11020 1844
rect 10874 1592 10930 1601
rect 10874 1527 10930 1536
rect 11164 800 11192 2042
rect 11716 800 11744 2790
rect 12084 2009 12112 4150
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12440 3392 12492 3398
rect 12544 3369 12572 4082
rect 12440 3334 12492 3340
rect 12530 3360 12586 3369
rect 12452 3126 12480 3334
rect 12530 3295 12586 3304
rect 12440 3120 12492 3126
rect 12440 3062 12492 3068
rect 12164 2576 12216 2582
rect 12164 2518 12216 2524
rect 12070 2000 12126 2009
rect 12070 1935 12126 1944
rect 12176 800 12204 2518
rect 12452 2514 12480 3062
rect 12636 2774 12664 5646
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12544 2746 12664 2774
rect 12544 2650 12572 2746
rect 12532 2644 12584 2650
rect 12532 2586 12584 2592
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12728 800 12756 3606
rect 12820 2446 12848 14214
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 13544 13320 13596 13326
rect 13544 13262 13596 13268
rect 13556 12434 13584 13262
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 13464 12406 13584 12434
rect 13268 11552 13320 11558
rect 13268 11494 13320 11500
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12912 8974 12940 9862
rect 12992 9716 13044 9722
rect 12992 9658 13044 9664
rect 12900 8968 12952 8974
rect 12900 8910 12952 8916
rect 12900 8832 12952 8838
rect 12900 8774 12952 8780
rect 12912 7886 12940 8774
rect 13004 8430 13032 9658
rect 12992 8424 13044 8430
rect 12992 8366 13044 8372
rect 13096 8090 13124 10610
rect 13280 10033 13308 11494
rect 13266 10024 13322 10033
rect 13266 9959 13322 9968
rect 13084 8084 13136 8090
rect 13084 8026 13136 8032
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7002 12940 7822
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13004 6882 13032 7686
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12912 6854 13032 6882
rect 12912 3942 12940 6854
rect 13096 5914 13124 7346
rect 13464 6882 13492 12406
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14200 11801 14228 12038
rect 14186 11792 14242 11801
rect 13820 11756 13872 11762
rect 14186 11727 14242 11736
rect 14280 11756 14332 11762
rect 13820 11698 13872 11704
rect 14280 11698 14332 11704
rect 13832 10810 13860 11698
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 14292 11286 14320 11698
rect 14280 11280 14332 11286
rect 14280 11222 14332 11228
rect 14384 11121 14412 12038
rect 14370 11112 14426 11121
rect 14370 11047 14426 11056
rect 14280 11008 14332 11014
rect 14280 10950 14332 10956
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 13832 10130 13860 10746
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 13820 10124 13872 10130
rect 13820 10066 13872 10072
rect 14292 10062 14320 10950
rect 14384 10266 14412 11047
rect 14372 10260 14424 10266
rect 14372 10202 14424 10208
rect 13544 10056 13596 10062
rect 13544 9998 13596 10004
rect 14280 10056 14332 10062
rect 14280 9998 14332 10004
rect 13556 9722 13584 9998
rect 14372 9920 14424 9926
rect 14372 9862 14424 9868
rect 13544 9716 13596 9722
rect 13544 9658 13596 9664
rect 13728 9512 13780 9518
rect 13728 9454 13780 9460
rect 13636 9444 13688 9450
rect 13636 9386 13688 9392
rect 13544 9172 13596 9178
rect 13544 9114 13596 9120
rect 13556 8838 13584 9114
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13648 8634 13676 9386
rect 13740 9178 13768 9454
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 13728 9172 13780 9178
rect 13728 9114 13780 9120
rect 14384 8634 14412 9862
rect 14476 9450 14504 16050
rect 14556 11552 14608 11558
rect 14556 11494 14608 11500
rect 14648 11552 14700 11558
rect 14648 11494 14700 11500
rect 14568 10742 14596 11494
rect 14660 11218 14688 11494
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14556 10736 14608 10742
rect 14556 10678 14608 10684
rect 14464 9444 14516 9450
rect 14464 9386 14516 9392
rect 14648 9376 14700 9382
rect 14648 9318 14700 9324
rect 14660 8906 14688 9318
rect 14648 8900 14700 8906
rect 14648 8842 14700 8848
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 13728 8424 13780 8430
rect 13728 8366 13780 8372
rect 13636 8016 13688 8022
rect 13636 7958 13688 7964
rect 13464 6854 13584 6882
rect 13452 6792 13504 6798
rect 13452 6734 13504 6740
rect 13464 6458 13492 6734
rect 13452 6452 13504 6458
rect 13452 6394 13504 6400
rect 13452 6316 13504 6322
rect 13452 6258 13504 6264
rect 13176 6248 13228 6254
rect 13176 6190 13228 6196
rect 13360 6248 13412 6254
rect 13360 6190 13412 6196
rect 13084 5908 13136 5914
rect 13084 5850 13136 5856
rect 13188 5370 13216 6190
rect 13372 5370 13400 6190
rect 13464 5914 13492 6258
rect 13452 5908 13504 5914
rect 13452 5850 13504 5856
rect 13176 5364 13228 5370
rect 13176 5306 13228 5312
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13360 4548 13412 4554
rect 13360 4490 13412 4496
rect 12992 4480 13044 4486
rect 12992 4422 13044 4428
rect 13004 4078 13032 4422
rect 13372 4214 13400 4490
rect 13268 4208 13320 4214
rect 13268 4150 13320 4156
rect 13360 4208 13412 4214
rect 13360 4150 13412 4156
rect 12992 4072 13044 4078
rect 12992 4014 13044 4020
rect 12900 3936 12952 3942
rect 12900 3878 12952 3884
rect 13176 3936 13228 3942
rect 13176 3878 13228 3884
rect 12808 2440 12860 2446
rect 12808 2382 12860 2388
rect 12808 2304 12860 2310
rect 12808 2246 12860 2252
rect 12820 1834 12848 2246
rect 12808 1828 12860 1834
rect 12808 1770 12860 1776
rect 12912 1630 12940 3878
rect 13188 3194 13216 3878
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 13280 2650 13308 4150
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13464 3194 13492 4082
rect 13556 4010 13584 6854
rect 13648 6390 13676 7958
rect 13740 7886 13768 8366
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13740 7546 13768 7822
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 14370 7168 14426 7177
rect 13945 7100 14253 7120
rect 14370 7103 14426 7112
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 13820 6656 13872 6662
rect 13820 6598 13872 6604
rect 13636 6384 13688 6390
rect 13636 6326 13688 6332
rect 13636 6248 13688 6254
rect 13636 6190 13688 6196
rect 13648 5234 13676 6190
rect 13728 5568 13780 5574
rect 13728 5510 13780 5516
rect 13636 5228 13688 5234
rect 13636 5170 13688 5176
rect 13648 4622 13676 5170
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13544 4004 13596 4010
rect 13544 3946 13596 3952
rect 13648 3534 13676 4558
rect 13740 4162 13768 5510
rect 13832 5302 13860 6598
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 13820 5296 13872 5302
rect 14188 5296 14240 5302
rect 13820 5238 13872 5244
rect 14186 5264 14188 5273
rect 14240 5264 14242 5273
rect 14186 5199 14242 5208
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 14292 4486 14320 5170
rect 14280 4480 14332 4486
rect 14280 4422 14332 4428
rect 13740 4134 13860 4162
rect 13728 4072 13780 4078
rect 13728 4014 13780 4020
rect 13636 3528 13688 3534
rect 13636 3470 13688 3476
rect 13740 3194 13768 4014
rect 13452 3188 13504 3194
rect 13452 3130 13504 3136
rect 13728 3188 13780 3194
rect 13728 3130 13780 3136
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13372 2990 13400 3062
rect 13728 3052 13780 3058
rect 13728 2994 13780 3000
rect 13360 2984 13412 2990
rect 13360 2926 13412 2932
rect 13360 2848 13412 2854
rect 13740 2825 13768 2994
rect 13360 2790 13412 2796
rect 13726 2816 13782 2825
rect 13268 2644 13320 2650
rect 13268 2586 13320 2592
rect 12900 1624 12952 1630
rect 12900 1566 12952 1572
rect 13372 1442 13400 2790
rect 13726 2751 13782 2760
rect 13280 1414 13400 1442
rect 13280 800 13308 1414
rect 13832 800 13860 4134
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 13912 3392 13964 3398
rect 13912 3334 13964 3340
rect 13924 2922 13952 3334
rect 14292 3126 14320 4422
rect 14384 3670 14412 7103
rect 14752 6458 14780 16546
rect 14924 13456 14976 13462
rect 14924 13398 14976 13404
rect 14832 12096 14884 12102
rect 14832 12038 14884 12044
rect 14844 11694 14872 12038
rect 14832 11688 14884 11694
rect 14832 11630 14884 11636
rect 14832 11144 14884 11150
rect 14832 11086 14884 11092
rect 14844 10674 14872 11086
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14740 6452 14792 6458
rect 14740 6394 14792 6400
rect 14832 6452 14884 6458
rect 14832 6394 14884 6400
rect 14844 6338 14872 6394
rect 14568 6310 14872 6338
rect 14936 6322 14964 13398
rect 15016 12640 15068 12646
rect 15016 12582 15068 12588
rect 15028 12238 15056 12582
rect 15016 12232 15068 12238
rect 15016 12174 15068 12180
rect 15028 9586 15056 12174
rect 15120 10266 15148 17206
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15212 14890 15240 16458
rect 15292 15564 15344 15570
rect 15292 15506 15344 15512
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15304 14074 15332 15506
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15292 14068 15344 14074
rect 15292 14010 15344 14016
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15290 13288 15346 13297
rect 15290 13223 15346 13232
rect 15200 12164 15252 12170
rect 15200 12106 15252 12112
rect 15212 11762 15240 12106
rect 15200 11756 15252 11762
rect 15200 11698 15252 11704
rect 15200 11620 15252 11626
rect 15200 11562 15252 11568
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15212 8650 15240 11562
rect 15304 10146 15332 13223
rect 15396 13190 15424 13806
rect 15384 13184 15436 13190
rect 15384 13126 15436 13132
rect 15396 11778 15424 13126
rect 15488 12442 15516 14554
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15476 12436 15528 12442
rect 15856 12434 15884 12718
rect 15856 12406 16068 12434
rect 15476 12378 15528 12384
rect 15396 11750 15976 11778
rect 15476 11688 15528 11694
rect 15476 11630 15528 11636
rect 15752 11688 15804 11694
rect 15752 11630 15804 11636
rect 15384 11008 15436 11014
rect 15384 10950 15436 10956
rect 15396 10742 15424 10950
rect 15384 10736 15436 10742
rect 15384 10678 15436 10684
rect 15304 10118 15424 10146
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9518 15332 9930
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 8838 15332 9454
rect 15292 8832 15344 8838
rect 15292 8774 15344 8780
rect 15212 8622 15332 8650
rect 15304 8498 15332 8622
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15304 8401 15332 8434
rect 15290 8392 15346 8401
rect 15290 8327 15346 8336
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6798 15240 7142
rect 15290 6896 15346 6905
rect 15290 6831 15346 6840
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 14924 6316 14976 6322
rect 14568 6118 14596 6310
rect 14924 6258 14976 6264
rect 14556 6112 14608 6118
rect 14556 6054 14608 6060
rect 14556 5772 14608 5778
rect 14556 5714 14608 5720
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 4282 14504 5510
rect 14568 5166 14596 5714
rect 14648 5568 14700 5574
rect 14648 5510 14700 5516
rect 14556 5160 14608 5166
rect 14556 5102 14608 5108
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14372 3664 14424 3670
rect 14372 3606 14424 3612
rect 14476 3233 14504 3674
rect 14462 3224 14518 3233
rect 14462 3159 14518 3168
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 13912 2916 13964 2922
rect 13912 2858 13964 2864
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 14660 2553 14688 5510
rect 14832 5296 14884 5302
rect 14830 5264 14832 5273
rect 14884 5264 14886 5273
rect 14830 5199 14886 5208
rect 14936 5250 14964 6258
rect 15106 5808 15162 5817
rect 15212 5778 15240 6734
rect 15304 6497 15332 6831
rect 15290 6488 15346 6497
rect 15290 6423 15346 6432
rect 15106 5743 15162 5752
rect 15200 5772 15252 5778
rect 15120 5710 15148 5743
rect 15200 5714 15252 5720
rect 15108 5704 15160 5710
rect 15108 5646 15160 5652
rect 14936 5234 15056 5250
rect 14936 5228 15068 5234
rect 14936 5222 15016 5228
rect 14844 4078 14872 5199
rect 14936 4690 14964 5222
rect 15016 5170 15068 5176
rect 14924 4684 14976 4690
rect 14924 4626 14976 4632
rect 15120 4146 15148 5646
rect 15396 4570 15424 10118
rect 15488 9722 15516 11630
rect 15568 10464 15620 10470
rect 15568 10406 15620 10412
rect 15660 10464 15712 10470
rect 15660 10406 15712 10412
rect 15580 10062 15608 10406
rect 15672 10198 15700 10406
rect 15764 10266 15792 11630
rect 15844 11620 15896 11626
rect 15844 11562 15896 11568
rect 15856 11286 15884 11562
rect 15844 11280 15896 11286
rect 15844 11222 15896 11228
rect 15948 11098 15976 11750
rect 15856 11070 15976 11098
rect 15856 10606 15884 11070
rect 15844 10600 15896 10606
rect 15844 10542 15896 10548
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15568 10056 15620 10062
rect 15568 9998 15620 10004
rect 15476 9716 15528 9722
rect 15476 9658 15528 9664
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15660 8832 15712 8838
rect 15660 8774 15712 8780
rect 15488 8430 15516 8774
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 7410 15516 8366
rect 15672 8362 15700 8774
rect 15660 8356 15712 8362
rect 15660 8298 15712 8304
rect 15568 7948 15620 7954
rect 15568 7890 15620 7896
rect 15476 7404 15528 7410
rect 15476 7346 15528 7352
rect 15580 6798 15608 7890
rect 15660 7812 15712 7818
rect 15660 7754 15712 7760
rect 15568 6792 15620 6798
rect 15568 6734 15620 6740
rect 15476 6656 15528 6662
rect 15476 6598 15528 6604
rect 15568 6656 15620 6662
rect 15568 6598 15620 6604
rect 15488 4826 15516 6598
rect 15580 5030 15608 6598
rect 15672 5710 15700 7754
rect 15856 7750 15884 10542
rect 15936 8560 15988 8566
rect 15936 8502 15988 8508
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15752 6792 15804 6798
rect 15752 6734 15804 6740
rect 15764 6662 15792 6734
rect 15844 6724 15896 6730
rect 15844 6666 15896 6672
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15752 6112 15804 6118
rect 15752 6054 15804 6060
rect 15764 5953 15792 6054
rect 15750 5944 15806 5953
rect 15750 5879 15806 5888
rect 15660 5704 15712 5710
rect 15660 5646 15712 5652
rect 15568 5024 15620 5030
rect 15568 4966 15620 4972
rect 15476 4820 15528 4826
rect 15476 4762 15528 4768
rect 15396 4542 15516 4570
rect 15384 4480 15436 4486
rect 15384 4422 15436 4428
rect 15396 4185 15424 4422
rect 15382 4176 15438 4185
rect 15108 4140 15160 4146
rect 15382 4111 15438 4120
rect 15108 4082 15160 4088
rect 14832 4072 14884 4078
rect 14832 4014 14884 4020
rect 14740 4004 14792 4010
rect 14740 3946 14792 3952
rect 14752 3738 14780 3946
rect 14740 3732 14792 3738
rect 14740 3674 14792 3680
rect 14740 3188 14792 3194
rect 14844 3176 14872 4014
rect 15488 3942 15516 4542
rect 15568 4208 15620 4214
rect 15568 4150 15620 4156
rect 15476 3936 15528 3942
rect 15476 3878 15528 3884
rect 15198 3632 15254 3641
rect 15198 3567 15254 3576
rect 15212 3534 15240 3567
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 14792 3148 14872 3176
rect 15200 3188 15252 3194
rect 14740 3130 14792 3136
rect 15200 3130 15252 3136
rect 14924 2916 14976 2922
rect 14924 2858 14976 2864
rect 14646 2544 14702 2553
rect 14646 2479 14702 2488
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 14188 2304 14240 2310
rect 14188 2246 14240 2252
rect 14200 2106 14228 2246
rect 14188 2100 14240 2106
rect 14188 2042 14240 2048
rect 14476 1170 14504 2382
rect 14384 1142 14504 1170
rect 14384 800 14412 1142
rect 14936 800 14964 2858
rect 15212 2514 15240 3130
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 15292 2304 15344 2310
rect 15292 2246 15344 2252
rect 15304 1970 15332 2246
rect 15292 1964 15344 1970
rect 15292 1906 15344 1912
rect 15488 800 15516 3334
rect 15580 2650 15608 4150
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 15672 3194 15700 3402
rect 15660 3188 15712 3194
rect 15660 3130 15712 3136
rect 15764 2650 15792 4082
rect 15856 2774 15884 6666
rect 15948 3913 15976 8502
rect 16040 7018 16068 12406
rect 16132 7886 16160 13942
rect 16224 11898 16252 19382
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 17328 16574 17356 20198
rect 18892 20058 18920 20402
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 19524 19848 19576 19854
rect 19524 19790 19576 19796
rect 19536 19514 19564 19790
rect 19524 19508 19576 19514
rect 19524 19450 19576 19456
rect 18420 19372 18472 19378
rect 18420 19314 18472 19320
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17236 16546 17356 16574
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17144 14346 17172 14826
rect 17132 14340 17184 14346
rect 17132 14282 17184 14288
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 17236 13326 17264 16546
rect 17972 16250 18000 17070
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17868 16108 17920 16114
rect 17868 16050 17920 16056
rect 17408 13864 17460 13870
rect 17408 13806 17460 13812
rect 17224 13320 17276 13326
rect 17224 13262 17276 13268
rect 17316 13252 17368 13258
rect 17316 13194 17368 13200
rect 17224 13184 17276 13190
rect 17224 13126 17276 13132
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16304 12096 16356 12102
rect 16304 12038 16356 12044
rect 16212 11892 16264 11898
rect 16212 11834 16264 11840
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16224 7546 16252 8842
rect 16212 7540 16264 7546
rect 16212 7482 16264 7488
rect 16040 6990 16252 7018
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 16040 6118 16068 6802
rect 16028 6112 16080 6118
rect 16028 6054 16080 6060
rect 16120 6112 16172 6118
rect 16120 6054 16172 6060
rect 16040 5778 16068 6054
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 16040 5302 16068 5714
rect 16028 5296 16080 5302
rect 16028 5238 16080 5244
rect 15934 3904 15990 3913
rect 15934 3839 15990 3848
rect 16132 3777 16160 6054
rect 16224 4214 16252 6990
rect 16316 6662 16344 12038
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 16580 11824 16632 11830
rect 16580 11766 16632 11772
rect 16592 11354 16620 11766
rect 16960 11558 16988 12854
rect 17040 12844 17092 12850
rect 17040 12786 17092 12792
rect 16948 11552 17000 11558
rect 16948 11494 17000 11500
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16684 11257 16712 11290
rect 16670 11248 16726 11257
rect 16670 11183 16726 11192
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16396 11008 16448 11014
rect 16396 10950 16448 10956
rect 16408 10690 16436 10950
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16960 10849 16988 11086
rect 16946 10840 17002 10849
rect 16946 10775 17002 10784
rect 17052 10690 17080 12786
rect 17132 12096 17184 12102
rect 17132 12038 17184 12044
rect 17144 11762 17172 12038
rect 17236 11830 17264 13126
rect 17224 11824 17276 11830
rect 17224 11766 17276 11772
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 17144 11218 17172 11698
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 17132 11212 17184 11218
rect 17132 11154 17184 11160
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 16408 10662 16620 10690
rect 16592 10266 16620 10662
rect 16960 10662 17080 10690
rect 16960 10470 16988 10662
rect 17040 10532 17092 10538
rect 17040 10474 17092 10480
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 16580 10260 16632 10266
rect 16580 10202 16632 10208
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 16960 9602 16988 10406
rect 17052 10266 17080 10474
rect 17040 10260 17092 10266
rect 17040 10202 17092 10208
rect 17144 10198 17172 10950
rect 17132 10192 17184 10198
rect 17132 10134 17184 10140
rect 17132 9920 17184 9926
rect 17132 9862 17184 9868
rect 16960 9574 17080 9602
rect 17052 9518 17080 9574
rect 16764 9512 16816 9518
rect 16764 9454 16816 9460
rect 16948 9512 17000 9518
rect 16948 9454 17000 9460
rect 17040 9512 17092 9518
rect 17040 9454 17092 9460
rect 16776 9042 16804 9454
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16408 8566 16436 8910
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 16960 8634 16988 9454
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16396 8560 16448 8566
rect 16396 8502 16448 8508
rect 17040 8288 17092 8294
rect 16394 8256 16450 8265
rect 17144 8276 17172 9862
rect 17236 8838 17264 11494
rect 17224 8832 17276 8838
rect 17224 8774 17276 8780
rect 17092 8248 17172 8276
rect 17040 8230 17092 8236
rect 16394 8191 16450 8200
rect 16408 7585 16436 8191
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16394 7576 16450 7585
rect 16544 7568 16852 7588
rect 16394 7511 16450 7520
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16396 6928 16448 6934
rect 16396 6870 16448 6876
rect 16304 6656 16356 6662
rect 16304 6598 16356 6604
rect 16408 5234 16436 6870
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 16856 6384 16908 6390
rect 16960 6372 16988 7278
rect 17144 6984 17172 8248
rect 17144 6956 17264 6984
rect 17040 6724 17092 6730
rect 17040 6666 17092 6672
rect 16908 6344 16988 6372
rect 16856 6326 16908 6332
rect 17052 5914 17080 6666
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 16396 5228 16448 5234
rect 16396 5170 16448 5176
rect 17040 5228 17092 5234
rect 17236 5216 17264 6956
rect 17092 5188 17264 5216
rect 17040 5170 17092 5176
rect 16856 5160 16908 5166
rect 16856 5102 16908 5108
rect 16868 4865 16896 5102
rect 16948 5024 17000 5030
rect 16948 4966 17000 4972
rect 16854 4856 16910 4865
rect 16854 4791 16910 4800
rect 16396 4616 16448 4622
rect 16396 4558 16448 4564
rect 16212 4208 16264 4214
rect 16212 4150 16264 4156
rect 16212 4072 16264 4078
rect 16212 4014 16264 4020
rect 16118 3768 16174 3777
rect 16224 3738 16252 4014
rect 16118 3703 16174 3712
rect 16212 3732 16264 3738
rect 16212 3674 16264 3680
rect 16304 3732 16356 3738
rect 16304 3674 16356 3680
rect 16028 3664 16080 3670
rect 16028 3606 16080 3612
rect 16040 3466 16068 3606
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16120 3460 16172 3466
rect 16120 3402 16172 3408
rect 16132 3194 16160 3402
rect 16316 3398 16344 3674
rect 16304 3392 16356 3398
rect 16210 3360 16266 3369
rect 16304 3334 16356 3340
rect 16210 3295 16266 3304
rect 16120 3188 16172 3194
rect 16120 3130 16172 3136
rect 16224 2922 16252 3295
rect 16302 3224 16358 3233
rect 16302 3159 16358 3168
rect 16316 3126 16344 3159
rect 16304 3120 16356 3126
rect 16304 3062 16356 3068
rect 16212 2916 16264 2922
rect 16212 2858 16264 2864
rect 15856 2746 16068 2774
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 15936 2440 15988 2446
rect 15936 2382 15988 2388
rect 15948 2038 15976 2382
rect 15936 2032 15988 2038
rect 15936 1974 15988 1980
rect 16040 800 16068 2746
rect 16408 2582 16436 4558
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 16488 4208 16540 4214
rect 16488 4150 16540 4156
rect 16500 3777 16528 4150
rect 16672 4140 16724 4146
rect 16672 4082 16724 4088
rect 16764 4140 16816 4146
rect 16764 4082 16816 4088
rect 16486 3768 16542 3777
rect 16486 3703 16542 3712
rect 16684 3602 16712 4082
rect 16776 4049 16804 4082
rect 16762 4040 16818 4049
rect 16762 3975 16818 3984
rect 16960 3738 16988 4966
rect 16948 3732 17000 3738
rect 16948 3674 17000 3680
rect 16672 3596 16724 3602
rect 16724 3556 16988 3584
rect 16672 3538 16724 3544
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 16856 3052 16908 3058
rect 16960 3040 16988 3556
rect 16908 3012 16988 3040
rect 16856 2994 16908 3000
rect 16396 2576 16448 2582
rect 16396 2518 16448 2524
rect 17052 2310 17080 5170
rect 17132 4752 17184 4758
rect 17132 4694 17184 4700
rect 17144 4486 17172 4694
rect 17224 4684 17276 4690
rect 17224 4626 17276 4632
rect 17132 4480 17184 4486
rect 17132 4422 17184 4428
rect 17236 4146 17264 4626
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 17222 3904 17278 3913
rect 17222 3839 17278 3848
rect 17132 3732 17184 3738
rect 17132 3674 17184 3680
rect 17040 2304 17092 2310
rect 17040 2246 17092 2252
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 16580 1148 16632 1154
rect 16580 1090 16632 1096
rect 16592 800 16620 1090
rect 17144 800 17172 3674
rect 17236 3602 17264 3839
rect 17224 3596 17276 3602
rect 17224 3538 17276 3544
rect 17236 2825 17264 3538
rect 17222 2816 17278 2825
rect 17222 2751 17278 2760
rect 17328 2514 17356 13194
rect 17420 9654 17448 13806
rect 17500 13320 17552 13326
rect 17500 13262 17552 13268
rect 17512 12238 17540 13262
rect 17684 12844 17736 12850
rect 17684 12786 17736 12792
rect 17592 12640 17644 12646
rect 17592 12582 17644 12588
rect 17500 12232 17552 12238
rect 17500 12174 17552 12180
rect 17500 11824 17552 11830
rect 17500 11766 17552 11772
rect 17512 11218 17540 11766
rect 17500 11212 17552 11218
rect 17500 11154 17552 11160
rect 17498 11112 17554 11121
rect 17498 11047 17554 11056
rect 17512 11014 17540 11047
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17500 10192 17552 10198
rect 17500 10134 17552 10140
rect 17512 9674 17540 10134
rect 17604 9994 17632 12582
rect 17696 11393 17724 12786
rect 17880 12646 17908 16050
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 13938 18000 14758
rect 18052 14544 18104 14550
rect 18052 14486 18104 14492
rect 18064 14414 18092 14486
rect 18052 14408 18104 14414
rect 18052 14350 18104 14356
rect 18144 14408 18196 14414
rect 18144 14350 18196 14356
rect 18156 14074 18184 14350
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 17960 13932 18012 13938
rect 17960 13874 18012 13880
rect 17868 12640 17920 12646
rect 17868 12582 17920 12588
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17868 12164 17920 12170
rect 17868 12106 17920 12112
rect 17788 11898 17816 12106
rect 17776 11892 17828 11898
rect 17776 11834 17828 11840
rect 17776 11756 17828 11762
rect 17776 11698 17828 11704
rect 17682 11384 17738 11393
rect 17682 11319 17738 11328
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17696 10169 17724 11154
rect 17682 10160 17738 10169
rect 17682 10095 17738 10104
rect 17592 9988 17644 9994
rect 17592 9930 17644 9936
rect 17684 9716 17736 9722
rect 17408 9648 17460 9654
rect 17512 9646 17632 9674
rect 17684 9658 17736 9664
rect 17408 9590 17460 9596
rect 17500 6792 17552 6798
rect 17500 6734 17552 6740
rect 17408 6656 17460 6662
rect 17408 6598 17460 6604
rect 17420 5914 17448 6598
rect 17408 5908 17460 5914
rect 17408 5850 17460 5856
rect 17408 5636 17460 5642
rect 17408 5578 17460 5584
rect 17420 5302 17448 5578
rect 17408 5296 17460 5302
rect 17408 5238 17460 5244
rect 17420 4214 17448 5238
rect 17512 4706 17540 6734
rect 17604 6662 17632 9646
rect 17696 8514 17724 9658
rect 17788 9382 17816 11698
rect 17880 11694 17908 12106
rect 17868 11688 17920 11694
rect 17972 11665 18000 13874
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 13326 18092 13806
rect 18052 13320 18104 13326
rect 18052 13262 18104 13268
rect 17868 11630 17920 11636
rect 17958 11656 18014 11665
rect 17880 11082 17908 11630
rect 17958 11591 18014 11600
rect 17960 11552 18012 11558
rect 17960 11494 18012 11500
rect 17868 11076 17920 11082
rect 17868 11018 17920 11024
rect 17880 9994 17908 11018
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17776 9376 17828 9382
rect 17776 9318 17828 9324
rect 17880 8974 17908 9930
rect 17868 8968 17920 8974
rect 17868 8910 17920 8916
rect 17880 8566 17908 8910
rect 17972 8566 18000 11494
rect 18064 10713 18092 13262
rect 18144 12640 18196 12646
rect 18144 12582 18196 12588
rect 18156 11762 18184 12582
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18142 11384 18198 11393
rect 18142 11319 18198 11328
rect 18156 11014 18184 11319
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18050 10704 18106 10713
rect 18050 10639 18106 10648
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17868 8560 17920 8566
rect 17696 8486 17816 8514
rect 17868 8502 17920 8508
rect 17960 8560 18012 8566
rect 18064 8537 18092 9522
rect 18248 8634 18276 16526
rect 18432 12714 18460 19314
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 19536 17270 19564 19314
rect 19524 17264 19576 17270
rect 19524 17206 19576 17212
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 19628 15910 19656 22199
rect 20442 21720 20498 21729
rect 20442 21655 20498 21664
rect 19706 21312 19762 21321
rect 19706 21247 19762 21256
rect 19720 20602 19748 21247
rect 20350 20904 20406 20913
rect 20350 20839 20406 20848
rect 19708 20596 19760 20602
rect 19708 20538 19760 20544
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 19892 19780 19944 19786
rect 19892 19722 19944 19728
rect 19904 19514 19932 19722
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20088 17338 20116 17614
rect 20076 17332 20128 17338
rect 20076 17274 20128 17280
rect 19616 15904 19668 15910
rect 19616 15846 19668 15852
rect 20076 15904 20128 15910
rect 20076 15846 20128 15852
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 18972 15496 19024 15502
rect 18972 15438 19024 15444
rect 18604 14544 18656 14550
rect 18604 14486 18656 14492
rect 18512 13932 18564 13938
rect 18512 13874 18564 13880
rect 18420 12708 18472 12714
rect 18420 12650 18472 12656
rect 18328 12640 18380 12646
rect 18328 12582 18380 12588
rect 18340 11830 18368 12582
rect 18524 12434 18552 13874
rect 18616 12866 18644 14486
rect 18880 13320 18932 13326
rect 18880 13262 18932 13268
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 12986 18736 13126
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 18616 12838 18736 12866
rect 18432 12406 18552 12434
rect 18328 11824 18380 11830
rect 18328 11766 18380 11772
rect 18328 11348 18380 11354
rect 18328 11290 18380 11296
rect 18340 11257 18368 11290
rect 18326 11248 18382 11257
rect 18326 11183 18382 11192
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18340 9489 18368 10678
rect 18326 9480 18382 9489
rect 18326 9415 18382 9424
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 17960 8502 18012 8508
rect 18050 8528 18106 8537
rect 17684 8356 17736 8362
rect 17684 8298 17736 8304
rect 17696 6866 17724 8298
rect 17684 6860 17736 6866
rect 17684 6802 17736 6808
rect 17592 6656 17644 6662
rect 17644 6616 17724 6644
rect 17592 6598 17644 6604
rect 17696 6066 17724 6616
rect 17788 6202 17816 8486
rect 17880 8090 17908 8502
rect 18050 8463 18106 8472
rect 17960 8424 18012 8430
rect 17960 8366 18012 8372
rect 17868 8084 17920 8090
rect 17868 8026 17920 8032
rect 17972 6662 18000 8366
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 18052 8016 18104 8022
rect 18050 7984 18052 7993
rect 18104 7984 18106 7993
rect 18050 7919 18106 7928
rect 18052 7880 18104 7886
rect 18052 7822 18104 7828
rect 18064 6905 18092 7822
rect 18050 6896 18106 6905
rect 18050 6831 18106 6840
rect 17960 6656 18012 6662
rect 18156 6633 18184 8026
rect 18326 7984 18382 7993
rect 18326 7919 18382 7928
rect 18236 7404 18288 7410
rect 18236 7346 18288 7352
rect 18248 6866 18276 7346
rect 18340 7041 18368 7919
rect 18326 7032 18382 7041
rect 18326 6967 18382 6976
rect 18236 6860 18288 6866
rect 18236 6802 18288 6808
rect 18328 6656 18380 6662
rect 17960 6598 18012 6604
rect 18142 6624 18198 6633
rect 18328 6598 18380 6604
rect 18142 6559 18198 6568
rect 17788 6174 18000 6202
rect 17696 6038 17908 6066
rect 17776 5908 17828 5914
rect 17776 5850 17828 5856
rect 17788 5794 17816 5850
rect 17604 5766 17816 5794
rect 17604 5574 17632 5766
rect 17682 5672 17738 5681
rect 17682 5607 17738 5616
rect 17592 5568 17644 5574
rect 17592 5510 17644 5516
rect 17696 5234 17724 5607
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17684 5228 17736 5234
rect 17684 5170 17736 5176
rect 17788 5098 17816 5510
rect 17776 5092 17828 5098
rect 17776 5034 17828 5040
rect 17774 4856 17830 4865
rect 17774 4791 17830 4800
rect 17512 4678 17632 4706
rect 17498 4584 17554 4593
rect 17498 4519 17554 4528
rect 17512 4486 17540 4519
rect 17500 4480 17552 4486
rect 17500 4422 17552 4428
rect 17408 4208 17460 4214
rect 17408 4150 17460 4156
rect 17498 4040 17554 4049
rect 17498 3975 17554 3984
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17420 3534 17448 3878
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17512 3398 17540 3975
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17604 3097 17632 4678
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17590 3088 17646 3097
rect 17590 3023 17646 3032
rect 17500 2984 17552 2990
rect 17500 2926 17552 2932
rect 17512 2650 17540 2926
rect 17500 2644 17552 2650
rect 17500 2586 17552 2592
rect 17512 2514 17540 2586
rect 17316 2508 17368 2514
rect 17316 2450 17368 2456
rect 17500 2508 17552 2514
rect 17500 2450 17552 2456
rect 17696 800 17724 4218
rect 17788 2990 17816 4791
rect 17880 4049 17908 6038
rect 17866 4040 17922 4049
rect 17866 3975 17922 3984
rect 17868 3936 17920 3942
rect 17868 3878 17920 3884
rect 17880 3602 17908 3878
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17880 3126 17908 3538
rect 17868 3120 17920 3126
rect 17868 3062 17920 3068
rect 17972 3058 18000 6174
rect 18050 5808 18106 5817
rect 18050 5743 18106 5752
rect 18064 3398 18092 5743
rect 18144 5704 18196 5710
rect 18142 5672 18144 5681
rect 18196 5672 18198 5681
rect 18142 5607 18198 5616
rect 18144 5568 18196 5574
rect 18144 5510 18196 5516
rect 18156 5370 18184 5510
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18236 5296 18288 5302
rect 18234 5264 18236 5273
rect 18288 5264 18290 5273
rect 18234 5199 18290 5208
rect 18234 5128 18290 5137
rect 18234 5063 18290 5072
rect 18248 4690 18276 5063
rect 18236 4684 18288 4690
rect 18236 4626 18288 4632
rect 18248 4570 18276 4626
rect 18156 4542 18276 4570
rect 18156 4282 18184 4542
rect 18236 4480 18288 4486
rect 18236 4422 18288 4428
rect 18144 4276 18196 4282
rect 18144 4218 18196 4224
rect 18052 3392 18104 3398
rect 18052 3334 18104 3340
rect 18248 3126 18276 4422
rect 18236 3120 18288 3126
rect 18236 3062 18288 3068
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 17776 2984 17828 2990
rect 17776 2926 17828 2932
rect 18144 2916 18196 2922
rect 18144 2858 18196 2864
rect 17774 2816 17830 2825
rect 17774 2751 17830 2760
rect 17788 2582 17816 2751
rect 17776 2576 17828 2582
rect 17776 2518 17828 2524
rect 18156 1154 18184 2858
rect 18340 2774 18368 6598
rect 18432 4826 18460 12406
rect 18604 12096 18656 12102
rect 18604 12038 18656 12044
rect 18616 11286 18644 12038
rect 18604 11280 18656 11286
rect 18604 11222 18656 11228
rect 18604 10600 18656 10606
rect 18708 10577 18736 12838
rect 18788 12844 18840 12850
rect 18788 12786 18840 12792
rect 18800 12442 18828 12786
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18786 12336 18842 12345
rect 18786 12271 18842 12280
rect 18800 11286 18828 12271
rect 18788 11280 18840 11286
rect 18788 11222 18840 11228
rect 18786 10840 18842 10849
rect 18786 10775 18842 10784
rect 18800 10742 18828 10775
rect 18788 10736 18840 10742
rect 18788 10678 18840 10684
rect 18604 10542 18656 10548
rect 18694 10568 18750 10577
rect 18616 9722 18644 10542
rect 18694 10503 18750 10512
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18892 9450 18920 13262
rect 18984 12073 19012 15438
rect 19708 15360 19760 15366
rect 19708 15302 19760 15308
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19064 14952 19116 14958
rect 19064 14894 19116 14900
rect 18970 12064 19026 12073
rect 18970 11999 19026 12008
rect 18970 11792 19026 11801
rect 18970 11727 19026 11736
rect 18984 11218 19012 11727
rect 18972 11212 19024 11218
rect 18972 11154 19024 11160
rect 18984 9761 19012 11154
rect 18970 9752 19026 9761
rect 18970 9687 19026 9696
rect 18880 9444 18932 9450
rect 18880 9386 18932 9392
rect 18892 9042 18920 9386
rect 18880 9036 18932 9042
rect 18880 8978 18932 8984
rect 18604 8900 18656 8906
rect 18604 8842 18656 8848
rect 18512 8492 18564 8498
rect 18512 8434 18564 8440
rect 18524 7342 18552 8434
rect 18616 7410 18644 8842
rect 18972 8492 19024 8498
rect 18972 8434 19024 8440
rect 18880 8424 18932 8430
rect 18880 8366 18932 8372
rect 18892 7546 18920 8366
rect 18880 7540 18932 7546
rect 18880 7482 18932 7488
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18512 7336 18564 7342
rect 18512 7278 18564 7284
rect 18512 7200 18564 7206
rect 18512 7142 18564 7148
rect 18524 5273 18552 7142
rect 18788 6996 18840 7002
rect 18788 6938 18840 6944
rect 18696 5568 18748 5574
rect 18696 5510 18748 5516
rect 18510 5264 18566 5273
rect 18510 5199 18566 5208
rect 18604 5228 18656 5234
rect 18604 5170 18656 5176
rect 18420 4820 18472 4826
rect 18420 4762 18472 4768
rect 18512 4480 18564 4486
rect 18512 4422 18564 4428
rect 18420 4208 18472 4214
rect 18420 4150 18472 4156
rect 18248 2746 18368 2774
rect 18144 1148 18196 1154
rect 18144 1090 18196 1096
rect 18248 800 18276 2746
rect 18432 2514 18460 4150
rect 18524 3194 18552 4422
rect 18616 4282 18644 5170
rect 18604 4276 18656 4282
rect 18604 4218 18656 4224
rect 18616 4185 18644 4218
rect 18602 4176 18658 4185
rect 18602 4111 18658 4120
rect 18602 3768 18658 3777
rect 18602 3703 18658 3712
rect 18616 3194 18644 3703
rect 18708 3641 18736 5510
rect 18800 4321 18828 6938
rect 18892 6798 18920 7482
rect 18984 7177 19012 8434
rect 19076 7886 19104 14894
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19628 14550 19656 14962
rect 19616 14544 19668 14550
rect 19616 14486 19668 14492
rect 19720 14482 19748 15302
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19800 14816 19852 14822
rect 19800 14758 19852 14764
rect 19708 14476 19760 14482
rect 19708 14418 19760 14424
rect 19524 14408 19576 14414
rect 19576 14356 19656 14362
rect 19524 14350 19656 14356
rect 19536 14334 19656 14350
rect 19524 14272 19576 14278
rect 19524 14214 19576 14220
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19536 13394 19564 14214
rect 19524 13388 19576 13394
rect 19524 13330 19576 13336
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19536 12238 19564 12582
rect 19524 12232 19576 12238
rect 19524 12174 19576 12180
rect 19524 11756 19576 11762
rect 19524 11698 19576 11704
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19154 11248 19210 11257
rect 19154 11183 19210 11192
rect 19168 10742 19196 11183
rect 19536 10742 19564 11698
rect 19156 10736 19208 10742
rect 19156 10678 19208 10684
rect 19524 10736 19576 10742
rect 19524 10678 19576 10684
rect 19536 10470 19564 10678
rect 19524 10464 19576 10470
rect 19524 10406 19576 10412
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19536 10062 19564 10406
rect 19628 10130 19656 14334
rect 19708 13864 19760 13870
rect 19708 13806 19760 13812
rect 19720 10810 19748 13806
rect 19812 13326 19840 14758
rect 19892 14408 19944 14414
rect 19892 14350 19944 14356
rect 19800 13320 19852 13326
rect 19904 13297 19932 14350
rect 19996 13530 20024 14962
rect 20088 14278 20116 15846
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 20076 13864 20128 13870
rect 20076 13806 20128 13812
rect 19984 13524 20036 13530
rect 19984 13466 20036 13472
rect 19800 13262 19852 13268
rect 19890 13288 19946 13297
rect 19890 13223 19946 13232
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19800 12164 19852 12170
rect 19800 12106 19852 12112
rect 19708 10804 19760 10810
rect 19708 10746 19760 10752
rect 19708 10464 19760 10470
rect 19708 10406 19760 10412
rect 19616 10124 19668 10130
rect 19616 10066 19668 10072
rect 19524 10056 19576 10062
rect 19524 9998 19576 10004
rect 19524 9920 19576 9926
rect 19524 9862 19576 9868
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19536 9110 19564 9862
rect 19720 9654 19748 10406
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19812 9330 19840 12106
rect 19720 9302 19840 9330
rect 19524 9104 19576 9110
rect 19524 9046 19576 9052
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19536 8498 19564 8910
rect 19720 8634 19748 9302
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 18970 7168 19026 7177
rect 18970 7103 19026 7112
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19352 6390 19380 6734
rect 19340 6384 19392 6390
rect 19340 6326 19392 6332
rect 19524 6316 19576 6322
rect 19524 6258 19576 6264
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 18970 5944 19026 5953
rect 19143 5936 19451 5956
rect 19026 5902 19104 5930
rect 18970 5879 19026 5888
rect 18892 5846 18920 5877
rect 18880 5840 18932 5846
rect 18878 5808 18880 5817
rect 18932 5808 18934 5817
rect 18878 5743 18934 5752
rect 18892 5710 18920 5743
rect 18880 5704 18932 5710
rect 18880 5646 18932 5652
rect 18972 4752 19024 4758
rect 18972 4694 19024 4700
rect 18880 4548 18932 4554
rect 18880 4490 18932 4496
rect 18786 4312 18842 4321
rect 18786 4247 18842 4256
rect 18892 4049 18920 4490
rect 18984 4146 19012 4694
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18878 4040 18934 4049
rect 18878 3975 18934 3984
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18694 3632 18750 3641
rect 18694 3567 18750 3576
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 18604 3188 18656 3194
rect 18604 3130 18656 3136
rect 18420 2508 18472 2514
rect 18420 2450 18472 2456
rect 18420 2372 18472 2378
rect 18420 2314 18472 2320
rect 18432 1873 18460 2314
rect 18418 1864 18474 1873
rect 18418 1799 18474 1808
rect 18800 800 18828 3878
rect 18892 3126 18920 3975
rect 18880 3120 18932 3126
rect 18880 3062 18932 3068
rect 18984 2990 19012 4082
rect 19076 3618 19104 5902
rect 19536 5166 19564 6258
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 19536 4690 19564 5102
rect 19524 4684 19576 4690
rect 19524 4626 19576 4632
rect 19628 4570 19656 8570
rect 19812 7698 19840 9114
rect 19904 8906 19932 13126
rect 19984 11552 20036 11558
rect 19984 11494 20036 11500
rect 19996 10810 20024 11494
rect 20088 11234 20116 13806
rect 20180 11370 20208 20198
rect 20364 20058 20392 20839
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20456 19446 20484 21655
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 21088 20460 21140 20466
rect 21088 20402 21140 20408
rect 20444 19440 20496 19446
rect 20444 19382 20496 19388
rect 20548 18970 20576 20402
rect 20810 20360 20866 20369
rect 20810 20295 20866 20304
rect 20720 20256 20772 20262
rect 20720 20198 20772 20204
rect 20732 19961 20760 20198
rect 20824 20058 20852 20295
rect 20812 20052 20864 20058
rect 20812 19994 20864 20000
rect 20718 19952 20774 19961
rect 20718 19887 20774 19896
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20628 19508 20680 19514
rect 20628 19450 20680 19456
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20260 18760 20312 18766
rect 20260 18702 20312 18708
rect 20272 18086 20300 18702
rect 20640 18601 20668 19450
rect 20720 19372 20772 19378
rect 20720 19314 20772 19320
rect 20626 18592 20682 18601
rect 20626 18527 20682 18536
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20536 18080 20588 18086
rect 20536 18022 20588 18028
rect 20548 17678 20576 18022
rect 20732 17882 20760 19314
rect 20824 18426 20852 19790
rect 21100 18970 21128 20402
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21272 19712 21324 19718
rect 21272 19654 21324 19660
rect 21284 19009 21312 19654
rect 21376 19417 21404 20198
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21270 19000 21326 19009
rect 21088 18964 21140 18970
rect 21270 18935 21326 18944
rect 21088 18906 21140 18912
rect 20996 18760 21048 18766
rect 20996 18702 21048 18708
rect 20812 18420 20864 18426
rect 20812 18362 20864 18368
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20904 18284 20956 18290
rect 20904 18226 20956 18232
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20718 17640 20774 17649
rect 20718 17575 20774 17584
rect 20732 17542 20760 17575
rect 20720 17536 20772 17542
rect 20720 17478 20772 17484
rect 20824 17354 20852 18226
rect 20732 17326 20852 17354
rect 20916 17338 20944 18226
rect 20904 17332 20956 17338
rect 20732 16266 20760 17326
rect 20904 17274 20956 17280
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20640 16250 20760 16266
rect 20824 16250 20852 17138
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 20628 16244 20760 16250
rect 20680 16238 20760 16244
rect 20812 16244 20864 16250
rect 20628 16186 20680 16192
rect 20812 16186 20864 16192
rect 20352 15496 20404 15502
rect 20352 15438 20404 15444
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20272 11898 20300 15302
rect 20364 14074 20392 15438
rect 20732 15162 20760 15438
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20640 14618 20668 14962
rect 20916 14890 20944 16526
rect 21008 16454 21036 18702
rect 21272 18624 21324 18630
rect 21272 18566 21324 18572
rect 21284 18057 21312 18566
rect 21364 18080 21416 18086
rect 21270 18048 21326 18057
rect 21364 18022 21416 18028
rect 21270 17983 21326 17992
rect 21088 17672 21140 17678
rect 21088 17614 21140 17620
rect 21100 16794 21128 17614
rect 21272 17536 21324 17542
rect 21272 17478 21324 17484
rect 21088 16788 21140 16794
rect 21088 16730 21140 16736
rect 21284 16697 21312 17478
rect 21376 17241 21404 18022
rect 21362 17232 21418 17241
rect 21362 17167 21418 17176
rect 21364 16992 21416 16998
rect 21364 16934 21416 16940
rect 21270 16688 21326 16697
rect 21270 16623 21326 16632
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21272 16448 21324 16454
rect 21272 16390 21324 16396
rect 21088 16108 21140 16114
rect 21088 16050 21140 16056
rect 21100 15706 21128 16050
rect 21284 15745 21312 16390
rect 21376 16289 21404 16934
rect 21362 16280 21418 16289
rect 21362 16215 21418 16224
rect 21364 15904 21416 15910
rect 21364 15846 21416 15852
rect 21270 15736 21326 15745
rect 21088 15700 21140 15706
rect 21270 15671 21326 15680
rect 21088 15642 21140 15648
rect 21088 15360 21140 15366
rect 21088 15302 21140 15308
rect 21272 15360 21324 15366
rect 21376 15337 21404 15846
rect 21272 15302 21324 15308
rect 21362 15328 21418 15337
rect 20904 14884 20956 14890
rect 20904 14826 20956 14832
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20444 14408 20496 14414
rect 20444 14350 20496 14356
rect 20352 14068 20404 14074
rect 20352 14010 20404 14016
rect 20350 13560 20406 13569
rect 20350 13495 20352 13504
rect 20404 13495 20406 13504
rect 20352 13466 20404 13472
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20260 11892 20312 11898
rect 20260 11834 20312 11840
rect 20364 11626 20392 12786
rect 20352 11620 20404 11626
rect 20352 11562 20404 11568
rect 20180 11342 20300 11370
rect 20088 11206 20208 11234
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19984 10804 20036 10810
rect 19984 10746 20036 10752
rect 20088 10538 20116 11086
rect 20076 10532 20128 10538
rect 20076 10474 20128 10480
rect 20088 9518 20116 10474
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 20088 8974 20116 9454
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 20076 8832 20128 8838
rect 20076 8774 20128 8780
rect 19812 7670 20024 7698
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19800 7200 19852 7206
rect 19800 7142 19852 7148
rect 19708 5228 19760 5234
rect 19708 5170 19760 5176
rect 19536 4542 19656 4570
rect 19536 3942 19564 4542
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 19076 3590 19380 3618
rect 19062 3360 19118 3369
rect 19062 3295 19118 3304
rect 18972 2984 19024 2990
rect 18972 2926 19024 2932
rect 18880 2440 18932 2446
rect 18878 2408 18880 2417
rect 18932 2408 18934 2417
rect 18878 2343 18934 2352
rect 18892 2009 18920 2343
rect 18878 2000 18934 2009
rect 18878 1935 18934 1944
rect 19076 1737 19104 3295
rect 19352 3194 19380 3590
rect 19524 3528 19576 3534
rect 19524 3470 19576 3476
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 19432 2984 19484 2990
rect 19430 2952 19432 2961
rect 19484 2952 19486 2961
rect 19430 2887 19486 2896
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 19432 2440 19484 2446
rect 19432 2382 19484 2388
rect 19340 1828 19392 1834
rect 19340 1770 19392 1776
rect 19062 1728 19118 1737
rect 19062 1663 19118 1672
rect 19352 800 19380 1770
rect 19444 1358 19472 2382
rect 19536 1601 19564 3470
rect 19628 2514 19656 4422
rect 19720 3754 19748 5170
rect 19812 4622 19840 7142
rect 19904 5370 19932 7482
rect 19892 5364 19944 5370
rect 19892 5306 19944 5312
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19720 3726 19840 3754
rect 19708 3528 19760 3534
rect 19708 3470 19760 3476
rect 19720 2650 19748 3470
rect 19812 3058 19840 3726
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19798 2952 19854 2961
rect 19798 2887 19854 2896
rect 19708 2644 19760 2650
rect 19708 2586 19760 2592
rect 19616 2508 19668 2514
rect 19616 2450 19668 2456
rect 19522 1592 19578 1601
rect 19522 1527 19578 1536
rect 19536 1426 19564 1527
rect 19524 1420 19576 1426
rect 19524 1362 19576 1368
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 202 0 258 800
rect 662 0 718 800
rect 1214 0 1270 800
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12162 0 12218 800
rect 12714 0 12770 800
rect 13266 0 13322 800
rect 13818 0 13874 800
rect 14370 0 14426 800
rect 14922 0 14978 800
rect 15474 0 15530 800
rect 16026 0 16082 800
rect 16578 0 16634 800
rect 17130 0 17186 800
rect 17682 0 17738 800
rect 18234 0 18290 800
rect 18786 0 18842 800
rect 19338 0 19394 800
rect 19444 241 19472 1294
rect 19812 1057 19840 2887
rect 19798 1048 19854 1057
rect 19798 983 19854 992
rect 19904 800 19932 3878
rect 19430 232 19486 241
rect 19430 167 19486 176
rect 19890 0 19946 800
rect 19996 762 20024 7670
rect 20088 7546 20116 8774
rect 20076 7540 20128 7546
rect 20076 7482 20128 7488
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20088 6610 20116 7346
rect 20180 6730 20208 11206
rect 20272 8838 20300 11342
rect 20352 10668 20404 10674
rect 20352 10610 20404 10616
rect 20364 10266 20392 10610
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20364 9586 20392 10066
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20350 8936 20406 8945
rect 20350 8871 20406 8880
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20272 7954 20300 8570
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20364 6882 20392 8871
rect 20272 6854 20392 6882
rect 20168 6724 20220 6730
rect 20168 6666 20220 6672
rect 20088 6582 20208 6610
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 20088 4690 20116 4966
rect 20076 4684 20128 4690
rect 20076 4626 20128 4632
rect 20180 4282 20208 6582
rect 20272 5250 20300 6854
rect 20350 6760 20406 6769
rect 20350 6695 20406 6704
rect 20364 6458 20392 6695
rect 20352 6452 20404 6458
rect 20352 6394 20404 6400
rect 20456 5370 20484 14350
rect 20548 12617 20576 14486
rect 21100 14414 21128 15302
rect 21284 14929 21312 15302
rect 21362 15263 21418 15272
rect 21270 14920 21326 14929
rect 21270 14855 21326 14864
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 21088 14408 21140 14414
rect 21284 14385 21312 14758
rect 21088 14350 21140 14356
rect 21270 14376 21326 14385
rect 20996 14340 21048 14346
rect 21270 14311 21326 14320
rect 20996 14282 21048 14288
rect 20628 14272 20680 14278
rect 20628 14214 20680 14220
rect 20640 13938 20668 14214
rect 20628 13932 20680 13938
rect 20628 13874 20680 13880
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20534 12608 20590 12617
rect 20534 12543 20590 12552
rect 20640 12102 20668 12786
rect 20732 12434 20760 13262
rect 20904 12640 20956 12646
rect 20904 12582 20956 12588
rect 20732 12406 20852 12434
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20640 10606 20668 12038
rect 20720 11076 20772 11082
rect 20720 11018 20772 11024
rect 20732 10810 20760 11018
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20628 10600 20680 10606
rect 20628 10542 20680 10548
rect 20718 10024 20774 10033
rect 20718 9959 20774 9968
rect 20732 9042 20760 9959
rect 20824 9178 20852 12406
rect 20916 11082 20944 12582
rect 21008 12238 21036 14282
rect 21272 14272 21324 14278
rect 21272 14214 21324 14220
rect 21284 13977 21312 14214
rect 21270 13968 21326 13977
rect 21270 13903 21326 13912
rect 21640 13864 21692 13870
rect 21640 13806 21692 13812
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 20904 11076 20956 11082
rect 20904 11018 20956 11024
rect 20904 10668 20956 10674
rect 20904 10610 20956 10616
rect 20916 9382 20944 10610
rect 21008 10606 21036 11290
rect 20996 10600 21048 10606
rect 20996 10542 21048 10548
rect 21008 10062 21036 10542
rect 20996 10056 21048 10062
rect 20996 9998 21048 10004
rect 20904 9376 20956 9382
rect 20904 9318 20956 9324
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20720 9036 20772 9042
rect 20720 8978 20772 8984
rect 20720 8288 20772 8294
rect 20720 8230 20772 8236
rect 20732 7886 20760 8230
rect 20720 7880 20772 7886
rect 20720 7822 20772 7828
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7546 20576 7686
rect 20536 7540 20588 7546
rect 20536 7482 20588 7488
rect 20824 7342 20852 9114
rect 20916 7546 20944 9318
rect 21100 8566 21128 13126
rect 21270 13016 21326 13025
rect 21270 12951 21326 12960
rect 21284 12442 21312 12951
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21456 11552 21508 11558
rect 21456 11494 21508 11500
rect 21364 9920 21416 9926
rect 21364 9862 21416 9868
rect 21376 8945 21404 9862
rect 21362 8936 21418 8945
rect 21362 8871 21418 8880
rect 21180 8832 21232 8838
rect 21180 8774 21232 8780
rect 21088 8560 21140 8566
rect 21088 8502 21140 8508
rect 21192 8265 21220 8774
rect 21178 8256 21234 8265
rect 21178 8191 21234 8200
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 20904 7540 20956 7546
rect 20904 7482 20956 7488
rect 21376 7478 21404 7686
rect 21364 7472 21416 7478
rect 20994 7440 21050 7449
rect 21364 7414 21416 7420
rect 20994 7375 20996 7384
rect 21048 7375 21050 7384
rect 20996 7346 21048 7352
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 21272 7268 21324 7274
rect 21272 7210 21324 7216
rect 20536 6792 20588 6798
rect 20536 6734 20588 6740
rect 20548 5710 20576 6734
rect 21284 6662 21312 7210
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20548 5250 20576 5646
rect 20272 5222 20392 5250
rect 20260 5160 20312 5166
rect 20260 5102 20312 5108
rect 20168 4276 20220 4282
rect 20168 4218 20220 4224
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 20088 1834 20116 3130
rect 20272 2854 20300 5102
rect 20364 3534 20392 5222
rect 20456 5222 20576 5250
rect 20456 4706 20484 5222
rect 20536 5160 20588 5166
rect 20536 5102 20588 5108
rect 20548 4826 20576 5102
rect 20536 4820 20588 4826
rect 20536 4762 20588 4768
rect 20456 4678 20576 4706
rect 20444 4276 20496 4282
rect 20444 4218 20496 4224
rect 20456 3602 20484 4218
rect 20548 4146 20576 4678
rect 20536 4140 20588 4146
rect 20536 4082 20588 4088
rect 20640 3738 20668 6394
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 20902 6352 20958 6361
rect 20628 3732 20680 3738
rect 20628 3674 20680 3680
rect 20444 3596 20496 3602
rect 20444 3538 20496 3544
rect 20352 3528 20404 3534
rect 20352 3470 20404 3476
rect 20628 3528 20680 3534
rect 20628 3470 20680 3476
rect 20536 3392 20588 3398
rect 20536 3334 20588 3340
rect 20548 3058 20576 3334
rect 20536 3052 20588 3058
rect 20536 2994 20588 3000
rect 20548 2961 20576 2994
rect 20534 2952 20590 2961
rect 20534 2887 20590 2896
rect 20260 2848 20312 2854
rect 20260 2790 20312 2796
rect 20272 2514 20300 2790
rect 20260 2508 20312 2514
rect 20260 2450 20312 2456
rect 20536 2440 20588 2446
rect 20534 2408 20536 2417
rect 20588 2408 20590 2417
rect 20534 2343 20590 2352
rect 20076 1828 20128 1834
rect 20076 1770 20128 1776
rect 20640 921 20668 3470
rect 20626 912 20682 921
rect 20364 870 20484 898
rect 20364 762 20392 870
rect 20456 800 20484 870
rect 20626 847 20682 856
rect 19996 734 20392 762
rect 20442 0 20498 800
rect 20732 762 20760 6326
rect 20902 6287 20958 6296
rect 21088 6316 21140 6322
rect 20812 6112 20864 6118
rect 20812 6054 20864 6060
rect 20824 5370 20852 6054
rect 20916 5710 20944 6287
rect 21088 6258 21140 6264
rect 21100 6225 21128 6258
rect 21086 6216 21142 6225
rect 21086 6151 21142 6160
rect 21180 6180 21232 6186
rect 21180 6122 21232 6128
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20904 5704 20956 5710
rect 20904 5646 20956 5652
rect 20812 5364 20864 5370
rect 20812 5306 20864 5312
rect 21008 5166 21036 5850
rect 21192 5642 21220 6122
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20996 5160 21048 5166
rect 20996 5102 21048 5108
rect 21100 2922 21128 5510
rect 21192 4690 21220 5578
rect 21180 4684 21232 4690
rect 21180 4626 21232 4632
rect 21284 4214 21312 6598
rect 21272 4208 21324 4214
rect 21272 4150 21324 4156
rect 21468 3942 21496 11494
rect 21548 7812 21600 7818
rect 21548 7754 21600 7760
rect 21456 3936 21508 3942
rect 21456 3878 21508 3884
rect 21088 2916 21140 2922
rect 21088 2858 21140 2864
rect 20916 870 21036 898
rect 20916 762 20944 870
rect 21008 800 21036 870
rect 21560 800 21588 7754
rect 21652 5914 21680 13806
rect 21732 8968 21784 8974
rect 21732 8910 21784 8916
rect 21640 5908 21692 5914
rect 21640 5850 21692 5856
rect 21744 4729 21772 8910
rect 22652 5840 22704 5846
rect 22652 5782 22704 5788
rect 21730 4720 21786 4729
rect 21730 4655 21786 4664
rect 22100 2100 22152 2106
rect 22100 2042 22152 2048
rect 22112 800 22140 2042
rect 22664 800 22692 5782
rect 20732 734 20944 762
rect 20994 0 21050 800
rect 21546 0 21602 800
rect 22098 0 22154 800
rect 22650 0 22706 800
<< via2 >>
rect 19246 22616 19302 22672
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 19614 22208 19670 22264
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 6550 17176 6606 17232
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 4986 12280 5042 12336
rect 1490 11500 1492 11520
rect 1492 11500 1544 11520
rect 1544 11500 1546 11520
rect 1490 11464 1546 11500
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3974 9016 4030 9072
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 2042 7384 2098 7440
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 2134 1808 2190 1864
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3698 2916 3754 2952
rect 3698 2896 3700 2916
rect 3700 2896 3752 2916
rect 3752 2896 3754 2916
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 2962 2352 3018 2408
rect 4618 3984 4674 4040
rect 4618 3032 4674 3088
rect 4618 2760 4674 2816
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 4802 2760 4858 2816
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 5354 6840 5410 6896
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 5630 8880 5686 8936
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6274 6724 6330 6760
rect 6274 6704 6276 6724
rect 6276 6704 6328 6724
rect 6328 6704 6330 6724
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 5998 5752 6054 5808
rect 5722 4664 5778 4720
rect 5538 4120 5594 4176
rect 4710 1672 4766 1728
rect 5538 1944 5594 2000
rect 5446 1536 5502 1592
rect 6550 5616 6606 5672
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6458 5244 6460 5264
rect 6460 5244 6512 5264
rect 6512 5244 6514 5264
rect 6458 5208 6514 5244
rect 7010 8336 7066 8392
rect 6918 7812 6974 7848
rect 6918 7792 6920 7812
rect 6920 7792 6972 7812
rect 6972 7792 6974 7812
rect 7010 6180 7066 6216
rect 7010 6160 7012 6180
rect 7012 6160 7064 6180
rect 7064 6160 7066 6180
rect 6550 5072 6606 5128
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6550 3576 6606 3632
rect 5814 2624 5870 2680
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6642 3440 6698 3496
rect 7102 4548 7158 4584
rect 7102 4528 7104 4548
rect 7104 4528 7156 4548
rect 7156 4528 7158 4548
rect 7010 3984 7066 4040
rect 7470 7928 7526 7984
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6826 2624 6882 2680
rect 6642 2488 6698 2544
rect 6826 2216 6882 2272
rect 8022 7268 8078 7304
rect 8022 7248 8024 7268
rect 8024 7248 8076 7268
rect 8076 7248 8078 7268
rect 7838 6432 7894 6488
rect 8114 4528 8170 4584
rect 7654 3712 7710 3768
rect 7562 3168 7618 3224
rect 8022 3712 8078 3768
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8390 2760 8446 2816
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 10230 10104 10286 10160
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 9632 7486 9688 7542
rect 9218 7384 9274 7440
rect 9126 6296 9182 6352
rect 9126 6024 9182 6080
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 9770 7112 9826 7168
rect 9586 6432 9642 6488
rect 9494 6296 9550 6352
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9126 3032 9182 3088
rect 9494 3052 9550 3088
rect 9494 3032 9496 3052
rect 9496 3032 9548 3052
rect 9548 3032 9550 3052
rect 9126 2760 9182 2816
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 8942 2488 8998 2544
rect 10414 9152 10470 9208
rect 10506 7520 10562 7576
rect 10414 5208 10470 5264
rect 10598 3168 10654 3224
rect 10966 7404 11022 7440
rect 10966 7384 10968 7404
rect 10968 7384 11020 7404
rect 11020 7384 11022 7404
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11886 9560 11942 9616
rect 11886 9288 11942 9344
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11794 6432 11850 6488
rect 11794 6024 11850 6080
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11978 9152 12034 9208
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 11794 3476 11796 3496
rect 11796 3476 11848 3496
rect 11848 3476 11850 3496
rect 11794 3440 11850 3476
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 10874 1536 10930 1592
rect 12530 3304 12586 3360
rect 12070 1944 12126 2000
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13266 9968 13322 10024
rect 14186 11736 14242 11792
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 14370 11056 14426 11112
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 14370 7112 14426 7168
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 14186 5244 14188 5264
rect 14188 5244 14240 5264
rect 14240 5244 14242 5264
rect 14186 5208 14242 5244
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 13726 2760 13782 2816
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 15290 13232 15346 13288
rect 15290 8336 15346 8392
rect 15290 6840 15346 6896
rect 14462 3168 14518 3224
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14830 5244 14832 5264
rect 14832 5244 14884 5264
rect 14884 5244 14886 5264
rect 14830 5208 14886 5244
rect 15106 5752 15162 5808
rect 15290 6432 15346 6488
rect 15750 5888 15806 5944
rect 15382 4120 15438 4176
rect 15198 3576 15254 3632
rect 14646 2488 14702 2544
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 15934 3848 15990 3904
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16670 11192 16726 11248
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16946 10784 17002 10840
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16394 8200 16450 8256
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16394 7520 16450 7576
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 16854 4800 16910 4856
rect 16118 3712 16174 3768
rect 16210 3304 16266 3360
rect 16302 3168 16358 3224
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 16486 3712 16542 3768
rect 16762 3984 16818 4040
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 17222 3848 17278 3904
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17222 2760 17278 2816
rect 17498 11056 17554 11112
rect 17682 11328 17738 11384
rect 17682 10104 17738 10160
rect 17958 11600 18014 11656
rect 18142 11328 18198 11384
rect 18050 10648 18106 10704
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 20442 21664 20498 21720
rect 19706 21256 19762 21312
rect 20350 20848 20406 20904
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 18326 11192 18382 11248
rect 18326 9424 18382 9480
rect 18050 8472 18106 8528
rect 18050 7964 18052 7984
rect 18052 7964 18104 7984
rect 18104 7964 18106 7984
rect 18050 7928 18106 7964
rect 18050 6840 18106 6896
rect 18326 7928 18382 7984
rect 18326 6976 18382 7032
rect 18142 6568 18198 6624
rect 17682 5616 17738 5672
rect 17774 4800 17830 4856
rect 17498 4528 17554 4584
rect 17498 3984 17554 4040
rect 17590 3032 17646 3088
rect 17866 3984 17922 4040
rect 18050 5752 18106 5808
rect 18142 5652 18144 5672
rect 18144 5652 18196 5672
rect 18196 5652 18198 5672
rect 18142 5616 18198 5652
rect 18234 5244 18236 5264
rect 18236 5244 18288 5264
rect 18288 5244 18290 5264
rect 18234 5208 18290 5244
rect 18234 5072 18290 5128
rect 17774 2760 17830 2816
rect 18786 12280 18842 12336
rect 18786 10784 18842 10840
rect 18694 10512 18750 10568
rect 18970 12008 19026 12064
rect 18970 11736 19026 11792
rect 18970 9696 19026 9752
rect 18510 5208 18566 5264
rect 18602 4120 18658 4176
rect 18602 3712 18658 3768
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19154 11192 19210 11248
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19890 13232 19946 13288
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 18970 7112 19026 7168
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 18970 5888 19026 5944
rect 18878 5788 18880 5808
rect 18880 5788 18932 5808
rect 18932 5788 18934 5808
rect 18878 5752 18934 5788
rect 18786 4256 18842 4312
rect 18878 3984 18934 4040
rect 18694 3576 18750 3632
rect 18418 1808 18474 1864
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 20810 20304 20866 20360
rect 20718 19896 20774 19952
rect 20626 18536 20682 18592
rect 21362 19352 21418 19408
rect 21270 18944 21326 19000
rect 20718 17584 20774 17640
rect 21270 17992 21326 18048
rect 21362 17176 21418 17232
rect 21270 16632 21326 16688
rect 21362 16224 21418 16280
rect 21270 15680 21326 15736
rect 20350 13524 20406 13560
rect 20350 13504 20352 13524
rect 20352 13504 20404 13524
rect 20404 13504 20406 13524
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 19062 3304 19118 3360
rect 18878 2388 18880 2408
rect 18880 2388 18932 2408
rect 18932 2388 18934 2408
rect 18878 2352 18934 2388
rect 18878 1944 18934 2000
rect 19430 2932 19432 2952
rect 19432 2932 19484 2952
rect 19484 2932 19486 2952
rect 19430 2896 19486 2932
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19062 1672 19118 1728
rect 19798 2896 19854 2952
rect 19522 1536 19578 1592
rect 19798 992 19854 1048
rect 19430 176 19486 232
rect 20350 8880 20406 8936
rect 20350 6704 20406 6760
rect 21362 15272 21418 15328
rect 21270 14864 21326 14920
rect 21270 14320 21326 14376
rect 20534 12552 20590 12608
rect 20718 9968 20774 10024
rect 21270 13912 21326 13968
rect 21270 12960 21326 13016
rect 21362 8880 21418 8936
rect 21178 8200 21234 8256
rect 20994 7404 21050 7440
rect 20994 7384 20996 7404
rect 20996 7384 21048 7404
rect 21048 7384 21050 7404
rect 20534 2896 20590 2952
rect 20534 2388 20536 2408
rect 20536 2388 20588 2408
rect 20588 2388 20590 2408
rect 20534 2352 20590 2388
rect 20626 856 20682 912
rect 20902 6296 20958 6352
rect 21086 6160 21142 6216
rect 21730 4664 21786 4720
<< metal3 >>
rect 19241 22674 19307 22677
rect 22200 22674 23000 22704
rect 19241 22672 23000 22674
rect 19241 22616 19246 22672
rect 19302 22616 23000 22672
rect 19241 22614 23000 22616
rect 19241 22611 19307 22614
rect 22200 22584 23000 22614
rect 19609 22266 19675 22269
rect 22200 22266 23000 22296
rect 19609 22264 23000 22266
rect 19609 22208 19614 22264
rect 19670 22208 23000 22264
rect 19609 22206 23000 22208
rect 19609 22203 19675 22206
rect 22200 22176 23000 22206
rect 20437 21722 20503 21725
rect 22200 21722 23000 21752
rect 20437 21720 23000 21722
rect 20437 21664 20442 21720
rect 20498 21664 23000 21720
rect 20437 21662 23000 21664
rect 20437 21659 20503 21662
rect 22200 21632 23000 21662
rect 19701 21314 19767 21317
rect 22200 21314 23000 21344
rect 19701 21312 23000 21314
rect 19701 21256 19706 21312
rect 19762 21256 23000 21312
rect 19701 21254 23000 21256
rect 19701 21251 19767 21254
rect 22200 21224 23000 21254
rect 20345 20906 20411 20909
rect 22200 20906 23000 20936
rect 20345 20904 23000 20906
rect 20345 20848 20350 20904
rect 20406 20848 23000 20904
rect 20345 20846 23000 20848
rect 20345 20843 20411 20846
rect 22200 20816 23000 20846
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 20639 16858 20640
rect 20805 20362 20871 20365
rect 22200 20362 23000 20392
rect 20805 20360 23000 20362
rect 20805 20304 20810 20360
rect 20866 20304 23000 20360
rect 20805 20302 23000 20304
rect 20805 20299 20871 20302
rect 22200 20272 23000 20302
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 20713 19954 20779 19957
rect 22200 19954 23000 19984
rect 20713 19952 23000 19954
rect 20713 19896 20718 19952
rect 20774 19896 23000 19952
rect 20713 19894 23000 19896
rect 20713 19891 20779 19894
rect 22200 19864 23000 19894
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 21357 19410 21423 19413
rect 22200 19410 23000 19440
rect 21357 19408 23000 19410
rect 21357 19352 21362 19408
rect 21418 19352 23000 19408
rect 21357 19350 23000 19352
rect 21357 19347 21423 19350
rect 22200 19320 23000 19350
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 21265 19002 21331 19005
rect 22200 19002 23000 19032
rect 21265 19000 23000 19002
rect 21265 18944 21270 19000
rect 21326 18944 23000 19000
rect 21265 18942 23000 18944
rect 21265 18939 21331 18942
rect 22200 18912 23000 18942
rect 20621 18594 20687 18597
rect 22200 18594 23000 18624
rect 20621 18592 23000 18594
rect 20621 18536 20626 18592
rect 20682 18536 23000 18592
rect 20621 18534 23000 18536
rect 20621 18531 20687 18534
rect 6142 18528 6462 18529
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 22200 18504 23000 18534
rect 16538 18463 16858 18464
rect 21265 18050 21331 18053
rect 22200 18050 23000 18080
rect 21265 18048 23000 18050
rect 21265 17992 21270 18048
rect 21326 17992 23000 18048
rect 21265 17990 23000 17992
rect 21265 17987 21331 17990
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 22200 17960 23000 17990
rect 19137 17919 19457 17920
rect 20713 17642 20779 17645
rect 22200 17642 23000 17672
rect 20713 17640 23000 17642
rect 20713 17584 20718 17640
rect 20774 17584 23000 17640
rect 20713 17582 23000 17584
rect 20713 17579 20779 17582
rect 22200 17552 23000 17582
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 17375 16858 17376
rect 6545 17234 6611 17237
rect 14958 17234 14964 17236
rect 6545 17232 14964 17234
rect 6545 17176 6550 17232
rect 6606 17176 14964 17232
rect 6545 17174 14964 17176
rect 6545 17171 6611 17174
rect 14958 17172 14964 17174
rect 15028 17172 15034 17236
rect 21357 17234 21423 17237
rect 22200 17234 23000 17264
rect 21357 17232 23000 17234
rect 21357 17176 21362 17232
rect 21418 17176 23000 17232
rect 21357 17174 23000 17176
rect 21357 17171 21423 17174
rect 22200 17144 23000 17174
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 21265 16690 21331 16693
rect 22200 16690 23000 16720
rect 21265 16688 23000 16690
rect 21265 16632 21270 16688
rect 21326 16632 23000 16688
rect 21265 16630 23000 16632
rect 21265 16627 21331 16630
rect 22200 16600 23000 16630
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 21357 16282 21423 16285
rect 22200 16282 23000 16312
rect 21357 16280 23000 16282
rect 21357 16224 21362 16280
rect 21418 16224 23000 16280
rect 21357 16222 23000 16224
rect 21357 16219 21423 16222
rect 22200 16192 23000 16222
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 21265 15738 21331 15741
rect 22200 15738 23000 15768
rect 21265 15736 23000 15738
rect 21265 15680 21270 15736
rect 21326 15680 23000 15736
rect 21265 15678 23000 15680
rect 21265 15675 21331 15678
rect 22200 15648 23000 15678
rect 21357 15330 21423 15333
rect 22200 15330 23000 15360
rect 21357 15328 23000 15330
rect 21357 15272 21362 15328
rect 21418 15272 23000 15328
rect 21357 15270 23000 15272
rect 21357 15267 21423 15270
rect 6142 15264 6462 15265
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 22200 15240 23000 15270
rect 16538 15199 16858 15200
rect 21265 14922 21331 14925
rect 22200 14922 23000 14952
rect 21265 14920 23000 14922
rect 21265 14864 21270 14920
rect 21326 14864 23000 14920
rect 21265 14862 23000 14864
rect 21265 14859 21331 14862
rect 22200 14832 23000 14862
rect 3543 14720 3863 14721
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 21265 14378 21331 14381
rect 22200 14378 23000 14408
rect 21265 14376 23000 14378
rect 21265 14320 21270 14376
rect 21326 14320 23000 14376
rect 21265 14318 23000 14320
rect 21265 14315 21331 14318
rect 22200 14288 23000 14318
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 14111 16858 14112
rect 21265 13970 21331 13973
rect 22200 13970 23000 14000
rect 21265 13968 23000 13970
rect 21265 13912 21270 13968
rect 21326 13912 23000 13968
rect 21265 13910 23000 13912
rect 21265 13907 21331 13910
rect 22200 13880 23000 13910
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 20345 13562 20411 13565
rect 22200 13562 23000 13592
rect 20345 13560 23000 13562
rect 20345 13504 20350 13560
rect 20406 13504 23000 13560
rect 20345 13502 23000 13504
rect 20345 13499 20411 13502
rect 22200 13472 23000 13502
rect 15285 13290 15351 13293
rect 19885 13290 19951 13293
rect 15285 13288 19951 13290
rect 15285 13232 15290 13288
rect 15346 13232 19890 13288
rect 19946 13232 19951 13288
rect 15285 13230 19951 13232
rect 15285 13227 15351 13230
rect 19885 13227 19951 13230
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 21265 13018 21331 13021
rect 22200 13018 23000 13048
rect 21265 13016 23000 13018
rect 21265 12960 21270 13016
rect 21326 12960 23000 13016
rect 21265 12958 23000 12960
rect 21265 12955 21331 12958
rect 22200 12928 23000 12958
rect 20529 12610 20595 12613
rect 22200 12610 23000 12640
rect 20529 12608 23000 12610
rect 20529 12552 20534 12608
rect 20590 12552 23000 12608
rect 20529 12550 23000 12552
rect 20529 12547 20595 12550
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 22200 12520 23000 12550
rect 19137 12479 19457 12480
rect 4981 12338 5047 12341
rect 18781 12338 18847 12341
rect 4981 12336 18847 12338
rect 4981 12280 4986 12336
rect 5042 12280 18786 12336
rect 18842 12280 18847 12336
rect 4981 12278 18847 12280
rect 4981 12275 5047 12278
rect 18781 12275 18847 12278
rect 18965 12066 19031 12069
rect 22200 12066 23000 12096
rect 18965 12064 23000 12066
rect 18965 12008 18970 12064
rect 19026 12008 23000 12064
rect 18965 12006 23000 12008
rect 18965 12003 19031 12006
rect 6142 12000 6462 12001
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 22200 11976 23000 12006
rect 16538 11935 16858 11936
rect 14181 11794 14247 11797
rect 18965 11794 19031 11797
rect 14181 11792 19031 11794
rect 14181 11736 14186 11792
rect 14242 11736 18970 11792
rect 19026 11736 19031 11792
rect 14181 11734 19031 11736
rect 14181 11731 14247 11734
rect 18965 11731 19031 11734
rect 17953 11658 18019 11661
rect 22200 11658 23000 11688
rect 17953 11656 23000 11658
rect 17953 11600 17958 11656
rect 18014 11600 23000 11656
rect 17953 11598 23000 11600
rect 17953 11595 18019 11598
rect 22200 11568 23000 11598
rect 0 11522 800 11552
rect 1485 11522 1551 11525
rect 0 11520 1551 11522
rect 0 11464 1490 11520
rect 1546 11464 1551 11520
rect 0 11462 1551 11464
rect 0 11432 800 11462
rect 1485 11459 1551 11462
rect 3543 11456 3863 11457
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 11391 19457 11392
rect 17677 11386 17743 11389
rect 18137 11386 18203 11389
rect 17677 11384 18203 11386
rect 17677 11328 17682 11384
rect 17738 11328 18142 11384
rect 18198 11328 18203 11384
rect 17677 11326 18203 11328
rect 17677 11323 17743 11326
rect 18137 11323 18203 11326
rect 16665 11250 16731 11253
rect 18321 11250 18387 11253
rect 16665 11248 18387 11250
rect 16665 11192 16670 11248
rect 16726 11192 18326 11248
rect 18382 11192 18387 11248
rect 16665 11190 18387 11192
rect 16665 11187 16731 11190
rect 18321 11187 18387 11190
rect 19149 11250 19215 11253
rect 22200 11250 23000 11280
rect 19149 11248 23000 11250
rect 19149 11192 19154 11248
rect 19210 11192 23000 11248
rect 19149 11190 23000 11192
rect 19149 11187 19215 11190
rect 22200 11160 23000 11190
rect 14365 11114 14431 11117
rect 17493 11114 17559 11117
rect 14365 11112 17559 11114
rect 14365 11056 14370 11112
rect 14426 11056 17498 11112
rect 17554 11056 17559 11112
rect 14365 11054 17559 11056
rect 14365 11051 14431 11054
rect 17493 11051 17559 11054
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 16941 10842 17007 10845
rect 18781 10842 18847 10845
rect 16941 10840 18847 10842
rect 16941 10784 16946 10840
rect 17002 10784 18786 10840
rect 18842 10784 18847 10840
rect 16941 10782 18847 10784
rect 16941 10779 17007 10782
rect 18781 10779 18847 10782
rect 18045 10706 18111 10709
rect 22200 10706 23000 10736
rect 18045 10704 23000 10706
rect 18045 10648 18050 10704
rect 18106 10648 23000 10704
rect 18045 10646 23000 10648
rect 18045 10643 18111 10646
rect 22200 10616 23000 10646
rect 18689 10570 18755 10573
rect 18689 10568 19626 10570
rect 18689 10512 18694 10568
rect 18750 10512 19626 10568
rect 18689 10510 19626 10512
rect 18689 10507 18755 10510
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 10303 19457 10304
rect 19566 10298 19626 10510
rect 22200 10298 23000 10328
rect 19566 10238 23000 10298
rect 22200 10208 23000 10238
rect 10225 10162 10291 10165
rect 17677 10162 17743 10165
rect 10225 10160 17743 10162
rect 10225 10104 10230 10160
rect 10286 10104 17682 10160
rect 17738 10104 17743 10160
rect 10225 10102 17743 10104
rect 10225 10099 10291 10102
rect 17677 10099 17743 10102
rect 13261 10026 13327 10029
rect 20713 10026 20779 10029
rect 13261 10024 20779 10026
rect 13261 9968 13266 10024
rect 13322 9968 20718 10024
rect 20774 9968 20779 10024
rect 13261 9966 20779 9968
rect 13261 9963 13327 9966
rect 20713 9963 20779 9966
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 18965 9754 19031 9757
rect 22200 9754 23000 9784
rect 18965 9752 23000 9754
rect 18965 9696 18970 9752
rect 19026 9696 23000 9752
rect 18965 9694 23000 9696
rect 18965 9691 19031 9694
rect 22200 9664 23000 9694
rect 11881 9618 11947 9621
rect 11838 9616 11947 9618
rect 11838 9560 11886 9616
rect 11942 9560 11947 9616
rect 11838 9555 11947 9560
rect 11838 9349 11898 9555
rect 18321 9482 18387 9485
rect 18321 9480 19626 9482
rect 18321 9424 18326 9480
rect 18382 9424 19626 9480
rect 18321 9422 19626 9424
rect 18321 9419 18387 9422
rect 11838 9344 11947 9349
rect 11838 9288 11886 9344
rect 11942 9288 11947 9344
rect 11838 9286 11947 9288
rect 19566 9346 19626 9422
rect 22200 9346 23000 9376
rect 19566 9286 23000 9346
rect 11881 9283 11947 9286
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 22200 9256 23000 9286
rect 19137 9215 19457 9216
rect 10409 9210 10475 9213
rect 11973 9210 12039 9213
rect 10409 9208 12039 9210
rect 10409 9152 10414 9208
rect 10470 9152 11978 9208
rect 12034 9152 12039 9208
rect 10409 9150 12039 9152
rect 10409 9147 10475 9150
rect 11973 9147 12039 9150
rect 3969 9074 4035 9077
rect 19742 9074 19748 9076
rect 3969 9072 19748 9074
rect 3969 9016 3974 9072
rect 4030 9016 19748 9072
rect 3969 9014 19748 9016
rect 3969 9011 4035 9014
rect 19742 9012 19748 9014
rect 19812 9012 19818 9076
rect 5625 8938 5691 8941
rect 20345 8938 20411 8941
rect 5625 8936 20411 8938
rect 5625 8880 5630 8936
rect 5686 8880 20350 8936
rect 20406 8880 20411 8936
rect 5625 8878 20411 8880
rect 5625 8875 5691 8878
rect 20345 8875 20411 8878
rect 21357 8938 21423 8941
rect 22200 8938 23000 8968
rect 21357 8936 23000 8938
rect 21357 8880 21362 8936
rect 21418 8880 23000 8936
rect 21357 8878 23000 8880
rect 21357 8875 21423 8878
rect 22200 8848 23000 8878
rect 6142 8736 6462 8737
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 18045 8530 18111 8533
rect 18045 8528 19810 8530
rect 18045 8472 18050 8528
rect 18106 8472 19810 8528
rect 18045 8470 19810 8472
rect 18045 8467 18111 8470
rect 7005 8394 7071 8397
rect 15285 8394 15351 8397
rect 19750 8394 19810 8470
rect 22200 8394 23000 8424
rect 7005 8392 15351 8394
rect 7005 8336 7010 8392
rect 7066 8336 15290 8392
rect 15346 8336 15351 8392
rect 7005 8334 15351 8336
rect 7005 8331 7071 8334
rect 15285 8331 15351 8334
rect 19014 8334 19626 8394
rect 19750 8334 23000 8394
rect 16389 8258 16455 8261
rect 19014 8258 19074 8334
rect 16389 8256 19074 8258
rect 16389 8200 16394 8256
rect 16450 8200 19074 8256
rect 16389 8198 19074 8200
rect 19566 8258 19626 8334
rect 22200 8304 23000 8334
rect 21173 8258 21239 8261
rect 19566 8256 21239 8258
rect 19566 8200 21178 8256
rect 21234 8200 21239 8256
rect 19566 8198 21239 8200
rect 16389 8195 16455 8198
rect 21173 8195 21239 8198
rect 3543 8192 3863 8193
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 7465 7986 7531 7989
rect 18045 7986 18111 7989
rect 7465 7984 18111 7986
rect 7465 7928 7470 7984
rect 7526 7928 18050 7984
rect 18106 7928 18111 7984
rect 7465 7926 18111 7928
rect 7465 7923 7531 7926
rect 18045 7923 18111 7926
rect 18321 7986 18387 7989
rect 22200 7986 23000 8016
rect 18321 7984 23000 7986
rect 18321 7928 18326 7984
rect 18382 7928 23000 7984
rect 18321 7926 23000 7928
rect 18321 7923 18387 7926
rect 22200 7896 23000 7926
rect 6913 7850 6979 7853
rect 6913 7848 17418 7850
rect 6913 7792 6918 7848
rect 6974 7792 17418 7848
rect 6913 7790 17418 7792
rect 6913 7787 6979 7790
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 10501 7578 10567 7581
rect 16389 7578 16455 7581
rect 9630 7576 10567 7578
rect 9630 7547 10506 7576
rect 9627 7542 10506 7547
rect 9627 7486 9632 7542
rect 9688 7520 10506 7542
rect 10562 7520 10567 7576
rect 9688 7518 10567 7520
rect 9688 7486 9693 7518
rect 10501 7515 10567 7518
rect 12390 7576 16455 7578
rect 12390 7520 16394 7576
rect 16450 7520 16455 7576
rect 12390 7518 16455 7520
rect 17358 7578 17418 7790
rect 22200 7578 23000 7608
rect 17358 7518 23000 7578
rect 9627 7481 9693 7486
rect 2037 7442 2103 7445
rect 9213 7442 9279 7445
rect 2037 7440 9279 7442
rect 2037 7384 2042 7440
rect 2098 7384 9218 7440
rect 9274 7384 9279 7440
rect 2037 7382 9279 7384
rect 2037 7379 2103 7382
rect 9213 7379 9279 7382
rect 10961 7442 11027 7445
rect 12390 7442 12450 7518
rect 16389 7515 16455 7518
rect 22200 7488 23000 7518
rect 20989 7442 21055 7445
rect 10961 7440 12450 7442
rect 10961 7384 10966 7440
rect 11022 7384 12450 7440
rect 10961 7382 12450 7384
rect 13494 7440 21055 7442
rect 13494 7384 20994 7440
rect 21050 7384 21055 7440
rect 13494 7382 21055 7384
rect 10961 7379 11027 7382
rect 8017 7306 8083 7309
rect 13494 7306 13554 7382
rect 20989 7379 21055 7382
rect 8017 7304 13554 7306
rect 8017 7248 8022 7304
rect 8078 7248 13554 7304
rect 8017 7246 13554 7248
rect 13678 7246 19626 7306
rect 8017 7243 8083 7246
rect 9765 7170 9831 7173
rect 13678 7170 13738 7246
rect 9765 7168 13738 7170
rect 9765 7112 9770 7168
rect 9826 7112 13738 7168
rect 9765 7110 13738 7112
rect 14365 7170 14431 7173
rect 18965 7170 19031 7173
rect 14365 7168 19031 7170
rect 14365 7112 14370 7168
rect 14426 7112 18970 7168
rect 19026 7112 19031 7168
rect 14365 7110 19031 7112
rect 9765 7107 9831 7110
rect 14365 7107 14431 7110
rect 18965 7107 19031 7110
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 18321 7034 18387 7037
rect 5582 6974 8586 7034
rect 5349 6898 5415 6901
rect 5582 6898 5642 6974
rect 5349 6896 5642 6898
rect 5349 6840 5354 6896
rect 5410 6840 5642 6896
rect 5349 6838 5642 6840
rect 8526 6898 8586 6974
rect 9262 6974 13738 7034
rect 9262 6898 9322 6974
rect 8526 6838 9322 6898
rect 13678 6898 13738 6974
rect 14414 7032 18387 7034
rect 14414 6976 18326 7032
rect 18382 6976 18387 7032
rect 14414 6974 18387 6976
rect 19566 7034 19626 7246
rect 22200 7034 23000 7064
rect 19566 6974 23000 7034
rect 14414 6898 14474 6974
rect 18321 6971 18387 6974
rect 22200 6944 23000 6974
rect 13678 6838 14474 6898
rect 15285 6898 15351 6901
rect 18045 6898 18111 6901
rect 15285 6896 18111 6898
rect 15285 6840 15290 6896
rect 15346 6840 18050 6896
rect 18106 6840 18111 6896
rect 15285 6838 18111 6840
rect 5349 6835 5415 6838
rect 15285 6835 15351 6838
rect 18045 6835 18111 6838
rect 6269 6762 6335 6765
rect 20345 6762 20411 6765
rect 6269 6760 20411 6762
rect 6269 6704 6274 6760
rect 6330 6704 20350 6760
rect 20406 6704 20411 6760
rect 6269 6702 20411 6704
rect 6269 6699 6335 6702
rect 20345 6699 20411 6702
rect 18137 6626 18203 6629
rect 22200 6626 23000 6656
rect 18137 6624 23000 6626
rect 18137 6568 18142 6624
rect 18198 6568 23000 6624
rect 18137 6566 23000 6568
rect 18137 6563 18203 6566
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 22200 6536 23000 6566
rect 16538 6495 16858 6496
rect 7833 6490 7899 6493
rect 9581 6490 9647 6493
rect 7833 6488 9647 6490
rect 7833 6432 7838 6488
rect 7894 6432 9586 6488
rect 9642 6432 9647 6488
rect 7833 6430 9647 6432
rect 7833 6427 7899 6430
rect 9581 6427 9647 6430
rect 11789 6490 11855 6493
rect 15285 6490 15351 6493
rect 11789 6488 15351 6490
rect 11789 6432 11794 6488
rect 11850 6432 15290 6488
rect 15346 6432 15351 6488
rect 11789 6430 15351 6432
rect 11789 6427 11855 6430
rect 15285 6427 15351 6430
rect 4654 6292 4660 6356
rect 4724 6354 4730 6356
rect 9121 6354 9187 6357
rect 4724 6352 9187 6354
rect 4724 6296 9126 6352
rect 9182 6296 9187 6352
rect 4724 6294 9187 6296
rect 4724 6292 4730 6294
rect 9121 6291 9187 6294
rect 9489 6354 9555 6357
rect 20897 6354 20963 6357
rect 9489 6352 20963 6354
rect 9489 6296 9494 6352
rect 9550 6296 20902 6352
rect 20958 6296 20963 6352
rect 9489 6294 20963 6296
rect 9489 6291 9555 6294
rect 20897 6291 20963 6294
rect 7005 6218 7071 6221
rect 21081 6218 21147 6221
rect 7005 6216 21147 6218
rect 7005 6160 7010 6216
rect 7066 6160 21086 6216
rect 21142 6160 21147 6216
rect 7005 6158 21147 6160
rect 7005 6155 7071 6158
rect 21081 6155 21147 6158
rect 9121 6082 9187 6085
rect 11789 6082 11855 6085
rect 22200 6082 23000 6112
rect 9121 6080 11855 6082
rect 9121 6024 9126 6080
rect 9182 6024 11794 6080
rect 11850 6024 11855 6080
rect 9121 6022 11855 6024
rect 9121 6019 9187 6022
rect 11789 6019 11855 6022
rect 19566 6022 23000 6082
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 5951 19457 5952
rect 15745 5946 15811 5949
rect 18965 5946 19031 5949
rect 14782 5886 15578 5946
rect 5993 5810 6059 5813
rect 14782 5810 14842 5886
rect 5993 5808 14842 5810
rect 5993 5752 5998 5808
rect 6054 5752 14842 5808
rect 5993 5750 14842 5752
rect 5993 5747 6059 5750
rect 14958 5748 14964 5812
rect 15028 5810 15034 5812
rect 15101 5810 15167 5813
rect 15028 5808 15167 5810
rect 15028 5752 15106 5808
rect 15162 5752 15167 5808
rect 15028 5750 15167 5752
rect 15518 5810 15578 5886
rect 15745 5944 19031 5946
rect 15745 5888 15750 5944
rect 15806 5888 18970 5944
rect 19026 5888 19031 5944
rect 15745 5886 19031 5888
rect 15745 5883 15811 5886
rect 18965 5883 19031 5886
rect 18045 5810 18111 5813
rect 15518 5808 18111 5810
rect 15518 5752 18050 5808
rect 18106 5752 18111 5808
rect 15518 5750 18111 5752
rect 15028 5748 15034 5750
rect 15101 5747 15167 5750
rect 18045 5747 18111 5750
rect 18873 5810 18939 5813
rect 19566 5810 19626 6022
rect 22200 5992 23000 6022
rect 18873 5808 19626 5810
rect 18873 5752 18878 5808
rect 18934 5752 19626 5808
rect 18873 5750 19626 5752
rect 18873 5747 18939 5750
rect 6545 5674 6611 5677
rect 17677 5674 17743 5677
rect 6545 5672 17743 5674
rect 6545 5616 6550 5672
rect 6606 5616 17682 5672
rect 17738 5616 17743 5672
rect 6545 5614 17743 5616
rect 6545 5611 6611 5614
rect 17677 5611 17743 5614
rect 18137 5674 18203 5677
rect 22200 5674 23000 5704
rect 18137 5672 23000 5674
rect 18137 5616 18142 5672
rect 18198 5616 23000 5672
rect 18137 5614 23000 5616
rect 18137 5611 18203 5614
rect 22200 5584 23000 5614
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 6453 5266 6519 5269
rect 10409 5266 10475 5269
rect 14181 5266 14247 5269
rect 6453 5264 14247 5266
rect 6453 5208 6458 5264
rect 6514 5208 10414 5264
rect 10470 5208 14186 5264
rect 14242 5208 14247 5264
rect 6453 5206 14247 5208
rect 6453 5203 6519 5206
rect 10409 5203 10475 5206
rect 14181 5203 14247 5206
rect 14825 5266 14891 5269
rect 18229 5266 18295 5269
rect 14825 5264 18295 5266
rect 14825 5208 14830 5264
rect 14886 5208 18234 5264
rect 18290 5208 18295 5264
rect 14825 5206 18295 5208
rect 14825 5203 14891 5206
rect 18229 5203 18295 5206
rect 18505 5266 18571 5269
rect 22200 5266 23000 5296
rect 18505 5264 23000 5266
rect 18505 5208 18510 5264
rect 18566 5208 23000 5264
rect 18505 5206 23000 5208
rect 18505 5203 18571 5206
rect 22200 5176 23000 5206
rect 6545 5130 6611 5133
rect 18229 5130 18295 5133
rect 6545 5128 18295 5130
rect 6545 5072 6550 5128
rect 6606 5072 18234 5128
rect 18290 5072 18295 5128
rect 6545 5070 18295 5072
rect 6545 5067 6611 5070
rect 18229 5067 18295 5070
rect 3543 4928 3863 4929
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 16849 4858 16915 4861
rect 17769 4858 17835 4861
rect 16849 4856 17835 4858
rect 16849 4800 16854 4856
rect 16910 4800 17774 4856
rect 17830 4800 17835 4856
rect 16849 4798 17835 4800
rect 16849 4795 16915 4798
rect 17769 4795 17835 4798
rect 5717 4722 5783 4725
rect 21725 4722 21791 4725
rect 22200 4722 23000 4752
rect 5717 4720 17556 4722
rect 5717 4664 5722 4720
rect 5778 4664 17556 4720
rect 5717 4662 17556 4664
rect 5717 4659 5783 4662
rect 17496 4589 17556 4662
rect 21725 4720 23000 4722
rect 21725 4664 21730 4720
rect 21786 4664 23000 4720
rect 21725 4662 23000 4664
rect 21725 4659 21791 4662
rect 22200 4632 23000 4662
rect 7097 4586 7163 4589
rect 8109 4586 8175 4589
rect 7097 4584 11898 4586
rect 7097 4528 7102 4584
rect 7158 4528 8114 4584
rect 8170 4528 11898 4584
rect 7097 4526 11898 4528
rect 7097 4523 7163 4526
rect 8109 4523 8175 4526
rect 11838 4450 11898 4526
rect 17493 4584 17559 4589
rect 17493 4528 17498 4584
rect 17554 4528 17559 4584
rect 17493 4523 17559 4528
rect 11838 4390 12450 4450
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 12390 4314 12450 4390
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 4319 16858 4320
rect 18781 4314 18847 4317
rect 22200 4314 23000 4344
rect 12390 4254 16314 4314
rect 5533 4178 5599 4181
rect 15377 4178 15443 4181
rect 5533 4176 15443 4178
rect 5533 4120 5538 4176
rect 5594 4120 15382 4176
rect 15438 4120 15443 4176
rect 5533 4118 15443 4120
rect 16254 4178 16314 4254
rect 18781 4312 23000 4314
rect 18781 4256 18786 4312
rect 18842 4256 23000 4312
rect 18781 4254 23000 4256
rect 18781 4251 18847 4254
rect 22200 4224 23000 4254
rect 18597 4178 18663 4181
rect 16254 4176 18663 4178
rect 16254 4120 18602 4176
rect 18658 4120 18663 4176
rect 16254 4118 18663 4120
rect 5533 4115 5599 4118
rect 15377 4115 15443 4118
rect 18597 4115 18663 4118
rect 4613 4044 4679 4045
rect 4613 4042 4660 4044
rect 4568 4040 4660 4042
rect 4568 3984 4618 4040
rect 4568 3982 4660 3984
rect 4613 3980 4660 3982
rect 4724 3980 4730 4044
rect 7005 4042 7071 4045
rect 16757 4042 16823 4045
rect 7005 4040 16823 4042
rect 7005 3984 7010 4040
rect 7066 3984 16762 4040
rect 16818 3984 16823 4040
rect 7005 3982 16823 3984
rect 4613 3979 4679 3980
rect 7005 3979 7071 3982
rect 16757 3979 16823 3982
rect 17493 4042 17559 4045
rect 17861 4042 17927 4045
rect 18873 4042 18939 4045
rect 17493 4040 18939 4042
rect 17493 3984 17498 4040
rect 17554 3984 17866 4040
rect 17922 3984 18878 4040
rect 18934 3984 18939 4040
rect 17493 3982 18939 3984
rect 17493 3979 17559 3982
rect 17861 3979 17927 3982
rect 18873 3979 18939 3982
rect 15929 3906 15995 3909
rect 17217 3906 17283 3909
rect 22200 3906 23000 3936
rect 15929 3904 17283 3906
rect 15929 3848 15934 3904
rect 15990 3848 17222 3904
rect 17278 3848 17283 3904
rect 15929 3846 17283 3848
rect 15929 3843 15995 3846
rect 17217 3843 17283 3846
rect 19566 3846 23000 3906
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 7649 3770 7715 3773
rect 8017 3770 8083 3773
rect 16113 3770 16179 3773
rect 7649 3768 8083 3770
rect 7649 3712 7654 3768
rect 7710 3712 8022 3768
rect 8078 3712 8083 3768
rect 7649 3710 8083 3712
rect 7649 3707 7715 3710
rect 8017 3707 8083 3710
rect 14966 3768 16179 3770
rect 14966 3712 16118 3768
rect 16174 3712 16179 3768
rect 14966 3710 16179 3712
rect 6545 3634 6611 3637
rect 14966 3634 15026 3710
rect 16113 3707 16179 3710
rect 16481 3770 16547 3773
rect 18597 3770 18663 3773
rect 16481 3768 18663 3770
rect 16481 3712 16486 3768
rect 16542 3712 18602 3768
rect 18658 3712 18663 3768
rect 16481 3710 18663 3712
rect 16481 3707 16547 3710
rect 18597 3707 18663 3710
rect 6545 3632 15026 3634
rect 6545 3576 6550 3632
rect 6606 3576 15026 3632
rect 6545 3574 15026 3576
rect 15193 3634 15259 3637
rect 18689 3634 18755 3637
rect 15193 3632 18755 3634
rect 15193 3576 15198 3632
rect 15254 3576 18694 3632
rect 18750 3576 18755 3632
rect 15193 3574 18755 3576
rect 6545 3571 6611 3574
rect 15193 3571 15259 3574
rect 18689 3571 18755 3574
rect 6637 3498 6703 3501
rect 11789 3498 11855 3501
rect 19566 3498 19626 3846
rect 22200 3816 23000 3846
rect 6637 3496 11855 3498
rect 6637 3440 6642 3496
rect 6698 3440 11794 3496
rect 11850 3440 11855 3496
rect 6637 3438 11855 3440
rect 6637 3435 6703 3438
rect 11789 3435 11855 3438
rect 12390 3438 19626 3498
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 7557 3226 7623 3229
rect 10593 3226 10659 3229
rect 7557 3224 10659 3226
rect 7557 3168 7562 3224
rect 7618 3168 10598 3224
rect 10654 3168 10659 3224
rect 7557 3166 10659 3168
rect 7557 3163 7623 3166
rect 10593 3163 10659 3166
rect 4613 3090 4679 3093
rect 9121 3090 9187 3093
rect 4613 3088 9187 3090
rect 4613 3032 4618 3088
rect 4674 3032 9126 3088
rect 9182 3032 9187 3088
rect 4613 3030 9187 3032
rect 4613 3027 4679 3030
rect 9121 3027 9187 3030
rect 9489 3090 9555 3093
rect 12390 3090 12450 3438
rect 12525 3362 12591 3365
rect 16205 3362 16271 3365
rect 12525 3360 16271 3362
rect 12525 3304 12530 3360
rect 12586 3304 16210 3360
rect 16266 3304 16271 3360
rect 12525 3302 16271 3304
rect 12525 3299 12591 3302
rect 16205 3299 16271 3302
rect 19057 3362 19123 3365
rect 22200 3362 23000 3392
rect 19057 3360 23000 3362
rect 19057 3304 19062 3360
rect 19118 3304 23000 3360
rect 19057 3302 23000 3304
rect 19057 3299 19123 3302
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 22200 3272 23000 3302
rect 16538 3231 16858 3232
rect 14457 3226 14523 3229
rect 16297 3226 16363 3229
rect 14457 3224 16363 3226
rect 14457 3168 14462 3224
rect 14518 3168 16302 3224
rect 16358 3168 16363 3224
rect 14457 3166 16363 3168
rect 14457 3163 14523 3166
rect 16297 3163 16363 3166
rect 17585 3090 17651 3093
rect 9489 3088 12450 3090
rect 9489 3032 9494 3088
rect 9550 3032 12450 3088
rect 9489 3030 12450 3032
rect 13494 3088 17651 3090
rect 13494 3032 17590 3088
rect 17646 3032 17651 3088
rect 13494 3030 17651 3032
rect 9489 3027 9555 3030
rect 3693 2954 3759 2957
rect 13494 2954 13554 3030
rect 17585 3027 17651 3030
rect 3693 2952 13554 2954
rect 3693 2896 3698 2952
rect 3754 2896 13554 2952
rect 3693 2894 13554 2896
rect 19425 2954 19491 2957
rect 19793 2956 19859 2957
rect 19742 2954 19748 2956
rect 19425 2952 19748 2954
rect 19812 2954 19859 2956
rect 20529 2954 20595 2957
rect 22200 2954 23000 2984
rect 19812 2952 19904 2954
rect 19425 2896 19430 2952
rect 19486 2896 19748 2952
rect 19854 2896 19904 2952
rect 19425 2894 19748 2896
rect 3693 2891 3759 2894
rect 19425 2891 19491 2894
rect 19742 2892 19748 2894
rect 19812 2894 19904 2896
rect 20529 2952 23000 2954
rect 20529 2896 20534 2952
rect 20590 2896 23000 2952
rect 20529 2894 23000 2896
rect 19812 2892 19859 2894
rect 19793 2891 19859 2892
rect 20529 2891 20595 2894
rect 22200 2864 23000 2894
rect 4613 2818 4679 2821
rect 4797 2818 4863 2821
rect 8385 2818 8451 2821
rect 4613 2816 8451 2818
rect 4613 2760 4618 2816
rect 4674 2760 4802 2816
rect 4858 2760 8390 2816
rect 8446 2760 8451 2816
rect 4613 2758 8451 2760
rect 4613 2755 4679 2758
rect 4797 2755 4863 2758
rect 8385 2755 8451 2758
rect 9121 2818 9187 2821
rect 13721 2818 13787 2821
rect 9121 2816 13787 2818
rect 9121 2760 9126 2816
rect 9182 2760 13726 2816
rect 13782 2760 13787 2816
rect 9121 2758 13787 2760
rect 9121 2755 9187 2758
rect 13721 2755 13787 2758
rect 17217 2818 17283 2821
rect 17769 2818 17835 2821
rect 17217 2816 17835 2818
rect 17217 2760 17222 2816
rect 17278 2760 17774 2816
rect 17830 2760 17835 2816
rect 17217 2758 17835 2760
rect 17217 2755 17283 2758
rect 17769 2755 17835 2758
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 5809 2682 5875 2685
rect 6821 2682 6887 2685
rect 5809 2680 6887 2682
rect 5809 2624 5814 2680
rect 5870 2624 6826 2680
rect 6882 2624 6887 2680
rect 5809 2622 6887 2624
rect 5809 2619 5875 2622
rect 6821 2619 6887 2622
rect 6637 2546 6703 2549
rect 8937 2546 9003 2549
rect 14641 2546 14707 2549
rect 6637 2544 9003 2546
rect 6637 2488 6642 2544
rect 6698 2488 8942 2544
rect 8998 2488 9003 2544
rect 6637 2486 9003 2488
rect 6637 2483 6703 2486
rect 8937 2483 9003 2486
rect 10734 2544 14707 2546
rect 10734 2488 14646 2544
rect 14702 2488 14707 2544
rect 10734 2486 14707 2488
rect 2957 2410 3023 2413
rect 10734 2410 10794 2486
rect 14641 2483 14707 2486
rect 18873 2410 18939 2413
rect 2957 2408 10794 2410
rect 2957 2352 2962 2408
rect 3018 2352 10794 2408
rect 2957 2350 10794 2352
rect 11102 2408 18939 2410
rect 11102 2352 18878 2408
rect 18934 2352 18939 2408
rect 11102 2350 18939 2352
rect 2957 2347 3023 2350
rect 6821 2274 6887 2277
rect 11102 2274 11162 2350
rect 18873 2347 18939 2350
rect 20529 2410 20595 2413
rect 22200 2410 23000 2440
rect 20529 2408 23000 2410
rect 20529 2352 20534 2408
rect 20590 2352 23000 2408
rect 20529 2350 23000 2352
rect 20529 2347 20595 2350
rect 22200 2320 23000 2350
rect 6821 2272 11162 2274
rect 6821 2216 6826 2272
rect 6882 2216 11162 2272
rect 6821 2214 11162 2216
rect 6821 2211 6887 2214
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 5533 2002 5599 2005
rect 12065 2002 12131 2005
rect 5533 2000 12131 2002
rect 5533 1944 5538 2000
rect 5594 1944 12070 2000
rect 12126 1944 12131 2000
rect 5533 1942 12131 1944
rect 5533 1939 5599 1942
rect 12065 1939 12131 1942
rect 18873 2002 18939 2005
rect 22200 2002 23000 2032
rect 18873 2000 23000 2002
rect 18873 1944 18878 2000
rect 18934 1944 23000 2000
rect 18873 1942 23000 1944
rect 18873 1939 18939 1942
rect 22200 1912 23000 1942
rect 2129 1866 2195 1869
rect 18413 1866 18479 1869
rect 2129 1864 18479 1866
rect 2129 1808 2134 1864
rect 2190 1808 18418 1864
rect 18474 1808 18479 1864
rect 2129 1806 18479 1808
rect 2129 1803 2195 1806
rect 18413 1803 18479 1806
rect 4705 1730 4771 1733
rect 19057 1730 19123 1733
rect 4705 1728 19123 1730
rect 4705 1672 4710 1728
rect 4766 1672 19062 1728
rect 19118 1672 19123 1728
rect 4705 1670 19123 1672
rect 4705 1667 4771 1670
rect 19057 1667 19123 1670
rect 5441 1594 5507 1597
rect 10869 1594 10935 1597
rect 5441 1592 10935 1594
rect 5441 1536 5446 1592
rect 5502 1536 10874 1592
rect 10930 1536 10935 1592
rect 5441 1534 10935 1536
rect 5441 1531 5507 1534
rect 10869 1531 10935 1534
rect 19517 1594 19583 1597
rect 22200 1594 23000 1624
rect 19517 1592 23000 1594
rect 19517 1536 19522 1592
rect 19578 1536 23000 1592
rect 19517 1534 23000 1536
rect 19517 1531 19583 1534
rect 22200 1504 23000 1534
rect 19793 1050 19859 1053
rect 22200 1050 23000 1080
rect 19793 1048 23000 1050
rect 19793 992 19798 1048
rect 19854 992 23000 1048
rect 19793 990 23000 992
rect 19793 987 19859 990
rect 22200 960 23000 990
rect 20621 914 20687 917
rect 20621 912 21282 914
rect 20621 856 20626 912
rect 20682 856 21282 912
rect 20621 854 21282 856
rect 20621 851 20687 854
rect 21222 642 21282 854
rect 22200 642 23000 672
rect 21222 582 23000 642
rect 22200 552 23000 582
rect 19425 234 19491 237
rect 22200 234 23000 264
rect 19425 232 23000 234
rect 19425 176 19430 232
rect 19486 176 23000 232
rect 19425 174 23000 176
rect 19425 171 19491 174
rect 22200 144 23000 174
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 14964 17172 15028 17236
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 19748 9012 19812 9076
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 4660 6292 4724 6356
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 14964 5748 15028 5812
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 4660 4040 4724 4044
rect 4660 3984 4674 4040
rect 4674 3984 4724 4040
rect 4660 3980 4724 3984
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 19748 2952 19812 2956
rect 19748 2896 19798 2952
rect 19798 2896 19812 2952
rect 19748 2892 19812 2896
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 13632 3863 14656
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 4659 6356 4725 6357
rect 4659 6292 4660 6356
rect 4724 6292 4725 6356
rect 4659 6291 4725 6292
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 4662 4045 4722 6291
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 4659 4044 4725 4045
rect 4659 3980 4660 4044
rect 4724 3980 4725 4044
rect 4659 3979 4725 3980
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 14963 17236 15029 17237
rect 14963 17172 14964 17236
rect 15028 17172 15029 17236
rect 14963 17171 15029 17172
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 14966 5813 15026 17171
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 14963 5812 15029 5813
rect 14963 5748 14964 5812
rect 15028 5748 15029 5812
rect 14963 5747 15029 5748
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19747 9076 19813 9077
rect 19747 9012 19748 9076
rect 19812 9012 19813 9076
rect 19747 9011 19813 9012
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19750 2957 19810 9011
rect 19747 2956 19813 2957
rect 19747 2892 19748 2956
rect 19812 2892 19813 2956
rect 19747 2891 19813 2892
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__74__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5152 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 1564 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 15272 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 12880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 18400 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 19504 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 6072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 6992 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 1564 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 5060 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2208 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 2392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 2024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_1.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_5.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15732 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_9.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 12512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_bottom_track_25.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 12328 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 11684 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_34.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 12696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_36.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_right_track_38.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output53_A
timestamp 1649977179
transform -1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output54_A
timestamp 1649977179
transform 1 0 1932 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1932 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16
timestamp 1649977179
transform 1 0 2576 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21
timestamp 1649977179
transform 1 0 3036 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 1649977179
transform 1 0 3496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44
timestamp 1649977179
transform 1 0 5152 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54
timestamp 1649977179
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59
timestamp 1649977179
transform 1 0 6532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64
timestamp 1649977179
transform 1 0 6992 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_82
timestamp 1649977179
transform 1 0 8648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_94
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_99
timestamp 1649977179
transform 1 0 10212 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 1649977179
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_121
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_132
timestamp 1649977179
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_138
timestamp 1649977179
transform 1 0 13800 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_145
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_149 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_159
timestamp 1649977179
transform 1 0 15732 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_171
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1649977179
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1649977179
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_6
timestamp 1649977179
transform 1 0 1656 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_11
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_16
timestamp 1649977179
transform 1 0 2576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_21
timestamp 1649977179
transform 1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1649977179
transform 1 0 3404 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_29
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_34
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_44
timestamp 1649977179
transform 1 0 5152 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_49
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_54
timestamp 1649977179
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_60
timestamp 1649977179
transform 1 0 6624 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_88
timestamp 1649977179
transform 1 0 9200 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_92
timestamp 1649977179
transform 1 0 9568 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 1649977179
transform 1 0 11224 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_117
timestamp 1649977179
transform 1 0 11868 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_135
timestamp 1649977179
transform 1 0 13524 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_146
timestamp 1649977179
transform 1 0 14536 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_165
timestamp 1649977179
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_178
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_184
timestamp 1649977179
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_196
timestamp 1649977179
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_221
timestamp 1649977179
transform 1 0 21436 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_6
timestamp 1649977179
transform 1 0 1656 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_10
timestamp 1649977179
transform 1 0 2024 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_14
timestamp 1649977179
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 1649977179
transform 1 0 2760 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_22
timestamp 1649977179
transform 1 0 3128 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_26
timestamp 1649977179
transform 1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_31
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_36
timestamp 1649977179
transform 1 0 4416 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_46
timestamp 1649977179
transform 1 0 5336 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_56
timestamp 1649977179
transform 1 0 6256 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_61
timestamp 1649977179
transform 1 0 6716 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_71
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_82
timestamp 1649977179
transform 1 0 8648 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_94
timestamp 1649977179
transform 1 0 9752 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_113
timestamp 1649977179
transform 1 0 11500 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_120
timestamp 1649977179
transform 1 0 12144 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_138
timestamp 1649977179
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_144
timestamp 1649977179
transform 1 0 14352 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_162
timestamp 1649977179
transform 1 0 16008 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 1649977179
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_194
timestamp 1649977179
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_5
timestamp 1649977179
transform 1 0 1564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_10
timestamp 1649977179
transform 1 0 2024 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_14
timestamp 1649977179
transform 1 0 2392 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_18
timestamp 1649977179
transform 1 0 2760 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_22
timestamp 1649977179
transform 1 0 3128 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_26
timestamp 1649977179
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 1649977179
transform 1 0 3864 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_34
timestamp 1649977179
transform 1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_44
timestamp 1649977179
transform 1 0 5152 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_49
timestamp 1649977179
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 1649977179
transform 1 0 6072 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_62
timestamp 1649977179
transform 1 0 6808 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_72
timestamp 1649977179
transform 1 0 7728 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_90
timestamp 1649977179
transform 1 0 9384 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_94
timestamp 1649977179
transform 1 0 9752 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_99
timestamp 1649977179
transform 1 0 10212 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_110
timestamp 1649977179
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_122
timestamp 1649977179
transform 1 0 12328 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_126
timestamp 1649977179
transform 1 0 12696 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_147
timestamp 1649977179
transform 1 0 14628 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_151
timestamp 1649977179
transform 1 0 14996 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_162
timestamp 1649977179
transform 1 0 16008 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 1649977179
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_185
timestamp 1649977179
transform 1 0 18124 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1649977179
transform 1 0 19780 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_221
timestamp 1649977179
transform 1 0 21436 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_8
timestamp 1649977179
transform 1 0 1840 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_12
timestamp 1649977179
transform 1 0 2208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_18
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_22
timestamp 1649977179
transform 1 0 3128 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_26
timestamp 1649977179
transform 1 0 3496 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_32
timestamp 1649977179
transform 1 0 4048 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_36
timestamp 1649977179
transform 1 0 4416 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_40
timestamp 1649977179
transform 1 0 4784 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_45
timestamp 1649977179
transform 1 0 5244 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_50
timestamp 1649977179
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_60
timestamp 1649977179
transform 1 0 6624 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1649977179
transform 1 0 7636 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_82
timestamp 1649977179
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_87
timestamp 1649977179
transform 1 0 9108 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1649977179
transform 1 0 9568 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_110
timestamp 1649977179
transform 1 0 11224 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_120
timestamp 1649977179
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_138
timestamp 1649977179
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_149
timestamp 1649977179
transform 1 0 14812 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_160
timestamp 1649977179
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_172
timestamp 1649977179
transform 1 0 16928 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_183
timestamp 1649977179
transform 1 0 17940 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_194
timestamp 1649977179
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_220
timestamp 1649977179
transform 1 0 21344 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_5 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_17 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2668 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_25
timestamp 1649977179
transform 1 0 3404 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_28 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_43
timestamp 1649977179
transform 1 0 5060 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_49
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 1649977179
transform 1 0 6072 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1649977179
transform 1 0 6532 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_64
timestamp 1649977179
transform 1 0 6992 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_82
timestamp 1649977179
transform 1 0 8648 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1649977179
transform 1 0 9568 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_110
timestamp 1649977179
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_119
timestamp 1649977179
transform 1 0 12052 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_148
timestamp 1649977179
transform 1 0 14720 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_166
timestamp 1649977179
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_178
timestamp 1649977179
transform 1 0 17480 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 1649977179
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_196
timestamp 1649977179
transform 1 0 19136 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 1649977179
transform 1 0 20148 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_218
timestamp 1649977179
transform 1 0 21160 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_37
timestamp 1649977179
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_46
timestamp 1649977179
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 1649977179
transform 1 0 5704 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_54
timestamp 1649977179
transform 1 0 6072 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_64
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_82
timestamp 1649977179
transform 1 0 8648 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_94
timestamp 1649977179
transform 1 0 9752 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_99
timestamp 1649977179
transform 1 0 10212 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_131
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_150
timestamp 1649977179
transform 1 0 14904 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_156
timestamp 1649977179
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_178
timestamp 1649977179
transform 1 0 17480 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1649977179
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_213
timestamp 1649977179
transform 1 0 20700 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_54
timestamp 1649977179
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 1649977179
transform 1 0 6624 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1649977179
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_75
timestamp 1649977179
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_110
timestamp 1649977179
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_128
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_139
timestamp 1649977179
transform 1 0 13892 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_145
timestamp 1649977179
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_163
timestamp 1649977179
transform 1 0 16100 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_186
timestamp 1649977179
transform 1 0 18216 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_204
timestamp 1649977179
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_215
timestamp 1649977179
transform 1 0 20884 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_49
timestamp 1649977179
transform 1 0 5612 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp 1649977179
transform 1 0 5888 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_57
timestamp 1649977179
transform 1 0 6348 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_62
timestamp 1649977179
transform 1 0 6808 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_72
timestamp 1649977179
transform 1 0 7728 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_82
timestamp 1649977179
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_94
timestamp 1649977179
transform 1 0 9752 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_100
timestamp 1649977179
transform 1 0 10304 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_118
timestamp 1649977179
transform 1 0 11960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_129
timestamp 1649977179
transform 1 0 12972 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 1649977179
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_151
timestamp 1649977179
transform 1 0 14996 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_162
timestamp 1649977179
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_173
timestamp 1649977179
transform 1 0 17020 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_184
timestamp 1649977179
transform 1 0 18032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 1649977179
transform 1 0 18952 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_201
timestamp 1649977179
transform 1 0 19596 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_219
timestamp 1649977179
transform 1 0 21252 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_61
timestamp 1649977179
transform 1 0 6716 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_66
timestamp 1649977179
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_71
timestamp 1649977179
transform 1 0 7636 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_76
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_104
timestamp 1649977179
transform 1 0 10672 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1649977179
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_119
timestamp 1649977179
transform 1 0 12052 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_155
timestamp 1649977179
transform 1 0 15364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 1649977179
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_188
timestamp 1649977179
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_198
timestamp 1649977179
transform 1 0 19320 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_209
timestamp 1649977179
transform 1 0 20332 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 1649977179
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_64
timestamp 1649977179
transform 1 0 6992 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_68
timestamp 1649977179
transform 1 0 7360 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_72
timestamp 1649977179
transform 1 0 7728 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_88
timestamp 1649977179
transform 1 0 9200 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_99
timestamp 1649977179
transform 1 0 10212 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_128
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 1649977179
transform 1 0 13800 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_164
timestamp 1649977179
transform 1 0 16192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_186
timestamp 1649977179
transform 1 0 18216 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_200
timestamp 1649977179
transform 1 0 19504 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_75
timestamp 1649977179
transform 1 0 8004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_92
timestamp 1649977179
transform 1 0 9568 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_110
timestamp 1649977179
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_121
timestamp 1649977179
transform 1 0 12236 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_126
timestamp 1649977179
transform 1 0 12696 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_150
timestamp 1649977179
transform 1 0 14904 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_163
timestamp 1649977179
transform 1 0 16100 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_185
timestamp 1649977179
transform 1 0 18124 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_196
timestamp 1649977179
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_202
timestamp 1649977179
transform 1 0 19688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_221
timestamp 1649977179
transform 1 0 21436 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_72
timestamp 1649977179
transform 1 0 7728 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 1649977179
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_101
timestamp 1649977179
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_105
timestamp 1649977179
transform 1 0 10764 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_116
timestamp 1649977179
transform 1 0 11776 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_120
timestamp 1649977179
transform 1 0 12144 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_157
timestamp 1649977179
transform 1 0 15548 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_175
timestamp 1649977179
transform 1 0 17204 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_183
timestamp 1649977179
transform 1 0 17940 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1649977179
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_216
timestamp 1649977179
transform 1 0 20976 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_92
timestamp 1649977179
transform 1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 1649977179
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_136
timestamp 1649977179
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_147
timestamp 1649977179
transform 1 0 14628 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_157
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_162
timestamp 1649977179
transform 1 0 16008 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_178
timestamp 1649977179
transform 1 0 17480 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_189
timestamp 1649977179
transform 1 0 18492 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_207
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_221
timestamp 1649977179
transform 1 0 21436 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_122
timestamp 1649977179
transform 1 0 12328 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_126
timestamp 1649977179
transform 1 0 12696 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_136
timestamp 1649977179
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_150
timestamp 1649977179
transform 1 0 14904 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_161
timestamp 1649977179
transform 1 0 15916 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_171
timestamp 1649977179
transform 1 0 16836 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_176
timestamp 1649977179
transform 1 0 17296 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1649977179
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_207
timestamp 1649977179
transform 1 0 20148 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_217
timestamp 1649977179
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_117
timestamp 1649977179
transform 1 0 11868 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_140
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_158
timestamp 1649977179
transform 1 0 15640 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_162
timestamp 1649977179
transform 1 0 16008 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_188
timestamp 1649977179
transform 1 0 18400 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_197
timestamp 1649977179
transform 1 0 19228 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_208
timestamp 1649977179
transform 1 0 20240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_219
timestamp 1649977179
transform 1 0 21252 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_124
timestamp 1649977179
transform 1 0 12512 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_128
timestamp 1649977179
transform 1 0 12880 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_144
timestamp 1649977179
transform 1 0 14352 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_164
timestamp 1649977179
transform 1 0 16192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_170
timestamp 1649977179
transform 1 0 16744 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_181
timestamp 1649977179
transform 1 0 17756 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_191
timestamp 1649977179
transform 1 0 18676 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_200
timestamp 1649977179
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_219
timestamp 1649977179
transform 1 0 21252 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_7
timestamp 1649977179
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_11
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_23
timestamp 1649977179
transform 1 0 3220 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_35
timestamp 1649977179
transform 1 0 4324 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_47
timestamp 1649977179
transform 1 0 5428 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 1649977179
transform 1 0 13340 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 1649977179
transform 1 0 14628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_154
timestamp 1649977179
transform 1 0 15272 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_172
timestamp 1649977179
transform 1 0 16928 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_182
timestamp 1649977179
transform 1 0 17848 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1649977179
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_204
timestamp 1649977179
transform 1 0 19872 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_214
timestamp 1649977179
transform 1 0 20792 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_143
timestamp 1649977179
transform 1 0 14260 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_147
timestamp 1649977179
transform 1 0 14628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_152
timestamp 1649977179
transform 1 0 15088 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_157
timestamp 1649977179
transform 1 0 15548 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_175
timestamp 1649977179
transform 1 0 17204 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_193
timestamp 1649977179
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_213
timestamp 1649977179
transform 1 0 20700 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_154
timestamp 1649977179
transform 1 0 15272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 1649977179
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_178
timestamp 1649977179
transform 1 0 17480 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_189
timestamp 1649977179
transform 1 0 18492 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_200
timestamp 1649977179
transform 1 0 19504 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_210
timestamp 1649977179
transform 1 0 20424 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 1649977179
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_20_161
timestamp 1649977179
transform 1 0 15916 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_179
timestamp 1649977179
transform 1 0 17572 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 1649977179
transform 1 0 18032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_194
timestamp 1649977179
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_211
timestamp 1649977179
transform 1 0 20516 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_116
timestamp 1649977179
transform 1 0 11776 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_128
timestamp 1649977179
transform 1 0 12880 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_140
timestamp 1649977179
transform 1 0 13984 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_152
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1649977179
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1649977179
transform 1 0 16836 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1649977179
transform 1 0 17204 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_180
timestamp 1649977179
transform 1 0 17664 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_186
timestamp 1649977179
transform 1 0 18216 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_191
timestamp 1649977179
transform 1 0 18676 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1649977179
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 1649977179
transform 1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_88
timestamp 1649977179
transform 1 0 9200 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_100
timestamp 1649977179
transform 1 0 10304 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_112
timestamp 1649977179
transform 1 0 11408 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_124
timestamp 1649977179
transform 1 0 12512 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_179
timestamp 1649977179
transform 1 0 17572 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_184
timestamp 1649977179
transform 1 0 18032 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 1649977179
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_202
timestamp 1649977179
transform 1 0 19688 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_207
timestamp 1649977179
transform 1 0 20148 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_212
timestamp 1649977179
transform 1 0 20608 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_216
timestamp 1649977179
transform 1 0 20976 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_23_92
timestamp 1649977179
transform 1 0 9568 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_104
timestamp 1649977179
transform 1 0 10672 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_117
timestamp 1649977179
transform 1 0 11868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_129
timestamp 1649977179
transform 1 0 12972 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_141
timestamp 1649977179
transform 1 0 14076 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_153
timestamp 1649977179
transform 1 0 15180 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_185
timestamp 1649977179
transform 1 0 18124 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_188
timestamp 1649977179
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_194
timestamp 1649977179
transform 1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1649977179
transform 1 0 20424 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_215
timestamp 1649977179
transform 1 0 20884 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_221
timestamp 1649977179
transform 1 0 21436 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_200
timestamp 1649977179
transform 1 0 19504 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 1649977179
transform 1 0 19964 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1649977179
transform 1 0 20424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1649977179
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_145
timestamp 1649977179
transform 1 0 14444 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_203
timestamp 1649977179
transform 1 0 19780 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_208
timestamp 1649977179
transform 1 0 20240 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_215
timestamp 1649977179
transform 1 0 20884 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_221
timestamp 1649977179
transform 1 0 21436 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_185
timestamp 1649977179
transform 1 0 18124 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_205
timestamp 1649977179
transform 1 0 19964 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1649977179
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_215
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_201
timestamp 1649977179
transform 1 0 19596 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1649977179
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_211
timestamp 1649977179
transform 1 0 20516 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_215
timestamp 1649977179
transform 1 0 20884 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_115
timestamp 1649977179
transform 1 0 11684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_127
timestamp 1649977179
transform 1 0 12788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_77
timestamp 1649977179
transform 1 0 8188 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_29_82
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_94
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_106
timestamp 1649977179
transform 1 0 10856 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_124
timestamp 1649977179
transform 1 0 12512 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_136
timestamp 1649977179
transform 1 0 13616 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_148
timestamp 1649977179
transform 1 0 14720 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1649977179
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_211
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_94
timestamp 1649977179
transform 1 0 9752 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_106
timestamp 1649977179
transform 1 0 10856 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_205
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_210
timestamp 1649977179
transform 1 0 20424 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_215
timestamp 1649977179
transform 1 0 20884 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_187
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_191
timestamp 1649977179
transform 1 0 18676 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_198
timestamp 1649977179
transform 1 0 19320 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_208
timestamp 1649977179
transform 1 0 20240 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_215
timestamp 1649977179
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_60
timestamp 1649977179
transform 1 0 6624 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_72
timestamp 1649977179
transform 1 0 7728 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_127
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_131
timestamp 1649977179
transform 1 0 13156 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_203
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_215
timestamp 1649977179
transform 1 0 20884 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_29
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_41
timestamp 1649977179
transform 1 0 4876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_49
timestamp 1649977179
transform 1 0 5612 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_71
timestamp 1649977179
transform 1 0 7636 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_83
timestamp 1649977179
transform 1 0 8740 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_85
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_97
timestamp 1649977179
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_141
timestamp 1649977179
transform 1 0 14076 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_153
timestamp 1649977179
transform 1 0 15180 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_165
timestamp 1649977179
transform 1 0 16284 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_175
timestamp 1649977179
transform 1 0 17204 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_183
timestamp 1649977179
transform 1 0 17940 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_194
timestamp 1649977179
transform 1 0 18952 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1649977179
transform 1 0 19228 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_203
timestamp 1649977179
transform 1 0 19780 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_209
timestamp 1649977179
transform 1 0 20332 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_215
timestamp 1649977179
transform 1 0 20884 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  _48_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6256 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _49_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18952 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _50_
timestamp 1649977179
transform -1 0 19504 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _51_
timestamp 1649977179
transform -1 0 20884 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _52_
timestamp 1649977179
transform -1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _53_
timestamp 1649977179
transform -1 0 20424 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _54_
timestamp 1649977179
transform -1 0 20424 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _55_
timestamp 1649977179
transform -1 0 19964 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _56_
timestamp 1649977179
transform -1 0 20884 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _57_
timestamp 1649977179
transform -1 0 20884 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _58_
timestamp 1649977179
transform -1 0 20884 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _59_
timestamp 1649977179
transform 1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _60_
timestamp 1649977179
transform -1 0 20424 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _61_
timestamp 1649977179
transform -1 0 20332 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _62_
timestamp 1649977179
transform -1 0 12512 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _63_
timestamp 1649977179
transform -1 0 20884 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _64_
timestamp 1649977179
transform -1 0 20424 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _65_
timestamp 1649977179
transform -1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _66_
timestamp 1649977179
transform -1 0 19780 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _67_
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _68_
timestamp 1649977179
transform -1 0 19320 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _69_
timestamp 1649977179
transform -1 0 6992 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _70_
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _71_
timestamp 1649977179
transform -1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _72_
timestamp 1649977179
transform -1 0 13340 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _73_
timestamp 1649977179
transform -1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _74_
timestamp 1649977179
transform -1 0 5152 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _75_
timestamp 1649977179
transform -1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _76_
timestamp 1649977179
transform -1 0 6624 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _77_
timestamp 1649977179
transform -1 0 5704 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _78_
timestamp 1649977179
transform -1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _79_
timestamp 1649977179
transform -1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _80_
timestamp 1649977179
transform 1 0 14996 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _81_
timestamp 1649977179
transform -1 0 10212 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _82_
timestamp 1649977179
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _83_
timestamp 1649977179
transform -1 0 5152 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _84_
timestamp 1649977179
transform -1 0 10304 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _85_
timestamp 1649977179
transform -1 0 11224 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _86_
timestamp 1649977179
transform -1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _87_
timestamp 1649977179
transform -1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _88_
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_bottom_track_1.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 16192 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_mem_bottom_track_1.prog_clk
timestamp 1649977179
transform 1 0 16376 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 18216 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 14996 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform -1 0 8648 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform 1 0 12420 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform -1 0 6624 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 20700 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 7912 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform -1 0 13616 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 17940 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform -1 0 8648 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform -1 0 18952 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform 1 0 18584 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform 1 0 15548 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform -1 0 20424 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform -1 0 8004 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 20332 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 17112 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform 1 0 16100 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform -1 0 6992 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform -1 0 9016 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform 1 0 20700 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform -1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform -1 0 7636 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform -1 0 17480 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform -1 0 12144 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform -1 0 20056 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform 1 0 20608 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform 1 0 13892 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform -1 0 9568 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform -1 0 6072 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform -1 0 7728 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform -1 0 21068 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform -1 0 13800 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 6072 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform 1 0 1564 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 17296 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 14812 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 17020 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform 1 0 16100 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 18032 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform 1 0 17756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 16744 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 18216 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 19964 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform 1 0 19412 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 21160 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 10028 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 8096 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 7268 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 6808 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 1656 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 4232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 4692 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform -1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform -1 0 5336 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform -1 0 5152 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform -1 0 6624 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 5612 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform -1 0 6992 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform -1 0 1656 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 2116 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 2576 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform -1 0 2576 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 3772 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform -1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19412 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform 1 0 20516 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform 1 0 19412 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform 1 0 19412 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input48
timestamp 1649977179
transform -1 0 18952 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input49
timestamp 1649977179
transform 1 0 20516 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input50
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 4416 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform -1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18032 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21252 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18400 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 20148 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19504 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_bottom_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 17572 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14628 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16376 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16744 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18400 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 19780 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 21436 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 19780 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 16284 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 16008 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 13800 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12052 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 8648 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7728 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7912 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 9568 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12328 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15732 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 16928 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13892 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13708 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12328 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11224 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_28.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_30.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8188 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 9200 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_32.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 10488 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 12236 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_34.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12512 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_36.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14720 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_right_track_38.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_1.mux_l2_in_0__108 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18676 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19412 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12052 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20424 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_5.mux_l2_in_0__110
timestamp 1649977179
transform 1 0 18584 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17664 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 13340 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19320 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_9.mux_l2_in_0__111
timestamp 1649977179
transform -1 0 15916 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18124 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 10212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 20516 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_bottom_track_25.mux_l2_in_0__109
timestamp 1649977179
transform -1 0 18952 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_bottom_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 19688 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_bottom_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7728 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_1_
timestamp 1649977179
transform -1 0 17480 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 15824 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_0_
timestamp 1649977179
transform 1 0 17664 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_0.mux_l2_in_1__112
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l2_in_1_
timestamp 1649977179
transform -1 0 16008 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_0.mux_l3_in_0_
timestamp 1649977179
transform 1 0 16192 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15548 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 20148 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l1_in_1_
timestamp 1649977179
transform -1 0 20332 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 20516 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_2.mux_l2_in_1__118
timestamp 1649977179
transform -1 0 6348 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 20884 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_2.mux_l3_in_0_
timestamp 1649977179
transform 1 0 20332 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l1_in_2_
timestamp 1649977179
transform -1 0 17940 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16928 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_4.mux_l2_in_1__105
timestamp 1649977179
transform -1 0 16376 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l2_in_1_
timestamp 1649977179
transform 1 0 18308 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 18952 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19136 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 17204 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_0_
timestamp 1649977179
transform 1 0 16192 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_6.mux_l2_in_1__106
timestamp 1649977179
transform -1 0 7728 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l2_in_1_
timestamp 1649977179
transform -1 0 15732 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 16008 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_8.mux_l1_in_1__107
timestamp 1649977179
transform -1 0 6256 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 13248 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13800 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_10.mux_l2_in_0__113
timestamp 1649977179
transform -1 0 6072 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11776 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_12.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_12.mux_l2_in_0__114
timestamp 1649977179
transform -1 0 6072 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9200 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9568 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_14.mux_l2_in_0__115
timestamp 1649977179
transform -1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9568 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_16.mux_l2_in_0__116
timestamp 1649977179
transform 1 0 12052 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11776 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l1_in_0_
timestamp 1649977179
transform -1 0 13708 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_18.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 15732 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14628 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14812 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16100 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_20.mux_l2_in_0__95
timestamp 1649977179
transform 1 0 17388 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20240 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l1_in_0_
timestamp 1649977179
transform -1 0 18032 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_22.mux_l2_in_0__96
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_22.mux_l2_in_0_
timestamp 1649977179
transform 1 0 18308 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18492 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13892 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_24.mux_l1_in_1__97
timestamp 1649977179
transform -1 0 6808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13892 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 20148 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_26.mux_l2_in_0_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_26.mux_l2_in_0__98
timestamp 1649977179
transform -1 0 6072 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 11684 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l1_in_0_
timestamp 1649977179
transform -1 0 7636 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_28.mux_l2_in_0__99
timestamp 1649977179
transform -1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_28.mux_l2_in_0_
timestamp 1649977179
transform -1 0 8648 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_28.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 8648 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_30.mux_l2_in_0__100
timestamp 1649977179
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_30.mux_l2_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_30.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 9752 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10212 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_32.mux_l2_in_0__101
timestamp 1649977179
transform -1 0 12696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_32.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12144 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_32.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 12236 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_34.mux_l2_in_0__102
timestamp 1649977179
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_34.mux_l2_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_34.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19780 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15916 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_36.mux_l2_in_0__103
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_36.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16284 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_36.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17756 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_right_track_38.mux_l2_in_0__104
timestamp 1649977179
transform 1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_right_track_38.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18492 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_right_track_38.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18676 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output53 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15088 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output54
timestamp 1649977179
transform -1 0 1748 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output55
timestamp 1649977179
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output56
timestamp 1649977179
transform 1 0 20516 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output57
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output58
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output59
timestamp 1649977179
transform 1 0 21068 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output60
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform 1 0 20516 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 19412 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 20148 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform 1 0 21068 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 12052 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform 1 0 19320 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 12512 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform 1 0 14076 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform 1 0 18584 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform -1 0 13800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 11776 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 17664 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 13432 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform 1 0 9844 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform 1 0 17664 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform 1 0 13432 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform 1 0 20884 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 14144
box -38 -48 1142 592
<< labels >>
rlabel metal2 s 5722 22200 5778 23000 6 SC_IN_TOP
port 0 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 SC_OUT_BOT
port 1 nsew signal tristate
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 2 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 3 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 3 nsew power input
rlabel metal2 s 202 0 258 800 6 bottom_left_grid_pin_1_
port 4 nsew signal input
rlabel metal2 s 17222 22200 17278 23000 6 ccff_head
port 5 nsew signal input
rlabel metal3 s 0 11432 800 11552 6 ccff_tail
port 6 nsew signal tristate
rlabel metal3 s 22200 3816 23000 3936 6 chanx_right_in[0]
port 7 nsew signal input
rlabel metal3 s 22200 8304 23000 8424 6 chanx_right_in[10]
port 8 nsew signal input
rlabel metal3 s 22200 8848 23000 8968 6 chanx_right_in[11]
port 9 nsew signal input
rlabel metal3 s 22200 9256 23000 9376 6 chanx_right_in[12]
port 10 nsew signal input
rlabel metal3 s 22200 9664 23000 9784 6 chanx_right_in[13]
port 11 nsew signal input
rlabel metal3 s 22200 10208 23000 10328 6 chanx_right_in[14]
port 12 nsew signal input
rlabel metal3 s 22200 10616 23000 10736 6 chanx_right_in[15]
port 13 nsew signal input
rlabel metal3 s 22200 11160 23000 11280 6 chanx_right_in[16]
port 14 nsew signal input
rlabel metal3 s 22200 11568 23000 11688 6 chanx_right_in[17]
port 15 nsew signal input
rlabel metal3 s 22200 11976 23000 12096 6 chanx_right_in[18]
port 16 nsew signal input
rlabel metal3 s 22200 12520 23000 12640 6 chanx_right_in[19]
port 17 nsew signal input
rlabel metal3 s 22200 4224 23000 4344 6 chanx_right_in[1]
port 18 nsew signal input
rlabel metal3 s 22200 4632 23000 4752 6 chanx_right_in[2]
port 19 nsew signal input
rlabel metal3 s 22200 5176 23000 5296 6 chanx_right_in[3]
port 20 nsew signal input
rlabel metal3 s 22200 5584 23000 5704 6 chanx_right_in[4]
port 21 nsew signal input
rlabel metal3 s 22200 5992 23000 6112 6 chanx_right_in[5]
port 22 nsew signal input
rlabel metal3 s 22200 6536 23000 6656 6 chanx_right_in[6]
port 23 nsew signal input
rlabel metal3 s 22200 6944 23000 7064 6 chanx_right_in[7]
port 24 nsew signal input
rlabel metal3 s 22200 7488 23000 7608 6 chanx_right_in[8]
port 25 nsew signal input
rlabel metal3 s 22200 7896 23000 8016 6 chanx_right_in[9]
port 26 nsew signal input
rlabel metal3 s 22200 12928 23000 13048 6 chanx_right_out[0]
port 27 nsew signal tristate
rlabel metal3 s 22200 17552 23000 17672 6 chanx_right_out[10]
port 28 nsew signal tristate
rlabel metal3 s 22200 17960 23000 18080 6 chanx_right_out[11]
port 29 nsew signal tristate
rlabel metal3 s 22200 18504 23000 18624 6 chanx_right_out[12]
port 30 nsew signal tristate
rlabel metal3 s 22200 18912 23000 19032 6 chanx_right_out[13]
port 31 nsew signal tristate
rlabel metal3 s 22200 19320 23000 19440 6 chanx_right_out[14]
port 32 nsew signal tristate
rlabel metal3 s 22200 19864 23000 19984 6 chanx_right_out[15]
port 33 nsew signal tristate
rlabel metal3 s 22200 20272 23000 20392 6 chanx_right_out[16]
port 34 nsew signal tristate
rlabel metal3 s 22200 20816 23000 20936 6 chanx_right_out[17]
port 35 nsew signal tristate
rlabel metal3 s 22200 21224 23000 21344 6 chanx_right_out[18]
port 36 nsew signal tristate
rlabel metal3 s 22200 21632 23000 21752 6 chanx_right_out[19]
port 37 nsew signal tristate
rlabel metal3 s 22200 13472 23000 13592 6 chanx_right_out[1]
port 38 nsew signal tristate
rlabel metal3 s 22200 13880 23000 14000 6 chanx_right_out[2]
port 39 nsew signal tristate
rlabel metal3 s 22200 14288 23000 14408 6 chanx_right_out[3]
port 40 nsew signal tristate
rlabel metal3 s 22200 14832 23000 14952 6 chanx_right_out[4]
port 41 nsew signal tristate
rlabel metal3 s 22200 15240 23000 15360 6 chanx_right_out[5]
port 42 nsew signal tristate
rlabel metal3 s 22200 15648 23000 15768 6 chanx_right_out[6]
port 43 nsew signal tristate
rlabel metal3 s 22200 16192 23000 16312 6 chanx_right_out[7]
port 44 nsew signal tristate
rlabel metal3 s 22200 16600 23000 16720 6 chanx_right_out[8]
port 45 nsew signal tristate
rlabel metal3 s 22200 17144 23000 17264 6 chanx_right_out[9]
port 46 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 chany_bottom_in[0]
port 47 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 chany_bottom_in[10]
port 48 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 chany_bottom_in[11]
port 49 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 chany_bottom_in[12]
port 50 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 chany_bottom_in[13]
port 51 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 chany_bottom_in[14]
port 52 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 chany_bottom_in[15]
port 53 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 chany_bottom_in[16]
port 54 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 chany_bottom_in[17]
port 55 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 chany_bottom_in[18]
port 56 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 chany_bottom_in[19]
port 57 nsew signal input
rlabel metal2 s 1214 0 1270 800 6 chany_bottom_in[1]
port 58 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 chany_bottom_in[2]
port 59 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 chany_bottom_in[3]
port 60 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 chany_bottom_in[4]
port 61 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 chany_bottom_in[5]
port 62 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 chany_bottom_in[6]
port 63 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 chany_bottom_in[7]
port 64 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 chany_bottom_in[8]
port 65 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 chany_bottom_in[9]
port 66 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 chany_bottom_out[0]
port 67 nsew signal tristate
rlabel metal2 s 17130 0 17186 800 6 chany_bottom_out[10]
port 68 nsew signal tristate
rlabel metal2 s 17682 0 17738 800 6 chany_bottom_out[11]
port 69 nsew signal tristate
rlabel metal2 s 18234 0 18290 800 6 chany_bottom_out[12]
port 70 nsew signal tristate
rlabel metal2 s 18786 0 18842 800 6 chany_bottom_out[13]
port 71 nsew signal tristate
rlabel metal2 s 19338 0 19394 800 6 chany_bottom_out[14]
port 72 nsew signal tristate
rlabel metal2 s 19890 0 19946 800 6 chany_bottom_out[15]
port 73 nsew signal tristate
rlabel metal2 s 20442 0 20498 800 6 chany_bottom_out[16]
port 74 nsew signal tristate
rlabel metal2 s 20994 0 21050 800 6 chany_bottom_out[17]
port 75 nsew signal tristate
rlabel metal2 s 21546 0 21602 800 6 chany_bottom_out[18]
port 76 nsew signal tristate
rlabel metal2 s 22098 0 22154 800 6 chany_bottom_out[19]
port 77 nsew signal tristate
rlabel metal2 s 12162 0 12218 800 6 chany_bottom_out[1]
port 78 nsew signal tristate
rlabel metal2 s 12714 0 12770 800 6 chany_bottom_out[2]
port 79 nsew signal tristate
rlabel metal2 s 13266 0 13322 800 6 chany_bottom_out[3]
port 80 nsew signal tristate
rlabel metal2 s 13818 0 13874 800 6 chany_bottom_out[4]
port 81 nsew signal tristate
rlabel metal2 s 14370 0 14426 800 6 chany_bottom_out[5]
port 82 nsew signal tristate
rlabel metal2 s 14922 0 14978 800 6 chany_bottom_out[6]
port 83 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 chany_bottom_out[7]
port 84 nsew signal tristate
rlabel metal2 s 16026 0 16082 800 6 chany_bottom_out[8]
port 85 nsew signal tristate
rlabel metal2 s 16578 0 16634 800 6 chany_bottom_out[9]
port 86 nsew signal tristate
rlabel metal3 s 22200 22176 23000 22296 6 prog_clk_0_E_in
port 87 nsew signal input
rlabel metal3 s 22200 144 23000 264 6 right_bottom_grid_pin_34_
port 88 nsew signal input
rlabel metal3 s 22200 552 23000 672 6 right_bottom_grid_pin_35_
port 89 nsew signal input
rlabel metal3 s 22200 960 23000 1080 6 right_bottom_grid_pin_36_
port 90 nsew signal input
rlabel metal3 s 22200 1504 23000 1624 6 right_bottom_grid_pin_37_
port 91 nsew signal input
rlabel metal3 s 22200 1912 23000 2032 6 right_bottom_grid_pin_38_
port 92 nsew signal input
rlabel metal3 s 22200 2320 23000 2440 6 right_bottom_grid_pin_39_
port 93 nsew signal input
rlabel metal3 s 22200 2864 23000 2984 6 right_bottom_grid_pin_40_
port 94 nsew signal input
rlabel metal3 s 22200 3272 23000 3392 6 right_bottom_grid_pin_41_
port 95 nsew signal input
rlabel metal3 s 22200 22584 23000 22704 6 right_top_grid_pin_1_
port 96 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
