magic
tech sky130A
magscale 1 2
timestamp 1650893844
<< viali >>
rect 5641 20553 5675 20587
rect 9137 20553 9171 20587
rect 13277 20553 13311 20587
rect 14197 20553 14231 20587
rect 15301 20553 15335 20587
rect 16773 20553 16807 20587
rect 17877 20553 17911 20587
rect 19349 20553 19383 20587
rect 19901 20553 19935 20587
rect 7941 20485 7975 20519
rect 9934 20485 9968 20519
rect 2329 20417 2363 20451
rect 4997 20417 5031 20451
rect 6745 20417 6779 20451
rect 8585 20417 8619 20451
rect 8953 20417 8987 20451
rect 11529 20417 11563 20451
rect 12725 20417 12759 20451
rect 13461 20417 13495 20451
rect 14381 20417 14415 20451
rect 14933 20417 14967 20451
rect 15485 20417 15519 20451
rect 16037 20417 16071 20451
rect 16957 20417 16991 20451
rect 17509 20417 17543 20451
rect 18061 20417 18095 20451
rect 18613 20417 18647 20451
rect 19533 20417 19567 20451
rect 20085 20417 20119 20451
rect 2053 20349 2087 20383
rect 3157 20349 3191 20383
rect 3433 20349 3467 20383
rect 3801 20349 3835 20383
rect 4077 20349 4111 20383
rect 5733 20349 5767 20383
rect 5917 20349 5951 20383
rect 6469 20349 6503 20383
rect 9689 20349 9723 20383
rect 21097 20349 21131 20383
rect 21373 20349 21407 20383
rect 14749 20281 14783 20315
rect 15853 20281 15887 20315
rect 17325 20281 17359 20315
rect 18429 20281 18463 20315
rect 5273 20213 5307 20247
rect 7389 20213 7423 20247
rect 11069 20213 11103 20247
rect 12173 20213 12207 20247
rect 12541 20213 12575 20247
rect 10057 20009 10091 20043
rect 15025 20009 15059 20043
rect 15577 20009 15611 20043
rect 16957 20009 16991 20043
rect 17417 20009 17451 20043
rect 18337 20009 18371 20043
rect 19809 20009 19843 20043
rect 13277 19941 13311 19975
rect 13737 19941 13771 19975
rect 2053 19873 2087 19907
rect 2881 19873 2915 19907
rect 9137 19873 9171 19907
rect 20729 19873 20763 19907
rect 2329 19805 2363 19839
rect 2605 19805 2639 19839
rect 5181 19805 5215 19839
rect 6662 19805 6696 19839
rect 6929 19805 6963 19839
rect 8585 19805 8619 19839
rect 11437 19805 11471 19839
rect 11713 19805 11747 19839
rect 12633 19805 12667 19839
rect 13553 19805 13587 19839
rect 14105 19805 14139 19839
rect 14565 19805 14599 19839
rect 15209 19805 15243 19839
rect 15761 19805 15795 19839
rect 16221 19805 16255 19839
rect 16497 19805 16531 19839
rect 17141 19805 17175 19839
rect 17601 19805 17635 19839
rect 18521 19805 18555 19839
rect 19349 19805 19383 19839
rect 19625 19805 19659 19839
rect 21373 19805 21407 19839
rect 4914 19737 4948 19771
rect 8340 19737 8374 19771
rect 11192 19737 11226 19771
rect 12357 19737 12391 19771
rect 3801 19669 3835 19703
rect 5549 19669 5583 19703
rect 7205 19669 7239 19703
rect 9321 19669 9355 19703
rect 9413 19669 9447 19703
rect 9781 19669 9815 19703
rect 14289 19669 14323 19703
rect 14749 19669 14783 19703
rect 16037 19669 16071 19703
rect 17969 19669 18003 19703
rect 18797 19669 18831 19703
rect 2605 19465 2639 19499
rect 5089 19465 5123 19499
rect 6745 19465 6779 19499
rect 7389 19465 7423 19499
rect 8125 19465 8159 19499
rect 9413 19465 9447 19499
rect 12817 19465 12851 19499
rect 13277 19465 13311 19499
rect 13921 19465 13955 19499
rect 15209 19465 15243 19499
rect 15669 19465 15703 19499
rect 15945 19465 15979 19499
rect 16681 19465 16715 19499
rect 17141 19465 17175 19499
rect 17601 19465 17635 19499
rect 18245 19465 18279 19499
rect 18521 19465 18555 19499
rect 19165 19465 19199 19499
rect 20269 19465 20303 19499
rect 20821 19465 20855 19499
rect 1961 19329 1995 19363
rect 3718 19329 3752 19363
rect 3985 19329 4019 19363
rect 4353 19329 4387 19363
rect 5457 19329 5491 19363
rect 6561 19329 6595 19363
rect 7481 19329 7515 19363
rect 8493 19329 8527 19363
rect 8585 19329 8619 19363
rect 10526 19329 10560 19363
rect 10793 19329 10827 19363
rect 11805 19329 11839 19363
rect 12449 19329 12483 19363
rect 13001 19329 13035 19363
rect 13461 19329 13495 19363
rect 13737 19329 13771 19363
rect 14841 19329 14875 19363
rect 15485 19329 15519 19363
rect 16129 19329 16163 19363
rect 16865 19329 16899 19363
rect 17325 19329 17359 19363
rect 17785 19329 17819 19363
rect 18061 19329 18095 19363
rect 18705 19329 18739 19363
rect 18981 19329 19015 19363
rect 19625 19329 19659 19363
rect 20085 19329 20119 19363
rect 20637 19329 20671 19363
rect 21373 19329 21407 19363
rect 2237 19261 2271 19295
rect 5549 19261 5583 19295
rect 5641 19261 5675 19295
rect 7297 19261 7331 19295
rect 8769 19261 8803 19295
rect 14565 19261 14599 19295
rect 14749 19261 14783 19295
rect 4537 19193 4571 19227
rect 19441 19193 19475 19227
rect 7849 19125 7883 19159
rect 11069 19125 11103 19159
rect 21189 19125 21223 19159
rect 1777 18921 1811 18955
rect 6745 18921 6779 18955
rect 8953 18921 8987 18955
rect 10609 18921 10643 18955
rect 16037 18921 16071 18955
rect 18613 18921 18647 18955
rect 21189 18921 21223 18955
rect 1501 18853 1535 18887
rect 3985 18853 4019 18887
rect 17877 18853 17911 18887
rect 18153 18853 18187 18887
rect 20545 18853 20579 18887
rect 2881 18785 2915 18819
rect 4537 18785 4571 18819
rect 4629 18785 4663 18819
rect 9505 18785 9539 18819
rect 9597 18785 9631 18819
rect 11989 18785 12023 18819
rect 2421 18717 2455 18751
rect 3801 18717 3835 18751
rect 5365 18717 5399 18751
rect 7021 18717 7055 18751
rect 8585 18717 8619 18751
rect 11253 18717 11287 18751
rect 12817 18717 12851 18751
rect 15761 18717 15795 18751
rect 16221 18717 16255 18751
rect 16773 18717 16807 18751
rect 17693 18717 17727 18751
rect 18337 18717 18371 18751
rect 18797 18717 18831 18751
rect 19257 18717 19291 18751
rect 19717 18717 19751 18751
rect 20729 18717 20763 18751
rect 21005 18717 21039 18751
rect 5610 18649 5644 18683
rect 9689 18649 9723 18683
rect 15516 18649 15550 18683
rect 2973 18581 3007 18615
rect 3065 18581 3099 18615
rect 3433 18581 3467 18615
rect 4721 18581 4755 18615
rect 5089 18581 5123 18615
rect 7665 18581 7699 18615
rect 7941 18581 7975 18615
rect 10057 18581 10091 18615
rect 12081 18581 12115 18615
rect 12173 18581 12207 18615
rect 12541 18581 12575 18615
rect 13461 18581 13495 18615
rect 14381 18581 14415 18615
rect 17417 18581 17451 18615
rect 19441 18581 19475 18615
rect 19901 18581 19935 18615
rect 1777 18377 1811 18411
rect 2697 18377 2731 18411
rect 3617 18377 3651 18411
rect 3985 18377 4019 18411
rect 4629 18377 4663 18411
rect 6561 18377 6595 18411
rect 10057 18377 10091 18411
rect 14933 18377 14967 18411
rect 16681 18377 16715 18411
rect 20177 18377 20211 18411
rect 21281 18377 21315 18411
rect 7472 18309 7506 18343
rect 12848 18309 12882 18343
rect 15945 18309 15979 18343
rect 2421 18241 2455 18275
rect 3341 18241 3375 18275
rect 4077 18241 4111 18275
rect 5742 18241 5776 18275
rect 6009 18241 6043 18275
rect 6377 18241 6411 18275
rect 9045 18241 9079 18275
rect 10333 18241 10367 18275
rect 13093 18241 13127 18275
rect 13737 18241 13771 18275
rect 13829 18241 13863 18275
rect 14565 18241 14599 18275
rect 15301 18241 15335 18275
rect 17794 18241 17828 18275
rect 18061 18241 18095 18275
rect 18337 18241 18371 18275
rect 19441 18241 19475 18275
rect 19901 18241 19935 18275
rect 20361 18241 20395 18275
rect 20821 18241 20855 18275
rect 21097 18241 21131 18275
rect 4169 18173 4203 18207
rect 7205 18173 7239 18207
rect 14013 18173 14047 18207
rect 15393 18173 15427 18207
rect 15577 18173 15611 18207
rect 19257 18105 19291 18139
rect 19717 18105 19751 18139
rect 20637 18105 20671 18139
rect 1501 18037 1535 18071
rect 8585 18037 8619 18071
rect 9689 18037 9723 18071
rect 10977 18037 11011 18071
rect 11713 18037 11747 18071
rect 13369 18037 13403 18071
rect 14381 18037 14415 18071
rect 18981 18037 19015 18071
rect 1593 17833 1627 17867
rect 10609 17833 10643 17867
rect 12265 17833 12299 17867
rect 14841 17833 14875 17867
rect 16497 17833 16531 17867
rect 19441 17833 19475 17867
rect 20637 17833 20671 17867
rect 21097 17833 21131 17867
rect 5641 17765 5675 17799
rect 18889 17765 18923 17799
rect 6193 17697 6227 17731
rect 7389 17697 7423 17731
rect 9229 17697 9263 17731
rect 13093 17697 13127 17731
rect 14289 17697 14323 17731
rect 15117 17697 15151 17731
rect 17693 17697 17727 17731
rect 18245 17697 18279 17731
rect 1409 17629 1443 17663
rect 2513 17629 2547 17663
rect 3433 17629 3467 17663
rect 5181 17629 5215 17663
rect 8585 17629 8619 17663
rect 10885 17629 10919 17663
rect 11152 17629 11186 17663
rect 12909 17629 12943 17663
rect 14473 17629 14507 17663
rect 16773 17629 16807 17663
rect 19257 17629 19291 17663
rect 20361 17629 20395 17663
rect 20821 17629 20855 17663
rect 21281 17629 21315 17663
rect 1869 17561 1903 17595
rect 4914 17561 4948 17595
rect 6101 17561 6135 17595
rect 7205 17561 7239 17595
rect 9496 17561 9530 17595
rect 13553 17561 13587 17595
rect 15362 17561 15396 17595
rect 18521 17561 18555 17595
rect 19717 17561 19751 17595
rect 2789 17493 2823 17527
rect 3801 17493 3835 17527
rect 6009 17493 6043 17527
rect 6837 17493 6871 17527
rect 7297 17493 7331 17527
rect 7941 17493 7975 17527
rect 12541 17493 12575 17527
rect 13001 17493 13035 17527
rect 14381 17493 14415 17527
rect 17417 17493 17451 17527
rect 18429 17493 18463 17527
rect 20177 17493 20211 17527
rect 1685 17289 1719 17323
rect 5365 17289 5399 17323
rect 6929 17289 6963 17323
rect 9045 17289 9079 17323
rect 10057 17289 10091 17323
rect 10793 17289 10827 17323
rect 11989 17289 12023 17323
rect 13001 17289 13035 17323
rect 14657 17289 14691 17323
rect 4270 17221 4304 17255
rect 8042 17221 8076 17255
rect 9597 17221 9631 17255
rect 21281 17221 21315 17255
rect 1869 17153 1903 17187
rect 2513 17153 2547 17187
rect 2605 17153 2639 17187
rect 5089 17153 5123 17187
rect 6009 17153 6043 17187
rect 6653 17153 6687 17187
rect 8861 17153 8895 17187
rect 9689 17153 9723 17187
rect 10701 17153 10735 17187
rect 11713 17153 11747 17187
rect 12357 17153 12391 17187
rect 13369 17153 13403 17187
rect 13461 17153 13495 17187
rect 14013 17153 14047 17187
rect 15301 17153 15335 17187
rect 16681 17153 16715 17187
rect 19093 17153 19127 17187
rect 19349 17153 19383 17187
rect 19901 17153 19935 17187
rect 20821 17153 20855 17187
rect 2697 17085 2731 17119
rect 4537 17085 4571 17119
rect 8309 17085 8343 17119
rect 9413 17085 9447 17119
rect 10977 17085 11011 17119
rect 12449 17085 12483 17119
rect 12633 17085 12667 17119
rect 13553 17085 13587 17119
rect 15117 17085 15151 17119
rect 15209 17085 15243 17119
rect 16129 17085 16163 17119
rect 3157 17017 3191 17051
rect 6469 17017 6503 17051
rect 15669 17017 15703 17051
rect 17601 17017 17635 17051
rect 17969 17017 18003 17051
rect 2145 16949 2179 16983
rect 4905 16949 4939 16983
rect 10333 16949 10367 16983
rect 11529 16949 11563 16983
rect 17325 16949 17359 16983
rect 20545 16949 20579 16983
rect 21005 16949 21039 16983
rect 3801 16745 3835 16779
rect 6285 16745 6319 16779
rect 7481 16745 7515 16779
rect 8493 16745 8527 16779
rect 15761 16745 15795 16779
rect 16865 16745 16899 16779
rect 19257 16745 19291 16779
rect 14105 16677 14139 16711
rect 4353 16609 4387 16643
rect 4905 16609 4939 16643
rect 7941 16609 7975 16643
rect 8125 16609 8159 16643
rect 10333 16609 10367 16643
rect 11897 16609 11931 16643
rect 12449 16609 12483 16643
rect 15485 16609 15519 16643
rect 16313 16609 16347 16643
rect 17141 16609 17175 16643
rect 18797 16609 18831 16643
rect 19717 16609 19751 16643
rect 19809 16609 19843 16643
rect 1409 16541 1443 16575
rect 2237 16541 2271 16575
rect 2697 16541 2731 16575
rect 3341 16541 3375 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 6561 16541 6595 16575
rect 10077 16541 10111 16575
rect 11805 16541 11839 16575
rect 12725 16541 12759 16575
rect 15229 16541 15263 16575
rect 17408 16541 17442 16575
rect 20269 16541 20303 16575
rect 20913 16541 20947 16575
rect 21373 16541 21407 16575
rect 5150 16473 5184 16507
rect 12633 16473 12667 16507
rect 16129 16473 16163 16507
rect 19625 16473 19659 16507
rect 1593 16405 1627 16439
rect 2053 16405 2087 16439
rect 7205 16405 7239 16439
rect 7849 16405 7883 16439
rect 8953 16405 8987 16439
rect 10609 16405 10643 16439
rect 11345 16405 11379 16439
rect 11713 16405 11747 16439
rect 13093 16405 13127 16439
rect 13369 16405 13403 16439
rect 16221 16405 16255 16439
rect 18521 16405 18555 16439
rect 21189 16405 21223 16439
rect 2145 16201 2179 16235
rect 3157 16201 3191 16235
rect 3709 16201 3743 16235
rect 5365 16201 5399 16235
rect 6377 16201 6411 16235
rect 8309 16201 8343 16235
rect 13461 16201 13495 16235
rect 13921 16201 13955 16235
rect 15301 16201 15335 16235
rect 15945 16201 15979 16235
rect 16681 16201 16715 16235
rect 19901 16201 19935 16235
rect 20177 16201 20211 16235
rect 20729 16201 20763 16235
rect 2605 16133 2639 16167
rect 6009 16133 6043 16167
rect 18788 16133 18822 16167
rect 1409 16065 1443 16099
rect 1961 16065 1995 16099
rect 3341 16065 3375 16099
rect 3985 16065 4019 16099
rect 5273 16065 5307 16099
rect 6745 16065 6779 16099
rect 7389 16065 7423 16099
rect 9597 16065 9631 16099
rect 10241 16065 10275 16099
rect 10885 16065 10919 16099
rect 12653 16065 12687 16099
rect 12909 16065 12943 16099
rect 13553 16065 13587 16099
rect 14565 16065 14599 16099
rect 17805 16065 17839 16099
rect 18061 16065 18095 16099
rect 18521 16065 18555 16099
rect 20361 16065 20395 16099
rect 5457 15997 5491 16031
rect 6837 15997 6871 16031
rect 6929 15997 6963 16031
rect 10333 15997 10367 16031
rect 10425 15997 10459 16031
rect 13277 15997 13311 16031
rect 14657 15997 14691 16031
rect 14749 15997 14783 16031
rect 15761 15997 15795 16031
rect 15853 15997 15887 16031
rect 2789 15929 2823 15963
rect 4905 15929 4939 15963
rect 14197 15929 14231 15963
rect 16313 15929 16347 15963
rect 21005 15929 21039 15963
rect 1593 15861 1627 15895
rect 4629 15861 4663 15895
rect 7573 15861 7607 15895
rect 9873 15861 9907 15895
rect 11529 15861 11563 15895
rect 2053 15657 2087 15691
rect 2697 15657 2731 15691
rect 3249 15657 3283 15691
rect 4353 15657 4387 15691
rect 8585 15657 8619 15691
rect 10333 15657 10367 15691
rect 13737 15657 13771 15691
rect 17141 15657 17175 15691
rect 18429 15657 18463 15691
rect 18889 15657 18923 15691
rect 20269 15589 20303 15623
rect 20637 15589 20671 15623
rect 5273 15521 5307 15555
rect 7941 15521 7975 15555
rect 8953 15521 8987 15555
rect 11897 15521 11931 15555
rect 13185 15521 13219 15555
rect 17877 15521 17911 15555
rect 19717 15521 19751 15555
rect 19901 15521 19935 15555
rect 1409 15453 1443 15487
rect 2237 15453 2271 15487
rect 2513 15453 2547 15487
rect 3065 15453 3099 15487
rect 3893 15453 3927 15487
rect 4997 15453 5031 15487
rect 7021 15453 7055 15487
rect 8401 15453 8435 15487
rect 10977 15453 11011 15487
rect 11805 15453 11839 15487
rect 12541 15453 12575 15487
rect 13369 15453 13403 15487
rect 15025 15453 15059 15487
rect 18705 15453 18739 15487
rect 9198 15385 9232 15419
rect 15669 15385 15703 15419
rect 17969 15385 18003 15419
rect 21005 15385 21039 15419
rect 1593 15317 1627 15351
rect 4077 15317 4111 15351
rect 7297 15317 7331 15351
rect 7665 15317 7699 15351
rect 7757 15317 7791 15351
rect 10793 15317 10827 15351
rect 11345 15317 11379 15351
rect 11713 15317 11747 15351
rect 12357 15317 12391 15351
rect 13277 15317 13311 15351
rect 14381 15317 14415 15351
rect 15301 15317 15335 15351
rect 18061 15317 18095 15351
rect 19257 15317 19291 15351
rect 19625 15317 19659 15351
rect 2053 15113 2087 15147
rect 4169 15113 4203 15147
rect 4629 15113 4663 15147
rect 6377 15113 6411 15147
rect 8493 15113 8527 15147
rect 9229 15113 9263 15147
rect 9597 15113 9631 15147
rect 10701 15113 10735 15147
rect 11161 15113 11195 15147
rect 11805 15113 11839 15147
rect 11897 15113 11931 15147
rect 12265 15113 12299 15147
rect 12541 15113 12575 15147
rect 13093 15113 13127 15147
rect 13461 15113 13495 15147
rect 15485 15113 15519 15147
rect 16681 15113 16715 15147
rect 17693 15113 17727 15147
rect 19441 15113 19475 15147
rect 21097 15113 21131 15147
rect 7380 15045 7414 15079
rect 9137 15045 9171 15079
rect 10057 15045 10091 15079
rect 10793 15045 10827 15079
rect 14372 15045 14406 15079
rect 1685 14977 1719 15011
rect 2237 14977 2271 15011
rect 2789 14977 2823 15011
rect 3045 14977 3079 15011
rect 5742 14977 5776 15011
rect 6009 14977 6043 15011
rect 6561 14977 6595 15011
rect 7113 14977 7147 15011
rect 12725 14977 12759 15011
rect 13553 14977 13587 15011
rect 14105 14977 14139 15011
rect 17049 14977 17083 15011
rect 18061 14977 18095 15011
rect 18328 14977 18362 15011
rect 19717 14977 19751 15011
rect 9045 14909 9079 14943
rect 10609 14909 10643 14943
rect 11713 14909 11747 14943
rect 13737 14909 13771 14943
rect 16221 14909 16255 14943
rect 17141 14909 17175 14943
rect 17233 14909 17267 14943
rect 20729 14841 20763 14875
rect 1501 14773 1535 14807
rect 20361 14773 20395 14807
rect 2053 14569 2087 14603
rect 5457 14569 5491 14603
rect 6377 14569 6411 14603
rect 8493 14569 8527 14603
rect 10149 14569 10183 14603
rect 12265 14569 12299 14603
rect 14105 14569 14139 14603
rect 18153 14569 18187 14603
rect 21005 14569 21039 14603
rect 20177 14501 20211 14535
rect 3341 14433 3375 14467
rect 5181 14433 5215 14467
rect 14657 14433 14691 14467
rect 17509 14433 17543 14467
rect 18429 14433 18463 14467
rect 21281 14433 21315 14467
rect 1685 14365 1719 14399
rect 2237 14365 2271 14399
rect 4914 14365 4948 14399
rect 6101 14365 6135 14399
rect 7757 14365 7791 14399
rect 9873 14365 9907 14399
rect 11529 14365 11563 14399
rect 13553 14365 13587 14399
rect 15761 14365 15795 14399
rect 17785 14365 17819 14399
rect 19257 14365 19291 14399
rect 20545 14365 20579 14399
rect 7490 14297 7524 14331
rect 9229 14297 9263 14331
rect 11262 14297 11296 14331
rect 14473 14297 14507 14331
rect 15117 14297 15151 14331
rect 16028 14297 16062 14331
rect 19901 14297 19935 14331
rect 1501 14229 1535 14263
rect 2697 14229 2731 14263
rect 3065 14229 3099 14263
rect 3157 14229 3191 14263
rect 3801 14229 3835 14263
rect 8033 14229 8067 14263
rect 14565 14229 14599 14263
rect 17141 14229 17175 14263
rect 17693 14229 17727 14263
rect 2329 14025 2363 14059
rect 3249 14025 3283 14059
rect 3985 14025 4019 14059
rect 6009 14025 6043 14059
rect 6929 14025 6963 14059
rect 7389 14025 7423 14059
rect 7941 14025 7975 14059
rect 8401 14025 8435 14059
rect 8953 14025 8987 14059
rect 10609 14025 10643 14059
rect 11529 14025 11563 14059
rect 12541 14025 12575 14059
rect 14381 14025 14415 14059
rect 16313 14025 16347 14059
rect 17417 14025 17451 14059
rect 19993 14025 20027 14059
rect 20729 14025 20763 14059
rect 21373 14025 21407 14059
rect 7297 13957 7331 13991
rect 11069 13957 11103 13991
rect 16957 13957 16991 13991
rect 17049 13957 17083 13991
rect 18828 13957 18862 13991
rect 1409 13889 1443 13923
rect 2605 13889 2639 13923
rect 3065 13889 3099 13923
rect 3893 13889 3927 13923
rect 4629 13889 4663 13923
rect 4885 13889 4919 13923
rect 6377 13889 6411 13923
rect 8309 13889 8343 13923
rect 10066 13889 10100 13923
rect 10333 13889 10367 13923
rect 11897 13889 11931 13923
rect 12725 13889 12759 13923
rect 13268 13889 13302 13923
rect 14933 13889 14967 13923
rect 15200 13889 15234 13923
rect 19349 13889 19383 13923
rect 20269 13889 20303 13923
rect 4169 13821 4203 13855
rect 7573 13821 7607 13855
rect 8585 13821 8619 13855
rect 11989 13821 12023 13855
rect 12081 13821 12115 13855
rect 13001 13821 13035 13855
rect 16865 13821 16899 13855
rect 19073 13821 19107 13855
rect 1593 13753 1627 13787
rect 2789 13753 2823 13787
rect 3525 13753 3559 13787
rect 17693 13685 17727 13719
rect 2513 13481 2547 13515
rect 7941 13481 7975 13515
rect 10149 13481 10183 13515
rect 10885 13481 10919 13515
rect 13737 13481 13771 13515
rect 16405 13481 16439 13515
rect 18153 13481 18187 13515
rect 21373 13481 21407 13515
rect 2789 13413 2823 13447
rect 4353 13413 4387 13447
rect 16129 13413 16163 13447
rect 20269 13413 20303 13447
rect 5733 13345 5767 13379
rect 6561 13345 6595 13379
rect 12449 13345 12483 13379
rect 13185 13345 13219 13379
rect 17601 13345 17635 13379
rect 1593 13277 1627 13311
rect 1869 13277 1903 13311
rect 2329 13277 2363 13311
rect 3433 13277 3467 13311
rect 3893 13277 3927 13311
rect 6377 13277 6411 13311
rect 7665 13277 7699 13311
rect 8585 13277 8619 13311
rect 9505 13277 9539 13311
rect 14749 13277 14783 13311
rect 17049 13277 17083 13311
rect 19257 13277 19291 13311
rect 5466 13209 5500 13243
rect 6469 13209 6503 13243
rect 9045 13209 9079 13243
rect 12173 13209 12207 13243
rect 13369 13209 13403 13243
rect 14105 13209 14139 13243
rect 15016 13209 15050 13243
rect 1409 13141 1443 13175
rect 2053 13141 2087 13175
rect 4077 13141 4111 13175
rect 6009 13141 6043 13175
rect 7021 13141 7055 13175
rect 13277 13141 13311 13175
rect 17693 13141 17727 13175
rect 17785 13141 17819 13175
rect 18613 13141 18647 13175
rect 19901 13141 19935 13175
rect 4261 12937 4295 12971
rect 4721 12937 4755 12971
rect 5641 12937 5675 12971
rect 8677 12937 8711 12971
rect 10333 12937 10367 12971
rect 10701 12937 10735 12971
rect 12909 12937 12943 12971
rect 14197 12937 14231 12971
rect 15577 12937 15611 12971
rect 18705 12937 18739 12971
rect 19993 12937 20027 12971
rect 1685 12869 1719 12903
rect 2605 12869 2639 12903
rect 4629 12869 4663 12903
rect 9198 12869 9232 12903
rect 11796 12869 11830 12903
rect 14565 12869 14599 12903
rect 1961 12801 1995 12835
rect 2881 12801 2915 12835
rect 3985 12801 4019 12835
rect 7021 12801 7055 12835
rect 7297 12801 7331 12835
rect 7564 12801 7598 12835
rect 13185 12801 13219 12835
rect 15209 12801 15243 12835
rect 15853 12801 15887 12835
rect 17325 12801 17359 12835
rect 17592 12801 17626 12835
rect 21106 12801 21140 12835
rect 21373 12801 21407 12835
rect 4813 12733 4847 12767
rect 5733 12733 5767 12767
rect 5917 12733 5951 12767
rect 8953 12733 8987 12767
rect 10977 12733 11011 12767
rect 11529 12733 11563 12767
rect 15025 12733 15059 12767
rect 15117 12733 15151 12767
rect 3065 12665 3099 12699
rect 2145 12597 2179 12631
rect 3341 12597 3375 12631
rect 5273 12597 5307 12631
rect 6377 12597 6411 12631
rect 13829 12597 13863 12631
rect 16681 12597 16715 12631
rect 19073 12597 19107 12631
rect 1409 12393 1443 12427
rect 2973 12393 3007 12427
rect 5825 12393 5859 12427
rect 14381 12393 14415 12427
rect 16681 12393 16715 12427
rect 17509 12393 17543 12427
rect 19257 12393 19291 12427
rect 2513 12325 2547 12359
rect 8309 12257 8343 12291
rect 15761 12257 15795 12291
rect 18153 12257 18187 12291
rect 19717 12257 19751 12291
rect 19809 12257 19843 12291
rect 1593 12189 1627 12223
rect 2053 12189 2087 12223
rect 2329 12189 2363 12223
rect 2789 12189 2823 12223
rect 3985 12189 4019 12223
rect 4445 12189 4479 12223
rect 7214 12189 7248 12223
rect 7481 12189 7515 12223
rect 11161 12189 11195 12223
rect 12909 12189 12943 12223
rect 16037 12189 16071 12223
rect 17049 12189 17083 12223
rect 19625 12189 19659 12223
rect 4690 12121 4724 12155
rect 10894 12121 10928 12155
rect 12664 12121 12698 12155
rect 15494 12121 15528 12155
rect 17969 12121 18003 12155
rect 18521 12121 18555 12155
rect 1869 12053 1903 12087
rect 3433 12053 3467 12087
rect 3801 12053 3835 12087
rect 6101 12053 6135 12087
rect 7757 12053 7791 12087
rect 8125 12053 8159 12087
rect 8217 12053 8251 12087
rect 9045 12053 9079 12087
rect 9781 12053 9815 12087
rect 11529 12053 11563 12087
rect 13185 12053 13219 12087
rect 13645 12053 13679 12087
rect 17877 12053 17911 12087
rect 1409 11849 1443 11883
rect 3433 11849 3467 11883
rect 8769 11849 8803 11883
rect 9781 11849 9815 11883
rect 10149 11849 10183 11883
rect 10701 11849 10735 11883
rect 11805 11849 11839 11883
rect 12173 11849 12207 11883
rect 15393 11849 15427 11883
rect 15853 11849 15887 11883
rect 21189 11849 21223 11883
rect 4844 11781 4878 11815
rect 5365 11781 5399 11815
rect 6745 11781 6779 11815
rect 7656 11781 7690 11815
rect 10793 11781 10827 11815
rect 18460 11781 18494 11815
rect 1593 11713 1627 11747
rect 1869 11713 1903 11747
rect 2329 11713 2363 11747
rect 2973 11713 3007 11747
rect 3249 11713 3283 11747
rect 5089 11713 5123 11747
rect 6009 11713 6043 11747
rect 6837 11713 6871 11747
rect 12265 11713 12299 11747
rect 13461 11713 13495 11747
rect 13737 11713 13771 11747
rect 14004 11713 14038 11747
rect 15761 11713 15795 11747
rect 16681 11713 16715 11747
rect 18981 11713 19015 11747
rect 20913 11713 20947 11747
rect 21373 11713 21407 11747
rect 6929 11645 6963 11679
rect 7389 11645 7423 11679
rect 9597 11645 9631 11679
rect 9689 11645 9723 11679
rect 10517 11645 10551 11679
rect 12357 11645 12391 11679
rect 15945 11645 15979 11679
rect 18705 11645 18739 11679
rect 2053 11577 2087 11611
rect 11161 11577 11195 11611
rect 17325 11577 17359 11611
rect 2513 11509 2547 11543
rect 2789 11509 2823 11543
rect 3709 11509 3743 11543
rect 6377 11509 6411 11543
rect 9045 11509 9079 11543
rect 12817 11509 12851 11543
rect 15117 11509 15151 11543
rect 19625 11509 19659 11543
rect 4353 11305 4387 11339
rect 6377 11305 6411 11339
rect 8033 11305 8067 11339
rect 8953 11305 8987 11339
rect 15117 11305 15151 11339
rect 18061 11305 18095 11339
rect 2697 11237 2731 11271
rect 3893 11237 3927 11271
rect 5365 11237 5399 11271
rect 13277 11237 13311 11271
rect 17049 11237 17083 11271
rect 1869 11169 1903 11203
rect 1961 11169 1995 11203
rect 3249 11169 3283 11203
rect 4813 11169 4847 11203
rect 4997 11169 5031 11203
rect 6009 11169 6043 11203
rect 7757 11169 7791 11203
rect 9505 11169 9539 11203
rect 14197 11169 14231 11203
rect 14381 11169 14415 11203
rect 17509 11169 17543 11203
rect 4077 11101 4111 11135
rect 4721 11101 4755 11135
rect 8217 11101 8251 11135
rect 9321 11101 9355 11135
rect 10149 11101 10183 11135
rect 11897 11101 11931 11135
rect 12164 11101 12198 11135
rect 14473 11101 14507 11135
rect 15669 11101 15703 11135
rect 3157 11033 3191 11067
rect 5733 11033 5767 11067
rect 7512 11033 7546 11067
rect 8493 11033 8527 11067
rect 9413 11033 9447 11067
rect 10394 11033 10428 11067
rect 13737 11033 13771 11067
rect 15936 11033 15970 11067
rect 17693 11033 17727 11067
rect 18337 11033 18371 11067
rect 2053 10965 2087 10999
rect 2421 10965 2455 10999
rect 3065 10965 3099 10999
rect 5825 10965 5859 10999
rect 11529 10965 11563 10999
rect 14841 10965 14875 10999
rect 17601 10965 17635 10999
rect 1685 10761 1719 10795
rect 2697 10761 2731 10795
rect 4353 10761 4387 10795
rect 4813 10761 4847 10795
rect 5365 10761 5399 10795
rect 6377 10761 6411 10795
rect 7573 10761 7607 10795
rect 10241 10761 10275 10795
rect 11805 10761 11839 10795
rect 14841 10761 14875 10795
rect 14933 10761 14967 10795
rect 15853 10761 15887 10795
rect 16313 10761 16347 10795
rect 3832 10693 3866 10727
rect 7849 10693 7883 10727
rect 12633 10693 12667 10727
rect 13154 10693 13188 10727
rect 2053 10625 2087 10659
rect 2145 10625 2179 10659
rect 4077 10625 4111 10659
rect 4721 10625 4755 10659
rect 6009 10625 6043 10659
rect 7205 10625 7239 10659
rect 11161 10625 11195 10659
rect 11897 10625 11931 10659
rect 15945 10625 15979 10659
rect 17805 10625 17839 10659
rect 18061 10625 18095 10659
rect 2329 10557 2363 10591
rect 4997 10557 5031 10591
rect 7021 10557 7055 10591
rect 7113 10557 7147 10591
rect 11713 10557 11747 10591
rect 12909 10557 12943 10591
rect 14749 10557 14783 10591
rect 15761 10557 15795 10591
rect 16681 10489 16715 10523
rect 9321 10421 9355 10455
rect 10517 10421 10551 10455
rect 12265 10421 12299 10455
rect 14289 10421 14323 10455
rect 15301 10421 15335 10455
rect 1869 10217 1903 10251
rect 3801 10217 3835 10251
rect 4813 10217 4847 10251
rect 5733 10217 5767 10251
rect 7481 10217 7515 10251
rect 9965 10217 9999 10251
rect 10885 10217 10919 10251
rect 13185 10217 13219 10251
rect 15393 10217 15427 10251
rect 16957 10217 16991 10251
rect 18337 10217 18371 10251
rect 1409 10149 1443 10183
rect 8953 10149 8987 10183
rect 3249 10081 3283 10115
rect 4445 10081 4479 10115
rect 9505 10081 9539 10115
rect 12633 10081 12667 10115
rect 12725 10081 12759 10115
rect 1593 10013 1627 10047
rect 4997 10013 5031 10047
rect 7021 10013 7055 10047
rect 8125 10013 8159 10047
rect 12173 10013 12207 10047
rect 12817 10013 12851 10047
rect 14749 10013 14783 10047
rect 17693 10013 17727 10047
rect 2982 9945 3016 9979
rect 4169 9945 4203 9979
rect 15669 9945 15703 9979
rect 4261 9877 4295 9911
rect 8401 9877 8435 9911
rect 9321 9877 9355 9911
rect 9413 9877 9447 9911
rect 2973 9673 3007 9707
rect 4169 9673 4203 9707
rect 12909 9673 12943 9707
rect 15301 9673 15335 9707
rect 10609 9605 10643 9639
rect 11796 9605 11830 9639
rect 13829 9605 13863 9639
rect 14289 9605 14323 9639
rect 1501 9537 1535 9571
rect 1961 9537 1995 9571
rect 3341 9537 3375 9571
rect 3985 9537 4019 9571
rect 4445 9537 4479 9571
rect 5273 9537 5307 9571
rect 5365 9537 5399 9571
rect 6653 9537 6687 9571
rect 7113 9537 7147 9571
rect 7380 9537 7414 9571
rect 8953 9537 8987 9571
rect 9220 9537 9254 9571
rect 11529 9537 11563 9571
rect 13185 9537 13219 9571
rect 14933 9537 14967 9571
rect 3433 9469 3467 9503
rect 3617 9469 3651 9503
rect 5457 9469 5491 9503
rect 1685 9401 1719 9435
rect 4629 9401 4663 9435
rect 5917 9401 5951 9435
rect 15577 9401 15611 9435
rect 2605 9333 2639 9367
rect 4905 9333 4939 9367
rect 6837 9333 6871 9367
rect 8493 9333 8527 9367
rect 10333 9333 10367 9367
rect 10977 9333 11011 9367
rect 8033 9129 8067 9163
rect 9689 9129 9723 9163
rect 10609 9129 10643 9163
rect 10977 9129 11011 9163
rect 3433 9061 3467 9095
rect 6285 9061 6319 9095
rect 4445 8993 4479 9027
rect 5457 8993 5491 9027
rect 6745 8993 6779 9027
rect 6837 8993 6871 9027
rect 7481 8993 7515 9027
rect 9137 8993 9171 9027
rect 9229 8993 9263 9027
rect 1409 8925 1443 8959
rect 2053 8925 2087 8959
rect 4629 8925 4663 8959
rect 5641 8925 5675 8959
rect 9965 8925 9999 8959
rect 2320 8857 2354 8891
rect 3801 8857 3835 8891
rect 6653 8857 6687 8891
rect 1593 8789 1627 8823
rect 4537 8789 4571 8823
rect 4997 8789 5031 8823
rect 5549 8789 5583 8823
rect 6009 8789 6043 8823
rect 7573 8789 7607 8823
rect 7665 8789 7699 8823
rect 8309 8789 8343 8823
rect 9321 8789 9355 8823
rect 11253 8789 11287 8823
rect 1409 8585 1443 8619
rect 2053 8585 2087 8619
rect 4905 8585 4939 8619
rect 5641 8585 5675 8619
rect 7021 8585 7055 8619
rect 7389 8585 7423 8619
rect 9689 8585 9723 8619
rect 1593 8449 1627 8483
rect 1869 8449 1903 8483
rect 2329 8449 2363 8483
rect 2973 8449 3007 8483
rect 3249 8449 3283 8483
rect 3516 8449 3550 8483
rect 6561 8449 6595 8483
rect 7481 8449 7515 8483
rect 9157 8449 9191 8483
rect 10333 8449 10367 8483
rect 5733 8381 5767 8415
rect 5917 8381 5951 8415
rect 7665 8381 7699 8415
rect 9413 8381 9447 8415
rect 2513 8313 2547 8347
rect 2789 8313 2823 8347
rect 5273 8313 5307 8347
rect 6377 8313 6411 8347
rect 8033 8313 8067 8347
rect 4629 8245 4663 8279
rect 1501 8041 1535 8075
rect 2237 8041 2271 8075
rect 8585 8041 8619 8075
rect 10609 8041 10643 8075
rect 18889 8041 18923 8075
rect 1961 7973 1995 8007
rect 3801 7973 3835 8007
rect 3341 7905 3375 7939
rect 4721 7905 4755 7939
rect 4813 7905 4847 7939
rect 5273 7905 5307 7939
rect 9505 7905 9539 7939
rect 1777 7837 1811 7871
rect 2421 7837 2455 7871
rect 3065 7837 3099 7871
rect 3985 7837 4019 7871
rect 4629 7837 4663 7871
rect 7205 7837 7239 7871
rect 9965 7837 9999 7871
rect 18705 7837 18739 7871
rect 19257 7837 19291 7871
rect 5540 7769 5574 7803
rect 7472 7769 7506 7803
rect 9321 7769 9355 7803
rect 2697 7701 2731 7735
rect 3157 7701 3191 7735
rect 4261 7701 4295 7735
rect 6653 7701 6687 7735
rect 8953 7701 8987 7735
rect 9413 7701 9447 7735
rect 2053 7497 2087 7531
rect 2513 7497 2547 7531
rect 5549 7497 5583 7531
rect 5917 7497 5951 7531
rect 9137 7497 9171 7531
rect 9597 7497 9631 7531
rect 10241 7497 10275 7531
rect 19441 7497 19475 7531
rect 3433 7429 3467 7463
rect 6644 7429 6678 7463
rect 1409 7361 1443 7395
rect 2237 7361 2271 7395
rect 2697 7361 2731 7395
rect 4169 7361 4203 7395
rect 4436 7361 4470 7395
rect 6377 7361 6411 7395
rect 8493 7361 8527 7395
rect 9505 7361 9539 7395
rect 19257 7361 19291 7395
rect 19717 7361 19751 7395
rect 3893 7293 3927 7327
rect 8585 7293 8619 7327
rect 8677 7293 8711 7327
rect 9689 7293 9723 7327
rect 1593 7225 1627 7259
rect 7757 7157 7791 7191
rect 8125 7157 8159 7191
rect 4169 6953 4203 6987
rect 6193 6953 6227 6987
rect 3249 6885 3283 6919
rect 8953 6885 8987 6919
rect 3801 6817 3835 6851
rect 4813 6817 4847 6851
rect 8217 6817 8251 6851
rect 1409 6749 1443 6783
rect 1869 6749 1903 6783
rect 2329 6749 2363 6783
rect 2789 6749 2823 6783
rect 3433 6749 3467 6783
rect 4537 6749 4571 6783
rect 5549 6749 5583 6783
rect 8033 6749 8067 6783
rect 19625 6749 19659 6783
rect 5181 6681 5215 6715
rect 1593 6613 1627 6647
rect 2053 6613 2087 6647
rect 2513 6613 2547 6647
rect 2973 6613 3007 6647
rect 4629 6613 4663 6647
rect 6745 6613 6779 6647
rect 7113 6613 7147 6647
rect 7665 6613 7699 6647
rect 8125 6613 8159 6647
rect 19809 6613 19843 6647
rect 1593 6409 1627 6443
rect 2513 6409 2547 6443
rect 2973 6409 3007 6443
rect 3801 6409 3835 6443
rect 6377 6409 6411 6443
rect 8309 6409 8343 6443
rect 20269 6409 20303 6443
rect 5733 6341 5767 6375
rect 1409 6273 1443 6307
rect 1869 6273 1903 6307
rect 2329 6273 2363 6307
rect 2789 6273 2823 6307
rect 3249 6273 3283 6307
rect 20085 6273 20119 6307
rect 6745 6205 6779 6239
rect 2053 6137 2087 6171
rect 3433 6137 3467 6171
rect 7941 6137 7975 6171
rect 4169 6069 4203 6103
rect 4721 6069 4755 6103
rect 5089 6069 5123 6103
rect 1593 5865 1627 5899
rect 4629 5865 4663 5899
rect 4997 5865 5031 5899
rect 5365 5865 5399 5899
rect 20729 5865 20763 5899
rect 2513 5797 2547 5831
rect 2973 5797 3007 5831
rect 3341 5797 3375 5831
rect 6377 5797 6411 5831
rect 21005 5797 21039 5831
rect 5641 5729 5675 5763
rect 1409 5661 1443 5695
rect 1869 5661 1903 5695
rect 2329 5661 2363 5695
rect 2789 5661 2823 5695
rect 6009 5661 6043 5695
rect 20545 5661 20579 5695
rect 21189 5661 21223 5695
rect 2053 5525 2087 5559
rect 3801 5525 3835 5559
rect 4261 5525 4295 5559
rect 20177 5525 20211 5559
rect 2053 5321 2087 5355
rect 2513 5321 2547 5355
rect 2881 5321 2915 5355
rect 4629 5321 4663 5355
rect 5365 5321 5399 5355
rect 5825 5321 5859 5355
rect 3157 5253 3191 5287
rect 4997 5253 5031 5287
rect 1409 5185 1443 5219
rect 1869 5185 1903 5219
rect 2329 5185 2363 5219
rect 4353 5185 4387 5219
rect 20821 5117 20855 5151
rect 1593 4981 1627 5015
rect 3525 4981 3559 5015
rect 3985 4981 4019 5015
rect 2053 4777 2087 4811
rect 3893 4777 3927 4811
rect 4169 4777 4203 4811
rect 2329 4709 2363 4743
rect 4537 4709 4571 4743
rect 3157 4641 3191 4675
rect 1409 4573 1443 4607
rect 1869 4573 1903 4607
rect 4905 4573 4939 4607
rect 1593 4437 1627 4471
rect 2789 4437 2823 4471
rect 3617 4233 3651 4267
rect 3985 4233 4019 4267
rect 1961 4097 1995 4131
rect 4721 4097 4755 4131
rect 2237 4029 2271 4063
rect 4353 4029 4387 4063
rect 2881 3961 2915 3995
rect 3249 3961 3283 3995
rect 2513 3893 2547 3927
rect 4169 3689 4203 3723
rect 3065 3621 3099 3655
rect 1961 3553 1995 3587
rect 2789 3553 2823 3587
rect 2237 3485 2271 3519
rect 4537 3485 4571 3519
rect 2605 3417 2639 3451
rect 3801 3349 3835 3383
rect 2605 3145 2639 3179
rect 1961 3009 1995 3043
rect 2697 3009 2731 3043
rect 3801 3009 3835 3043
rect 2237 2941 2271 2975
rect 4169 2941 4203 2975
rect 4537 2873 4571 2907
rect 3065 2805 3099 2839
rect 3433 2805 3467 2839
rect 2697 2601 2731 2635
rect 3157 2601 3191 2635
rect 4077 2601 4111 2635
rect 1961 2465 1995 2499
rect 2237 2397 2271 2431
rect 2605 2397 2639 2431
rect 4905 2397 4939 2431
rect 11897 2397 11931 2431
rect 12173 2397 12207 2431
rect 3249 2329 3283 2363
rect 4169 2329 4203 2363
rect 4537 2329 4571 2363
rect 11713 2261 11747 2295
<< metal1 >>
rect 2774 21292 2780 21344
rect 2832 21332 2838 21344
rect 9122 21332 9128 21344
rect 2832 21304 9128 21332
rect 2832 21292 2838 21304
rect 9122 21292 9128 21304
rect 9180 21292 9186 21344
rect 5626 20884 5632 20936
rect 5684 20924 5690 20936
rect 6178 20924 6184 20936
rect 5684 20896 6184 20924
rect 5684 20884 5690 20896
rect 6178 20884 6184 20896
rect 6236 20884 6242 20936
rect 3970 20816 3976 20868
rect 4028 20856 4034 20868
rect 6822 20856 6828 20868
rect 4028 20828 6828 20856
rect 4028 20816 4034 20828
rect 6822 20816 6828 20828
rect 6880 20816 6886 20868
rect 11238 20816 11244 20868
rect 11296 20856 11302 20868
rect 16114 20856 16120 20868
rect 11296 20828 16120 20856
rect 11296 20816 11302 20828
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 8386 20748 8392 20800
rect 8444 20788 8450 20800
rect 8938 20788 8944 20800
rect 8444 20760 8944 20788
rect 8444 20748 8450 20760
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 11698 20748 11704 20800
rect 11756 20788 11762 20800
rect 12802 20788 12808 20800
rect 11756 20760 12808 20788
rect 11756 20748 11762 20760
rect 12802 20748 12808 20760
rect 12860 20748 12866 20800
rect 1104 20698 21896 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21896 20698
rect 1104 20624 21896 20646
rect 3418 20544 3424 20596
rect 3476 20584 3482 20596
rect 3970 20584 3976 20596
rect 3476 20556 3976 20584
rect 3476 20544 3482 20556
rect 3970 20544 3976 20556
rect 4028 20544 4034 20596
rect 5629 20587 5687 20593
rect 5629 20553 5641 20587
rect 5675 20584 5687 20587
rect 8478 20584 8484 20596
rect 5675 20556 8484 20584
rect 5675 20553 5687 20556
rect 5629 20547 5687 20553
rect 8478 20544 8484 20556
rect 8536 20544 8542 20596
rect 9122 20584 9128 20596
rect 9083 20556 9128 20584
rect 9122 20544 9128 20556
rect 9180 20544 9186 20596
rect 12986 20584 12992 20596
rect 10980 20556 12992 20584
rect 2038 20476 2044 20528
rect 2096 20476 2102 20528
rect 7929 20519 7987 20525
rect 2746 20488 6868 20516
rect 842 20408 848 20460
rect 900 20448 906 20460
rect 2056 20448 2084 20476
rect 2317 20451 2375 20457
rect 2317 20448 2329 20451
rect 900 20420 2329 20448
rect 900 20408 906 20420
rect 2317 20417 2329 20420
rect 2363 20417 2375 20451
rect 2317 20411 2375 20417
rect 2041 20383 2099 20389
rect 2041 20349 2053 20383
rect 2087 20349 2099 20383
rect 2041 20343 2099 20349
rect 2056 20312 2084 20343
rect 2746 20312 2774 20488
rect 2958 20408 2964 20460
rect 3016 20448 3022 20460
rect 4985 20451 5043 20457
rect 3016 20420 3372 20448
rect 3016 20408 3022 20420
rect 3344 20392 3372 20420
rect 4985 20417 4997 20451
rect 5031 20448 5043 20451
rect 6730 20448 6736 20460
rect 5031 20420 5856 20448
rect 5031 20417 5043 20420
rect 4985 20411 5043 20417
rect 5828 20392 5856 20420
rect 5920 20420 6736 20448
rect 3145 20383 3203 20389
rect 3145 20349 3157 20383
rect 3191 20349 3203 20383
rect 3145 20343 3203 20349
rect 2056 20284 2774 20312
rect 3160 20312 3188 20343
rect 3326 20340 3332 20392
rect 3384 20380 3390 20392
rect 3421 20383 3479 20389
rect 3421 20380 3433 20383
rect 3384 20352 3433 20380
rect 3384 20340 3390 20352
rect 3421 20349 3433 20352
rect 3467 20349 3479 20383
rect 3421 20343 3479 20349
rect 3789 20383 3847 20389
rect 3789 20349 3801 20383
rect 3835 20380 3847 20383
rect 3970 20380 3976 20392
rect 3835 20352 3976 20380
rect 3835 20349 3847 20352
rect 3789 20343 3847 20349
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4065 20383 4123 20389
rect 4065 20349 4077 20383
rect 4111 20380 4123 20383
rect 5534 20380 5540 20392
rect 4111 20352 5540 20380
rect 4111 20349 4123 20352
rect 4065 20343 4123 20349
rect 5534 20340 5540 20352
rect 5592 20340 5598 20392
rect 5718 20380 5724 20392
rect 5679 20352 5724 20380
rect 5718 20340 5724 20352
rect 5776 20340 5782 20392
rect 5810 20340 5816 20392
rect 5868 20340 5874 20392
rect 5920 20389 5948 20420
rect 6730 20408 6736 20420
rect 6788 20408 6794 20460
rect 6840 20448 6868 20488
rect 7929 20485 7941 20519
rect 7975 20516 7987 20519
rect 9922 20519 9980 20525
rect 9922 20516 9934 20519
rect 7975 20488 9934 20516
rect 7975 20485 7987 20488
rect 7929 20479 7987 20485
rect 9922 20485 9934 20488
rect 9968 20485 9980 20519
rect 9922 20479 9980 20485
rect 8294 20448 8300 20460
rect 6840 20420 8300 20448
rect 8294 20408 8300 20420
rect 8352 20408 8358 20460
rect 8573 20451 8631 20457
rect 8573 20417 8585 20451
rect 8619 20448 8631 20451
rect 8662 20448 8668 20460
rect 8619 20420 8668 20448
rect 8619 20417 8631 20420
rect 8573 20411 8631 20417
rect 8662 20408 8668 20420
rect 8720 20408 8726 20460
rect 8938 20448 8944 20460
rect 8899 20420 8944 20448
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 9490 20408 9496 20460
rect 9548 20448 9554 20460
rect 10980 20448 11008 20556
rect 12986 20544 12992 20556
rect 13044 20544 13050 20596
rect 13078 20544 13084 20596
rect 13136 20584 13142 20596
rect 13265 20587 13323 20593
rect 13265 20584 13277 20587
rect 13136 20556 13277 20584
rect 13136 20544 13142 20556
rect 13265 20553 13277 20556
rect 13311 20553 13323 20587
rect 13265 20547 13323 20553
rect 13538 20544 13544 20596
rect 13596 20584 13602 20596
rect 14185 20587 14243 20593
rect 14185 20584 14197 20587
rect 13596 20556 14197 20584
rect 13596 20544 13602 20556
rect 14185 20553 14197 20556
rect 14231 20553 14243 20587
rect 14185 20547 14243 20553
rect 14458 20544 14464 20596
rect 14516 20584 14522 20596
rect 15289 20587 15347 20593
rect 15289 20584 15301 20587
rect 14516 20556 15301 20584
rect 14516 20544 14522 20556
rect 15289 20553 15301 20556
rect 15335 20553 15347 20587
rect 15289 20547 15347 20553
rect 15838 20544 15844 20596
rect 15896 20584 15902 20596
rect 16761 20587 16819 20593
rect 16761 20584 16773 20587
rect 15896 20556 16773 20584
rect 15896 20544 15902 20556
rect 16761 20553 16773 20556
rect 16807 20553 16819 20587
rect 16761 20547 16819 20553
rect 17218 20544 17224 20596
rect 17276 20584 17282 20596
rect 17865 20587 17923 20593
rect 17865 20584 17877 20587
rect 17276 20556 17877 20584
rect 17276 20544 17282 20556
rect 17865 20553 17877 20556
rect 17911 20553 17923 20587
rect 17865 20547 17923 20553
rect 18598 20544 18604 20596
rect 18656 20584 18662 20596
rect 19337 20587 19395 20593
rect 19337 20584 19349 20587
rect 18656 20556 19349 20584
rect 18656 20544 18662 20556
rect 19337 20553 19349 20556
rect 19383 20553 19395 20587
rect 19337 20547 19395 20553
rect 19426 20544 19432 20596
rect 19484 20584 19490 20596
rect 19889 20587 19947 20593
rect 19889 20584 19901 20587
rect 19484 20556 19901 20584
rect 19484 20544 19490 20556
rect 19889 20553 19901 20556
rect 19935 20553 19947 20587
rect 19889 20547 19947 20553
rect 12618 20476 12624 20528
rect 12676 20516 12682 20528
rect 15930 20516 15936 20528
rect 12676 20488 15936 20516
rect 12676 20476 12682 20488
rect 15930 20476 15936 20488
rect 15988 20476 15994 20528
rect 17586 20516 17592 20528
rect 16040 20488 17592 20516
rect 9548 20420 11008 20448
rect 9548 20408 9554 20420
rect 11054 20408 11060 20460
rect 11112 20448 11118 20460
rect 11517 20451 11575 20457
rect 11517 20448 11529 20451
rect 11112 20420 11529 20448
rect 11112 20408 11118 20420
rect 11517 20417 11529 20420
rect 11563 20417 11575 20451
rect 12710 20448 12716 20460
rect 12671 20420 12716 20448
rect 11517 20411 11575 20417
rect 12710 20408 12716 20420
rect 12768 20408 12774 20460
rect 13446 20448 13452 20460
rect 13407 20420 13452 20448
rect 13446 20408 13452 20420
rect 13504 20408 13510 20460
rect 14369 20451 14427 20457
rect 14369 20417 14381 20451
rect 14415 20448 14427 20451
rect 14921 20451 14979 20457
rect 14415 20420 14872 20448
rect 14415 20417 14427 20420
rect 14369 20411 14427 20417
rect 5905 20383 5963 20389
rect 5905 20349 5917 20383
rect 5951 20349 5963 20383
rect 5905 20343 5963 20349
rect 6457 20383 6515 20389
rect 6457 20349 6469 20383
rect 6503 20380 6515 20383
rect 9398 20380 9404 20392
rect 6503 20352 9404 20380
rect 6503 20349 6515 20352
rect 6457 20343 6515 20349
rect 9398 20340 9404 20352
rect 9456 20340 9462 20392
rect 9582 20340 9588 20392
rect 9640 20380 9646 20392
rect 9677 20383 9735 20389
rect 9677 20380 9689 20383
rect 9640 20352 9689 20380
rect 9640 20340 9646 20352
rect 9677 20349 9689 20352
rect 9723 20349 9735 20383
rect 9677 20343 9735 20349
rect 13630 20312 13636 20324
rect 3160 20284 9674 20312
rect 5258 20244 5264 20256
rect 5219 20216 5264 20244
rect 5258 20204 5264 20216
rect 5316 20204 5322 20256
rect 6638 20204 6644 20256
rect 6696 20244 6702 20256
rect 7377 20247 7435 20253
rect 7377 20244 7389 20247
rect 6696 20216 7389 20244
rect 6696 20204 6702 20216
rect 7377 20213 7389 20216
rect 7423 20213 7435 20247
rect 9646 20244 9674 20284
rect 10888 20284 13636 20312
rect 10888 20244 10916 20284
rect 13630 20272 13636 20284
rect 13688 20272 13694 20324
rect 13998 20272 14004 20324
rect 14056 20312 14062 20324
rect 14737 20315 14795 20321
rect 14737 20312 14749 20315
rect 14056 20284 14749 20312
rect 14056 20272 14062 20284
rect 14737 20281 14749 20284
rect 14783 20281 14795 20315
rect 14737 20275 14795 20281
rect 11054 20244 11060 20256
rect 9646 20216 10916 20244
rect 11015 20216 11060 20244
rect 7377 20207 7435 20213
rect 11054 20204 11060 20216
rect 11112 20204 11118 20256
rect 12158 20244 12164 20256
rect 12119 20216 12164 20244
rect 12158 20204 12164 20216
rect 12216 20204 12222 20256
rect 12250 20204 12256 20256
rect 12308 20244 12314 20256
rect 12529 20247 12587 20253
rect 12529 20244 12541 20247
rect 12308 20216 12541 20244
rect 12308 20204 12314 20216
rect 12529 20213 12541 20216
rect 12575 20213 12587 20247
rect 14844 20244 14872 20420
rect 14921 20417 14933 20451
rect 14967 20417 14979 20451
rect 15470 20448 15476 20460
rect 15431 20420 15476 20448
rect 14921 20411 14979 20417
rect 14936 20380 14964 20411
rect 15470 20408 15476 20420
rect 15528 20408 15534 20460
rect 16040 20457 16068 20488
rect 17586 20476 17592 20488
rect 17644 20476 17650 20528
rect 21082 20516 21088 20528
rect 17880 20488 19472 20516
rect 16025 20451 16083 20457
rect 16025 20417 16037 20451
rect 16071 20417 16083 20451
rect 16025 20411 16083 20417
rect 16945 20451 17003 20457
rect 16945 20417 16957 20451
rect 16991 20448 17003 20451
rect 17497 20451 17555 20457
rect 16991 20420 17448 20448
rect 16991 20417 17003 20420
rect 16945 20411 17003 20417
rect 17218 20380 17224 20392
rect 14936 20352 17224 20380
rect 17218 20340 17224 20352
rect 17276 20340 17282 20392
rect 17420 20380 17448 20420
rect 17497 20417 17509 20451
rect 17543 20448 17555 20451
rect 17880 20448 17908 20488
rect 18046 20448 18052 20460
rect 17543 20420 17908 20448
rect 18007 20420 18052 20448
rect 17543 20417 17555 20420
rect 17497 20411 17555 20417
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 18598 20448 18604 20460
rect 18559 20420 18604 20448
rect 18598 20408 18604 20420
rect 18656 20408 18662 20460
rect 17954 20380 17960 20392
rect 17420 20352 17960 20380
rect 17954 20340 17960 20352
rect 18012 20340 18018 20392
rect 19444 20380 19472 20488
rect 19536 20488 21088 20516
rect 19536 20457 19564 20488
rect 21082 20476 21088 20488
rect 21140 20476 21146 20528
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20417 19579 20451
rect 19521 20411 19579 20417
rect 20073 20451 20131 20457
rect 20073 20417 20085 20451
rect 20119 20448 20131 20451
rect 20806 20448 20812 20460
rect 20119 20420 20812 20448
rect 20119 20417 20131 20420
rect 20073 20411 20131 20417
rect 20806 20408 20812 20420
rect 20864 20408 20870 20460
rect 20530 20380 20536 20392
rect 19444 20352 20536 20380
rect 20530 20340 20536 20352
rect 20588 20340 20594 20392
rect 20990 20340 20996 20392
rect 21048 20380 21054 20392
rect 21085 20383 21143 20389
rect 21085 20380 21097 20383
rect 21048 20352 21097 20380
rect 21048 20340 21054 20352
rect 21085 20349 21097 20352
rect 21131 20349 21143 20383
rect 21085 20343 21143 20349
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20380 21419 20383
rect 21450 20380 21456 20392
rect 21407 20352 21456 20380
rect 21407 20349 21419 20352
rect 21361 20343 21419 20349
rect 21450 20340 21456 20352
rect 21508 20380 21514 20392
rect 22738 20380 22744 20392
rect 21508 20352 22744 20380
rect 21508 20340 21514 20352
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 14918 20272 14924 20324
rect 14976 20312 14982 20324
rect 15841 20315 15899 20321
rect 15841 20312 15853 20315
rect 14976 20284 15853 20312
rect 14976 20272 14982 20284
rect 15841 20281 15853 20284
rect 15887 20281 15899 20315
rect 15841 20275 15899 20281
rect 16298 20272 16304 20324
rect 16356 20312 16362 20324
rect 17313 20315 17371 20321
rect 17313 20312 17325 20315
rect 16356 20284 17325 20312
rect 16356 20272 16362 20284
rect 17313 20281 17325 20284
rect 17359 20281 17371 20315
rect 17313 20275 17371 20281
rect 17678 20272 17684 20324
rect 17736 20312 17742 20324
rect 18417 20315 18475 20321
rect 18417 20312 18429 20315
rect 17736 20284 18429 20312
rect 17736 20272 17742 20284
rect 18417 20281 18429 20284
rect 18463 20281 18475 20315
rect 18417 20275 18475 20281
rect 18506 20244 18512 20256
rect 14844 20216 18512 20244
rect 12529 20207 12587 20213
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 8570 20040 8576 20052
rect 2884 20012 8576 20040
rect 2884 19913 2912 20012
rect 8570 20000 8576 20012
rect 8628 20000 8634 20052
rect 9674 20000 9680 20052
rect 9732 20040 9738 20052
rect 10045 20043 10103 20049
rect 10045 20040 10057 20043
rect 9732 20012 10057 20040
rect 9732 20000 9738 20012
rect 10045 20009 10057 20012
rect 10091 20040 10103 20043
rect 10091 20012 11744 20040
rect 10091 20009 10103 20012
rect 10045 20003 10103 20009
rect 8754 19932 8760 19984
rect 8812 19972 8818 19984
rect 8812 19944 10088 19972
rect 8812 19932 8818 19944
rect 10060 19916 10088 19944
rect 2041 19907 2099 19913
rect 2041 19873 2053 19907
rect 2087 19904 2099 19907
rect 2869 19907 2927 19913
rect 2087 19876 2774 19904
rect 2087 19873 2099 19876
rect 2041 19867 2099 19873
rect 1210 19796 1216 19848
rect 1268 19836 1274 19848
rect 1578 19836 1584 19848
rect 1268 19808 1584 19836
rect 1268 19796 1274 19808
rect 1578 19796 1584 19808
rect 1636 19836 1642 19848
rect 2317 19839 2375 19845
rect 2317 19836 2329 19839
rect 1636 19808 2329 19836
rect 1636 19796 1642 19808
rect 2317 19805 2329 19808
rect 2363 19805 2375 19839
rect 2317 19799 2375 19805
rect 2498 19796 2504 19848
rect 2556 19836 2562 19848
rect 2593 19839 2651 19845
rect 2593 19836 2605 19839
rect 2556 19808 2605 19836
rect 2556 19796 2562 19808
rect 2593 19805 2605 19808
rect 2639 19805 2651 19839
rect 2746 19836 2774 19876
rect 2869 19873 2881 19907
rect 2915 19873 2927 19907
rect 5442 19904 5448 19916
rect 2869 19867 2927 19873
rect 5092 19876 5448 19904
rect 5092 19836 5120 19876
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 8662 19864 8668 19916
rect 8720 19904 8726 19916
rect 9125 19907 9183 19913
rect 9125 19904 9137 19907
rect 8720 19876 9137 19904
rect 8720 19864 8726 19876
rect 9125 19873 9137 19876
rect 9171 19873 9183 19907
rect 9125 19867 9183 19873
rect 10042 19864 10048 19916
rect 10100 19864 10106 19916
rect 2746 19808 5120 19836
rect 2593 19799 2651 19805
rect 5166 19796 5172 19848
rect 5224 19836 5230 19848
rect 5224 19808 5269 19836
rect 5224 19796 5230 19808
rect 5534 19796 5540 19848
rect 5592 19796 5598 19848
rect 6638 19796 6644 19848
rect 6696 19845 6702 19848
rect 6696 19836 6708 19845
rect 6914 19836 6920 19848
rect 6696 19808 6741 19836
rect 6875 19808 6920 19836
rect 6696 19799 6708 19808
rect 6696 19796 6702 19799
rect 6914 19796 6920 19808
rect 6972 19796 6978 19848
rect 8573 19839 8631 19845
rect 8573 19805 8585 19839
rect 8619 19836 8631 19839
rect 9214 19836 9220 19848
rect 8619 19808 9220 19836
rect 8619 19805 8631 19808
rect 8573 19799 8631 19805
rect 9214 19796 9220 19808
rect 9272 19836 9278 19848
rect 9582 19836 9588 19848
rect 9272 19808 9588 19836
rect 9272 19796 9278 19808
rect 9582 19796 9588 19808
rect 9640 19836 9646 19848
rect 10778 19836 10784 19848
rect 9640 19808 10784 19836
rect 9640 19796 9646 19808
rect 10778 19796 10784 19808
rect 10836 19836 10842 19848
rect 11716 19845 11744 20012
rect 13446 20000 13452 20052
rect 13504 20040 13510 20052
rect 15013 20043 15071 20049
rect 15013 20040 15025 20043
rect 13504 20012 15025 20040
rect 13504 20000 13510 20012
rect 15013 20009 15025 20012
rect 15059 20009 15071 20043
rect 15013 20003 15071 20009
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15565 20043 15623 20049
rect 15565 20040 15577 20043
rect 15436 20012 15577 20040
rect 15436 20000 15442 20012
rect 15565 20009 15577 20012
rect 15611 20009 15623 20043
rect 16942 20040 16948 20052
rect 16903 20012 16948 20040
rect 15565 20003 15623 20009
rect 16942 20000 16948 20012
rect 17000 20000 17006 20052
rect 17218 20000 17224 20052
rect 17276 20040 17282 20052
rect 17405 20043 17463 20049
rect 17405 20040 17417 20043
rect 17276 20012 17417 20040
rect 17276 20000 17282 20012
rect 17405 20009 17417 20012
rect 17451 20009 17463 20043
rect 17405 20003 17463 20009
rect 18138 20000 18144 20052
rect 18196 20040 18202 20052
rect 18325 20043 18383 20049
rect 18325 20040 18337 20043
rect 18196 20012 18337 20040
rect 18196 20000 18202 20012
rect 18325 20009 18337 20012
rect 18371 20009 18383 20043
rect 18325 20003 18383 20009
rect 19518 20000 19524 20052
rect 19576 20040 19582 20052
rect 19797 20043 19855 20049
rect 19797 20040 19809 20043
rect 19576 20012 19809 20040
rect 19576 20000 19582 20012
rect 19797 20009 19809 20012
rect 19843 20009 19855 20043
rect 19797 20003 19855 20009
rect 11790 19932 11796 19984
rect 11848 19972 11854 19984
rect 13265 19975 13323 19981
rect 13265 19972 13277 19975
rect 11848 19944 13277 19972
rect 11848 19932 11854 19944
rect 13265 19941 13277 19944
rect 13311 19941 13323 19975
rect 13265 19935 13323 19941
rect 13725 19975 13783 19981
rect 13725 19941 13737 19975
rect 13771 19972 13783 19975
rect 19610 19972 19616 19984
rect 13771 19944 19616 19972
rect 13771 19941 13783 19944
rect 13725 19935 13783 19941
rect 19610 19932 19616 19944
rect 19668 19932 19674 19984
rect 13906 19864 13912 19916
rect 13964 19904 13970 19916
rect 13964 19876 17540 19904
rect 13964 19864 13970 19876
rect 11425 19839 11483 19845
rect 11425 19836 11437 19839
rect 10836 19808 11437 19836
rect 10836 19796 10842 19808
rect 11425 19805 11437 19808
rect 11471 19805 11483 19839
rect 11425 19799 11483 19805
rect 11701 19839 11759 19845
rect 11701 19805 11713 19839
rect 11747 19805 11759 19839
rect 11701 19799 11759 19805
rect 11882 19796 11888 19848
rect 11940 19836 11946 19848
rect 12621 19839 12679 19845
rect 12621 19836 12633 19839
rect 11940 19808 12633 19836
rect 11940 19796 11946 19808
rect 12621 19805 12633 19808
rect 12667 19805 12679 19839
rect 12621 19799 12679 19805
rect 13170 19796 13176 19848
rect 13228 19836 13234 19848
rect 13541 19839 13599 19845
rect 13541 19836 13553 19839
rect 13228 19808 13553 19836
rect 13228 19796 13234 19808
rect 13541 19805 13553 19808
rect 13587 19805 13599 19839
rect 13541 19799 13599 19805
rect 14093 19839 14151 19845
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14550 19836 14556 19848
rect 14511 19808 14556 19836
rect 14093 19799 14151 19805
rect 4154 19728 4160 19780
rect 4212 19768 4218 19780
rect 4902 19771 4960 19777
rect 4902 19768 4914 19771
rect 4212 19740 4914 19768
rect 4212 19728 4218 19740
rect 4902 19737 4914 19740
rect 4948 19737 4960 19771
rect 5552 19768 5580 19796
rect 8328 19771 8386 19777
rect 5552 19740 6500 19768
rect 4902 19731 4960 19737
rect 3789 19703 3847 19709
rect 3789 19669 3801 19703
rect 3835 19700 3847 19703
rect 3970 19700 3976 19712
rect 3835 19672 3976 19700
rect 3835 19669 3847 19672
rect 3789 19663 3847 19669
rect 3970 19660 3976 19672
rect 4028 19660 4034 19712
rect 5534 19700 5540 19712
rect 5495 19672 5540 19700
rect 5534 19660 5540 19672
rect 5592 19660 5598 19712
rect 6472 19700 6500 19740
rect 8328 19737 8340 19771
rect 8374 19768 8386 19771
rect 11180 19771 11238 19777
rect 8374 19740 10364 19768
rect 8374 19737 8386 19740
rect 8328 19731 8386 19737
rect 6638 19700 6644 19712
rect 6472 19672 6644 19700
rect 6638 19660 6644 19672
rect 6696 19660 6702 19712
rect 7190 19700 7196 19712
rect 7151 19672 7196 19700
rect 7190 19660 7196 19672
rect 7248 19660 7254 19712
rect 8478 19660 8484 19712
rect 8536 19700 8542 19712
rect 8846 19700 8852 19712
rect 8536 19672 8852 19700
rect 8536 19660 8542 19672
rect 8846 19660 8852 19672
rect 8904 19660 8910 19712
rect 9306 19700 9312 19712
rect 9267 19672 9312 19700
rect 9306 19660 9312 19672
rect 9364 19660 9370 19712
rect 9401 19703 9459 19709
rect 9401 19669 9413 19703
rect 9447 19700 9459 19703
rect 9582 19700 9588 19712
rect 9447 19672 9588 19700
rect 9447 19669 9459 19672
rect 9401 19663 9459 19669
rect 9582 19660 9588 19672
rect 9640 19660 9646 19712
rect 9766 19700 9772 19712
rect 9727 19672 9772 19700
rect 9766 19660 9772 19672
rect 9824 19660 9830 19712
rect 10336 19700 10364 19740
rect 11180 19737 11192 19771
rect 11226 19768 11238 19771
rect 12158 19768 12164 19780
rect 11226 19740 12164 19768
rect 11226 19737 11238 19740
rect 11180 19731 11238 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 12345 19771 12403 19777
rect 12345 19768 12357 19771
rect 12268 19740 12357 19768
rect 12268 19700 12296 19740
rect 12345 19737 12357 19740
rect 12391 19737 12403 19771
rect 12345 19731 12403 19737
rect 13446 19728 13452 19780
rect 13504 19768 13510 19780
rect 14108 19768 14136 19799
rect 14550 19796 14556 19808
rect 14608 19796 14614 19848
rect 15197 19839 15255 19845
rect 15197 19836 15209 19839
rect 14752 19808 15209 19836
rect 13504 19740 14136 19768
rect 13504 19728 13510 19740
rect 14274 19700 14280 19712
rect 10336 19672 12296 19700
rect 14235 19672 14280 19700
rect 14274 19660 14280 19672
rect 14332 19660 14338 19712
rect 14752 19709 14780 19808
rect 15197 19805 15209 19808
rect 15243 19805 15255 19839
rect 15197 19799 15255 19805
rect 15749 19839 15807 19845
rect 15749 19805 15761 19839
rect 15795 19805 15807 19839
rect 15749 19799 15807 19805
rect 15764 19768 15792 19799
rect 15930 19796 15936 19848
rect 15988 19836 15994 19848
rect 16209 19839 16267 19845
rect 16209 19836 16221 19839
rect 15988 19808 16221 19836
rect 15988 19796 15994 19808
rect 16209 19805 16221 19808
rect 16255 19836 16267 19839
rect 16390 19836 16396 19848
rect 16255 19808 16396 19836
rect 16255 19805 16267 19808
rect 16209 19799 16267 19805
rect 16390 19796 16396 19808
rect 16448 19796 16454 19848
rect 16482 19796 16488 19848
rect 16540 19836 16546 19848
rect 17126 19836 17132 19848
rect 16540 19808 16585 19836
rect 17087 19808 17132 19836
rect 16540 19796 16546 19808
rect 17126 19796 17132 19808
rect 17184 19796 17190 19848
rect 17512 19832 17540 19876
rect 17862 19864 17868 19916
rect 17920 19904 17926 19916
rect 19702 19904 19708 19916
rect 17920 19876 19708 19904
rect 17920 19864 17926 19876
rect 19702 19864 19708 19876
rect 19760 19864 19766 19916
rect 20714 19904 20720 19916
rect 20675 19876 20720 19904
rect 20714 19864 20720 19876
rect 20772 19864 20778 19916
rect 17589 19839 17647 19845
rect 17589 19832 17601 19839
rect 17512 19805 17601 19832
rect 17635 19805 17647 19839
rect 17512 19804 17647 19805
rect 17589 19799 17647 19804
rect 18509 19839 18567 19845
rect 18509 19805 18521 19839
rect 18555 19836 18567 19839
rect 19058 19836 19064 19848
rect 18555 19808 19064 19836
rect 18555 19805 18567 19808
rect 18509 19799 18567 19805
rect 19058 19796 19064 19808
rect 19116 19796 19122 19848
rect 19334 19836 19340 19848
rect 19295 19808 19340 19836
rect 19334 19796 19340 19808
rect 19392 19796 19398 19848
rect 19613 19839 19671 19845
rect 19613 19805 19625 19839
rect 19659 19836 19671 19839
rect 20162 19836 20168 19848
rect 19659 19808 20168 19836
rect 19659 19805 19671 19808
rect 19613 19799 19671 19805
rect 20162 19796 20168 19808
rect 20220 19796 20226 19848
rect 21358 19836 21364 19848
rect 21271 19808 21364 19836
rect 21358 19796 21364 19808
rect 21416 19836 21422 19848
rect 22278 19836 22284 19848
rect 21416 19808 22284 19836
rect 21416 19796 21422 19808
rect 22278 19796 22284 19808
rect 22336 19796 22342 19848
rect 19426 19768 19432 19780
rect 15764 19740 19432 19768
rect 19426 19728 19432 19740
rect 19484 19728 19490 19780
rect 14737 19703 14795 19709
rect 14737 19669 14749 19703
rect 14783 19669 14795 19703
rect 16022 19700 16028 19712
rect 15983 19672 16028 19700
rect 14737 19663 14795 19669
rect 16022 19660 16028 19672
rect 16080 19660 16086 19712
rect 17126 19660 17132 19712
rect 17184 19700 17190 19712
rect 17862 19700 17868 19712
rect 17184 19672 17868 19700
rect 17184 19660 17190 19672
rect 17862 19660 17868 19672
rect 17920 19660 17926 19712
rect 17957 19703 18015 19709
rect 17957 19669 17969 19703
rect 18003 19700 18015 19703
rect 18138 19700 18144 19712
rect 18003 19672 18144 19700
rect 18003 19669 18015 19672
rect 17957 19663 18015 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 18782 19700 18788 19712
rect 18743 19672 18788 19700
rect 18782 19660 18788 19672
rect 18840 19660 18846 19712
rect 1104 19610 21896 19632
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21896 19610
rect 1104 19536 21896 19558
rect 2593 19499 2651 19505
rect 2593 19465 2605 19499
rect 2639 19496 2651 19499
rect 2866 19496 2872 19508
rect 2639 19468 2872 19496
rect 2639 19465 2651 19468
rect 2593 19459 2651 19465
rect 2866 19456 2872 19468
rect 2924 19456 2930 19508
rect 4062 19456 4068 19508
rect 4120 19496 4126 19508
rect 5077 19499 5135 19505
rect 5077 19496 5089 19499
rect 4120 19468 5089 19496
rect 4120 19456 4126 19468
rect 5077 19465 5089 19468
rect 5123 19465 5135 19499
rect 5077 19459 5135 19465
rect 5442 19456 5448 19508
rect 5500 19496 5506 19508
rect 6733 19499 6791 19505
rect 5500 19468 6500 19496
rect 5500 19456 5506 19468
rect 4982 19428 4988 19440
rect 1964 19400 4988 19428
rect 1964 19369 1992 19400
rect 4982 19388 4988 19400
rect 5040 19388 5046 19440
rect 5350 19388 5356 19440
rect 5408 19428 5414 19440
rect 6472 19428 6500 19468
rect 6733 19465 6745 19499
rect 6779 19496 6791 19499
rect 7006 19496 7012 19508
rect 6779 19468 7012 19496
rect 6779 19465 6791 19468
rect 6733 19459 6791 19465
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7282 19496 7288 19508
rect 7116 19468 7288 19496
rect 7116 19428 7144 19468
rect 7282 19456 7288 19468
rect 7340 19456 7346 19508
rect 7377 19499 7435 19505
rect 7377 19465 7389 19499
rect 7423 19496 7435 19499
rect 8113 19499 8171 19505
rect 8113 19496 8125 19499
rect 7423 19468 8125 19496
rect 7423 19465 7435 19468
rect 7377 19459 7435 19465
rect 8113 19465 8125 19468
rect 8159 19465 8171 19499
rect 8113 19459 8171 19465
rect 8662 19456 8668 19508
rect 8720 19496 8726 19508
rect 9401 19499 9459 19505
rect 9401 19496 9413 19499
rect 8720 19468 9413 19496
rect 8720 19456 8726 19468
rect 9401 19465 9413 19468
rect 9447 19465 9459 19499
rect 11882 19496 11888 19508
rect 9401 19459 9459 19465
rect 9508 19468 11888 19496
rect 5408 19400 5764 19428
rect 6472 19400 7144 19428
rect 5408 19388 5414 19400
rect 1949 19363 2007 19369
rect 1949 19329 1961 19363
rect 1995 19329 2007 19363
rect 1949 19323 2007 19329
rect 2038 19320 2044 19372
rect 2096 19360 2102 19372
rect 3706 19363 3764 19369
rect 3706 19360 3718 19363
rect 2096 19332 3718 19360
rect 2096 19320 2102 19332
rect 3706 19329 3718 19332
rect 3752 19329 3764 19363
rect 3706 19323 3764 19329
rect 3973 19363 4031 19369
rect 3973 19329 3985 19363
rect 4019 19360 4031 19363
rect 4341 19363 4399 19369
rect 4019 19332 4292 19360
rect 4019 19329 4031 19332
rect 3973 19323 4031 19329
rect 934 19252 940 19304
rect 992 19292 998 19304
rect 1118 19292 1124 19304
rect 992 19264 1124 19292
rect 992 19252 998 19264
rect 1118 19252 1124 19264
rect 1176 19292 1182 19304
rect 2225 19295 2283 19301
rect 2225 19292 2237 19295
rect 1176 19264 2237 19292
rect 1176 19252 1182 19264
rect 2225 19261 2237 19264
rect 2271 19261 2283 19295
rect 4264 19292 4292 19332
rect 4341 19329 4353 19363
rect 4387 19360 4399 19363
rect 4430 19360 4436 19372
rect 4387 19332 4436 19360
rect 4387 19329 4399 19332
rect 4341 19323 4399 19329
rect 4430 19320 4436 19332
rect 4488 19320 4494 19372
rect 5074 19320 5080 19372
rect 5132 19360 5138 19372
rect 5445 19363 5503 19369
rect 5445 19360 5457 19363
rect 5132 19332 5457 19360
rect 5132 19320 5138 19332
rect 5445 19329 5457 19332
rect 5491 19329 5503 19363
rect 5445 19323 5503 19329
rect 5166 19292 5172 19304
rect 4264 19264 5172 19292
rect 2225 19255 2283 19261
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 5537 19295 5595 19301
rect 5537 19292 5549 19295
rect 5460 19264 5549 19292
rect 5460 19236 5488 19264
rect 5537 19261 5549 19264
rect 5583 19261 5595 19295
rect 5537 19255 5595 19261
rect 5629 19295 5687 19301
rect 5629 19261 5641 19295
rect 5675 19261 5687 19295
rect 5736 19292 5764 19400
rect 7190 19388 7196 19440
rect 7248 19428 7254 19440
rect 9508 19428 9536 19468
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12805 19499 12863 19505
rect 12805 19496 12817 19499
rect 12544 19468 12817 19496
rect 7248 19400 9536 19428
rect 7248 19388 7254 19400
rect 5810 19320 5816 19372
rect 5868 19360 5874 19372
rect 6086 19360 6092 19372
rect 5868 19332 6092 19360
rect 5868 19320 5874 19332
rect 6086 19320 6092 19332
rect 6144 19320 6150 19372
rect 6546 19360 6552 19372
rect 6507 19332 6552 19360
rect 6546 19320 6552 19332
rect 6604 19320 6610 19372
rect 7190 19292 7196 19304
rect 5736 19264 7196 19292
rect 5629 19255 5687 19261
rect 566 19184 572 19236
rect 624 19224 630 19236
rect 2498 19224 2504 19236
rect 624 19196 2504 19224
rect 624 19184 630 19196
rect 2498 19184 2504 19196
rect 2556 19184 2562 19236
rect 4522 19224 4528 19236
rect 4483 19196 4528 19224
rect 4522 19184 4528 19196
rect 4580 19184 4586 19236
rect 5442 19184 5448 19236
rect 5500 19184 5506 19236
rect 4614 19116 4620 19168
rect 4672 19156 4678 19168
rect 5644 19156 5672 19255
rect 7190 19252 7196 19264
rect 7248 19252 7254 19304
rect 7300 19301 7328 19400
rect 9950 19388 9956 19440
rect 10008 19428 10014 19440
rect 10008 19400 12296 19428
rect 10008 19388 10014 19400
rect 7466 19360 7472 19372
rect 7427 19332 7472 19360
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 8481 19363 8539 19369
rect 8481 19329 8493 19363
rect 8527 19329 8539 19363
rect 8481 19323 8539 19329
rect 7285 19295 7343 19301
rect 7285 19261 7297 19295
rect 7331 19261 7343 19295
rect 7285 19255 7343 19261
rect 7374 19252 7380 19304
rect 7432 19292 7438 19304
rect 8496 19292 8524 19323
rect 8570 19320 8576 19372
rect 8628 19360 8634 19372
rect 8628 19332 8673 19360
rect 8628 19320 8634 19332
rect 8846 19320 8852 19372
rect 8904 19360 8910 19372
rect 9582 19360 9588 19372
rect 8904 19332 9588 19360
rect 8904 19320 8910 19332
rect 9582 19320 9588 19332
rect 9640 19320 9646 19372
rect 10502 19360 10508 19372
rect 10560 19369 10566 19372
rect 10472 19332 10508 19360
rect 10502 19320 10508 19332
rect 10560 19323 10572 19369
rect 10778 19360 10784 19372
rect 10739 19332 10784 19360
rect 10560 19320 10566 19323
rect 10778 19320 10784 19332
rect 10836 19320 10842 19372
rect 11146 19320 11152 19372
rect 11204 19360 11210 19372
rect 11793 19363 11851 19369
rect 11793 19360 11805 19363
rect 11204 19332 11805 19360
rect 11204 19320 11210 19332
rect 11793 19329 11805 19332
rect 11839 19329 11851 19363
rect 12268 19360 12296 19400
rect 12342 19388 12348 19440
rect 12400 19428 12406 19440
rect 12544 19428 12572 19468
rect 12805 19465 12817 19468
rect 12851 19465 12863 19499
rect 12805 19459 12863 19465
rect 13265 19499 13323 19505
rect 13265 19465 13277 19499
rect 13311 19465 13323 19499
rect 13906 19496 13912 19508
rect 13867 19468 13912 19496
rect 13265 19459 13323 19465
rect 13280 19428 13308 19459
rect 13906 19456 13912 19468
rect 13964 19456 13970 19508
rect 15197 19499 15255 19505
rect 15197 19465 15209 19499
rect 15243 19496 15255 19499
rect 15657 19499 15715 19505
rect 15243 19468 15608 19496
rect 15243 19465 15255 19468
rect 15197 19459 15255 19465
rect 12400 19400 12572 19428
rect 12636 19400 13308 19428
rect 12400 19388 12406 19400
rect 12268 19332 12388 19360
rect 11793 19323 11851 19329
rect 7432 19264 8524 19292
rect 8757 19295 8815 19301
rect 7432 19252 7438 19264
rect 8757 19261 8769 19295
rect 8803 19292 8815 19295
rect 9674 19292 9680 19304
rect 8803 19264 9680 19292
rect 8803 19261 8815 19264
rect 8757 19255 8815 19261
rect 9674 19252 9680 19264
rect 9732 19252 9738 19304
rect 12360 19224 12388 19332
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 12636 19224 12664 19400
rect 12986 19360 12992 19372
rect 12947 19332 12992 19360
rect 12986 19320 12992 19332
rect 13044 19320 13050 19372
rect 13449 19363 13507 19369
rect 13449 19360 13461 19363
rect 13096 19332 13461 19360
rect 12894 19252 12900 19304
rect 12952 19292 12958 19304
rect 13096 19292 13124 19332
rect 13449 19329 13461 19332
rect 13495 19329 13507 19363
rect 13722 19360 13728 19372
rect 13683 19332 13728 19360
rect 13449 19323 13507 19329
rect 13722 19320 13728 19332
rect 13780 19320 13786 19372
rect 14826 19360 14832 19372
rect 14787 19332 14832 19360
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 15473 19363 15531 19369
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 12952 19264 13124 19292
rect 14553 19295 14611 19301
rect 12952 19252 12958 19264
rect 14553 19261 14565 19295
rect 14599 19261 14611 19295
rect 14734 19292 14740 19304
rect 14695 19264 14740 19292
rect 14553 19255 14611 19261
rect 12360 19196 12664 19224
rect 12802 19184 12808 19236
rect 12860 19224 12866 19236
rect 14458 19224 14464 19236
rect 12860 19196 14464 19224
rect 12860 19184 12866 19196
rect 14458 19184 14464 19196
rect 14516 19184 14522 19236
rect 14568 19224 14596 19255
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 15497 19292 15525 19323
rect 15252 19264 15525 19292
rect 15252 19252 15258 19264
rect 15286 19224 15292 19236
rect 14568 19196 15292 19224
rect 15286 19184 15292 19196
rect 15344 19184 15350 19236
rect 15580 19224 15608 19468
rect 15657 19465 15669 19499
rect 15703 19465 15715 19499
rect 15657 19459 15715 19465
rect 15672 19428 15700 19459
rect 15746 19456 15752 19508
rect 15804 19496 15810 19508
rect 15933 19499 15991 19505
rect 15933 19496 15945 19499
rect 15804 19468 15945 19496
rect 15804 19456 15810 19468
rect 15933 19465 15945 19468
rect 15979 19465 15991 19499
rect 16669 19499 16727 19505
rect 15933 19459 15991 19465
rect 16040 19468 16620 19496
rect 16040 19428 16068 19468
rect 15672 19400 16068 19428
rect 16592 19428 16620 19468
rect 16669 19465 16681 19499
rect 16715 19496 16727 19499
rect 16942 19496 16948 19508
rect 16715 19468 16948 19496
rect 16715 19465 16727 19468
rect 16669 19459 16727 19465
rect 16942 19456 16948 19468
rect 17000 19456 17006 19508
rect 17129 19499 17187 19505
rect 17129 19465 17141 19499
rect 17175 19496 17187 19499
rect 17310 19496 17316 19508
rect 17175 19468 17316 19496
rect 17175 19465 17187 19468
rect 17129 19459 17187 19465
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 17586 19496 17592 19508
rect 17547 19468 17592 19496
rect 17586 19456 17592 19468
rect 17644 19456 17650 19508
rect 18233 19499 18291 19505
rect 18233 19465 18245 19499
rect 18279 19465 18291 19499
rect 18506 19496 18512 19508
rect 18467 19468 18512 19496
rect 18233 19459 18291 19465
rect 16592 19400 17816 19428
rect 16114 19360 16120 19372
rect 16075 19332 16120 19360
rect 16114 19320 16120 19332
rect 16172 19320 16178 19372
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17313 19363 17371 19369
rect 16908 19332 16953 19360
rect 16908 19320 16914 19332
rect 17313 19329 17325 19363
rect 17359 19360 17371 19363
rect 17402 19360 17408 19372
rect 17359 19332 17408 19360
rect 17359 19329 17371 19332
rect 17313 19323 17371 19329
rect 17402 19320 17408 19332
rect 17460 19320 17466 19372
rect 17788 19369 17816 19400
rect 17773 19363 17831 19369
rect 17773 19329 17785 19363
rect 17819 19329 17831 19363
rect 18049 19363 18107 19369
rect 18049 19360 18061 19363
rect 17773 19323 17831 19329
rect 17926 19332 18061 19360
rect 17926 19224 17954 19332
rect 18049 19329 18061 19332
rect 18095 19329 18107 19363
rect 18248 19360 18276 19459
rect 18506 19456 18512 19468
rect 18564 19456 18570 19508
rect 19153 19499 19211 19505
rect 19153 19465 19165 19499
rect 19199 19496 19211 19499
rect 19886 19496 19892 19508
rect 19199 19468 19892 19496
rect 19199 19465 19211 19468
rect 19153 19459 19211 19465
rect 19886 19456 19892 19468
rect 19944 19456 19950 19508
rect 19978 19456 19984 19508
rect 20036 19496 20042 19508
rect 20257 19499 20315 19505
rect 20257 19496 20269 19499
rect 20036 19468 20269 19496
rect 20036 19456 20042 19468
rect 20257 19465 20269 19468
rect 20303 19465 20315 19499
rect 20257 19459 20315 19465
rect 20438 19456 20444 19508
rect 20496 19496 20502 19508
rect 20809 19499 20867 19505
rect 20809 19496 20821 19499
rect 20496 19468 20821 19496
rect 20496 19456 20502 19468
rect 20809 19465 20821 19468
rect 20855 19465 20867 19499
rect 20809 19459 20867 19465
rect 18322 19388 18328 19440
rect 18380 19428 18386 19440
rect 18380 19400 19012 19428
rect 18380 19388 18386 19400
rect 18984 19369 19012 19400
rect 19518 19388 19524 19440
rect 19576 19428 19582 19440
rect 19576 19400 20116 19428
rect 19576 19388 19582 19400
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 18248 19332 18705 19360
rect 18049 19323 18107 19329
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 18969 19363 19027 19369
rect 18969 19329 18981 19363
rect 19015 19329 19027 19363
rect 18969 19323 19027 19329
rect 19426 19320 19432 19372
rect 19484 19320 19490 19372
rect 19610 19360 19616 19372
rect 19571 19332 19616 19360
rect 19610 19320 19616 19332
rect 19668 19320 19674 19372
rect 20088 19369 20116 19400
rect 20073 19363 20131 19369
rect 20073 19329 20085 19363
rect 20119 19329 20131 19363
rect 20622 19360 20628 19372
rect 20583 19332 20628 19360
rect 20073 19323 20131 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 21361 19363 21419 19369
rect 21361 19329 21373 19363
rect 21407 19360 21419 19363
rect 21726 19360 21732 19372
rect 21407 19332 21732 19360
rect 21407 19329 21419 19332
rect 21361 19323 21419 19329
rect 21726 19320 21732 19332
rect 21784 19320 21790 19372
rect 19444 19233 19472 19320
rect 15580 19196 17954 19224
rect 19429 19227 19487 19233
rect 19429 19193 19441 19227
rect 19475 19193 19487 19227
rect 19429 19187 19487 19193
rect 7834 19156 7840 19168
rect 4672 19128 5672 19156
rect 7795 19128 7840 19156
rect 4672 19116 4678 19128
rect 7834 19116 7840 19128
rect 7892 19116 7898 19168
rect 10410 19116 10416 19168
rect 10468 19156 10474 19168
rect 10870 19156 10876 19168
rect 10468 19128 10876 19156
rect 10468 19116 10474 19128
rect 10870 19116 10876 19128
rect 10928 19156 10934 19168
rect 11057 19159 11115 19165
rect 11057 19156 11069 19159
rect 10928 19128 11069 19156
rect 10928 19116 10934 19128
rect 11057 19125 11069 19128
rect 11103 19125 11115 19159
rect 11057 19119 11115 19125
rect 14274 19116 14280 19168
rect 14332 19156 14338 19168
rect 15838 19156 15844 19168
rect 14332 19128 15844 19156
rect 14332 19116 14338 19128
rect 15838 19116 15844 19128
rect 15896 19116 15902 19168
rect 21174 19156 21180 19168
rect 21135 19128 21180 19156
rect 21174 19116 21180 19128
rect 21232 19116 21238 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1765 18955 1823 18961
rect 1765 18921 1777 18955
rect 1811 18952 1823 18955
rect 4154 18952 4160 18964
rect 1811 18924 4160 18952
rect 1811 18921 1823 18924
rect 1765 18915 1823 18921
rect 4154 18912 4160 18924
rect 4212 18912 4218 18964
rect 5534 18952 5540 18964
rect 4632 18924 5540 18952
rect 1489 18887 1547 18893
rect 1489 18853 1501 18887
rect 1535 18884 1547 18887
rect 3694 18884 3700 18896
rect 1535 18856 3700 18884
rect 1535 18853 1547 18856
rect 1489 18847 1547 18853
rect 3694 18844 3700 18856
rect 3752 18844 3758 18896
rect 3878 18844 3884 18896
rect 3936 18884 3942 18896
rect 3973 18887 4031 18893
rect 3973 18884 3985 18887
rect 3936 18856 3985 18884
rect 3936 18844 3942 18856
rect 3973 18853 3985 18856
rect 4019 18853 4031 18887
rect 4632 18884 4660 18924
rect 5534 18912 5540 18924
rect 5592 18912 5598 18964
rect 6730 18952 6736 18964
rect 6691 18924 6736 18952
rect 6730 18912 6736 18924
rect 6788 18912 6794 18964
rect 8478 18912 8484 18964
rect 8536 18952 8542 18964
rect 8941 18955 8999 18961
rect 8941 18952 8953 18955
rect 8536 18924 8953 18952
rect 8536 18912 8542 18924
rect 8941 18921 8953 18924
rect 8987 18921 8999 18955
rect 10226 18952 10232 18964
rect 8941 18915 8999 18921
rect 9416 18924 10232 18952
rect 3973 18847 4031 18853
rect 4540 18856 4660 18884
rect 2866 18816 2872 18828
rect 2827 18788 2872 18816
rect 2866 18776 2872 18788
rect 2924 18776 2930 18828
rect 4540 18825 4568 18856
rect 4798 18844 4804 18896
rect 4856 18884 4862 18896
rect 4856 18856 5396 18884
rect 4856 18844 4862 18856
rect 4525 18819 4583 18825
rect 4525 18816 4537 18819
rect 3620 18788 4537 18816
rect 2409 18751 2467 18757
rect 2409 18717 2421 18751
rect 2455 18748 2467 18751
rect 3620 18748 3648 18788
rect 4525 18785 4537 18788
rect 4571 18785 4583 18819
rect 4525 18779 4583 18785
rect 4617 18819 4675 18825
rect 4617 18785 4629 18819
rect 4663 18816 4675 18819
rect 5258 18816 5264 18828
rect 4663 18788 5264 18816
rect 4663 18785 4675 18788
rect 4617 18779 4675 18785
rect 5258 18776 5264 18788
rect 5316 18776 5322 18828
rect 5368 18816 5396 18856
rect 7558 18844 7564 18896
rect 7616 18884 7622 18896
rect 9416 18884 9444 18924
rect 10226 18912 10232 18924
rect 10284 18912 10290 18964
rect 10502 18912 10508 18964
rect 10560 18952 10566 18964
rect 10597 18955 10655 18961
rect 10597 18952 10609 18955
rect 10560 18924 10609 18952
rect 10560 18912 10566 18924
rect 10597 18921 10609 18924
rect 10643 18921 10655 18955
rect 10597 18915 10655 18921
rect 10962 18912 10968 18964
rect 11020 18952 11026 18964
rect 15378 18952 15384 18964
rect 11020 18924 15384 18952
rect 11020 18912 11026 18924
rect 15378 18912 15384 18924
rect 15436 18912 15442 18964
rect 15470 18912 15476 18964
rect 15528 18952 15534 18964
rect 16025 18955 16083 18961
rect 16025 18952 16037 18955
rect 15528 18924 16037 18952
rect 15528 18912 15534 18924
rect 16025 18921 16037 18924
rect 16071 18921 16083 18955
rect 16025 18915 16083 18921
rect 18046 18912 18052 18964
rect 18104 18952 18110 18964
rect 18601 18955 18659 18961
rect 18601 18952 18613 18955
rect 18104 18924 18613 18952
rect 18104 18912 18110 18924
rect 18601 18921 18613 18924
rect 18647 18921 18659 18955
rect 18601 18915 18659 18921
rect 20898 18912 20904 18964
rect 20956 18952 20962 18964
rect 21177 18955 21235 18961
rect 21177 18952 21189 18955
rect 20956 18924 21189 18952
rect 20956 18912 20962 18924
rect 21177 18921 21189 18924
rect 21223 18921 21235 18955
rect 21177 18915 21235 18921
rect 11054 18884 11060 18896
rect 7616 18856 9444 18884
rect 9508 18856 11060 18884
rect 7616 18844 7622 18856
rect 5368 18788 5488 18816
rect 3786 18748 3792 18760
rect 2455 18720 3648 18748
rect 3747 18720 3792 18748
rect 2455 18717 2467 18720
rect 2409 18711 2467 18717
rect 3786 18708 3792 18720
rect 3844 18708 3850 18760
rect 5166 18708 5172 18760
rect 5224 18748 5230 18760
rect 5353 18751 5411 18757
rect 5353 18748 5365 18751
rect 5224 18720 5365 18748
rect 5224 18708 5230 18720
rect 5353 18717 5365 18720
rect 5399 18717 5411 18751
rect 5460 18748 5488 18788
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 9508 18825 9536 18856
rect 11054 18844 11060 18856
rect 11112 18844 11118 18896
rect 13814 18884 13820 18896
rect 11900 18856 13820 18884
rect 9493 18819 9551 18825
rect 8352 18788 8708 18816
rect 8352 18776 8358 18788
rect 5994 18748 6000 18760
rect 5460 18720 6000 18748
rect 5353 18711 5411 18717
rect 5994 18708 6000 18720
rect 6052 18708 6058 18760
rect 7006 18748 7012 18760
rect 6967 18720 7012 18748
rect 7006 18708 7012 18720
rect 7064 18708 7070 18760
rect 8202 18708 8208 18760
rect 8260 18748 8266 18760
rect 8573 18751 8631 18757
rect 8573 18748 8585 18751
rect 8260 18720 8585 18748
rect 8260 18708 8266 18720
rect 8573 18717 8585 18720
rect 8619 18717 8631 18751
rect 8680 18748 8708 18788
rect 9493 18785 9505 18819
rect 9539 18785 9551 18819
rect 9493 18779 9551 18785
rect 9585 18819 9643 18825
rect 9585 18785 9597 18819
rect 9631 18816 9643 18819
rect 9766 18816 9772 18828
rect 9631 18788 9772 18816
rect 9631 18785 9643 18788
rect 9585 18779 9643 18785
rect 9766 18776 9772 18788
rect 9824 18776 9830 18828
rect 11900 18816 11928 18856
rect 13814 18844 13820 18856
rect 13872 18844 13878 18896
rect 15746 18844 15752 18896
rect 15804 18844 15810 18896
rect 17865 18887 17923 18893
rect 17865 18853 17877 18887
rect 17911 18853 17923 18887
rect 17865 18847 17923 18853
rect 11072 18788 11928 18816
rect 11977 18819 12035 18825
rect 11072 18748 11100 18788
rect 11977 18785 11989 18819
rect 12023 18816 12035 18819
rect 12434 18816 12440 18828
rect 12023 18788 12440 18816
rect 12023 18785 12035 18788
rect 11977 18779 12035 18785
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 15764 18816 15792 18844
rect 15764 18788 17816 18816
rect 11238 18748 11244 18760
rect 8680 18720 11100 18748
rect 11199 18720 11244 18748
rect 8573 18711 8631 18717
rect 11238 18708 11244 18720
rect 11296 18708 11302 18760
rect 12618 18708 12624 18760
rect 12676 18748 12682 18760
rect 12805 18751 12863 18757
rect 12805 18748 12817 18751
rect 12676 18720 12817 18748
rect 12676 18708 12682 18720
rect 12805 18717 12817 18720
rect 12851 18717 12863 18751
rect 12805 18711 12863 18717
rect 15102 18708 15108 18760
rect 15160 18748 15166 18760
rect 15749 18751 15807 18757
rect 15749 18748 15761 18751
rect 15160 18720 15761 18748
rect 15160 18708 15166 18720
rect 15749 18717 15761 18720
rect 15795 18717 15807 18751
rect 15749 18711 15807 18717
rect 2682 18640 2688 18692
rect 2740 18680 2746 18692
rect 5598 18683 5656 18689
rect 5598 18680 5610 18683
rect 2740 18652 5610 18680
rect 2740 18640 2746 18652
rect 5598 18649 5610 18652
rect 5644 18649 5656 18683
rect 9490 18680 9496 18692
rect 5598 18643 5656 18649
rect 7484 18652 9496 18680
rect 2958 18612 2964 18624
rect 2919 18584 2964 18612
rect 2958 18572 2964 18584
rect 3016 18572 3022 18624
rect 3053 18615 3111 18621
rect 3053 18581 3065 18615
rect 3099 18612 3111 18615
rect 3234 18612 3240 18624
rect 3099 18584 3240 18612
rect 3099 18581 3111 18584
rect 3053 18575 3111 18581
rect 3234 18572 3240 18584
rect 3292 18572 3298 18624
rect 3418 18612 3424 18624
rect 3379 18584 3424 18612
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 3694 18572 3700 18624
rect 3752 18612 3758 18624
rect 4430 18612 4436 18624
rect 3752 18584 4436 18612
rect 3752 18572 3758 18584
rect 4430 18572 4436 18584
rect 4488 18572 4494 18624
rect 4706 18572 4712 18624
rect 4764 18612 4770 18624
rect 5077 18615 5135 18621
rect 4764 18584 4809 18612
rect 4764 18572 4770 18584
rect 5077 18581 5089 18615
rect 5123 18612 5135 18615
rect 7484 18612 7512 18652
rect 9490 18640 9496 18652
rect 9548 18640 9554 18692
rect 9677 18683 9735 18689
rect 9677 18649 9689 18683
rect 9723 18680 9735 18683
rect 11054 18680 11060 18692
rect 9723 18652 11060 18680
rect 9723 18649 9735 18652
rect 9677 18643 9735 18649
rect 11054 18640 11060 18652
rect 11112 18640 11118 18692
rect 15504 18683 15562 18689
rect 15504 18649 15516 18683
rect 15550 18680 15562 18683
rect 15764 18680 15792 18711
rect 15838 18708 15844 18760
rect 15896 18748 15902 18760
rect 16209 18751 16267 18757
rect 16209 18748 16221 18751
rect 15896 18720 16221 18748
rect 15896 18708 15902 18720
rect 16209 18717 16221 18720
rect 16255 18717 16267 18751
rect 16209 18711 16267 18717
rect 16298 18708 16304 18760
rect 16356 18748 16362 18760
rect 16761 18751 16819 18757
rect 16761 18748 16773 18751
rect 16356 18720 16773 18748
rect 16356 18708 16362 18720
rect 16761 18717 16773 18720
rect 16807 18717 16819 18751
rect 17678 18748 17684 18760
rect 17639 18720 17684 18748
rect 16761 18711 16819 18717
rect 17678 18708 17684 18720
rect 17736 18708 17742 18760
rect 17126 18680 17132 18692
rect 15550 18652 15700 18680
rect 15764 18652 17132 18680
rect 15550 18649 15562 18652
rect 15504 18643 15562 18649
rect 7650 18612 7656 18624
rect 5123 18584 7512 18612
rect 7611 18584 7656 18612
rect 5123 18581 5135 18584
rect 5077 18575 5135 18581
rect 7650 18572 7656 18584
rect 7708 18572 7714 18624
rect 7926 18612 7932 18624
rect 7887 18584 7932 18612
rect 7926 18572 7932 18584
rect 7984 18572 7990 18624
rect 10045 18615 10103 18621
rect 10045 18581 10057 18615
rect 10091 18612 10103 18615
rect 11698 18612 11704 18624
rect 10091 18584 11704 18612
rect 10091 18581 10103 18584
rect 10045 18575 10103 18581
rect 11698 18572 11704 18584
rect 11756 18572 11762 18624
rect 12066 18612 12072 18624
rect 12027 18584 12072 18612
rect 12066 18572 12072 18584
rect 12124 18572 12130 18624
rect 12158 18572 12164 18624
rect 12216 18612 12222 18624
rect 12526 18612 12532 18624
rect 12216 18584 12261 18612
rect 12487 18584 12532 18612
rect 12216 18572 12222 18584
rect 12526 18572 12532 18584
rect 12584 18572 12590 18624
rect 12802 18572 12808 18624
rect 12860 18612 12866 18624
rect 13449 18615 13507 18621
rect 13449 18612 13461 18615
rect 12860 18584 13461 18612
rect 12860 18572 12866 18584
rect 13449 18581 13461 18584
rect 13495 18581 13507 18615
rect 13449 18575 13507 18581
rect 13998 18572 14004 18624
rect 14056 18612 14062 18624
rect 14369 18615 14427 18621
rect 14369 18612 14381 18615
rect 14056 18584 14381 18612
rect 14056 18572 14062 18584
rect 14369 18581 14381 18584
rect 14415 18581 14427 18615
rect 15672 18612 15700 18652
rect 17126 18640 17132 18652
rect 17184 18680 17190 18692
rect 17586 18680 17592 18692
rect 17184 18652 17592 18680
rect 17184 18640 17190 18652
rect 17586 18640 17592 18652
rect 17644 18640 17650 18692
rect 17788 18680 17816 18788
rect 17880 18748 17908 18847
rect 17954 18844 17960 18896
rect 18012 18884 18018 18896
rect 18141 18887 18199 18893
rect 18141 18884 18153 18887
rect 18012 18856 18153 18884
rect 18012 18844 18018 18856
rect 18141 18853 18153 18856
rect 18187 18853 18199 18887
rect 18141 18847 18199 18853
rect 20533 18887 20591 18893
rect 20533 18853 20545 18887
rect 20579 18884 20591 18887
rect 21818 18884 21824 18896
rect 20579 18856 21824 18884
rect 20579 18853 20591 18856
rect 20533 18847 20591 18853
rect 21818 18844 21824 18856
rect 21876 18844 21882 18896
rect 21174 18816 21180 18828
rect 18800 18788 21180 18816
rect 18800 18757 18828 18788
rect 21174 18776 21180 18788
rect 21232 18776 21238 18828
rect 18325 18751 18383 18757
rect 18325 18748 18337 18751
rect 17880 18720 18337 18748
rect 18325 18717 18337 18720
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18785 18751 18843 18757
rect 18785 18717 18797 18751
rect 18831 18717 18843 18751
rect 18785 18711 18843 18717
rect 18874 18708 18880 18760
rect 18932 18748 18938 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18932 18720 19257 18748
rect 18932 18708 18938 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 20993 18751 21051 18757
rect 20993 18717 21005 18751
rect 21039 18748 21051 18751
rect 21634 18748 21640 18760
rect 21039 18720 21640 18748
rect 21039 18717 21051 18720
rect 20993 18711 21051 18717
rect 18414 18680 18420 18692
rect 17788 18652 18420 18680
rect 18414 18640 18420 18652
rect 18472 18640 18478 18692
rect 18506 18640 18512 18692
rect 18564 18680 18570 18692
rect 19720 18680 19748 18711
rect 18564 18652 19748 18680
rect 20732 18680 20760 18711
rect 21634 18708 21640 18720
rect 21692 18708 21698 18760
rect 21818 18680 21824 18692
rect 20732 18652 21824 18680
rect 18564 18640 18570 18652
rect 21818 18640 21824 18652
rect 21876 18640 21882 18692
rect 17405 18615 17463 18621
rect 17405 18612 17417 18615
rect 15672 18584 17417 18612
rect 14369 18575 14427 18581
rect 17405 18581 17417 18584
rect 17451 18581 17463 18615
rect 17405 18575 17463 18581
rect 19429 18615 19487 18621
rect 19429 18581 19441 18615
rect 19475 18612 19487 18615
rect 19794 18612 19800 18624
rect 19475 18584 19800 18612
rect 19475 18581 19487 18584
rect 19429 18575 19487 18581
rect 19794 18572 19800 18584
rect 19852 18572 19858 18624
rect 19889 18615 19947 18621
rect 19889 18581 19901 18615
rect 19935 18612 19947 18615
rect 20254 18612 20260 18624
rect 19935 18584 20260 18612
rect 19935 18581 19947 18584
rect 19889 18575 19947 18581
rect 20254 18572 20260 18584
rect 20312 18572 20318 18624
rect 1104 18522 21896 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21896 18522
rect 1104 18448 21896 18470
rect 1765 18411 1823 18417
rect 1765 18377 1777 18411
rect 1811 18408 1823 18411
rect 2038 18408 2044 18420
rect 1811 18380 2044 18408
rect 1811 18377 1823 18380
rect 1765 18371 1823 18377
rect 2038 18368 2044 18380
rect 2096 18368 2102 18420
rect 2682 18408 2688 18420
rect 2643 18380 2688 18408
rect 2682 18368 2688 18380
rect 2740 18368 2746 18420
rect 2958 18368 2964 18420
rect 3016 18408 3022 18420
rect 3605 18411 3663 18417
rect 3605 18408 3617 18411
rect 3016 18380 3617 18408
rect 3016 18368 3022 18380
rect 3605 18377 3617 18380
rect 3651 18377 3663 18411
rect 3605 18371 3663 18377
rect 3973 18411 4031 18417
rect 3973 18377 3985 18411
rect 4019 18408 4031 18411
rect 4154 18408 4160 18420
rect 4019 18380 4160 18408
rect 4019 18377 4031 18380
rect 3973 18371 4031 18377
rect 4154 18368 4160 18380
rect 4212 18368 4218 18420
rect 4614 18408 4620 18420
rect 4575 18380 4620 18408
rect 4614 18368 4620 18380
rect 4672 18368 4678 18420
rect 5810 18368 5816 18420
rect 5868 18408 5874 18420
rect 6549 18411 6607 18417
rect 5868 18380 6224 18408
rect 5868 18368 5874 18380
rect 4632 18340 4660 18368
rect 3344 18312 4660 18340
rect 3344 18281 3372 18312
rect 5166 18300 5172 18352
rect 5224 18340 5230 18352
rect 5224 18312 6040 18340
rect 5224 18300 5230 18312
rect 2409 18275 2467 18281
rect 2409 18241 2421 18275
rect 2455 18272 2467 18275
rect 3329 18275 3387 18281
rect 2455 18244 2774 18272
rect 2455 18241 2467 18244
rect 2409 18235 2467 18241
rect 2746 18204 2774 18244
rect 3329 18241 3341 18275
rect 3375 18241 3387 18275
rect 3329 18235 3387 18241
rect 3510 18232 3516 18284
rect 3568 18272 3574 18284
rect 3878 18272 3884 18284
rect 3568 18244 3884 18272
rect 3568 18232 3574 18244
rect 3878 18232 3884 18244
rect 3936 18232 3942 18284
rect 4065 18275 4123 18281
rect 4065 18241 4077 18275
rect 4111 18272 4123 18275
rect 4798 18272 4804 18284
rect 4111 18244 4804 18272
rect 4111 18241 4123 18244
rect 4065 18235 4123 18241
rect 4798 18232 4804 18244
rect 4856 18232 4862 18284
rect 5718 18232 5724 18284
rect 5776 18281 5782 18284
rect 6012 18281 6040 18312
rect 5776 18272 5788 18281
rect 5997 18275 6055 18281
rect 5776 18244 5821 18272
rect 5776 18235 5788 18244
rect 5997 18241 6009 18275
rect 6043 18241 6055 18275
rect 6196 18272 6224 18380
rect 6549 18377 6561 18411
rect 6595 18408 6607 18411
rect 6822 18408 6828 18420
rect 6595 18380 6828 18408
rect 6595 18377 6607 18380
rect 6549 18371 6607 18377
rect 6822 18368 6828 18380
rect 6880 18368 6886 18420
rect 7098 18368 7104 18420
rect 7156 18408 7162 18420
rect 8294 18408 8300 18420
rect 7156 18380 8300 18408
rect 7156 18368 7162 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8478 18368 8484 18420
rect 8536 18408 8542 18420
rect 9582 18408 9588 18420
rect 8536 18380 9588 18408
rect 8536 18368 8542 18380
rect 9582 18368 9588 18380
rect 9640 18368 9646 18420
rect 10042 18408 10048 18420
rect 10003 18380 10048 18408
rect 10042 18368 10048 18380
rect 10100 18368 10106 18420
rect 14734 18368 14740 18420
rect 14792 18408 14798 18420
rect 14921 18411 14979 18417
rect 14921 18408 14933 18411
rect 14792 18380 14933 18408
rect 14792 18368 14798 18380
rect 14921 18377 14933 18380
rect 14967 18377 14979 18411
rect 14921 18371 14979 18377
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 16298 18408 16304 18420
rect 15344 18380 16304 18408
rect 15344 18368 15350 18380
rect 16298 18368 16304 18380
rect 16356 18408 16362 18420
rect 16669 18411 16727 18417
rect 16669 18408 16681 18411
rect 16356 18380 16681 18408
rect 16356 18368 16362 18380
rect 16669 18377 16681 18380
rect 16715 18377 16727 18411
rect 16669 18371 16727 18377
rect 18598 18368 18604 18420
rect 18656 18408 18662 18420
rect 20165 18411 20223 18417
rect 20165 18408 20177 18411
rect 18656 18380 20177 18408
rect 18656 18368 18662 18380
rect 20165 18377 20177 18380
rect 20211 18377 20223 18411
rect 21266 18408 21272 18420
rect 21227 18380 21272 18408
rect 20165 18371 20223 18377
rect 21266 18368 21272 18380
rect 21324 18368 21330 18420
rect 7460 18343 7518 18349
rect 7460 18309 7472 18343
rect 7506 18340 7518 18343
rect 11790 18340 11796 18352
rect 7506 18312 11796 18340
rect 7506 18309 7518 18312
rect 7460 18303 7518 18309
rect 11790 18300 11796 18312
rect 11848 18300 11854 18352
rect 12250 18340 12256 18352
rect 11900 18312 12256 18340
rect 6365 18275 6423 18281
rect 6365 18272 6377 18275
rect 6196 18244 6377 18272
rect 5997 18235 6055 18241
rect 6365 18241 6377 18244
rect 6411 18241 6423 18275
rect 6365 18235 6423 18241
rect 5776 18232 5782 18235
rect 4157 18207 4215 18213
rect 2746 18176 4016 18204
rect 3988 18148 4016 18176
rect 4157 18173 4169 18207
rect 4203 18173 4215 18207
rect 6012 18204 6040 18235
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 9033 18275 9091 18281
rect 6512 18244 8984 18272
rect 6512 18232 6518 18244
rect 6914 18204 6920 18216
rect 6012 18176 6920 18204
rect 4157 18167 4215 18173
rect 2498 18096 2504 18148
rect 2556 18136 2562 18148
rect 3786 18136 3792 18148
rect 2556 18108 3792 18136
rect 2556 18096 2562 18108
rect 3786 18096 3792 18108
rect 3844 18096 3850 18148
rect 3970 18096 3976 18148
rect 4028 18136 4034 18148
rect 4172 18136 4200 18167
rect 6914 18164 6920 18176
rect 6972 18204 6978 18216
rect 7193 18207 7251 18213
rect 7193 18204 7205 18207
rect 6972 18176 7205 18204
rect 6972 18164 6978 18176
rect 7193 18173 7205 18176
rect 7239 18173 7251 18207
rect 8956 18204 8984 18244
rect 9033 18241 9045 18275
rect 9079 18272 9091 18275
rect 9766 18272 9772 18284
rect 9079 18244 9772 18272
rect 9079 18241 9091 18244
rect 9033 18235 9091 18241
rect 9766 18232 9772 18244
rect 9824 18232 9830 18284
rect 10321 18275 10379 18281
rect 10321 18241 10333 18275
rect 10367 18272 10379 18275
rect 10410 18272 10416 18284
rect 10367 18244 10416 18272
rect 10367 18241 10379 18244
rect 10321 18235 10379 18241
rect 10410 18232 10416 18244
rect 10468 18232 10474 18284
rect 11900 18204 11928 18312
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 12710 18300 12716 18352
rect 12768 18300 12774 18352
rect 12836 18343 12894 18349
rect 12836 18309 12848 18343
rect 12882 18340 12894 18343
rect 13538 18340 13544 18352
rect 12882 18312 13544 18340
rect 12882 18309 12894 18312
rect 12836 18303 12894 18309
rect 13538 18300 13544 18312
rect 13596 18340 13602 18352
rect 13998 18340 14004 18352
rect 13596 18312 14004 18340
rect 13596 18300 13602 18312
rect 13998 18300 14004 18312
rect 14056 18300 14062 18352
rect 14458 18300 14464 18352
rect 14516 18340 14522 18352
rect 15933 18343 15991 18349
rect 15933 18340 15945 18343
rect 14516 18312 15945 18340
rect 14516 18300 14522 18312
rect 15933 18309 15945 18312
rect 15979 18309 15991 18343
rect 15933 18303 15991 18309
rect 16390 18300 16396 18352
rect 16448 18340 16454 18352
rect 17494 18340 17500 18352
rect 16448 18312 17500 18340
rect 16448 18300 16454 18312
rect 17494 18300 17500 18312
rect 17552 18300 17558 18352
rect 17586 18300 17592 18352
rect 17644 18340 17650 18352
rect 17644 18312 18092 18340
rect 17644 18300 17650 18312
rect 12728 18272 12756 18300
rect 8956 18176 11928 18204
rect 11992 18244 12756 18272
rect 13081 18275 13139 18281
rect 7193 18167 7251 18173
rect 11992 18136 12020 18244
rect 13081 18241 13093 18275
rect 13127 18272 13139 18275
rect 13262 18272 13268 18284
rect 13127 18244 13268 18272
rect 13127 18241 13139 18244
rect 13081 18235 13139 18241
rect 13262 18232 13268 18244
rect 13320 18232 13326 18284
rect 13630 18232 13636 18284
rect 13688 18272 13694 18284
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13688 18244 13737 18272
rect 13688 18232 13694 18244
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 13872 18244 13917 18272
rect 13872 18232 13878 18244
rect 14090 18232 14096 18284
rect 14148 18272 14154 18284
rect 14553 18275 14611 18281
rect 14553 18272 14565 18275
rect 14148 18244 14565 18272
rect 14148 18232 14154 18244
rect 14553 18241 14565 18244
rect 14599 18241 14611 18275
rect 14553 18235 14611 18241
rect 15289 18275 15347 18281
rect 15289 18241 15301 18275
rect 15335 18272 15347 18275
rect 15746 18272 15752 18284
rect 15335 18244 15752 18272
rect 15335 18241 15347 18244
rect 15289 18235 15347 18241
rect 13998 18204 14004 18216
rect 13959 18176 14004 18204
rect 13998 18164 14004 18176
rect 14056 18164 14062 18216
rect 4028 18108 4200 18136
rect 8128 18108 12020 18136
rect 4028 18096 4034 18108
rect 1489 18071 1547 18077
rect 1489 18037 1501 18071
rect 1535 18068 1547 18071
rect 2866 18068 2872 18080
rect 1535 18040 2872 18068
rect 1535 18037 1547 18040
rect 1489 18031 1547 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 3418 18028 3424 18080
rect 3476 18068 3482 18080
rect 6822 18068 6828 18080
rect 3476 18040 6828 18068
rect 3476 18028 3482 18040
rect 6822 18028 6828 18040
rect 6880 18028 6886 18080
rect 7190 18028 7196 18080
rect 7248 18068 7254 18080
rect 8128 18068 8156 18108
rect 7248 18040 8156 18068
rect 7248 18028 7254 18040
rect 8202 18028 8208 18080
rect 8260 18068 8266 18080
rect 8573 18071 8631 18077
rect 8573 18068 8585 18071
rect 8260 18040 8585 18068
rect 8260 18028 8266 18040
rect 8573 18037 8585 18040
rect 8619 18037 8631 18071
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 8573 18031 8631 18037
rect 9674 18028 9680 18040
rect 9732 18028 9738 18080
rect 10962 18068 10968 18080
rect 10923 18040 10968 18068
rect 10962 18028 10968 18040
rect 11020 18028 11026 18080
rect 11701 18071 11759 18077
rect 11701 18037 11713 18071
rect 11747 18068 11759 18071
rect 12434 18068 12440 18080
rect 11747 18040 12440 18068
rect 11747 18037 11759 18040
rect 11701 18031 11759 18037
rect 12434 18028 12440 18040
rect 12492 18068 12498 18080
rect 13078 18068 13084 18080
rect 12492 18040 13084 18068
rect 12492 18028 12498 18040
rect 13078 18028 13084 18040
rect 13136 18028 13142 18080
rect 13354 18068 13360 18080
rect 13315 18040 13360 18068
rect 13354 18028 13360 18040
rect 13412 18028 13418 18080
rect 14366 18068 14372 18080
rect 14327 18040 14372 18068
rect 14366 18028 14372 18040
rect 14424 18028 14430 18080
rect 14568 18068 14596 18235
rect 15746 18232 15752 18244
rect 15804 18232 15810 18284
rect 16482 18232 16488 18284
rect 16540 18272 16546 18284
rect 18064 18281 18092 18312
rect 17782 18275 17840 18281
rect 17782 18272 17794 18275
rect 16540 18244 17794 18272
rect 16540 18232 16546 18244
rect 17782 18241 17794 18244
rect 17828 18241 17840 18275
rect 17782 18235 17840 18241
rect 18049 18275 18107 18281
rect 18049 18241 18061 18275
rect 18095 18241 18107 18275
rect 18322 18272 18328 18284
rect 18283 18244 18328 18272
rect 18049 18235 18107 18241
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 18414 18232 18420 18284
rect 18472 18272 18478 18284
rect 19429 18275 19487 18281
rect 19429 18272 19441 18275
rect 18472 18244 19441 18272
rect 18472 18232 18478 18244
rect 19429 18241 19441 18244
rect 19475 18241 19487 18275
rect 19429 18235 19487 18241
rect 15378 18204 15384 18216
rect 15339 18176 15384 18204
rect 15378 18164 15384 18176
rect 15436 18164 15442 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 16500 18204 16528 18232
rect 15611 18176 16528 18204
rect 19444 18204 19472 18235
rect 19794 18232 19800 18284
rect 19852 18272 19858 18284
rect 19889 18275 19947 18281
rect 19889 18272 19901 18275
rect 19852 18244 19901 18272
rect 19852 18232 19858 18244
rect 19889 18241 19901 18244
rect 19935 18241 19947 18275
rect 20346 18272 20352 18284
rect 20307 18244 20352 18272
rect 19889 18235 19947 18241
rect 20346 18232 20352 18244
rect 20404 18232 20410 18284
rect 20806 18272 20812 18284
rect 20767 18244 20812 18272
rect 20806 18232 20812 18244
rect 20864 18232 20870 18284
rect 21085 18275 21143 18281
rect 21085 18241 21097 18275
rect 21131 18272 21143 18275
rect 21542 18272 21548 18284
rect 21131 18244 21548 18272
rect 21131 18241 21143 18244
rect 21085 18235 21143 18241
rect 21542 18232 21548 18244
rect 21600 18232 21606 18284
rect 21174 18204 21180 18216
rect 19444 18176 21180 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 21174 18164 21180 18176
rect 21232 18164 21238 18216
rect 18046 18096 18052 18148
rect 18104 18136 18110 18148
rect 19245 18139 19303 18145
rect 19245 18136 19257 18139
rect 18104 18108 19257 18136
rect 18104 18096 18110 18108
rect 19245 18105 19257 18108
rect 19291 18105 19303 18139
rect 19702 18136 19708 18148
rect 19663 18108 19708 18136
rect 19245 18099 19303 18105
rect 19702 18096 19708 18108
rect 19760 18096 19766 18148
rect 20622 18136 20628 18148
rect 20583 18108 20628 18136
rect 20622 18096 20628 18108
rect 20680 18096 20686 18148
rect 18782 18068 18788 18080
rect 14568 18040 18788 18068
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 18966 18068 18972 18080
rect 18927 18040 18972 18068
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1581 17867 1639 17873
rect 1581 17833 1593 17867
rect 1627 17864 1639 17867
rect 5534 17864 5540 17876
rect 1627 17836 5540 17864
rect 1627 17833 1639 17836
rect 1581 17827 1639 17833
rect 5534 17824 5540 17836
rect 5592 17824 5598 17876
rect 5994 17824 6000 17876
rect 6052 17864 6058 17876
rect 10318 17864 10324 17876
rect 6052 17836 10324 17864
rect 6052 17824 6058 17836
rect 10318 17824 10324 17836
rect 10376 17824 10382 17876
rect 10597 17867 10655 17873
rect 10597 17833 10609 17867
rect 10643 17864 10655 17867
rect 11238 17864 11244 17876
rect 10643 17836 11244 17864
rect 10643 17833 10655 17836
rect 10597 17827 10655 17833
rect 11238 17824 11244 17836
rect 11296 17824 11302 17876
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 12618 17864 12624 17876
rect 12299 17836 12624 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 14826 17864 14832 17876
rect 14787 17836 14832 17864
rect 14826 17824 14832 17836
rect 14884 17824 14890 17876
rect 16482 17864 16488 17876
rect 14936 17836 16488 17864
rect 2866 17756 2872 17808
rect 2924 17796 2930 17808
rect 4154 17796 4160 17808
rect 2924 17768 4160 17796
rect 2924 17756 2930 17768
rect 4154 17756 4160 17768
rect 4212 17756 4218 17808
rect 5442 17756 5448 17808
rect 5500 17796 5506 17808
rect 5629 17799 5687 17805
rect 5629 17796 5641 17799
rect 5500 17768 5641 17796
rect 5500 17756 5506 17768
rect 5629 17765 5641 17768
rect 5675 17765 5687 17799
rect 5629 17759 5687 17765
rect 7282 17756 7288 17808
rect 7340 17796 7346 17808
rect 14734 17796 14740 17808
rect 7340 17768 8432 17796
rect 7340 17756 7346 17768
rect 5994 17688 6000 17740
rect 6052 17728 6058 17740
rect 6181 17731 6239 17737
rect 6181 17728 6193 17731
rect 6052 17700 6193 17728
rect 6052 17688 6058 17700
rect 6181 17697 6193 17700
rect 6227 17697 6239 17731
rect 6181 17691 6239 17697
rect 7006 17688 7012 17740
rect 7064 17728 7070 17740
rect 7377 17731 7435 17737
rect 7377 17728 7389 17731
rect 7064 17700 7389 17728
rect 7064 17688 7070 17700
rect 7377 17697 7389 17700
rect 7423 17697 7435 17731
rect 8404 17728 8432 17768
rect 11900 17768 14740 17796
rect 8938 17728 8944 17740
rect 8404 17700 8944 17728
rect 7377 17691 7435 17697
rect 8938 17688 8944 17700
rect 8996 17688 9002 17740
rect 9214 17728 9220 17740
rect 9175 17700 9220 17728
rect 9214 17688 9220 17700
rect 9272 17688 9278 17740
rect 750 17620 756 17672
rect 808 17660 814 17672
rect 1397 17663 1455 17669
rect 1397 17660 1409 17663
rect 808 17632 1409 17660
rect 808 17620 814 17632
rect 1397 17629 1409 17632
rect 1443 17660 1455 17663
rect 1486 17660 1492 17672
rect 1443 17632 1492 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1486 17620 1492 17632
rect 1544 17620 1550 17672
rect 2501 17663 2559 17669
rect 2501 17629 2513 17663
rect 2547 17660 2559 17663
rect 2682 17660 2688 17672
rect 2547 17632 2688 17660
rect 2547 17629 2559 17632
rect 2501 17623 2559 17629
rect 2682 17620 2688 17632
rect 2740 17620 2746 17672
rect 3421 17663 3479 17669
rect 3421 17629 3433 17663
rect 3467 17660 3479 17663
rect 5166 17660 5172 17672
rect 3467 17632 3832 17660
rect 5127 17632 5172 17660
rect 3467 17629 3479 17632
rect 3421 17623 3479 17629
rect 1857 17595 1915 17601
rect 1857 17561 1869 17595
rect 1903 17592 1915 17595
rect 2866 17592 2872 17604
rect 1903 17564 2872 17592
rect 1903 17561 1915 17564
rect 1857 17555 1915 17561
rect 2866 17552 2872 17564
rect 2924 17552 2930 17604
rect 2774 17484 2780 17536
rect 2832 17524 2838 17536
rect 3804 17533 3832 17632
rect 5166 17620 5172 17632
rect 5224 17620 5230 17672
rect 6546 17660 6552 17672
rect 5276 17632 6552 17660
rect 3878 17552 3884 17604
rect 3936 17592 3942 17604
rect 4902 17595 4960 17601
rect 4902 17592 4914 17595
rect 3936 17564 4914 17592
rect 3936 17552 3942 17564
rect 4902 17561 4914 17564
rect 4948 17561 4960 17595
rect 4902 17555 4960 17561
rect 3789 17527 3847 17533
rect 2832 17496 2877 17524
rect 2832 17484 2838 17496
rect 3789 17493 3801 17527
rect 3835 17524 3847 17527
rect 4338 17524 4344 17536
rect 3835 17496 4344 17524
rect 3835 17493 3847 17496
rect 3789 17487 3847 17493
rect 4338 17484 4344 17496
rect 4396 17484 4402 17536
rect 4430 17484 4436 17536
rect 4488 17524 4494 17536
rect 5276 17524 5304 17632
rect 6546 17620 6552 17632
rect 6604 17620 6610 17672
rect 8478 17620 8484 17672
rect 8536 17660 8542 17672
rect 8573 17663 8631 17669
rect 8573 17660 8585 17663
rect 8536 17632 8585 17660
rect 8536 17620 8542 17632
rect 8573 17629 8585 17632
rect 8619 17629 8631 17663
rect 9232 17660 9260 17688
rect 11146 17669 11152 17672
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 9232 17632 10885 17660
rect 8573 17623 8631 17629
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 11140 17660 11152 17669
rect 11107 17632 11152 17660
rect 10873 17623 10931 17629
rect 11140 17623 11152 17632
rect 11146 17620 11152 17623
rect 11204 17620 11210 17672
rect 5626 17552 5632 17604
rect 5684 17592 5690 17604
rect 6089 17595 6147 17601
rect 6089 17592 6101 17595
rect 5684 17564 6101 17592
rect 5684 17552 5690 17564
rect 6089 17561 6101 17564
rect 6135 17561 6147 17595
rect 6089 17555 6147 17561
rect 7193 17595 7251 17601
rect 7193 17561 7205 17595
rect 7239 17592 7251 17595
rect 9484 17595 9542 17601
rect 7239 17564 9444 17592
rect 7239 17561 7251 17564
rect 7193 17555 7251 17561
rect 4488 17496 5304 17524
rect 4488 17484 4494 17496
rect 5902 17484 5908 17536
rect 5960 17524 5966 17536
rect 5997 17527 6055 17533
rect 5997 17524 6009 17527
rect 5960 17496 6009 17524
rect 5960 17484 5966 17496
rect 5997 17493 6009 17496
rect 6043 17493 6055 17527
rect 5997 17487 6055 17493
rect 6730 17484 6736 17536
rect 6788 17524 6794 17536
rect 6825 17527 6883 17533
rect 6825 17524 6837 17527
rect 6788 17496 6837 17524
rect 6788 17484 6794 17496
rect 6825 17493 6837 17496
rect 6871 17493 6883 17527
rect 6825 17487 6883 17493
rect 7282 17484 7288 17536
rect 7340 17524 7346 17536
rect 7340 17496 7385 17524
rect 7340 17484 7346 17496
rect 7466 17484 7472 17536
rect 7524 17524 7530 17536
rect 7929 17527 7987 17533
rect 7929 17524 7941 17527
rect 7524 17496 7941 17524
rect 7524 17484 7530 17496
rect 7929 17493 7941 17496
rect 7975 17493 7987 17527
rect 9416 17524 9444 17564
rect 9484 17561 9496 17595
rect 9530 17592 9542 17595
rect 9674 17592 9680 17604
rect 9530 17564 9680 17592
rect 9530 17561 9542 17564
rect 9484 17555 9542 17561
rect 9674 17552 9680 17564
rect 9732 17552 9738 17604
rect 9858 17552 9864 17604
rect 9916 17592 9922 17604
rect 11900 17592 11928 17768
rect 14734 17756 14740 17768
rect 14792 17756 14798 17808
rect 13078 17728 13084 17740
rect 13039 17700 13084 17728
rect 13078 17688 13084 17700
rect 13136 17688 13142 17740
rect 14277 17731 14335 17737
rect 14277 17697 14289 17731
rect 14323 17728 14335 17731
rect 14936 17728 14964 17836
rect 16482 17824 16488 17836
rect 16540 17824 16546 17876
rect 19429 17867 19487 17873
rect 17236 17836 19380 17864
rect 15102 17728 15108 17740
rect 14323 17700 14964 17728
rect 15063 17700 15108 17728
rect 14323 17697 14335 17700
rect 14277 17691 14335 17697
rect 15102 17688 15108 17700
rect 15160 17688 15166 17740
rect 12897 17663 12955 17669
rect 12897 17629 12909 17663
rect 12943 17660 12955 17663
rect 13354 17660 13360 17672
rect 12943 17632 13360 17660
rect 12943 17629 12955 17632
rect 12897 17623 12955 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 14458 17660 14464 17672
rect 14419 17632 14464 17660
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 15838 17660 15844 17672
rect 14568 17632 15844 17660
rect 9916 17564 11928 17592
rect 9916 17552 9922 17564
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 13541 17595 13599 17601
rect 13541 17592 13553 17595
rect 12216 17564 13553 17592
rect 12216 17552 12222 17564
rect 13541 17561 13553 17564
rect 13587 17561 13599 17595
rect 13541 17555 13599 17561
rect 13630 17552 13636 17604
rect 13688 17592 13694 17604
rect 14568 17592 14596 17632
rect 15838 17620 15844 17632
rect 15896 17620 15902 17672
rect 16761 17663 16819 17669
rect 16761 17629 16773 17663
rect 16807 17660 16819 17663
rect 16942 17660 16948 17672
rect 16807 17632 16948 17660
rect 16807 17629 16819 17632
rect 16761 17623 16819 17629
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 13688 17564 14596 17592
rect 13688 17552 13694 17564
rect 14642 17552 14648 17604
rect 14700 17592 14706 17604
rect 15350 17595 15408 17601
rect 15350 17592 15362 17595
rect 14700 17564 15362 17592
rect 14700 17552 14706 17564
rect 15350 17561 15362 17564
rect 15396 17561 15408 17595
rect 15350 17555 15408 17561
rect 10502 17524 10508 17536
rect 9416 17496 10508 17524
rect 7929 17487 7987 17493
rect 10502 17484 10508 17496
rect 10560 17484 10566 17536
rect 12529 17527 12587 17533
rect 12529 17493 12541 17527
rect 12575 17524 12587 17527
rect 12618 17524 12624 17536
rect 12575 17496 12624 17524
rect 12575 17493 12587 17496
rect 12529 17487 12587 17493
rect 12618 17484 12624 17496
rect 12676 17484 12682 17536
rect 12989 17527 13047 17533
rect 12989 17493 13001 17527
rect 13035 17524 13047 17527
rect 13078 17524 13084 17536
rect 13035 17496 13084 17524
rect 13035 17493 13047 17496
rect 12989 17487 13047 17493
rect 13078 17484 13084 17496
rect 13136 17484 13142 17536
rect 14369 17527 14427 17533
rect 14369 17493 14381 17527
rect 14415 17524 14427 17527
rect 15010 17524 15016 17536
rect 14415 17496 15016 17524
rect 14415 17493 14427 17496
rect 14369 17487 14427 17493
rect 15010 17484 15016 17496
rect 15068 17484 15074 17536
rect 15102 17484 15108 17536
rect 15160 17524 15166 17536
rect 17236 17524 17264 17836
rect 18877 17799 18935 17805
rect 18877 17765 18889 17799
rect 18923 17796 18935 17799
rect 18923 17768 19288 17796
rect 18923 17765 18935 17768
rect 18877 17759 18935 17765
rect 17586 17688 17592 17740
rect 17644 17728 17650 17740
rect 17681 17731 17739 17737
rect 17681 17728 17693 17731
rect 17644 17700 17693 17728
rect 17644 17688 17650 17700
rect 17681 17697 17693 17700
rect 17727 17697 17739 17731
rect 17681 17691 17739 17697
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 18233 17731 18291 17737
rect 18233 17728 18245 17731
rect 18012 17700 18245 17728
rect 18012 17688 18018 17700
rect 18233 17697 18245 17700
rect 18279 17728 18291 17731
rect 18322 17728 18328 17740
rect 18279 17700 18328 17728
rect 18279 17697 18291 17700
rect 18233 17691 18291 17697
rect 18322 17688 18328 17700
rect 18380 17688 18386 17740
rect 19260 17669 19288 17768
rect 19245 17663 19303 17669
rect 19245 17629 19257 17663
rect 19291 17629 19303 17663
rect 19352 17660 19380 17836
rect 19429 17833 19441 17867
rect 19475 17864 19487 17867
rect 20346 17864 20352 17876
rect 19475 17836 20352 17864
rect 19475 17833 19487 17836
rect 19429 17827 19487 17833
rect 20346 17824 20352 17836
rect 20404 17824 20410 17876
rect 20530 17824 20536 17876
rect 20588 17864 20594 17876
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 20588 17836 20637 17864
rect 20588 17824 20594 17836
rect 20625 17833 20637 17836
rect 20671 17833 20683 17867
rect 20625 17827 20683 17833
rect 20898 17824 20904 17876
rect 20956 17864 20962 17876
rect 21085 17867 21143 17873
rect 21085 17864 21097 17867
rect 20956 17836 21097 17864
rect 20956 17824 20962 17836
rect 21085 17833 21097 17836
rect 21131 17833 21143 17867
rect 21085 17827 21143 17833
rect 19886 17688 19892 17740
rect 19944 17728 19950 17740
rect 19944 17700 20852 17728
rect 19944 17688 19950 17700
rect 20346 17660 20352 17672
rect 19352 17632 20352 17660
rect 19245 17623 19303 17629
rect 20346 17620 20352 17632
rect 20404 17620 20410 17672
rect 20824 17669 20852 17700
rect 20809 17663 20867 17669
rect 20809 17629 20821 17663
rect 20855 17629 20867 17663
rect 20809 17623 20867 17629
rect 21269 17663 21327 17669
rect 21269 17629 21281 17663
rect 21315 17629 21327 17663
rect 21269 17623 21327 17629
rect 18509 17595 18567 17601
rect 18509 17561 18521 17595
rect 18555 17592 18567 17595
rect 19705 17595 19763 17601
rect 19705 17592 19717 17595
rect 18555 17564 19717 17592
rect 18555 17561 18567 17564
rect 18509 17555 18567 17561
rect 19705 17561 19717 17564
rect 19751 17561 19763 17595
rect 19705 17555 19763 17561
rect 20070 17552 20076 17604
rect 20128 17592 20134 17604
rect 21284 17592 21312 17623
rect 20128 17564 21312 17592
rect 20128 17552 20134 17564
rect 17402 17524 17408 17536
rect 15160 17496 17264 17524
rect 17363 17496 17408 17524
rect 15160 17484 15166 17496
rect 17402 17484 17408 17496
rect 17460 17484 17466 17536
rect 18414 17524 18420 17536
rect 18375 17496 18420 17524
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18598 17484 18604 17536
rect 18656 17524 18662 17536
rect 20165 17527 20223 17533
rect 20165 17524 20177 17527
rect 18656 17496 20177 17524
rect 18656 17484 18662 17496
rect 20165 17493 20177 17496
rect 20211 17493 20223 17527
rect 20165 17487 20223 17493
rect 1104 17434 21896 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21896 17434
rect 1104 17360 21896 17382
rect 1670 17320 1676 17332
rect 1631 17292 1676 17320
rect 1670 17280 1676 17292
rect 1728 17280 1734 17332
rect 5258 17320 5264 17332
rect 1872 17292 5264 17320
rect 1872 17193 1900 17292
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 5353 17323 5411 17329
rect 5353 17289 5365 17323
rect 5399 17320 5411 17323
rect 5718 17320 5724 17332
rect 5399 17292 5724 17320
rect 5399 17289 5411 17292
rect 5353 17283 5411 17289
rect 5718 17280 5724 17292
rect 5776 17280 5782 17332
rect 5902 17280 5908 17332
rect 5960 17320 5966 17332
rect 6638 17320 6644 17332
rect 5960 17292 6644 17320
rect 5960 17280 5966 17292
rect 6638 17280 6644 17292
rect 6696 17280 6702 17332
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17320 6975 17323
rect 7006 17320 7012 17332
rect 6963 17292 7012 17320
rect 6963 17289 6975 17292
rect 6917 17283 6975 17289
rect 7006 17280 7012 17292
rect 7064 17280 7070 17332
rect 9033 17323 9091 17329
rect 7383 17292 8984 17320
rect 2774 17212 2780 17264
rect 2832 17252 2838 17264
rect 4258 17255 4316 17261
rect 4258 17252 4270 17255
rect 2832 17224 4270 17252
rect 2832 17212 2838 17224
rect 4258 17221 4270 17224
rect 4304 17221 4316 17255
rect 7383 17252 7411 17292
rect 4258 17215 4316 17221
rect 5085 17224 7411 17252
rect 1857 17187 1915 17193
rect 1857 17153 1869 17187
rect 1903 17153 1915 17187
rect 1857 17147 1915 17153
rect 2222 17144 2228 17196
rect 2280 17184 2286 17196
rect 2501 17187 2559 17193
rect 2501 17184 2513 17187
rect 2280 17156 2513 17184
rect 2280 17144 2286 17156
rect 2501 17153 2513 17156
rect 2547 17153 2559 17187
rect 2501 17147 2559 17153
rect 2593 17187 2651 17193
rect 2593 17153 2605 17187
rect 2639 17184 2651 17187
rect 3418 17184 3424 17196
rect 2639 17156 3424 17184
rect 2639 17153 2651 17156
rect 2593 17147 2651 17153
rect 3418 17144 3424 17156
rect 3476 17144 3482 17196
rect 4798 17184 4804 17196
rect 3528 17156 4804 17184
rect 2682 17116 2688 17128
rect 2643 17088 2688 17116
rect 2682 17076 2688 17088
rect 2740 17116 2746 17128
rect 2740 17076 2774 17116
rect 3050 17076 3056 17128
rect 3108 17116 3114 17128
rect 3528 17116 3556 17156
rect 4798 17144 4804 17156
rect 4856 17144 4862 17196
rect 5085 17193 5113 17224
rect 7926 17212 7932 17264
rect 7984 17252 7990 17264
rect 8030 17255 8088 17261
rect 8030 17252 8042 17255
rect 7984 17224 8042 17252
rect 7984 17212 7990 17224
rect 8030 17221 8042 17224
rect 8076 17221 8088 17255
rect 8956 17252 8984 17292
rect 9033 17289 9045 17323
rect 9079 17320 9091 17323
rect 9306 17320 9312 17332
rect 9079 17292 9312 17320
rect 9079 17289 9091 17292
rect 9033 17283 9091 17289
rect 9306 17280 9312 17292
rect 9364 17280 9370 17332
rect 9950 17320 9956 17332
rect 9416 17292 9956 17320
rect 9416 17252 9444 17292
rect 9950 17280 9956 17292
rect 10008 17280 10014 17332
rect 10045 17323 10103 17329
rect 10045 17289 10057 17323
rect 10091 17320 10103 17323
rect 10781 17323 10839 17329
rect 10781 17320 10793 17323
rect 10091 17292 10793 17320
rect 10091 17289 10103 17292
rect 10045 17283 10103 17289
rect 10781 17289 10793 17292
rect 10827 17289 10839 17323
rect 10781 17283 10839 17289
rect 11977 17323 12035 17329
rect 11977 17289 11989 17323
rect 12023 17320 12035 17323
rect 12066 17320 12072 17332
rect 12023 17292 12072 17320
rect 12023 17289 12035 17292
rect 11977 17283 12035 17289
rect 12066 17280 12072 17292
rect 12124 17280 12130 17332
rect 12989 17323 13047 17329
rect 12406 17292 12664 17320
rect 8956 17224 9444 17252
rect 9585 17255 9643 17261
rect 8030 17215 8088 17221
rect 9585 17221 9597 17255
rect 9631 17252 9643 17255
rect 12406 17252 12434 17292
rect 9631 17224 12434 17252
rect 12636 17252 12664 17292
rect 12989 17289 13001 17323
rect 13035 17320 13047 17323
rect 13078 17320 13084 17332
rect 13035 17292 13084 17320
rect 13035 17289 13047 17292
rect 12989 17283 13047 17289
rect 13078 17280 13084 17292
rect 13136 17280 13142 17332
rect 14642 17320 14648 17332
rect 14603 17292 14648 17320
rect 14642 17280 14648 17292
rect 14700 17280 14706 17332
rect 15194 17280 15200 17332
rect 15252 17320 15258 17332
rect 20714 17320 20720 17332
rect 15252 17292 20720 17320
rect 15252 17280 15258 17292
rect 20714 17280 20720 17292
rect 20772 17280 20778 17332
rect 12636 17224 16804 17252
rect 9631 17221 9643 17224
rect 9585 17215 9643 17221
rect 5077 17187 5135 17193
rect 5077 17153 5089 17187
rect 5123 17153 5135 17187
rect 5994 17184 6000 17196
rect 5907 17156 6000 17184
rect 5077 17147 5135 17153
rect 5994 17144 6000 17156
rect 6052 17184 6058 17196
rect 6270 17184 6276 17196
rect 6052 17156 6276 17184
rect 6052 17144 6058 17156
rect 6270 17144 6276 17156
rect 6328 17144 6334 17196
rect 6638 17184 6644 17196
rect 6599 17156 6644 17184
rect 6638 17144 6644 17156
rect 6696 17144 6702 17196
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17184 8907 17187
rect 9306 17184 9312 17196
rect 8895 17156 9312 17184
rect 8895 17153 8907 17156
rect 8849 17147 8907 17153
rect 9306 17144 9312 17156
rect 9364 17144 9370 17196
rect 9674 17184 9680 17196
rect 9635 17156 9680 17184
rect 9674 17144 9680 17156
rect 9732 17144 9738 17196
rect 10042 17144 10048 17196
rect 10100 17184 10106 17196
rect 10689 17187 10747 17193
rect 10689 17184 10701 17187
rect 10100 17156 10701 17184
rect 10100 17144 10106 17156
rect 10689 17153 10701 17156
rect 10735 17153 10747 17187
rect 10689 17147 10747 17153
rect 11701 17187 11759 17193
rect 11701 17153 11713 17187
rect 11747 17153 11759 17187
rect 11701 17147 11759 17153
rect 3108 17088 3556 17116
rect 4525 17119 4583 17125
rect 3108 17076 3114 17088
rect 4525 17085 4537 17119
rect 4571 17116 4583 17119
rect 4890 17116 4896 17128
rect 4571 17088 4896 17116
rect 4571 17085 4583 17088
rect 4525 17079 4583 17085
rect 4890 17076 4896 17088
rect 4948 17116 4954 17128
rect 5166 17116 5172 17128
rect 4948 17088 5172 17116
rect 4948 17076 4954 17088
rect 5166 17076 5172 17088
rect 5224 17076 5230 17128
rect 8294 17076 8300 17128
rect 8352 17116 8358 17128
rect 9214 17116 9220 17128
rect 8352 17088 9220 17116
rect 8352 17076 8358 17088
rect 9214 17076 9220 17088
rect 9272 17076 9278 17128
rect 9401 17119 9459 17125
rect 9401 17085 9413 17119
rect 9447 17085 9459 17119
rect 9858 17116 9864 17128
rect 9401 17079 9459 17085
rect 9646 17088 9864 17116
rect 2746 17048 2774 17076
rect 3145 17051 3203 17057
rect 3145 17048 3157 17051
rect 2746 17020 3157 17048
rect 3145 17017 3157 17020
rect 3191 17017 3203 17051
rect 6457 17051 6515 17057
rect 6457 17048 6469 17051
rect 3145 17011 3203 17017
rect 4632 17020 6469 17048
rect 1854 16940 1860 16992
rect 1912 16980 1918 16992
rect 2133 16983 2191 16989
rect 2133 16980 2145 16983
rect 1912 16952 2145 16980
rect 1912 16940 1918 16952
rect 2133 16949 2145 16952
rect 2179 16949 2191 16983
rect 2133 16943 2191 16949
rect 2406 16940 2412 16992
rect 2464 16980 2470 16992
rect 4632 16980 4660 17020
rect 6457 17017 6469 17020
rect 6503 17017 6515 17051
rect 9416 17048 9444 17079
rect 9646 17048 9674 17088
rect 9858 17076 9864 17088
rect 9916 17076 9922 17128
rect 10965 17119 11023 17125
rect 10965 17085 10977 17119
rect 11011 17116 11023 17119
rect 11238 17116 11244 17128
rect 11011 17088 11244 17116
rect 11011 17085 11023 17088
rect 10965 17079 11023 17085
rect 11238 17076 11244 17088
rect 11296 17076 11302 17128
rect 11716 17048 11744 17147
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12345 17187 12403 17193
rect 12345 17184 12357 17187
rect 11848 17156 12357 17184
rect 11848 17144 11854 17156
rect 12345 17153 12357 17156
rect 12391 17153 12403 17187
rect 13354 17184 13360 17196
rect 13315 17156 13360 17184
rect 12345 17147 12403 17153
rect 13354 17144 13360 17156
rect 13412 17144 13418 17196
rect 13449 17187 13507 17193
rect 13449 17153 13461 17187
rect 13495 17184 13507 17187
rect 13630 17184 13636 17196
rect 13495 17156 13636 17184
rect 13495 17153 13507 17156
rect 13449 17147 13507 17153
rect 13630 17144 13636 17156
rect 13688 17144 13694 17196
rect 14001 17187 14059 17193
rect 14001 17153 14013 17187
rect 14047 17153 14059 17187
rect 15286 17184 15292 17196
rect 15247 17156 15292 17184
rect 14001 17147 14059 17153
rect 12250 17076 12256 17128
rect 12308 17116 12314 17128
rect 12437 17119 12495 17125
rect 12437 17116 12449 17119
rect 12308 17088 12449 17116
rect 12308 17076 12314 17088
rect 12437 17085 12449 17088
rect 12483 17085 12495 17119
rect 12437 17079 12495 17085
rect 12621 17119 12679 17125
rect 12621 17085 12633 17119
rect 12667 17116 12679 17119
rect 13538 17116 13544 17128
rect 12667 17088 13544 17116
rect 12667 17085 12679 17088
rect 12621 17079 12679 17085
rect 13538 17076 13544 17088
rect 13596 17076 13602 17128
rect 14016 17116 14044 17147
rect 15286 17144 15292 17156
rect 15344 17144 15350 17196
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15528 17156 16681 17184
rect 15528 17144 15534 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16776 17184 16804 17224
rect 17126 17212 17132 17264
rect 17184 17252 17190 17264
rect 21269 17255 21327 17261
rect 21269 17252 21281 17255
rect 17184 17224 19380 17252
rect 17184 17212 17190 17224
rect 18598 17184 18604 17196
rect 16776 17156 18604 17184
rect 16669 17147 16727 17153
rect 18598 17144 18604 17156
rect 18656 17144 18662 17196
rect 19352 17193 19380 17224
rect 20732 17224 21281 17252
rect 19081 17187 19139 17193
rect 19081 17153 19093 17187
rect 19127 17184 19139 17187
rect 19337 17187 19395 17193
rect 19127 17156 19288 17184
rect 19127 17153 19139 17156
rect 19081 17147 19139 17153
rect 14274 17116 14280 17128
rect 14016 17088 14280 17116
rect 14274 17076 14280 17088
rect 14332 17116 14338 17128
rect 15105 17119 15163 17125
rect 15105 17116 15117 17119
rect 14332 17088 15117 17116
rect 14332 17076 14338 17088
rect 15105 17085 15117 17088
rect 15151 17085 15163 17119
rect 15105 17079 15163 17085
rect 15197 17119 15255 17125
rect 15197 17085 15209 17119
rect 15243 17116 15255 17119
rect 15562 17116 15568 17128
rect 15243 17088 15568 17116
rect 15243 17085 15255 17088
rect 15197 17079 15255 17085
rect 13078 17048 13084 17060
rect 9416 17020 9674 17048
rect 9876 17020 11652 17048
rect 11716 17020 13084 17048
rect 6457 17011 6515 17017
rect 2464 16952 4660 16980
rect 2464 16940 2470 16952
rect 4798 16940 4804 16992
rect 4856 16980 4862 16992
rect 4893 16983 4951 16989
rect 4893 16980 4905 16983
rect 4856 16952 4905 16980
rect 4856 16940 4862 16952
rect 4893 16949 4905 16952
rect 4939 16949 4951 16983
rect 4893 16943 4951 16949
rect 5166 16940 5172 16992
rect 5224 16980 5230 16992
rect 9876 16980 9904 17020
rect 5224 16952 9904 16980
rect 5224 16940 5230 16952
rect 9950 16940 9956 16992
rect 10008 16980 10014 16992
rect 10321 16983 10379 16989
rect 10321 16980 10333 16983
rect 10008 16952 10333 16980
rect 10008 16940 10014 16952
rect 10321 16949 10333 16952
rect 10367 16949 10379 16983
rect 10321 16943 10379 16949
rect 10686 16940 10692 16992
rect 10744 16980 10750 16992
rect 11517 16983 11575 16989
rect 11517 16980 11529 16983
rect 10744 16952 11529 16980
rect 10744 16940 10750 16952
rect 11517 16949 11529 16952
rect 11563 16949 11575 16983
rect 11624 16980 11652 17020
rect 13078 17008 13084 17020
rect 13136 17008 13142 17060
rect 15120 17048 15148 17079
rect 15562 17076 15568 17088
rect 15620 17076 15626 17128
rect 16114 17116 16120 17128
rect 16075 17088 16120 17116
rect 16114 17076 16120 17088
rect 16172 17076 16178 17128
rect 16206 17076 16212 17128
rect 16264 17116 16270 17128
rect 19260 17116 19288 17156
rect 19337 17153 19349 17187
rect 19383 17153 19395 17187
rect 19886 17184 19892 17196
rect 19847 17156 19892 17184
rect 19337 17147 19395 17153
rect 19886 17144 19892 17156
rect 19944 17144 19950 17196
rect 20622 17116 20628 17128
rect 16264 17088 17724 17116
rect 19260 17088 20628 17116
rect 16264 17076 16270 17088
rect 15120 17020 15240 17048
rect 14366 16980 14372 16992
rect 11624 16952 14372 16980
rect 11517 16943 11575 16949
rect 14366 16940 14372 16952
rect 14424 16940 14430 16992
rect 15212 16980 15240 17020
rect 15378 17008 15384 17060
rect 15436 17048 15442 17060
rect 15657 17051 15715 17057
rect 15657 17048 15669 17051
rect 15436 17020 15669 17048
rect 15436 17008 15442 17020
rect 15657 17017 15669 17020
rect 15703 17017 15715 17051
rect 15657 17011 15715 17017
rect 15838 17008 15844 17060
rect 15896 17048 15902 17060
rect 17589 17051 17647 17057
rect 17589 17048 17601 17051
rect 15896 17020 17601 17048
rect 15896 17008 15902 17020
rect 17589 17017 17601 17020
rect 17635 17017 17647 17051
rect 17589 17011 17647 17017
rect 16298 16980 16304 16992
rect 15212 16952 16304 16980
rect 16298 16940 16304 16952
rect 16356 16940 16362 16992
rect 16574 16940 16580 16992
rect 16632 16980 16638 16992
rect 17313 16983 17371 16989
rect 17313 16980 17325 16983
rect 16632 16952 17325 16980
rect 16632 16940 16638 16952
rect 17313 16949 17325 16952
rect 17359 16949 17371 16983
rect 17696 16980 17724 17088
rect 20622 17076 20628 17088
rect 20680 17076 20686 17128
rect 17954 17048 17960 17060
rect 17915 17020 17960 17048
rect 17954 17008 17960 17020
rect 18012 17008 18018 17060
rect 20732 17048 20760 17224
rect 21269 17221 21281 17224
rect 21315 17221 21327 17255
rect 21269 17215 21327 17221
rect 20809 17187 20867 17193
rect 20809 17153 20821 17187
rect 20855 17153 20867 17187
rect 20809 17147 20867 17153
rect 19352 17020 20760 17048
rect 19352 16980 19380 17020
rect 20824 16992 20852 17147
rect 20530 16980 20536 16992
rect 17696 16952 19380 16980
rect 20491 16952 20536 16980
rect 17313 16943 17371 16949
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 20806 16940 20812 16992
rect 20864 16940 20870 16992
rect 20990 16980 20996 16992
rect 20951 16952 20996 16980
rect 20990 16940 20996 16952
rect 21048 16940 21054 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 3418 16736 3424 16788
rect 3476 16776 3482 16788
rect 3789 16779 3847 16785
rect 3789 16776 3801 16779
rect 3476 16748 3801 16776
rect 3476 16736 3482 16748
rect 3789 16745 3801 16748
rect 3835 16745 3847 16779
rect 5166 16776 5172 16788
rect 3789 16739 3847 16745
rect 4724 16748 5172 16776
rect 2774 16668 2780 16720
rect 2832 16708 2838 16720
rect 4430 16708 4436 16720
rect 2832 16680 4436 16708
rect 2832 16668 2838 16680
rect 4430 16668 4436 16680
rect 4488 16668 4494 16720
rect 4338 16640 4344 16652
rect 4299 16612 4344 16640
rect 4338 16600 4344 16612
rect 4396 16600 4402 16652
rect 4724 16640 4752 16748
rect 5166 16736 5172 16748
rect 5224 16736 5230 16788
rect 6270 16776 6276 16788
rect 6231 16748 6276 16776
rect 6270 16736 6276 16748
rect 6328 16736 6334 16788
rect 7282 16736 7288 16788
rect 7340 16776 7346 16788
rect 7469 16779 7527 16785
rect 7469 16776 7481 16779
rect 7340 16748 7481 16776
rect 7340 16736 7346 16748
rect 7469 16745 7481 16748
rect 7515 16745 7527 16779
rect 7469 16739 7527 16745
rect 7742 16736 7748 16788
rect 7800 16776 7806 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 7800 16748 8493 16776
rect 7800 16736 7806 16748
rect 8481 16745 8493 16748
rect 8527 16776 8539 16779
rect 8527 16748 9168 16776
rect 8527 16745 8539 16748
rect 8481 16739 8539 16745
rect 9140 16708 9168 16748
rect 9214 16736 9220 16788
rect 9272 16776 9278 16788
rect 9272 16748 10364 16776
rect 9272 16736 9278 16748
rect 9306 16708 9312 16720
rect 9140 16680 9312 16708
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 4890 16640 4896 16652
rect 4448 16612 4752 16640
rect 4851 16612 4896 16640
rect 1397 16575 1455 16581
rect 1397 16541 1409 16575
rect 1443 16572 1455 16575
rect 1946 16572 1952 16584
rect 1443 16544 1952 16572
rect 1443 16541 1455 16544
rect 1397 16535 1455 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16541 2283 16575
rect 2225 16535 2283 16541
rect 2685 16575 2743 16581
rect 2685 16541 2697 16575
rect 2731 16572 2743 16575
rect 2958 16572 2964 16584
rect 2731 16544 2964 16572
rect 2731 16541 2743 16544
rect 2685 16535 2743 16541
rect 2240 16504 2268 16535
rect 2958 16532 2964 16544
rect 3016 16532 3022 16584
rect 3329 16575 3387 16581
rect 3329 16541 3341 16575
rect 3375 16572 3387 16575
rect 3878 16572 3884 16584
rect 3375 16544 3884 16572
rect 3375 16541 3387 16544
rect 3329 16535 3387 16541
rect 3878 16532 3884 16544
rect 3936 16532 3942 16584
rect 4154 16572 4160 16584
rect 4115 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4249 16575 4307 16581
rect 4249 16541 4261 16575
rect 4295 16572 4307 16575
rect 4448 16572 4476 16612
rect 4890 16600 4896 16612
rect 4948 16600 4954 16652
rect 7926 16640 7932 16652
rect 6380 16612 6684 16640
rect 7887 16612 7932 16640
rect 4295 16544 4476 16572
rect 4295 16541 4307 16544
rect 4249 16535 4307 16541
rect 4522 16532 4528 16584
rect 4580 16572 4586 16584
rect 6380 16572 6408 16612
rect 6546 16572 6552 16584
rect 4580 16544 6408 16572
rect 6507 16544 6552 16572
rect 4580 16532 4586 16544
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 6656 16572 6684 16612
rect 7926 16600 7932 16612
rect 7984 16600 7990 16652
rect 8110 16640 8116 16652
rect 8071 16612 8116 16640
rect 8110 16600 8116 16612
rect 8168 16600 8174 16652
rect 10336 16649 10364 16748
rect 12636 16748 13216 16776
rect 12636 16708 12664 16748
rect 11716 16680 12664 16708
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 11146 16600 11152 16652
rect 11204 16640 11210 16652
rect 11716 16640 11744 16680
rect 12710 16668 12716 16720
rect 12768 16668 12774 16720
rect 13188 16708 13216 16748
rect 13262 16736 13268 16788
rect 13320 16776 13326 16788
rect 15746 16776 15752 16788
rect 13320 16748 15516 16776
rect 15707 16748 15752 16776
rect 13320 16736 13326 16748
rect 13998 16708 14004 16720
rect 13188 16680 14004 16708
rect 13998 16668 14004 16680
rect 14056 16668 14062 16720
rect 14093 16711 14151 16717
rect 14093 16677 14105 16711
rect 14139 16708 14151 16711
rect 14274 16708 14280 16720
rect 14139 16680 14280 16708
rect 14139 16677 14151 16680
rect 14093 16671 14151 16677
rect 14274 16668 14280 16680
rect 14332 16668 14338 16720
rect 11882 16640 11888 16652
rect 11204 16612 11744 16640
rect 11843 16612 11888 16640
rect 11204 16600 11210 16612
rect 8386 16572 8392 16584
rect 6656 16544 8392 16572
rect 8386 16532 8392 16544
rect 8444 16572 8450 16584
rect 8662 16572 8668 16584
rect 8444 16544 8668 16572
rect 8444 16532 8450 16544
rect 8662 16532 8668 16544
rect 8720 16532 8726 16584
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 9674 16572 9680 16584
rect 8812 16544 9680 16572
rect 8812 16532 8818 16544
rect 9674 16532 9680 16544
rect 9732 16532 9738 16584
rect 10065 16575 10123 16581
rect 10065 16541 10077 16575
rect 10111 16572 10123 16575
rect 10962 16572 10968 16584
rect 10111 16544 10968 16572
rect 10111 16541 10123 16544
rect 10065 16535 10123 16541
rect 10962 16532 10968 16544
rect 11020 16532 11026 16584
rect 11716 16572 11744 16612
rect 11882 16600 11888 16612
rect 11940 16600 11946 16652
rect 12437 16643 12495 16649
rect 12437 16609 12449 16643
rect 12483 16640 12495 16643
rect 12728 16640 12756 16668
rect 12483 16612 12756 16640
rect 12483 16609 12495 16612
rect 12437 16603 12495 16609
rect 13354 16600 13360 16652
rect 13412 16640 13418 16652
rect 13538 16640 13544 16652
rect 13412 16612 13544 16640
rect 13412 16600 13418 16612
rect 13538 16600 13544 16612
rect 13596 16600 13602 16652
rect 15488 16649 15516 16748
rect 15746 16736 15752 16748
rect 15804 16736 15810 16788
rect 16853 16779 16911 16785
rect 16853 16745 16865 16779
rect 16899 16776 16911 16779
rect 17034 16776 17040 16788
rect 16899 16748 17040 16776
rect 16899 16745 16911 16748
rect 16853 16739 16911 16745
rect 17034 16736 17040 16748
rect 17092 16776 17098 16788
rect 17092 16748 18092 16776
rect 17092 16736 17098 16748
rect 18064 16708 18092 16748
rect 18414 16736 18420 16788
rect 18472 16776 18478 16788
rect 19245 16779 19303 16785
rect 19245 16776 19257 16779
rect 18472 16748 19257 16776
rect 18472 16736 18478 16748
rect 19245 16745 19257 16748
rect 19291 16745 19303 16779
rect 19245 16739 19303 16745
rect 21266 16708 21272 16720
rect 18064 16680 21272 16708
rect 15473 16643 15531 16649
rect 15473 16609 15485 16643
rect 15519 16609 15531 16643
rect 16298 16640 16304 16652
rect 16259 16612 16304 16640
rect 15473 16603 15531 16609
rect 16298 16600 16304 16612
rect 16356 16600 16362 16652
rect 17126 16640 17132 16652
rect 17087 16612 17132 16640
rect 17126 16600 17132 16612
rect 17184 16600 17190 16652
rect 18782 16640 18788 16652
rect 18743 16612 18788 16640
rect 18782 16600 18788 16612
rect 18840 16600 18846 16652
rect 19720 16649 19748 16680
rect 21266 16668 21272 16680
rect 21324 16668 21330 16720
rect 19705 16643 19763 16649
rect 19705 16609 19717 16643
rect 19751 16609 19763 16643
rect 19705 16603 19763 16609
rect 19797 16643 19855 16649
rect 19797 16609 19809 16643
rect 19843 16609 19855 16643
rect 19797 16603 19855 16609
rect 11793 16575 11851 16581
rect 11793 16572 11805 16575
rect 11716 16544 11805 16572
rect 11793 16541 11805 16544
rect 11839 16541 11851 16575
rect 11793 16535 11851 16541
rect 12526 16532 12532 16584
rect 12584 16572 12590 16584
rect 12713 16575 12771 16581
rect 12713 16572 12725 16575
rect 12584 16544 12725 16572
rect 12584 16532 12590 16544
rect 12713 16541 12725 16544
rect 12759 16541 12771 16575
rect 15217 16575 15275 16581
rect 12713 16535 12771 16541
rect 13004 16544 14596 16572
rect 952 16476 2268 16504
rect 952 16448 980 16476
rect 4338 16464 4344 16516
rect 4396 16504 4402 16516
rect 5138 16507 5196 16513
rect 5138 16504 5150 16507
rect 4396 16476 5150 16504
rect 4396 16464 4402 16476
rect 5138 16473 5150 16476
rect 5184 16473 5196 16507
rect 10686 16504 10692 16516
rect 5138 16467 5196 16473
rect 5276 16476 10692 16504
rect 934 16396 940 16448
rect 992 16396 998 16448
rect 1578 16436 1584 16448
rect 1539 16408 1584 16436
rect 1578 16396 1584 16408
rect 1636 16396 1642 16448
rect 2038 16436 2044 16448
rect 1999 16408 2044 16436
rect 2038 16396 2044 16408
rect 2096 16396 2102 16448
rect 3418 16396 3424 16448
rect 3476 16436 3482 16448
rect 4062 16436 4068 16448
rect 3476 16408 4068 16436
rect 3476 16396 3482 16408
rect 4062 16396 4068 16408
rect 4120 16396 4126 16448
rect 4430 16396 4436 16448
rect 4488 16436 4494 16448
rect 5276 16436 5304 16476
rect 10686 16464 10692 16476
rect 10744 16464 10750 16516
rect 10778 16464 10784 16516
rect 10836 16504 10842 16516
rect 12618 16504 12624 16516
rect 10836 16476 11744 16504
rect 12579 16476 12624 16504
rect 10836 16464 10842 16476
rect 7190 16436 7196 16448
rect 4488 16408 5304 16436
rect 7151 16408 7196 16436
rect 4488 16396 4494 16408
rect 7190 16396 7196 16408
rect 7248 16396 7254 16448
rect 7834 16436 7840 16448
rect 7795 16408 7840 16436
rect 7834 16396 7840 16408
rect 7892 16396 7898 16448
rect 8941 16439 8999 16445
rect 8941 16405 8953 16439
rect 8987 16436 8999 16439
rect 9858 16436 9864 16448
rect 8987 16408 9864 16436
rect 8987 16405 8999 16408
rect 8941 16399 8999 16405
rect 9858 16396 9864 16408
rect 9916 16396 9922 16448
rect 10318 16396 10324 16448
rect 10376 16436 10382 16448
rect 10597 16439 10655 16445
rect 10597 16436 10609 16439
rect 10376 16408 10609 16436
rect 10376 16396 10382 16408
rect 10597 16405 10609 16408
rect 10643 16405 10655 16439
rect 10597 16399 10655 16405
rect 11238 16396 11244 16448
rect 11296 16436 11302 16448
rect 11716 16445 11744 16476
rect 12618 16464 12624 16476
rect 12676 16464 12682 16516
rect 11333 16439 11391 16445
rect 11333 16436 11345 16439
rect 11296 16408 11345 16436
rect 11296 16396 11302 16408
rect 11333 16405 11345 16408
rect 11379 16405 11391 16439
rect 11333 16399 11391 16405
rect 11701 16439 11759 16445
rect 11701 16405 11713 16439
rect 11747 16436 11759 16439
rect 13004 16436 13032 16544
rect 13722 16504 13728 16516
rect 13096 16476 13728 16504
rect 13096 16445 13124 16476
rect 13722 16464 13728 16476
rect 13780 16464 13786 16516
rect 14568 16504 14596 16544
rect 15217 16541 15229 16575
rect 15263 16572 15275 16575
rect 16574 16572 16580 16584
rect 15263 16544 16580 16572
rect 15263 16541 15275 16544
rect 15217 16535 15275 16541
rect 16574 16532 16580 16544
rect 16632 16532 16638 16584
rect 17402 16581 17408 16584
rect 17396 16572 17408 16581
rect 17363 16544 17408 16572
rect 17396 16535 17408 16544
rect 17402 16532 17408 16535
rect 17460 16532 17466 16584
rect 19812 16572 19840 16603
rect 20257 16575 20315 16581
rect 20257 16572 20269 16575
rect 18524 16544 20269 16572
rect 16117 16507 16175 16513
rect 16117 16504 16129 16507
rect 14568 16476 16129 16504
rect 16117 16473 16129 16476
rect 16163 16504 16175 16507
rect 17218 16504 17224 16516
rect 16163 16476 17224 16504
rect 16163 16473 16175 16476
rect 16117 16467 16175 16473
rect 17218 16464 17224 16476
rect 17276 16464 17282 16516
rect 11747 16408 13032 16436
rect 13081 16439 13139 16445
rect 11747 16405 11759 16408
rect 11701 16399 11759 16405
rect 13081 16405 13093 16439
rect 13127 16405 13139 16439
rect 13354 16436 13360 16448
rect 13315 16408 13360 16436
rect 13081 16399 13139 16405
rect 13354 16396 13360 16408
rect 13412 16396 13418 16448
rect 13998 16396 14004 16448
rect 14056 16436 14062 16448
rect 16209 16439 16267 16445
rect 16209 16436 16221 16439
rect 14056 16408 16221 16436
rect 14056 16396 14062 16408
rect 16209 16405 16221 16408
rect 16255 16436 16267 16439
rect 16390 16436 16396 16448
rect 16255 16408 16396 16436
rect 16255 16405 16267 16408
rect 16209 16399 16267 16405
rect 16390 16396 16396 16408
rect 16448 16396 16454 16448
rect 18524 16445 18552 16544
rect 20257 16541 20269 16544
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20622 16532 20628 16584
rect 20680 16572 20686 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20680 16544 20913 16572
rect 20680 16532 20686 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 20990 16532 20996 16584
rect 21048 16572 21054 16584
rect 21361 16575 21419 16581
rect 21361 16572 21373 16575
rect 21048 16544 21373 16572
rect 21048 16532 21054 16544
rect 21361 16541 21373 16544
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 19613 16507 19671 16513
rect 19613 16473 19625 16507
rect 19659 16504 19671 16507
rect 19794 16504 19800 16516
rect 19659 16476 19800 16504
rect 19659 16473 19671 16476
rect 19613 16467 19671 16473
rect 19794 16464 19800 16476
rect 19852 16464 19858 16516
rect 18509 16439 18567 16445
rect 18509 16405 18521 16439
rect 18555 16405 18567 16439
rect 18509 16399 18567 16405
rect 21082 16396 21088 16448
rect 21140 16436 21146 16448
rect 21177 16439 21235 16445
rect 21177 16436 21189 16439
rect 21140 16408 21189 16436
rect 21140 16396 21146 16408
rect 21177 16405 21189 16408
rect 21223 16405 21235 16439
rect 21177 16399 21235 16405
rect 1104 16346 21896 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21896 16346
rect 1104 16272 21896 16294
rect 2130 16232 2136 16244
rect 2091 16204 2136 16232
rect 2130 16192 2136 16204
rect 2188 16192 2194 16244
rect 3142 16232 3148 16244
rect 3103 16204 3148 16232
rect 3142 16192 3148 16204
rect 3200 16192 3206 16244
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 4522 16232 4528 16244
rect 3743 16204 4528 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 4522 16192 4528 16204
rect 4580 16192 4586 16244
rect 5353 16235 5411 16241
rect 5353 16201 5365 16235
rect 5399 16232 5411 16235
rect 6365 16235 6423 16241
rect 6365 16232 6377 16235
rect 5399 16204 6377 16232
rect 5399 16201 5411 16204
rect 5353 16195 5411 16201
rect 6365 16201 6377 16204
rect 6411 16201 6423 16235
rect 8294 16232 8300 16244
rect 6365 16195 6423 16201
rect 6564 16204 8156 16232
rect 8255 16204 8300 16232
rect 198 16124 204 16176
rect 256 16164 262 16176
rect 2593 16167 2651 16173
rect 2593 16164 2605 16167
rect 256 16136 2605 16164
rect 256 16124 262 16136
rect 2593 16133 2605 16136
rect 2639 16133 2651 16167
rect 5994 16164 6000 16176
rect 5955 16136 6000 16164
rect 2593 16127 2651 16133
rect 5994 16124 6000 16136
rect 6052 16164 6058 16176
rect 6564 16164 6592 16204
rect 6052 16136 6592 16164
rect 8128 16164 8156 16204
rect 8294 16192 8300 16204
rect 8352 16192 8358 16244
rect 10778 16232 10784 16244
rect 8404 16204 10784 16232
rect 8404 16164 8432 16204
rect 10778 16192 10784 16204
rect 10836 16192 10842 16244
rect 11054 16192 11060 16244
rect 11112 16232 11118 16244
rect 13354 16232 13360 16244
rect 11112 16204 13360 16232
rect 11112 16192 11118 16204
rect 13354 16192 13360 16204
rect 13412 16192 13418 16244
rect 13449 16235 13507 16241
rect 13449 16201 13461 16235
rect 13495 16232 13507 16235
rect 13722 16232 13728 16244
rect 13495 16204 13728 16232
rect 13495 16201 13507 16204
rect 13449 16195 13507 16201
rect 13722 16192 13728 16204
rect 13780 16192 13786 16244
rect 13909 16235 13967 16241
rect 13909 16201 13921 16235
rect 13955 16232 13967 16235
rect 14550 16232 14556 16244
rect 13955 16204 14556 16232
rect 13955 16201 13967 16204
rect 13909 16195 13967 16201
rect 14550 16192 14556 16204
rect 14608 16192 14614 16244
rect 15289 16235 15347 16241
rect 15289 16201 15301 16235
rect 15335 16232 15347 16235
rect 15838 16232 15844 16244
rect 15335 16204 15844 16232
rect 15335 16201 15347 16204
rect 15289 16195 15347 16201
rect 15838 16192 15844 16204
rect 15896 16192 15902 16244
rect 15933 16235 15991 16241
rect 15933 16201 15945 16235
rect 15979 16232 15991 16235
rect 16114 16232 16120 16244
rect 15979 16204 16120 16232
rect 15979 16201 15991 16204
rect 15933 16195 15991 16201
rect 16114 16192 16120 16204
rect 16172 16192 16178 16244
rect 16669 16235 16727 16241
rect 16669 16201 16681 16235
rect 16715 16232 16727 16235
rect 16942 16232 16948 16244
rect 16715 16204 16948 16232
rect 16715 16201 16727 16204
rect 16669 16195 16727 16201
rect 12434 16164 12440 16176
rect 8128 16136 8432 16164
rect 9600 16136 12440 16164
rect 6052 16124 6058 16136
rect 1397 16099 1455 16105
rect 1397 16065 1409 16099
rect 1443 16096 1455 16099
rect 1670 16096 1676 16108
rect 1443 16068 1676 16096
rect 1443 16065 1455 16068
rect 1397 16059 1455 16065
rect 1670 16056 1676 16068
rect 1728 16056 1734 16108
rect 1762 16056 1768 16108
rect 1820 16096 1826 16108
rect 1949 16099 2007 16105
rect 1949 16096 1961 16099
rect 1820 16068 1961 16096
rect 1820 16056 1826 16068
rect 1949 16065 1961 16068
rect 1995 16065 2007 16099
rect 1949 16059 2007 16065
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16065 3387 16099
rect 3970 16096 3976 16108
rect 3931 16068 3976 16096
rect 3329 16059 3387 16065
rect 3344 16028 3372 16059
rect 3970 16056 3976 16068
rect 4028 16056 4034 16108
rect 4062 16056 4068 16108
rect 4120 16096 4126 16108
rect 5261 16099 5319 16105
rect 5261 16096 5273 16099
rect 4120 16068 5273 16096
rect 4120 16056 4126 16068
rect 5261 16065 5273 16068
rect 5307 16065 5319 16099
rect 5261 16059 5319 16065
rect 6733 16099 6791 16105
rect 6733 16065 6745 16099
rect 6779 16096 6791 16099
rect 6779 16068 7052 16096
rect 6779 16065 6791 16068
rect 6733 16059 6791 16065
rect 4430 16028 4436 16040
rect 3344 16000 4436 16028
rect 4430 15988 4436 16000
rect 4488 15988 4494 16040
rect 5442 16028 5448 16040
rect 5403 16000 5448 16028
rect 5442 15988 5448 16000
rect 5500 15988 5506 16040
rect 5534 15988 5540 16040
rect 5592 16028 5598 16040
rect 6825 16031 6883 16037
rect 6825 16028 6837 16031
rect 5592 16000 6837 16028
rect 5592 15988 5598 16000
rect 6825 15997 6837 16000
rect 6871 15997 6883 16031
rect 6825 15991 6883 15997
rect 6917 16031 6975 16037
rect 6917 15997 6929 16031
rect 6963 15997 6975 16031
rect 6917 15991 6975 15997
rect 2777 15963 2835 15969
rect 2777 15929 2789 15963
rect 2823 15960 2835 15963
rect 4798 15960 4804 15972
rect 2823 15932 4804 15960
rect 2823 15929 2835 15932
rect 2777 15923 2835 15929
rect 4798 15920 4804 15932
rect 4856 15920 4862 15972
rect 4893 15963 4951 15969
rect 4893 15929 4905 15963
rect 4939 15960 4951 15963
rect 4939 15932 6040 15960
rect 4939 15929 4951 15932
rect 4893 15923 4951 15929
rect 1578 15892 1584 15904
rect 1539 15864 1584 15892
rect 1578 15852 1584 15864
rect 1636 15852 1642 15904
rect 4614 15892 4620 15904
rect 4575 15864 4620 15892
rect 4614 15852 4620 15864
rect 4672 15852 4678 15904
rect 6012 15892 6040 15932
rect 6086 15920 6092 15972
rect 6144 15960 6150 15972
rect 6932 15960 6960 15991
rect 7024 15972 7052 16068
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7377 16099 7435 16105
rect 7377 16096 7389 16099
rect 7156 16068 7389 16096
rect 7156 16056 7162 16068
rect 7377 16065 7389 16068
rect 7423 16065 7435 16099
rect 7377 16059 7435 16065
rect 8294 16056 8300 16108
rect 8352 16096 8358 16108
rect 9600 16105 9628 16136
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 15470 16164 15476 16176
rect 13464 16136 15476 16164
rect 9585 16099 9643 16105
rect 9585 16096 9597 16099
rect 8352 16068 9597 16096
rect 8352 16056 8358 16068
rect 9585 16065 9597 16068
rect 9631 16065 9643 16099
rect 9585 16059 9643 16065
rect 10229 16099 10287 16105
rect 10229 16065 10241 16099
rect 10275 16096 10287 16099
rect 10873 16099 10931 16105
rect 10873 16096 10885 16099
rect 10275 16068 10885 16096
rect 10275 16065 10287 16068
rect 10229 16059 10287 16065
rect 10873 16065 10885 16068
rect 10919 16065 10931 16099
rect 10873 16059 10931 16065
rect 12641 16099 12699 16105
rect 12641 16065 12653 16099
rect 12687 16096 12699 16099
rect 12802 16096 12808 16108
rect 12687 16068 12808 16096
rect 12687 16065 12699 16068
rect 12641 16059 12699 16065
rect 12802 16056 12808 16068
rect 12860 16056 12866 16108
rect 12897 16099 12955 16105
rect 12897 16065 12909 16099
rect 12943 16096 12955 16099
rect 12986 16096 12992 16108
rect 12943 16068 12992 16096
rect 12943 16065 12955 16068
rect 12897 16059 12955 16065
rect 12986 16056 12992 16068
rect 13044 16096 13050 16108
rect 13354 16096 13360 16108
rect 13044 16068 13360 16096
rect 13044 16056 13050 16068
rect 13354 16056 13360 16068
rect 13412 16056 13418 16108
rect 10318 16028 10324 16040
rect 10279 16000 10324 16028
rect 10318 15988 10324 16000
rect 10376 15988 10382 16040
rect 10410 15988 10416 16040
rect 10468 16028 10474 16040
rect 13265 16031 13323 16037
rect 10468 16000 10513 16028
rect 10468 15988 10474 16000
rect 13265 15997 13277 16031
rect 13311 16028 13323 16031
rect 13464 16028 13492 16136
rect 15470 16124 15476 16136
rect 15528 16124 15534 16176
rect 13541 16099 13599 16105
rect 13541 16065 13553 16099
rect 13587 16096 13599 16099
rect 13814 16096 13820 16108
rect 13587 16068 13820 16096
rect 13587 16065 13599 16068
rect 13541 16059 13599 16065
rect 13814 16056 13820 16068
rect 13872 16056 13878 16108
rect 14553 16099 14611 16105
rect 14553 16065 14565 16099
rect 14599 16096 14611 16099
rect 16684 16096 16712 16195
rect 16942 16192 16948 16204
rect 17000 16192 17006 16244
rect 19886 16232 19892 16244
rect 17052 16204 18736 16232
rect 19847 16204 19892 16232
rect 14599 16068 15700 16096
rect 14599 16065 14611 16068
rect 14553 16059 14611 16065
rect 13311 16000 13492 16028
rect 13311 15997 13323 16000
rect 13265 15991 13323 15997
rect 13906 15988 13912 16040
rect 13964 16028 13970 16040
rect 14274 16028 14280 16040
rect 13964 16000 14280 16028
rect 13964 15988 13970 16000
rect 14274 15988 14280 16000
rect 14332 16028 14338 16040
rect 14645 16031 14703 16037
rect 14645 16028 14657 16031
rect 14332 16000 14657 16028
rect 14332 15988 14338 16000
rect 14645 15997 14657 16000
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 14792 16000 14837 16028
rect 14792 15988 14798 16000
rect 6144 15932 6960 15960
rect 6144 15920 6150 15932
rect 7006 15920 7012 15972
rect 7064 15920 7070 15972
rect 7098 15920 7104 15972
rect 7156 15960 7162 15972
rect 7156 15932 11652 15960
rect 7156 15920 7162 15932
rect 7282 15892 7288 15904
rect 6012 15864 7288 15892
rect 7282 15852 7288 15864
rect 7340 15852 7346 15904
rect 7561 15895 7619 15901
rect 7561 15861 7573 15895
rect 7607 15892 7619 15895
rect 9582 15892 9588 15904
rect 7607 15864 9588 15892
rect 7607 15861 7619 15864
rect 7561 15855 7619 15861
rect 9582 15852 9588 15864
rect 9640 15852 9646 15904
rect 9861 15895 9919 15901
rect 9861 15861 9873 15895
rect 9907 15892 9919 15895
rect 10134 15892 10140 15904
rect 9907 15864 10140 15892
rect 9907 15861 9919 15864
rect 9861 15855 9919 15861
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 11146 15852 11152 15904
rect 11204 15892 11210 15904
rect 11517 15895 11575 15901
rect 11517 15892 11529 15895
rect 11204 15864 11529 15892
rect 11204 15852 11210 15864
rect 11517 15861 11529 15864
rect 11563 15861 11575 15895
rect 11624 15892 11652 15932
rect 13354 15920 13360 15972
rect 13412 15960 13418 15972
rect 14185 15963 14243 15969
rect 14185 15960 14197 15963
rect 13412 15932 14197 15960
rect 13412 15920 13418 15932
rect 14185 15929 14197 15932
rect 14231 15929 14243 15963
rect 14185 15923 14243 15929
rect 13630 15892 13636 15904
rect 11624 15864 13636 15892
rect 11517 15855 11575 15861
rect 13630 15852 13636 15864
rect 13688 15852 13694 15904
rect 15672 15892 15700 16068
rect 15764 16068 16712 16096
rect 15764 16037 15792 16068
rect 15749 16031 15807 16037
rect 15749 15997 15761 16031
rect 15795 15997 15807 16031
rect 15749 15991 15807 15997
rect 15841 16031 15899 16037
rect 15841 15997 15853 16031
rect 15887 16028 15899 16031
rect 16942 16028 16948 16040
rect 15887 16000 16948 16028
rect 15887 15997 15899 16000
rect 15841 15991 15899 15997
rect 16942 15988 16948 16000
rect 17000 15988 17006 16040
rect 16301 15963 16359 15969
rect 16301 15929 16313 15963
rect 16347 15960 16359 15963
rect 17052 15960 17080 16204
rect 17126 16124 17132 16176
rect 17184 16164 17190 16176
rect 17184 16136 18092 16164
rect 17184 16124 17190 16136
rect 18064 16105 18092 16136
rect 17793 16099 17851 16105
rect 17793 16065 17805 16099
rect 17839 16096 17851 16099
rect 18049 16099 18107 16105
rect 17839 16068 18000 16096
rect 17839 16065 17851 16068
rect 17793 16059 17851 16065
rect 17972 16028 18000 16068
rect 18049 16065 18061 16099
rect 18095 16096 18107 16099
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 18095 16068 18521 16096
rect 18095 16065 18107 16068
rect 18049 16059 18107 16065
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18708 16096 18736 16204
rect 19886 16192 19892 16204
rect 19944 16192 19950 16244
rect 20165 16235 20223 16241
rect 20165 16201 20177 16235
rect 20211 16201 20223 16235
rect 20165 16195 20223 16201
rect 20717 16235 20775 16241
rect 20717 16201 20729 16235
rect 20763 16232 20775 16235
rect 20898 16232 20904 16244
rect 20763 16204 20904 16232
rect 20763 16201 20775 16204
rect 20717 16195 20775 16201
rect 18776 16167 18834 16173
rect 18776 16133 18788 16167
rect 18822 16164 18834 16167
rect 18966 16164 18972 16176
rect 18822 16136 18972 16164
rect 18822 16133 18834 16136
rect 18776 16127 18834 16133
rect 18966 16124 18972 16136
rect 19024 16124 19030 16176
rect 19058 16124 19064 16176
rect 19116 16164 19122 16176
rect 20180 16164 20208 16195
rect 20898 16192 20904 16204
rect 20956 16192 20962 16244
rect 19116 16136 20208 16164
rect 19116 16124 19122 16136
rect 18708 16068 19564 16096
rect 18509 16059 18567 16065
rect 19536 16028 19564 16068
rect 20254 16056 20260 16108
rect 20312 16096 20318 16108
rect 20349 16099 20407 16105
rect 20349 16096 20361 16099
rect 20312 16068 20361 16096
rect 20312 16056 20318 16068
rect 20349 16065 20361 16068
rect 20395 16065 20407 16099
rect 20349 16059 20407 16065
rect 21726 16028 21732 16040
rect 17972 16000 18552 16028
rect 19536 16000 21732 16028
rect 16347 15932 17080 15960
rect 16347 15929 16359 15932
rect 16301 15923 16359 15929
rect 17034 15892 17040 15904
rect 15672 15864 17040 15892
rect 17034 15852 17040 15864
rect 17092 15852 17098 15904
rect 18524 15892 18552 16000
rect 21726 15988 21732 16000
rect 21784 15988 21790 16040
rect 20622 15920 20628 15972
rect 20680 15960 20686 15972
rect 20993 15963 21051 15969
rect 20993 15960 21005 15963
rect 20680 15932 21005 15960
rect 20680 15920 20686 15932
rect 20993 15929 21005 15932
rect 21039 15929 21051 15963
rect 20993 15923 21051 15929
rect 19978 15892 19984 15904
rect 18524 15864 19984 15892
rect 19978 15852 19984 15864
rect 20036 15852 20042 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 1486 15648 1492 15700
rect 1544 15688 1550 15700
rect 2041 15691 2099 15697
rect 2041 15688 2053 15691
rect 1544 15660 2053 15688
rect 1544 15648 1550 15660
rect 2041 15657 2053 15660
rect 2087 15657 2099 15691
rect 2041 15651 2099 15657
rect 2590 15648 2596 15700
rect 2648 15688 2654 15700
rect 2685 15691 2743 15697
rect 2685 15688 2697 15691
rect 2648 15660 2697 15688
rect 2648 15648 2654 15660
rect 2685 15657 2697 15660
rect 2731 15657 2743 15691
rect 3234 15688 3240 15700
rect 3195 15660 3240 15688
rect 2685 15651 2743 15657
rect 3234 15648 3240 15660
rect 3292 15648 3298 15700
rect 4338 15688 4344 15700
rect 4299 15660 4344 15688
rect 4338 15648 4344 15660
rect 4396 15648 4402 15700
rect 8294 15688 8300 15700
rect 7024 15660 8300 15688
rect 3234 15552 3240 15564
rect 2240 15524 3240 15552
rect 1394 15484 1400 15496
rect 1355 15456 1400 15484
rect 1394 15444 1400 15456
rect 1452 15444 1458 15496
rect 2240 15493 2268 15524
rect 3234 15512 3240 15524
rect 3292 15512 3298 15564
rect 4890 15512 4896 15564
rect 4948 15552 4954 15564
rect 5166 15552 5172 15564
rect 4948 15524 5172 15552
rect 4948 15512 4954 15524
rect 5166 15512 5172 15524
rect 5224 15552 5230 15564
rect 5261 15555 5319 15561
rect 5261 15552 5273 15555
rect 5224 15524 5273 15552
rect 5224 15512 5230 15524
rect 5261 15521 5273 15524
rect 5307 15521 5319 15555
rect 5261 15515 5319 15521
rect 2225 15487 2283 15493
rect 2225 15453 2237 15487
rect 2271 15453 2283 15487
rect 2225 15447 2283 15453
rect 2501 15487 2559 15493
rect 2501 15453 2513 15487
rect 2547 15453 2559 15487
rect 2501 15447 2559 15453
rect 2130 15376 2136 15428
rect 2188 15416 2194 15428
rect 2516 15416 2544 15447
rect 2958 15444 2964 15496
rect 3016 15484 3022 15496
rect 3053 15487 3111 15493
rect 3053 15484 3065 15487
rect 3016 15456 3065 15484
rect 3016 15444 3022 15456
rect 3053 15453 3065 15456
rect 3099 15453 3111 15487
rect 3878 15484 3884 15496
rect 3839 15456 3884 15484
rect 3053 15447 3111 15453
rect 3878 15444 3884 15456
rect 3936 15444 3942 15496
rect 4982 15484 4988 15496
rect 4895 15456 4988 15484
rect 4982 15444 4988 15456
rect 5040 15484 5046 15496
rect 5442 15484 5448 15496
rect 5040 15456 5448 15484
rect 5040 15444 5046 15456
rect 5442 15444 5448 15456
rect 5500 15444 5506 15496
rect 5718 15444 5724 15496
rect 5776 15484 5782 15496
rect 6086 15484 6092 15496
rect 5776 15456 6092 15484
rect 5776 15444 5782 15456
rect 6086 15444 6092 15456
rect 6144 15444 6150 15496
rect 7024 15493 7052 15660
rect 8294 15648 8300 15660
rect 8352 15648 8358 15700
rect 8570 15688 8576 15700
rect 8531 15660 8576 15688
rect 8570 15648 8576 15660
rect 8628 15648 8634 15700
rect 9306 15648 9312 15700
rect 9364 15688 9370 15700
rect 10321 15691 10379 15697
rect 9364 15660 10272 15688
rect 9364 15648 9370 15660
rect 8386 15580 8392 15632
rect 8444 15580 8450 15632
rect 10244 15620 10272 15660
rect 10321 15657 10333 15691
rect 10367 15688 10379 15691
rect 10410 15688 10416 15700
rect 10367 15660 10416 15688
rect 10367 15657 10379 15660
rect 10321 15651 10379 15657
rect 10410 15648 10416 15660
rect 10468 15648 10474 15700
rect 10778 15648 10784 15700
rect 10836 15688 10842 15700
rect 12526 15688 12532 15700
rect 10836 15660 12532 15688
rect 10836 15648 10842 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 13722 15688 13728 15700
rect 13683 15660 13728 15688
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 17126 15688 17132 15700
rect 17087 15660 17132 15688
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 18417 15691 18475 15697
rect 18417 15657 18429 15691
rect 18463 15688 18475 15691
rect 18506 15688 18512 15700
rect 18463 15660 18512 15688
rect 18463 15657 18475 15660
rect 18417 15651 18475 15657
rect 18506 15648 18512 15660
rect 18564 15648 18570 15700
rect 18877 15691 18935 15697
rect 18877 15657 18889 15691
rect 18923 15688 18935 15691
rect 20070 15688 20076 15700
rect 18923 15660 20076 15688
rect 18923 15657 18935 15660
rect 18877 15651 18935 15657
rect 20070 15648 20076 15660
rect 20128 15648 20134 15700
rect 15562 15620 15568 15632
rect 10244 15592 11100 15620
rect 7929 15555 7987 15561
rect 7929 15521 7941 15555
rect 7975 15552 7987 15555
rect 8404 15552 8432 15580
rect 10428 15564 10456 15592
rect 8941 15555 8999 15561
rect 8941 15552 8953 15555
rect 7975 15524 8340 15552
rect 8404 15524 8953 15552
rect 7975 15521 7987 15524
rect 7929 15515 7987 15521
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 2188 15388 2544 15416
rect 2188 15376 2194 15388
rect 4154 15376 4160 15428
rect 4212 15416 4218 15428
rect 4798 15416 4804 15428
rect 4212 15388 4804 15416
rect 4212 15376 4218 15388
rect 4798 15376 4804 15388
rect 4856 15416 4862 15428
rect 7834 15416 7840 15428
rect 4856 15388 7840 15416
rect 4856 15376 4862 15388
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 8312 15416 8340 15524
rect 8941 15521 8953 15524
rect 8987 15521 8999 15555
rect 8941 15515 8999 15521
rect 10410 15512 10416 15564
rect 10468 15512 10474 15564
rect 8389 15487 8447 15493
rect 8389 15453 8401 15487
rect 8435 15484 8447 15487
rect 8662 15484 8668 15496
rect 8435 15456 8668 15484
rect 8435 15453 8447 15456
rect 8389 15447 8447 15453
rect 8662 15444 8668 15456
rect 8720 15444 8726 15496
rect 10778 15484 10784 15496
rect 9324 15456 10784 15484
rect 8478 15416 8484 15428
rect 8312 15388 8484 15416
rect 8478 15376 8484 15388
rect 8536 15376 8542 15428
rect 8570 15376 8576 15428
rect 8628 15416 8634 15428
rect 9186 15419 9244 15425
rect 9186 15416 9198 15419
rect 8628 15388 9198 15416
rect 8628 15376 8634 15388
rect 9186 15385 9198 15388
rect 9232 15385 9244 15419
rect 9186 15379 9244 15385
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 4065 15351 4123 15357
rect 4065 15317 4077 15351
rect 4111 15348 4123 15351
rect 4522 15348 4528 15360
rect 4111 15320 4528 15348
rect 4111 15317 4123 15320
rect 4065 15311 4123 15317
rect 4522 15308 4528 15320
rect 4580 15308 4586 15360
rect 6914 15308 6920 15360
rect 6972 15348 6978 15360
rect 7285 15351 7343 15357
rect 7285 15348 7297 15351
rect 6972 15320 7297 15348
rect 6972 15308 6978 15320
rect 7285 15317 7297 15320
rect 7331 15317 7343 15351
rect 7285 15311 7343 15317
rect 7374 15308 7380 15360
rect 7432 15348 7438 15360
rect 7653 15351 7711 15357
rect 7653 15348 7665 15351
rect 7432 15320 7665 15348
rect 7432 15308 7438 15320
rect 7653 15317 7665 15320
rect 7699 15317 7711 15351
rect 7653 15311 7711 15317
rect 7742 15308 7748 15360
rect 7800 15348 7806 15360
rect 7800 15320 7845 15348
rect 7800 15308 7806 15320
rect 8294 15308 8300 15360
rect 8352 15348 8358 15360
rect 9324 15348 9352 15456
rect 10778 15444 10784 15456
rect 10836 15444 10842 15496
rect 10870 15444 10876 15496
rect 10928 15484 10934 15496
rect 10965 15487 11023 15493
rect 10965 15484 10977 15487
rect 10928 15456 10977 15484
rect 10928 15444 10934 15456
rect 10965 15453 10977 15456
rect 11011 15453 11023 15487
rect 11072 15484 11100 15592
rect 13096 15592 15568 15620
rect 11146 15512 11152 15564
rect 11204 15552 11210 15564
rect 11882 15552 11888 15564
rect 11204 15524 11888 15552
rect 11204 15512 11210 15524
rect 11882 15512 11888 15524
rect 11940 15512 11946 15564
rect 13096 15552 13124 15592
rect 15562 15580 15568 15592
rect 15620 15580 15626 15632
rect 17218 15580 17224 15632
rect 17276 15620 17282 15632
rect 20257 15623 20315 15629
rect 20257 15620 20269 15623
rect 17276 15592 20269 15620
rect 17276 15580 17282 15592
rect 12406 15524 13124 15552
rect 13173 15555 13231 15561
rect 11793 15487 11851 15493
rect 11793 15484 11805 15487
rect 11072 15456 11805 15484
rect 10965 15447 11023 15453
rect 11793 15453 11805 15456
rect 11839 15484 11851 15487
rect 12406 15484 12434 15524
rect 13173 15521 13185 15555
rect 13219 15552 13231 15555
rect 14642 15552 14648 15564
rect 13219 15524 14648 15552
rect 13219 15521 13231 15524
rect 13173 15515 13231 15521
rect 14642 15512 14648 15524
rect 14700 15552 14706 15564
rect 17865 15555 17923 15561
rect 14700 15524 15056 15552
rect 14700 15512 14706 15524
rect 12526 15484 12532 15496
rect 11839 15456 12434 15484
rect 12487 15456 12532 15484
rect 11839 15453 11851 15456
rect 11793 15447 11851 15453
rect 12526 15444 12532 15456
rect 12584 15444 12590 15496
rect 13354 15484 13360 15496
rect 13315 15456 13360 15484
rect 13354 15444 13360 15456
rect 13412 15444 13418 15496
rect 15028 15493 15056 15524
rect 17865 15521 17877 15555
rect 17911 15552 17923 15555
rect 19426 15552 19432 15564
rect 17911 15524 19432 15552
rect 17911 15521 17923 15524
rect 17865 15515 17923 15521
rect 19426 15512 19432 15524
rect 19484 15512 19490 15564
rect 19720 15561 19748 15592
rect 20257 15589 20269 15592
rect 20303 15620 20315 15623
rect 20625 15623 20683 15629
rect 20625 15620 20637 15623
rect 20303 15592 20637 15620
rect 20303 15589 20315 15592
rect 20257 15583 20315 15589
rect 20625 15589 20637 15592
rect 20671 15589 20683 15623
rect 20625 15583 20683 15589
rect 19705 15555 19763 15561
rect 19705 15521 19717 15555
rect 19751 15521 19763 15555
rect 19886 15552 19892 15564
rect 19847 15524 19892 15552
rect 19705 15515 19763 15521
rect 19886 15512 19892 15524
rect 19944 15512 19950 15564
rect 15013 15487 15071 15493
rect 15013 15453 15025 15487
rect 15059 15453 15071 15487
rect 15013 15447 15071 15453
rect 18230 15444 18236 15496
rect 18288 15484 18294 15496
rect 18693 15487 18751 15493
rect 18693 15484 18705 15487
rect 18288 15456 18705 15484
rect 18288 15444 18294 15456
rect 18693 15453 18705 15456
rect 18739 15453 18751 15487
rect 18693 15447 18751 15453
rect 9766 15376 9772 15428
rect 9824 15416 9830 15428
rect 9824 15388 12388 15416
rect 9824 15376 9830 15388
rect 8352 15320 9352 15348
rect 8352 15308 8358 15320
rect 9674 15308 9680 15360
rect 9732 15348 9738 15360
rect 10781 15351 10839 15357
rect 10781 15348 10793 15351
rect 9732 15320 10793 15348
rect 9732 15308 9738 15320
rect 10781 15317 10793 15320
rect 10827 15317 10839 15351
rect 10781 15311 10839 15317
rect 11054 15308 11060 15360
rect 11112 15348 11118 15360
rect 11333 15351 11391 15357
rect 11333 15348 11345 15351
rect 11112 15320 11345 15348
rect 11112 15308 11118 15320
rect 11333 15317 11345 15320
rect 11379 15317 11391 15351
rect 11333 15311 11391 15317
rect 11701 15351 11759 15357
rect 11701 15317 11713 15351
rect 11747 15348 11759 15351
rect 11974 15348 11980 15360
rect 11747 15320 11980 15348
rect 11747 15317 11759 15320
rect 11701 15311 11759 15317
rect 11974 15308 11980 15320
rect 12032 15308 12038 15360
rect 12360 15357 12388 15388
rect 12434 15376 12440 15428
rect 12492 15416 12498 15428
rect 15657 15419 15715 15425
rect 15657 15416 15669 15419
rect 12492 15388 15669 15416
rect 12492 15376 12498 15388
rect 15657 15385 15669 15388
rect 15703 15385 15715 15419
rect 15657 15379 15715 15385
rect 17957 15419 18015 15425
rect 17957 15385 17969 15419
rect 18003 15416 18015 15419
rect 20993 15419 21051 15425
rect 20993 15416 21005 15419
rect 18003 15388 19288 15416
rect 18003 15385 18015 15388
rect 17957 15379 18015 15385
rect 12345 15351 12403 15357
rect 12345 15317 12357 15351
rect 12391 15317 12403 15351
rect 13262 15348 13268 15360
rect 13223 15320 13268 15348
rect 12345 15311 12403 15317
rect 13262 15308 13268 15320
rect 13320 15308 13326 15360
rect 14366 15348 14372 15360
rect 14327 15320 14372 15348
rect 14366 15308 14372 15320
rect 14424 15308 14430 15360
rect 15102 15308 15108 15360
rect 15160 15348 15166 15360
rect 15289 15351 15347 15357
rect 15289 15348 15301 15351
rect 15160 15320 15301 15348
rect 15160 15308 15166 15320
rect 15289 15317 15301 15320
rect 15335 15317 15347 15351
rect 18046 15348 18052 15360
rect 18007 15320 18052 15348
rect 15289 15311 15347 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 19260 15357 19288 15388
rect 19628 15388 21005 15416
rect 19628 15360 19656 15388
rect 20993 15385 21005 15388
rect 21039 15385 21051 15419
rect 20993 15379 21051 15385
rect 19245 15351 19303 15357
rect 19245 15317 19257 15351
rect 19291 15317 19303 15351
rect 19610 15348 19616 15360
rect 19571 15320 19616 15348
rect 19245 15311 19303 15317
rect 19610 15308 19616 15320
rect 19668 15308 19674 15360
rect 1104 15258 21896 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21896 15258
rect 1104 15184 21896 15206
rect 1486 15104 1492 15156
rect 1544 15144 1550 15156
rect 2041 15147 2099 15153
rect 2041 15144 2053 15147
rect 1544 15116 2053 15144
rect 1544 15104 1550 15116
rect 2041 15113 2053 15116
rect 2087 15113 2099 15147
rect 2041 15107 2099 15113
rect 3970 15104 3976 15156
rect 4028 15144 4034 15156
rect 4157 15147 4215 15153
rect 4157 15144 4169 15147
rect 4028 15116 4169 15144
rect 4028 15104 4034 15116
rect 4157 15113 4169 15116
rect 4203 15113 4215 15147
rect 4157 15107 4215 15113
rect 4617 15147 4675 15153
rect 4617 15113 4629 15147
rect 4663 15144 4675 15147
rect 4982 15144 4988 15156
rect 4663 15116 4988 15144
rect 4663 15113 4675 15116
rect 4617 15107 4675 15113
rect 4982 15104 4988 15116
rect 5040 15104 5046 15156
rect 5258 15104 5264 15156
rect 5316 15144 5322 15156
rect 6365 15147 6423 15153
rect 6365 15144 6377 15147
rect 5316 15116 6377 15144
rect 5316 15104 5322 15116
rect 6365 15113 6377 15116
rect 6411 15113 6423 15147
rect 8478 15144 8484 15156
rect 8439 15116 8484 15144
rect 6365 15107 6423 15113
rect 8478 15104 8484 15116
rect 8536 15104 8542 15156
rect 9030 15104 9036 15156
rect 9088 15144 9094 15156
rect 9217 15147 9275 15153
rect 9217 15144 9229 15147
rect 9088 15116 9229 15144
rect 9088 15104 9094 15116
rect 9217 15113 9229 15116
rect 9263 15144 9275 15147
rect 9306 15144 9312 15156
rect 9263 15116 9312 15144
rect 9263 15113 9275 15116
rect 9217 15107 9275 15113
rect 9306 15104 9312 15116
rect 9364 15104 9370 15156
rect 9585 15147 9643 15153
rect 9585 15113 9597 15147
rect 9631 15144 9643 15147
rect 10318 15144 10324 15156
rect 9631 15116 10324 15144
rect 9631 15113 9643 15116
rect 9585 15107 9643 15113
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 10689 15147 10747 15153
rect 10689 15113 10701 15147
rect 10735 15144 10747 15147
rect 11054 15144 11060 15156
rect 10735 15116 11060 15144
rect 10735 15113 10747 15116
rect 10689 15107 10747 15113
rect 11054 15104 11060 15116
rect 11112 15104 11118 15156
rect 11149 15147 11207 15153
rect 11149 15113 11161 15147
rect 11195 15144 11207 15147
rect 11793 15147 11851 15153
rect 11793 15144 11805 15147
rect 11195 15116 11805 15144
rect 11195 15113 11207 15116
rect 11149 15107 11207 15113
rect 11793 15113 11805 15116
rect 11839 15113 11851 15147
rect 11793 15107 11851 15113
rect 11882 15104 11888 15156
rect 11940 15144 11946 15156
rect 12253 15147 12311 15153
rect 11940 15116 11985 15144
rect 11940 15104 11946 15116
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 12529 15147 12587 15153
rect 12299 15116 12434 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 5166 15076 5172 15088
rect 2792 15048 5172 15076
rect 1210 14968 1216 15020
rect 1268 15008 1274 15020
rect 2792 15017 2820 15048
rect 5166 15036 5172 15048
rect 5224 15076 5230 15088
rect 7368 15079 7426 15085
rect 5224 15048 7144 15076
rect 5224 15036 5230 15048
rect 1673 15011 1731 15017
rect 1673 15008 1685 15011
rect 1268 14980 1685 15008
rect 1268 14968 1274 14980
rect 1673 14977 1685 14980
rect 1719 14977 1731 15011
rect 1673 14971 1731 14977
rect 2225 15011 2283 15017
rect 2225 14977 2237 15011
rect 2271 14977 2283 15011
rect 2225 14971 2283 14977
rect 2777 15011 2835 15017
rect 2777 14977 2789 15011
rect 2823 14977 2835 15011
rect 2777 14971 2835 14977
rect 1486 14804 1492 14816
rect 1447 14776 1492 14804
rect 1486 14764 1492 14776
rect 1544 14764 1550 14816
rect 2240 14804 2268 14971
rect 2866 14968 2872 15020
rect 2924 15008 2930 15020
rect 3033 15011 3091 15017
rect 3033 15008 3045 15011
rect 2924 14980 3045 15008
rect 2924 14968 2930 14980
rect 3033 14977 3045 14980
rect 3079 14977 3091 15011
rect 3033 14971 3091 14977
rect 5442 14968 5448 15020
rect 5500 15008 5506 15020
rect 6012 15017 6040 15048
rect 7116 15020 7144 15048
rect 7368 15045 7380 15079
rect 7414 15076 7426 15079
rect 7650 15076 7656 15088
rect 7414 15048 7656 15076
rect 7414 15045 7426 15048
rect 7368 15039 7426 15045
rect 7650 15036 7656 15048
rect 7708 15036 7714 15088
rect 9125 15079 9183 15085
rect 9125 15045 9137 15079
rect 9171 15076 9183 15079
rect 9674 15076 9680 15088
rect 9171 15048 9680 15076
rect 9171 15045 9183 15048
rect 9125 15039 9183 15045
rect 9674 15036 9680 15048
rect 9732 15036 9738 15088
rect 10042 15076 10048 15088
rect 10003 15048 10048 15076
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 10781 15079 10839 15085
rect 10781 15045 10793 15079
rect 10827 15076 10839 15079
rect 11238 15076 11244 15088
rect 10827 15048 11244 15076
rect 10827 15045 10839 15048
rect 10781 15039 10839 15045
rect 11238 15036 11244 15048
rect 11296 15036 11302 15088
rect 11698 15036 11704 15088
rect 11756 15076 11762 15088
rect 12406 15076 12434 15116
rect 12529 15113 12541 15147
rect 12575 15144 12587 15147
rect 12894 15144 12900 15156
rect 12575 15116 12900 15144
rect 12575 15113 12587 15116
rect 12529 15107 12587 15113
rect 12894 15104 12900 15116
rect 12952 15104 12958 15156
rect 13081 15147 13139 15153
rect 13081 15113 13093 15147
rect 13127 15144 13139 15147
rect 13262 15144 13268 15156
rect 13127 15116 13268 15144
rect 13127 15113 13139 15116
rect 13081 15107 13139 15113
rect 13262 15104 13268 15116
rect 13320 15104 13326 15156
rect 13449 15147 13507 15153
rect 13449 15113 13461 15147
rect 13495 15144 13507 15147
rect 13538 15144 13544 15156
rect 13495 15116 13544 15144
rect 13495 15113 13507 15116
rect 13449 15107 13507 15113
rect 13538 15104 13544 15116
rect 13596 15144 13602 15156
rect 15102 15144 15108 15156
rect 13596 15116 15108 15144
rect 13596 15104 13602 15116
rect 15102 15104 15108 15116
rect 15160 15104 15166 15156
rect 15470 15144 15476 15156
rect 15431 15116 15476 15144
rect 15470 15104 15476 15116
rect 15528 15104 15534 15156
rect 16669 15147 16727 15153
rect 16669 15113 16681 15147
rect 16715 15144 16727 15147
rect 16942 15144 16948 15156
rect 16715 15116 16948 15144
rect 16715 15113 16727 15116
rect 16669 15107 16727 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17681 15147 17739 15153
rect 17681 15144 17693 15147
rect 17052 15116 17693 15144
rect 11756 15048 12020 15076
rect 12406 15048 12940 15076
rect 11756 15036 11762 15048
rect 5730 15011 5788 15017
rect 5730 15008 5742 15011
rect 5500 14980 5742 15008
rect 5500 14968 5506 14980
rect 5730 14977 5742 14980
rect 5776 14977 5788 15011
rect 5730 14971 5788 14977
rect 5997 15011 6055 15017
rect 5997 14977 6009 15011
rect 6043 14977 6055 15011
rect 5997 14971 6055 14977
rect 6549 15011 6607 15017
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 7098 15008 7104 15020
rect 7011 14980 7104 15008
rect 6549 14971 6607 14977
rect 6564 14940 6592 14971
rect 7098 14968 7104 14980
rect 7156 14968 7162 15020
rect 11992 15008 12020 15048
rect 12713 15011 12771 15017
rect 12713 15008 12725 15011
rect 7217 14980 9168 15008
rect 7217 14940 7245 14980
rect 9030 14940 9036 14952
rect 6564 14912 7245 14940
rect 8991 14912 9036 14940
rect 9030 14900 9036 14912
rect 9088 14900 9094 14952
rect 9140 14940 9168 14980
rect 10428 14980 11836 15008
rect 11992 14980 12725 15008
rect 10428 14940 10456 14980
rect 10594 14940 10600 14952
rect 9140 14912 10456 14940
rect 10555 14912 10600 14940
rect 10594 14900 10600 14912
rect 10652 14900 10658 14952
rect 11701 14943 11759 14949
rect 11701 14909 11713 14943
rect 11747 14909 11759 14943
rect 11808 14940 11836 14980
rect 12713 14977 12725 14980
rect 12759 14977 12771 15011
rect 12912 15008 12940 15048
rect 12986 15036 12992 15088
rect 13044 15076 13050 15088
rect 14366 15085 14372 15088
rect 14360 15076 14372 15085
rect 13044 15048 14136 15076
rect 14327 15048 14372 15076
rect 13044 15036 13050 15048
rect 13354 15008 13360 15020
rect 12912 14980 13360 15008
rect 12713 14971 12771 14977
rect 13354 14968 13360 14980
rect 13412 14968 13418 15020
rect 13541 15011 13599 15017
rect 13541 14977 13553 15011
rect 13587 15008 13599 15011
rect 13630 15008 13636 15020
rect 13587 14980 13636 15008
rect 13587 14977 13599 14980
rect 13541 14971 13599 14977
rect 13630 14968 13636 14980
rect 13688 14968 13694 15020
rect 14108 15017 14136 15048
rect 14360 15039 14372 15048
rect 14366 15036 14372 15039
rect 14424 15036 14430 15088
rect 17052 15076 17080 15116
rect 17681 15113 17693 15116
rect 17727 15144 17739 15147
rect 19426 15144 19432 15156
rect 17727 15116 19334 15144
rect 19387 15116 19432 15144
rect 17727 15113 17739 15116
rect 17681 15107 17739 15113
rect 16868 15048 17080 15076
rect 14093 15011 14151 15017
rect 14093 14977 14105 15011
rect 14139 14977 14151 15011
rect 14734 15008 14740 15020
rect 14093 14971 14151 14977
rect 14200 14980 14740 15008
rect 12342 14940 12348 14952
rect 11808 14912 12348 14940
rect 11701 14903 11759 14909
rect 11716 14872 11744 14903
rect 12342 14900 12348 14912
rect 12400 14900 12406 14952
rect 13722 14940 13728 14952
rect 13683 14912 13728 14940
rect 13722 14900 13728 14912
rect 13780 14940 13786 14952
rect 14200 14940 14228 14980
rect 14734 14968 14740 14980
rect 14792 14968 14798 15020
rect 13780 14912 14228 14940
rect 16209 14943 16267 14949
rect 13780 14900 13786 14912
rect 16209 14909 16221 14943
rect 16255 14909 16267 14943
rect 16209 14903 16267 14909
rect 12894 14872 12900 14884
rect 11716 14844 12900 14872
rect 12894 14832 12900 14844
rect 12952 14832 12958 14884
rect 16224 14872 16252 14903
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 16868 14940 16896 15048
rect 17126 15036 17132 15088
rect 17184 15076 17190 15088
rect 19306 15076 19334 15116
rect 19426 15104 19432 15116
rect 19484 15104 19490 15156
rect 21085 15147 21143 15153
rect 21085 15113 21097 15147
rect 21131 15144 21143 15147
rect 21266 15144 21272 15156
rect 21131 15116 21272 15144
rect 21131 15113 21143 15116
rect 21085 15107 21143 15113
rect 21266 15104 21272 15116
rect 21324 15104 21330 15156
rect 20622 15076 20628 15088
rect 17184 15048 18092 15076
rect 19306 15048 20628 15076
rect 17184 15036 17190 15048
rect 17034 15008 17040 15020
rect 16995 14980 17040 15008
rect 17034 14968 17040 14980
rect 17092 15008 17098 15020
rect 17092 14980 17448 15008
rect 17092 14968 17098 14980
rect 17129 14943 17187 14949
rect 17129 14940 17141 14943
rect 16448 14912 17141 14940
rect 16448 14900 16454 14912
rect 17129 14909 17141 14912
rect 17175 14909 17187 14943
rect 17129 14903 17187 14909
rect 17218 14900 17224 14952
rect 17276 14940 17282 14952
rect 17420 14940 17448 14980
rect 17494 14968 17500 15020
rect 17552 15008 17558 15020
rect 17954 15008 17960 15020
rect 17552 14980 17960 15008
rect 17552 14968 17558 14980
rect 17954 14968 17960 14980
rect 18012 14968 18018 15020
rect 18064 15017 18092 15048
rect 20622 15036 20628 15048
rect 20680 15036 20686 15088
rect 18049 15011 18107 15017
rect 18049 14977 18061 15011
rect 18095 14977 18107 15011
rect 18049 14971 18107 14977
rect 18316 15011 18374 15017
rect 18316 14977 18328 15011
rect 18362 15008 18374 15011
rect 18362 14980 19380 15008
rect 18362 14977 18374 14980
rect 18316 14971 18374 14977
rect 19352 14940 19380 14980
rect 19426 14968 19432 15020
rect 19484 15008 19490 15020
rect 19705 15011 19763 15017
rect 19705 15008 19717 15011
rect 19484 14980 19717 15008
rect 19484 14968 19490 14980
rect 19705 14977 19717 14980
rect 19751 14977 19763 15011
rect 19705 14971 19763 14977
rect 20530 14940 20536 14952
rect 17276 14912 17321 14940
rect 17420 14912 17908 14940
rect 19352 14912 20536 14940
rect 17276 14900 17282 14912
rect 17770 14872 17776 14884
rect 16224 14844 17776 14872
rect 17770 14832 17776 14844
rect 17828 14832 17834 14884
rect 4154 14804 4160 14816
rect 2240 14776 4160 14804
rect 4154 14764 4160 14776
rect 4212 14764 4218 14816
rect 4338 14764 4344 14816
rect 4396 14804 4402 14816
rect 7374 14804 7380 14816
rect 4396 14776 7380 14804
rect 4396 14764 4402 14776
rect 7374 14764 7380 14776
rect 7432 14764 7438 14816
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 17494 14804 17500 14816
rect 8444 14776 17500 14804
rect 8444 14764 8450 14776
rect 17494 14764 17500 14776
rect 17552 14764 17558 14816
rect 17880 14804 17908 14912
rect 20530 14900 20536 14912
rect 20588 14900 20594 14952
rect 20717 14875 20775 14881
rect 20717 14872 20729 14875
rect 18984 14844 20729 14872
rect 18984 14804 19012 14844
rect 20717 14841 20729 14844
rect 20763 14841 20775 14875
rect 20717 14835 20775 14841
rect 17880 14776 19012 14804
rect 19058 14764 19064 14816
rect 19116 14804 19122 14816
rect 20349 14807 20407 14813
rect 20349 14804 20361 14807
rect 19116 14776 20361 14804
rect 19116 14764 19122 14776
rect 20349 14773 20361 14776
rect 20395 14773 20407 14807
rect 20349 14767 20407 14773
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 2041 14603 2099 14609
rect 2041 14569 2053 14603
rect 2087 14600 2099 14603
rect 2314 14600 2320 14612
rect 2087 14572 2320 14600
rect 2087 14569 2099 14572
rect 2041 14563 2099 14569
rect 2314 14560 2320 14572
rect 2372 14560 2378 14612
rect 5442 14600 5448 14612
rect 5403 14572 5448 14600
rect 5442 14560 5448 14572
rect 5500 14560 5506 14612
rect 5902 14560 5908 14612
rect 5960 14600 5966 14612
rect 6365 14603 6423 14609
rect 6365 14600 6377 14603
rect 5960 14572 6377 14600
rect 5960 14560 5966 14572
rect 6365 14569 6377 14572
rect 6411 14600 6423 14603
rect 6546 14600 6552 14612
rect 6411 14572 6552 14600
rect 6411 14569 6423 14572
rect 6365 14563 6423 14569
rect 6546 14560 6552 14572
rect 6604 14560 6610 14612
rect 8294 14560 8300 14612
rect 8352 14600 8358 14612
rect 8481 14603 8539 14609
rect 8481 14600 8493 14603
rect 8352 14572 8493 14600
rect 8352 14560 8358 14572
rect 8481 14569 8493 14572
rect 8527 14569 8539 14603
rect 8481 14563 8539 14569
rect 10137 14603 10195 14609
rect 10137 14569 10149 14603
rect 10183 14600 10195 14603
rect 10594 14600 10600 14612
rect 10183 14572 10600 14600
rect 10183 14569 10195 14572
rect 10137 14563 10195 14569
rect 2866 14492 2872 14544
rect 2924 14532 2930 14544
rect 2924 14504 4016 14532
rect 2924 14492 2930 14504
rect 3329 14467 3387 14473
rect 3329 14433 3341 14467
rect 3375 14464 3387 14467
rect 3786 14464 3792 14476
rect 3375 14436 3792 14464
rect 3375 14433 3387 14436
rect 3329 14427 3387 14433
rect 3786 14424 3792 14436
rect 3844 14424 3850 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 2225 14399 2283 14405
rect 2225 14365 2237 14399
rect 2271 14396 2283 14399
rect 2406 14396 2412 14408
rect 2271 14368 2412 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 1688 14328 1716 14359
rect 2406 14356 2412 14368
rect 2464 14356 2470 14408
rect 2746 14368 3924 14396
rect 2746 14328 2774 14368
rect 1688 14300 2774 14328
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 2685 14263 2743 14269
rect 2685 14260 2697 14263
rect 2372 14232 2697 14260
rect 2372 14220 2378 14232
rect 2685 14229 2697 14232
rect 2731 14229 2743 14263
rect 3050 14260 3056 14272
rect 3011 14232 3056 14260
rect 2685 14223 2743 14229
rect 3050 14220 3056 14232
rect 3108 14220 3114 14272
rect 3142 14220 3148 14272
rect 3200 14260 3206 14272
rect 3786 14260 3792 14272
rect 3200 14232 3245 14260
rect 3747 14232 3792 14260
rect 3200 14220 3206 14232
rect 3786 14220 3792 14232
rect 3844 14220 3850 14272
rect 3896 14260 3924 14368
rect 3988 14328 4016 14504
rect 5166 14464 5172 14476
rect 5127 14436 5172 14464
rect 5166 14424 5172 14436
rect 5224 14424 5230 14476
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 4902 14399 4960 14405
rect 4902 14396 4914 14399
rect 4672 14368 4914 14396
rect 4672 14356 4678 14368
rect 4902 14365 4914 14368
rect 4948 14365 4960 14399
rect 4902 14359 4960 14365
rect 5718 14356 5724 14408
rect 5776 14396 5782 14408
rect 5994 14396 6000 14408
rect 5776 14368 6000 14396
rect 5776 14356 5782 14368
rect 5994 14356 6000 14368
rect 6052 14396 6058 14408
rect 6089 14399 6147 14405
rect 6089 14396 6101 14399
rect 6052 14368 6101 14396
rect 6052 14356 6058 14368
rect 6089 14365 6101 14368
rect 6135 14365 6147 14399
rect 6089 14359 6147 14365
rect 7098 14356 7104 14408
rect 7156 14396 7162 14408
rect 7745 14399 7803 14405
rect 7745 14396 7757 14399
rect 7156 14368 7757 14396
rect 7156 14356 7162 14368
rect 7745 14365 7757 14368
rect 7791 14365 7803 14399
rect 7745 14359 7803 14365
rect 9861 14399 9919 14405
rect 9861 14365 9873 14399
rect 9907 14396 9919 14399
rect 10152 14396 10180 14563
rect 10594 14560 10600 14572
rect 10652 14600 10658 14612
rect 12066 14600 12072 14612
rect 10652 14572 12072 14600
rect 10652 14560 10658 14572
rect 12066 14560 12072 14572
rect 12124 14560 12130 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12434 14600 12440 14612
rect 12299 14572 12440 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12434 14560 12440 14572
rect 12492 14560 12498 14612
rect 13814 14560 13820 14612
rect 13872 14600 13878 14612
rect 14093 14603 14151 14609
rect 14093 14600 14105 14603
rect 13872 14572 14105 14600
rect 13872 14560 13878 14572
rect 14093 14569 14105 14572
rect 14139 14569 14151 14603
rect 14093 14563 14151 14569
rect 16022 14560 16028 14612
rect 16080 14600 16086 14612
rect 18141 14603 18199 14609
rect 16080 14572 16712 14600
rect 16080 14560 16086 14572
rect 16684 14532 16712 14572
rect 18141 14569 18153 14603
rect 18187 14600 18199 14603
rect 18874 14600 18880 14612
rect 18187 14572 18880 14600
rect 18187 14569 18199 14572
rect 18141 14563 18199 14569
rect 18874 14560 18880 14572
rect 18932 14560 18938 14612
rect 20993 14603 21051 14609
rect 20993 14569 21005 14603
rect 21039 14600 21051 14603
rect 21910 14600 21916 14612
rect 21039 14572 21916 14600
rect 21039 14569 21051 14572
rect 20993 14563 21051 14569
rect 21910 14560 21916 14572
rect 21968 14560 21974 14612
rect 20165 14535 20223 14541
rect 20165 14532 20177 14535
rect 16684 14504 20177 14532
rect 20165 14501 20177 14504
rect 20211 14501 20223 14535
rect 20165 14495 20223 14501
rect 14642 14464 14648 14476
rect 14603 14436 14648 14464
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 17494 14464 17500 14476
rect 17455 14436 17500 14464
rect 17494 14424 17500 14436
rect 17552 14464 17558 14476
rect 17552 14436 17908 14464
rect 17552 14424 17558 14436
rect 11517 14399 11575 14405
rect 11517 14396 11529 14399
rect 9907 14368 10180 14396
rect 11164 14368 11529 14396
rect 9907 14365 9919 14368
rect 9861 14359 9919 14365
rect 11164 14340 11192 14368
rect 11517 14365 11529 14368
rect 11563 14396 11575 14399
rect 12986 14396 12992 14408
rect 11563 14368 12992 14396
rect 11563 14365 11575 14368
rect 11517 14359 11575 14365
rect 12986 14356 12992 14368
rect 13044 14356 13050 14408
rect 13541 14399 13599 14405
rect 13541 14365 13553 14399
rect 13587 14396 13599 14399
rect 15194 14396 15200 14408
rect 13587 14368 15200 14396
rect 13587 14365 13599 14368
rect 13541 14359 13599 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 15749 14399 15807 14405
rect 15749 14365 15761 14399
rect 15795 14396 15807 14399
rect 17126 14396 17132 14408
rect 15795 14368 17132 14396
rect 15795 14365 15807 14368
rect 15749 14359 15807 14365
rect 17126 14356 17132 14368
rect 17184 14356 17190 14408
rect 17770 14396 17776 14408
rect 17731 14368 17776 14396
rect 17770 14356 17776 14368
rect 17828 14356 17834 14408
rect 17880 14396 17908 14436
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 18417 14467 18475 14473
rect 18417 14464 18429 14467
rect 18104 14436 18429 14464
rect 18104 14424 18110 14436
rect 18417 14433 18429 14436
rect 18463 14433 18475 14467
rect 18417 14427 18475 14433
rect 18690 14424 18696 14476
rect 18748 14464 18754 14476
rect 21269 14467 21327 14473
rect 21269 14464 21281 14467
rect 18748 14436 21281 14464
rect 18748 14424 18754 14436
rect 21269 14433 21281 14436
rect 21315 14433 21327 14467
rect 21269 14427 21327 14433
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 17880 14368 19257 14396
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 20530 14396 20536 14408
rect 20491 14368 20536 14396
rect 19245 14359 19303 14365
rect 20530 14356 20536 14368
rect 20588 14356 20594 14408
rect 6546 14328 6552 14340
rect 3988 14300 6552 14328
rect 6546 14288 6552 14300
rect 6604 14288 6610 14340
rect 7466 14288 7472 14340
rect 7524 14337 7530 14340
rect 7524 14328 7536 14337
rect 9217 14331 9275 14337
rect 7524 14300 7569 14328
rect 7524 14291 7536 14300
rect 9217 14297 9229 14331
rect 9263 14328 9275 14331
rect 9263 14300 11100 14328
rect 9263 14297 9275 14300
rect 9217 14291 9275 14297
rect 7524 14288 7530 14291
rect 5442 14260 5448 14272
rect 3896 14232 5448 14260
rect 5442 14220 5448 14232
rect 5500 14220 5506 14272
rect 8018 14260 8024 14272
rect 7979 14232 8024 14260
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 11072 14260 11100 14300
rect 11146 14288 11152 14340
rect 11204 14288 11210 14340
rect 11238 14288 11244 14340
rect 11296 14337 11302 14340
rect 11296 14328 11308 14337
rect 14461 14331 14519 14337
rect 11296 14300 11341 14328
rect 11296 14291 11308 14300
rect 14461 14297 14473 14331
rect 14507 14328 14519 14331
rect 15105 14331 15163 14337
rect 15105 14328 15117 14331
rect 14507 14300 15117 14328
rect 14507 14297 14519 14300
rect 14461 14291 14519 14297
rect 15105 14297 15117 14300
rect 15151 14297 15163 14331
rect 15105 14291 15163 14297
rect 16016 14331 16074 14337
rect 16016 14297 16028 14331
rect 16062 14328 16074 14331
rect 19889 14331 19947 14337
rect 19889 14328 19901 14331
rect 16062 14300 19901 14328
rect 16062 14297 16074 14300
rect 16016 14291 16074 14297
rect 19889 14297 19901 14300
rect 19935 14297 19947 14331
rect 19889 14291 19947 14297
rect 11296 14288 11302 14291
rect 11790 14260 11796 14272
rect 11072 14232 11796 14260
rect 11790 14220 11796 14232
rect 11848 14220 11854 14272
rect 14550 14260 14556 14272
rect 14511 14232 14556 14260
rect 14550 14220 14556 14232
rect 14608 14220 14614 14272
rect 17126 14260 17132 14272
rect 17087 14232 17132 14260
rect 17126 14220 17132 14232
rect 17184 14220 17190 14272
rect 17402 14220 17408 14272
rect 17460 14260 17466 14272
rect 17681 14263 17739 14269
rect 17681 14260 17693 14263
rect 17460 14232 17693 14260
rect 17460 14220 17466 14232
rect 17681 14229 17693 14232
rect 17727 14229 17739 14263
rect 17681 14223 17739 14229
rect 1104 14170 21896 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21896 14170
rect 1104 14096 21896 14118
rect 2317 14059 2375 14065
rect 2317 14025 2329 14059
rect 2363 14056 2375 14059
rect 3050 14056 3056 14068
rect 2363 14028 3056 14056
rect 2363 14025 2375 14028
rect 2317 14019 2375 14025
rect 3050 14016 3056 14028
rect 3108 14016 3114 14068
rect 3237 14059 3295 14065
rect 3237 14025 3249 14059
rect 3283 14056 3295 14059
rect 3973 14059 4031 14065
rect 3973 14056 3985 14059
rect 3283 14028 3985 14056
rect 3283 14025 3295 14028
rect 3237 14019 3295 14025
rect 3973 14025 3985 14028
rect 4019 14025 4031 14059
rect 5534 14056 5540 14068
rect 3973 14019 4031 14025
rect 4540 14028 5540 14056
rect 4540 13988 4568 14028
rect 5534 14016 5540 14028
rect 5592 14016 5598 14068
rect 5994 14056 6000 14068
rect 5955 14028 6000 14056
rect 5994 14016 6000 14028
rect 6052 14016 6058 14068
rect 6546 14016 6552 14068
rect 6604 14056 6610 14068
rect 6917 14059 6975 14065
rect 6917 14056 6929 14059
rect 6604 14028 6929 14056
rect 6604 14016 6610 14028
rect 6917 14025 6929 14028
rect 6963 14025 6975 14059
rect 6917 14019 6975 14025
rect 7377 14059 7435 14065
rect 7377 14025 7389 14059
rect 7423 14056 7435 14059
rect 7929 14059 7987 14065
rect 7929 14056 7941 14059
rect 7423 14028 7941 14056
rect 7423 14025 7435 14028
rect 7377 14019 7435 14025
rect 7929 14025 7941 14028
rect 7975 14025 7987 14059
rect 8386 14056 8392 14068
rect 8347 14028 8392 14056
rect 7929 14019 7987 14025
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 8941 14059 8999 14065
rect 8941 14025 8953 14059
rect 8987 14056 8999 14059
rect 9122 14056 9128 14068
rect 8987 14028 9128 14056
rect 8987 14025 8999 14028
rect 8941 14019 8999 14025
rect 9122 14016 9128 14028
rect 9180 14016 9186 14068
rect 10502 14016 10508 14068
rect 10560 14056 10566 14068
rect 10597 14059 10655 14065
rect 10597 14056 10609 14059
rect 10560 14028 10609 14056
rect 10560 14016 10566 14028
rect 10597 14025 10609 14028
rect 10643 14025 10655 14059
rect 10597 14019 10655 14025
rect 11517 14059 11575 14065
rect 11517 14025 11529 14059
rect 11563 14056 11575 14059
rect 11882 14056 11888 14068
rect 11563 14028 11888 14056
rect 11563 14025 11575 14028
rect 11517 14019 11575 14025
rect 11882 14016 11888 14028
rect 11940 14016 11946 14068
rect 11974 14016 11980 14068
rect 12032 14056 12038 14068
rect 12529 14059 12587 14065
rect 12529 14056 12541 14059
rect 12032 14028 12541 14056
rect 12032 14016 12038 14028
rect 12529 14025 12541 14028
rect 12575 14025 12587 14059
rect 12529 14019 12587 14025
rect 13078 14016 13084 14068
rect 13136 14056 13142 14068
rect 13630 14056 13636 14068
rect 13136 14028 13636 14056
rect 13136 14016 13142 14028
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 14369 14059 14427 14065
rect 14369 14025 14381 14059
rect 14415 14056 14427 14059
rect 14642 14056 14648 14068
rect 14415 14028 14648 14056
rect 14415 14025 14427 14028
rect 14369 14019 14427 14025
rect 14642 14016 14648 14028
rect 14700 14016 14706 14068
rect 16301 14059 16359 14065
rect 16301 14025 16313 14059
rect 16347 14056 16359 14059
rect 17402 14056 17408 14068
rect 16347 14028 17264 14056
rect 17363 14028 17408 14056
rect 16347 14025 16359 14028
rect 16301 14019 16359 14025
rect 5718 13988 5724 14000
rect 2976 13960 4568 13988
rect 4632 13960 5724 13988
rect 1397 13923 1455 13929
rect 1397 13889 1409 13923
rect 1443 13920 1455 13923
rect 1762 13920 1768 13932
rect 1443 13892 1768 13920
rect 1443 13889 1455 13892
rect 1397 13883 1455 13889
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 2774 13920 2780 13932
rect 2639 13892 2780 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 2774 13880 2780 13892
rect 2832 13880 2838 13932
rect 2976 13852 3004 13960
rect 3050 13880 3056 13932
rect 3108 13920 3114 13932
rect 3881 13923 3939 13929
rect 3108 13892 3648 13920
rect 3108 13880 3114 13892
rect 2792 13824 3004 13852
rect 1578 13784 1584 13796
rect 1539 13756 1584 13784
rect 1578 13744 1584 13756
rect 1636 13744 1642 13796
rect 2792 13793 2820 13824
rect 3142 13812 3148 13864
rect 3200 13852 3206 13864
rect 3620 13852 3648 13892
rect 3881 13889 3893 13923
rect 3927 13920 3939 13923
rect 4338 13920 4344 13932
rect 3927 13892 4344 13920
rect 3927 13889 3939 13892
rect 3881 13883 3939 13889
rect 4338 13880 4344 13892
rect 4396 13880 4402 13932
rect 4632 13929 4660 13960
rect 5718 13948 5724 13960
rect 5776 13948 5782 14000
rect 7285 13991 7343 13997
rect 7285 13957 7297 13991
rect 7331 13988 7343 13991
rect 8478 13988 8484 14000
rect 7331 13960 8484 13988
rect 7331 13957 7343 13960
rect 7285 13951 7343 13957
rect 8478 13948 8484 13960
rect 8536 13948 8542 14000
rect 10226 13948 10232 14000
rect 10284 13988 10290 14000
rect 11057 13991 11115 13997
rect 11057 13988 11069 13991
rect 10284 13960 11069 13988
rect 10284 13948 10290 13960
rect 11057 13957 11069 13960
rect 11103 13988 11115 13991
rect 11103 13960 12756 13988
rect 11103 13957 11115 13960
rect 11057 13951 11115 13957
rect 4617 13923 4675 13929
rect 4617 13889 4629 13923
rect 4663 13889 4675 13923
rect 4617 13883 4675 13889
rect 4706 13880 4712 13932
rect 4764 13920 4770 13932
rect 4873 13923 4931 13929
rect 4873 13920 4885 13923
rect 4764 13892 4885 13920
rect 4764 13880 4770 13892
rect 4873 13889 4885 13892
rect 4919 13889 4931 13923
rect 4873 13883 4931 13889
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 6365 13923 6423 13929
rect 6365 13920 6377 13923
rect 5224 13892 6377 13920
rect 5224 13880 5230 13892
rect 6365 13889 6377 13892
rect 6411 13889 6423 13923
rect 6365 13883 6423 13889
rect 7006 13880 7012 13932
rect 7064 13920 7070 13932
rect 8297 13923 8355 13929
rect 8297 13920 8309 13923
rect 7064 13892 8309 13920
rect 7064 13880 7070 13892
rect 8297 13889 8309 13892
rect 8343 13889 8355 13923
rect 10042 13920 10048 13932
rect 10100 13929 10106 13932
rect 10012 13892 10048 13920
rect 8297 13883 8355 13889
rect 10042 13880 10048 13892
rect 10100 13883 10112 13929
rect 10321 13923 10379 13929
rect 10321 13889 10333 13923
rect 10367 13920 10379 13923
rect 11146 13920 11152 13932
rect 10367 13892 11152 13920
rect 10367 13889 10379 13892
rect 10321 13883 10379 13889
rect 10100 13880 10106 13883
rect 11146 13880 11152 13892
rect 11204 13880 11210 13932
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 12434 13920 12440 13932
rect 11931 13892 12440 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 12728 13929 12756 13960
rect 12986 13948 12992 14000
rect 13044 13988 13050 14000
rect 16945 13991 17003 13997
rect 13044 13960 14964 13988
rect 13044 13948 13050 13960
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13889 12771 13923
rect 12713 13883 12771 13889
rect 13256 13923 13314 13929
rect 13256 13889 13268 13923
rect 13302 13920 13314 13923
rect 13814 13920 13820 13932
rect 13302 13892 13820 13920
rect 13302 13889 13314 13892
rect 13256 13883 13314 13889
rect 13814 13880 13820 13892
rect 13872 13880 13878 13932
rect 14936 13929 14964 13960
rect 16945 13957 16957 13991
rect 16991 13957 17003 13991
rect 16945 13951 17003 13957
rect 17037 13991 17095 13997
rect 17037 13957 17049 13991
rect 17083 13957 17095 13991
rect 17236 13988 17264 14028
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 17586 14016 17592 14068
rect 17644 14056 17650 14068
rect 19978 14056 19984 14068
rect 17644 14028 19472 14056
rect 19939 14028 19984 14056
rect 17644 14016 17650 14028
rect 17494 13988 17500 14000
rect 17236 13960 17500 13988
rect 17037 13951 17095 13957
rect 14921 13923 14979 13929
rect 14921 13889 14933 13923
rect 14967 13889 14979 13923
rect 14921 13883 14979 13889
rect 15188 13923 15246 13929
rect 15188 13889 15200 13923
rect 15234 13920 15246 13923
rect 16390 13920 16396 13932
rect 15234 13892 16396 13920
rect 15234 13889 15246 13892
rect 15188 13883 15246 13889
rect 16390 13880 16396 13892
rect 16448 13880 16454 13932
rect 16960 13864 16988 13951
rect 17052 13864 17080 13951
rect 17494 13948 17500 13960
rect 17552 13948 17558 14000
rect 18816 13991 18874 13997
rect 18816 13957 18828 13991
rect 18862 13988 18874 13991
rect 19058 13988 19064 14000
rect 18862 13960 19064 13988
rect 18862 13957 18874 13960
rect 18816 13951 18874 13957
rect 19058 13948 19064 13960
rect 19116 13948 19122 14000
rect 17126 13880 17132 13932
rect 17184 13920 17190 13932
rect 19337 13923 19395 13929
rect 19337 13920 19349 13923
rect 17184 13892 19349 13920
rect 17184 13880 17190 13892
rect 19337 13889 19349 13892
rect 19383 13889 19395 13923
rect 19444 13920 19472 14028
rect 19978 14016 19984 14028
rect 20036 14016 20042 14068
rect 20717 14059 20775 14065
rect 20717 14025 20729 14059
rect 20763 14056 20775 14059
rect 21174 14056 21180 14068
rect 20763 14028 21180 14056
rect 20763 14025 20775 14028
rect 20717 14019 20775 14025
rect 21174 14016 21180 14028
rect 21232 14016 21238 14068
rect 21358 14056 21364 14068
rect 21319 14028 21364 14056
rect 21358 14016 21364 14028
rect 21416 14016 21422 14068
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19444 13892 20269 13920
rect 19337 13883 19395 13889
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 3200 13824 3556 13852
rect 3620 13824 3924 13852
rect 3200 13812 3206 13824
rect 3528 13793 3556 13824
rect 2777 13787 2835 13793
rect 2777 13753 2789 13787
rect 2823 13753 2835 13787
rect 2777 13747 2835 13753
rect 3513 13787 3571 13793
rect 3513 13753 3525 13787
rect 3559 13753 3571 13787
rect 3896 13784 3924 13824
rect 3970 13812 3976 13864
rect 4028 13852 4034 13864
rect 4157 13855 4215 13861
rect 4157 13852 4169 13855
rect 4028 13824 4169 13852
rect 4028 13812 4034 13824
rect 4157 13821 4169 13824
rect 4203 13821 4215 13855
rect 4157 13815 4215 13821
rect 4246 13812 4252 13864
rect 4304 13812 4310 13864
rect 7558 13852 7564 13864
rect 7519 13824 7564 13852
rect 7558 13812 7564 13824
rect 7616 13812 7622 13864
rect 8573 13855 8631 13861
rect 8573 13821 8585 13855
rect 8619 13821 8631 13855
rect 8573 13815 8631 13821
rect 4264 13784 4292 13812
rect 3896 13756 4292 13784
rect 8588 13784 8616 13815
rect 11054 13812 11060 13864
rect 11112 13852 11118 13864
rect 11977 13855 12035 13861
rect 11977 13852 11989 13855
rect 11112 13824 11989 13852
rect 11112 13812 11118 13824
rect 11977 13821 11989 13824
rect 12023 13821 12035 13855
rect 11977 13815 12035 13821
rect 12066 13812 12072 13864
rect 12124 13852 12130 13864
rect 12124 13824 12169 13852
rect 12124 13812 12130 13824
rect 12342 13812 12348 13864
rect 12400 13852 12406 13864
rect 12989 13855 13047 13861
rect 12989 13852 13001 13855
rect 12400 13824 13001 13852
rect 12400 13812 12406 13824
rect 12989 13821 13001 13824
rect 13035 13821 13047 13855
rect 16853 13855 16911 13861
rect 16853 13852 16865 13855
rect 12989 13815 13047 13821
rect 16776 13824 16865 13852
rect 16776 13796 16804 13824
rect 16853 13821 16865 13824
rect 16899 13821 16911 13855
rect 16853 13815 16911 13821
rect 16942 13812 16948 13864
rect 17000 13812 17006 13864
rect 17034 13812 17040 13864
rect 17092 13812 17098 13864
rect 19058 13852 19064 13864
rect 19019 13824 19064 13852
rect 19058 13812 19064 13824
rect 19116 13812 19122 13864
rect 8662 13784 8668 13796
rect 8588 13756 8668 13784
rect 3513 13747 3571 13753
rect 8662 13744 8668 13756
rect 8720 13744 8726 13796
rect 16758 13744 16764 13796
rect 16816 13744 16822 13796
rect 3878 13676 3884 13728
rect 3936 13716 3942 13728
rect 6822 13716 6828 13728
rect 3936 13688 6828 13716
rect 3936 13676 3942 13688
rect 6822 13676 6828 13688
rect 6880 13676 6886 13728
rect 17586 13676 17592 13728
rect 17644 13716 17650 13728
rect 17681 13719 17739 13725
rect 17681 13716 17693 13719
rect 17644 13688 17693 13716
rect 17644 13676 17650 13688
rect 17681 13685 17693 13688
rect 17727 13685 17739 13719
rect 17681 13679 17739 13685
rect 1104 13626 21896 13648
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13512 2559 13515
rect 2958 13512 2964 13524
rect 2547 13484 2964 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 2958 13472 2964 13484
rect 3016 13472 3022 13524
rect 4706 13512 4712 13524
rect 3344 13484 4712 13512
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 3344 13444 3372 13484
rect 4706 13472 4712 13484
rect 4764 13472 4770 13524
rect 6730 13512 6736 13524
rect 4816 13484 6736 13512
rect 4338 13444 4344 13456
rect 2823 13416 3372 13444
rect 3436 13416 4344 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 1578 13308 1584 13320
rect 1539 13280 1584 13308
rect 1578 13268 1584 13280
rect 1636 13268 1642 13320
rect 1854 13308 1860 13320
rect 1815 13280 1860 13308
rect 1854 13268 1860 13280
rect 1912 13268 1918 13320
rect 2317 13311 2375 13317
rect 2317 13277 2329 13311
rect 2363 13308 2375 13311
rect 2590 13308 2596 13320
rect 2363 13280 2596 13308
rect 2363 13277 2375 13280
rect 2317 13271 2375 13277
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 3436 13317 3464 13416
rect 4338 13404 4344 13416
rect 4396 13404 4402 13456
rect 4816 13444 4844 13484
rect 6730 13472 6736 13484
rect 6788 13472 6794 13524
rect 7929 13515 7987 13521
rect 7929 13481 7941 13515
rect 7975 13512 7987 13515
rect 8570 13512 8576 13524
rect 7975 13484 8576 13512
rect 7975 13481 7987 13484
rect 7929 13475 7987 13481
rect 8570 13472 8576 13484
rect 8628 13472 8634 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10137 13515 10195 13521
rect 10137 13512 10149 13515
rect 10100 13484 10149 13512
rect 10100 13472 10106 13484
rect 10137 13481 10149 13484
rect 10183 13481 10195 13515
rect 10137 13475 10195 13481
rect 10873 13515 10931 13521
rect 10873 13481 10885 13515
rect 10919 13512 10931 13515
rect 11146 13512 11152 13524
rect 10919 13484 11152 13512
rect 10919 13481 10931 13484
rect 10873 13475 10931 13481
rect 11146 13472 11152 13484
rect 11204 13472 11210 13524
rect 13725 13515 13783 13521
rect 13725 13481 13737 13515
rect 13771 13512 13783 13515
rect 14550 13512 14556 13524
rect 13771 13484 14556 13512
rect 13771 13481 13783 13484
rect 13725 13475 13783 13481
rect 14550 13472 14556 13484
rect 14608 13472 14614 13524
rect 16390 13512 16396 13524
rect 16351 13484 16396 13512
rect 16390 13472 16396 13484
rect 16448 13472 16454 13524
rect 18141 13515 18199 13521
rect 18141 13481 18153 13515
rect 18187 13512 18199 13515
rect 20806 13512 20812 13524
rect 18187 13484 20812 13512
rect 18187 13481 18199 13484
rect 18141 13475 18199 13481
rect 20806 13472 20812 13484
rect 20864 13472 20870 13524
rect 21361 13515 21419 13521
rect 21361 13481 21373 13515
rect 21407 13512 21419 13515
rect 21450 13512 21456 13524
rect 21407 13484 21456 13512
rect 21407 13481 21419 13484
rect 21361 13475 21419 13481
rect 21450 13472 21456 13484
rect 21508 13472 21514 13524
rect 4448 13416 4844 13444
rect 3510 13336 3516 13388
rect 3568 13376 3574 13388
rect 4448 13376 4476 13416
rect 7558 13404 7564 13456
rect 7616 13444 7622 13456
rect 16117 13447 16175 13453
rect 7616 13416 9536 13444
rect 7616 13404 7622 13416
rect 5718 13376 5724 13388
rect 3568 13348 4476 13376
rect 5679 13348 5724 13376
rect 3568 13336 3574 13348
rect 5718 13336 5724 13348
rect 5776 13336 5782 13388
rect 6546 13376 6552 13388
rect 6507 13348 6552 13376
rect 6546 13336 6552 13348
rect 6604 13336 6610 13388
rect 8662 13376 8668 13388
rect 7668 13348 8668 13376
rect 3421 13311 3479 13317
rect 3421 13277 3433 13311
rect 3467 13277 3479 13311
rect 3421 13271 3479 13277
rect 3881 13311 3939 13317
rect 3881 13277 3893 13311
rect 3927 13308 3939 13311
rect 3970 13308 3976 13320
rect 3927 13280 3976 13308
rect 3927 13277 3939 13280
rect 3881 13271 3939 13277
rect 3970 13268 3976 13280
rect 4028 13268 4034 13320
rect 5626 13308 5632 13320
rect 4080 13280 5632 13308
rect 1397 13175 1455 13181
rect 1397 13141 1409 13175
rect 1443 13172 1455 13175
rect 1486 13172 1492 13184
rect 1443 13144 1492 13172
rect 1443 13141 1455 13144
rect 1397 13135 1455 13141
rect 1486 13132 1492 13144
rect 1544 13132 1550 13184
rect 2041 13175 2099 13181
rect 2041 13141 2053 13175
rect 2087 13172 2099 13175
rect 2406 13172 2412 13184
rect 2087 13144 2412 13172
rect 2087 13141 2099 13144
rect 2041 13135 2099 13141
rect 2406 13132 2412 13144
rect 2464 13132 2470 13184
rect 4080 13181 4108 13280
rect 5626 13268 5632 13280
rect 5684 13268 5690 13320
rect 6365 13311 6423 13317
rect 6365 13277 6377 13311
rect 6411 13308 6423 13311
rect 7006 13308 7012 13320
rect 6411 13280 7012 13308
rect 6411 13277 6423 13280
rect 6365 13271 6423 13277
rect 7006 13268 7012 13280
rect 7064 13308 7070 13320
rect 7466 13308 7472 13320
rect 7064 13280 7472 13308
rect 7064 13268 7070 13280
rect 7466 13268 7472 13280
rect 7524 13268 7530 13320
rect 7668 13317 7696 13348
rect 8662 13336 8668 13348
rect 8720 13336 8726 13388
rect 7653 13311 7711 13317
rect 7653 13277 7665 13311
rect 7699 13277 7711 13311
rect 7653 13271 7711 13277
rect 8573 13311 8631 13317
rect 8573 13277 8585 13311
rect 8619 13308 8631 13311
rect 9122 13308 9128 13320
rect 8619 13280 9128 13308
rect 8619 13277 8631 13280
rect 8573 13271 8631 13277
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 9508 13317 9536 13416
rect 16117 13413 16129 13447
rect 16163 13413 16175 13447
rect 16117 13407 16175 13413
rect 20257 13447 20315 13453
rect 20257 13413 20269 13447
rect 20303 13444 20315 13447
rect 20346 13444 20352 13456
rect 20303 13416 20352 13444
rect 20303 13413 20315 13416
rect 20257 13407 20315 13413
rect 12434 13336 12440 13388
rect 12492 13376 12498 13388
rect 13173 13379 13231 13385
rect 12492 13348 12537 13376
rect 12492 13336 12498 13348
rect 13173 13345 13185 13379
rect 13219 13376 13231 13379
rect 13814 13376 13820 13388
rect 13219 13348 13820 13376
rect 13219 13345 13231 13348
rect 13173 13339 13231 13345
rect 13814 13336 13820 13348
rect 13872 13376 13878 13388
rect 13872 13348 14872 13376
rect 13872 13336 13878 13348
rect 9493 13311 9551 13317
rect 9493 13277 9505 13311
rect 9539 13308 9551 13311
rect 10318 13308 10324 13320
rect 9539 13280 10324 13308
rect 9539 13277 9551 13280
rect 9493 13271 9551 13277
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 12342 13268 12348 13320
rect 12400 13308 12406 13320
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 12400 13280 14749 13308
rect 12400 13268 12406 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14844 13308 14872 13348
rect 16132 13308 16160 13407
rect 20346 13404 20352 13416
rect 20404 13404 20410 13456
rect 17589 13379 17647 13385
rect 17589 13345 17601 13379
rect 17635 13376 17647 13379
rect 18690 13376 18696 13388
rect 17635 13348 18696 13376
rect 17635 13345 17647 13348
rect 17589 13339 17647 13345
rect 18690 13336 18696 13348
rect 18748 13376 18754 13388
rect 18748 13348 19288 13376
rect 18748 13336 18754 13348
rect 16758 13308 16764 13320
rect 14844 13280 15884 13308
rect 16132 13280 16764 13308
rect 14737 13271 14795 13277
rect 5350 13200 5356 13252
rect 5408 13240 5414 13252
rect 5454 13243 5512 13249
rect 5454 13240 5466 13243
rect 5408 13212 5466 13240
rect 5408 13200 5414 13212
rect 5454 13209 5466 13212
rect 5500 13209 5512 13243
rect 5454 13203 5512 13209
rect 6457 13243 6515 13249
rect 6457 13209 6469 13243
rect 6503 13240 6515 13243
rect 6503 13212 8432 13240
rect 6503 13209 6515 13212
rect 6457 13203 6515 13209
rect 4065 13175 4123 13181
rect 4065 13141 4077 13175
rect 4111 13141 4123 13175
rect 4065 13135 4123 13141
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 5997 13175 6055 13181
rect 5997 13172 6009 13175
rect 4764 13144 6009 13172
rect 4764 13132 4770 13144
rect 5997 13141 6009 13144
rect 6043 13141 6055 13175
rect 5997 13135 6055 13141
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 7834 13172 7840 13184
rect 7055 13144 7840 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 7834 13132 7840 13144
rect 7892 13132 7898 13184
rect 8404 13172 8432 13212
rect 8478 13200 8484 13252
rect 8536 13240 8542 13252
rect 9033 13243 9091 13249
rect 9033 13240 9045 13243
rect 8536 13212 9045 13240
rect 8536 13200 8542 13212
rect 9033 13209 9045 13212
rect 9079 13209 9091 13243
rect 9033 13203 9091 13209
rect 11238 13200 11244 13252
rect 11296 13240 11302 13252
rect 12161 13243 12219 13249
rect 12161 13240 12173 13243
rect 11296 13212 12173 13240
rect 11296 13200 11302 13212
rect 12161 13209 12173 13212
rect 12207 13240 12219 13243
rect 12526 13240 12532 13252
rect 12207 13212 12532 13240
rect 12207 13209 12219 13212
rect 12161 13203 12219 13209
rect 12526 13200 12532 13212
rect 12584 13200 12590 13252
rect 13354 13240 13360 13252
rect 13315 13212 13360 13240
rect 13354 13200 13360 13212
rect 13412 13240 13418 13252
rect 14093 13243 14151 13249
rect 14093 13240 14105 13243
rect 13412 13212 14105 13240
rect 13412 13200 13418 13212
rect 14093 13209 14105 13212
rect 14139 13209 14151 13243
rect 14093 13203 14151 13209
rect 15004 13243 15062 13249
rect 15004 13209 15016 13243
rect 15050 13240 15062 13243
rect 15746 13240 15752 13252
rect 15050 13212 15752 13240
rect 15050 13209 15062 13212
rect 15004 13203 15062 13209
rect 15746 13200 15752 13212
rect 15804 13200 15810 13252
rect 15856 13240 15884 13280
rect 16758 13268 16764 13280
rect 16816 13308 16822 13320
rect 19260 13317 19288 13348
rect 17037 13311 17095 13317
rect 17037 13308 17049 13311
rect 16816 13280 17049 13308
rect 16816 13268 16822 13280
rect 17037 13277 17049 13280
rect 17083 13277 17095 13311
rect 17037 13271 17095 13277
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 19978 13240 19984 13252
rect 15856 13212 19984 13240
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 9766 13172 9772 13184
rect 8404 13144 9772 13172
rect 9766 13132 9772 13144
rect 9824 13132 9830 13184
rect 12250 13132 12256 13184
rect 12308 13172 12314 13184
rect 13265 13175 13323 13181
rect 13265 13172 13277 13175
rect 12308 13144 13277 13172
rect 12308 13132 12314 13144
rect 13265 13141 13277 13144
rect 13311 13141 13323 13175
rect 17678 13172 17684 13184
rect 17639 13144 17684 13172
rect 13265 13135 13323 13141
rect 17678 13132 17684 13144
rect 17736 13132 17742 13184
rect 17773 13175 17831 13181
rect 17773 13141 17785 13175
rect 17819 13172 17831 13175
rect 18046 13172 18052 13184
rect 17819 13144 18052 13172
rect 17819 13141 17831 13144
rect 17773 13135 17831 13141
rect 18046 13132 18052 13144
rect 18104 13132 18110 13184
rect 18601 13175 18659 13181
rect 18601 13141 18613 13175
rect 18647 13172 18659 13175
rect 19610 13172 19616 13184
rect 18647 13144 19616 13172
rect 18647 13141 18659 13144
rect 18601 13135 18659 13141
rect 19610 13132 19616 13144
rect 19668 13132 19674 13184
rect 19886 13172 19892 13184
rect 19847 13144 19892 13172
rect 19886 13132 19892 13144
rect 19944 13132 19950 13184
rect 1104 13082 21896 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21896 13082
rect 1104 13008 21896 13030
rect 1578 12928 1584 12980
rect 1636 12968 1642 12980
rect 4249 12971 4307 12977
rect 4249 12968 4261 12971
rect 1636 12940 4261 12968
rect 1636 12928 1642 12940
rect 4249 12937 4261 12940
rect 4295 12937 4307 12971
rect 4706 12968 4712 12980
rect 4667 12940 4712 12968
rect 4249 12931 4307 12937
rect 4706 12928 4712 12940
rect 4764 12928 4770 12980
rect 5629 12971 5687 12977
rect 5629 12937 5641 12971
rect 5675 12968 5687 12971
rect 8018 12968 8024 12980
rect 5675 12940 8024 12968
rect 5675 12937 5687 12940
rect 5629 12931 5687 12937
rect 8018 12928 8024 12940
rect 8076 12928 8082 12980
rect 8662 12968 8668 12980
rect 8623 12940 8668 12968
rect 8662 12928 8668 12940
rect 8720 12928 8726 12980
rect 10318 12968 10324 12980
rect 10279 12940 10324 12968
rect 10318 12928 10324 12940
rect 10376 12928 10382 12980
rect 10689 12971 10747 12977
rect 10689 12937 10701 12971
rect 10735 12968 10747 12971
rect 12158 12968 12164 12980
rect 10735 12940 12164 12968
rect 10735 12937 10747 12940
rect 10689 12931 10747 12937
rect 12158 12928 12164 12940
rect 12216 12928 12222 12980
rect 12894 12968 12900 12980
rect 12855 12940 12900 12968
rect 12894 12928 12900 12940
rect 12952 12928 12958 12980
rect 14185 12971 14243 12977
rect 14185 12937 14197 12971
rect 14231 12968 14243 12971
rect 14274 12968 14280 12980
rect 14231 12940 14280 12968
rect 14231 12937 14243 12940
rect 14185 12931 14243 12937
rect 14274 12928 14280 12940
rect 14332 12928 14338 12980
rect 15565 12971 15623 12977
rect 15565 12937 15577 12971
rect 15611 12968 15623 12971
rect 18138 12968 18144 12980
rect 15611 12940 18144 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 18138 12928 18144 12940
rect 18196 12928 18202 12980
rect 18690 12968 18696 12980
rect 18651 12940 18696 12968
rect 18690 12928 18696 12940
rect 18748 12928 18754 12980
rect 19978 12968 19984 12980
rect 19939 12940 19984 12968
rect 19978 12928 19984 12940
rect 20036 12928 20042 12980
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 2222 12900 2228 12912
rect 1719 12872 2228 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2222 12860 2228 12872
rect 2280 12860 2286 12912
rect 2593 12903 2651 12909
rect 2593 12869 2605 12903
rect 2639 12900 2651 12903
rect 4062 12900 4068 12912
rect 2639 12872 4068 12900
rect 2639 12869 2651 12872
rect 2593 12863 2651 12869
rect 4062 12860 4068 12872
rect 4120 12860 4126 12912
rect 4617 12903 4675 12909
rect 4617 12869 4629 12903
rect 4663 12900 4675 12903
rect 5166 12900 5172 12912
rect 4663 12872 5172 12900
rect 4663 12869 4675 12872
rect 4617 12863 4675 12869
rect 5166 12860 5172 12872
rect 5224 12860 5230 12912
rect 5718 12860 5724 12912
rect 5776 12900 5782 12912
rect 5776 12872 7328 12900
rect 5776 12860 5782 12872
rect 1949 12835 2007 12841
rect 1949 12801 1961 12835
rect 1995 12832 2007 12835
rect 2682 12832 2688 12844
rect 1995 12804 2688 12832
rect 1995 12801 2007 12804
rect 1949 12795 2007 12801
rect 2682 12792 2688 12804
rect 2740 12792 2746 12844
rect 2869 12835 2927 12841
rect 2869 12801 2881 12835
rect 2915 12832 2927 12835
rect 3510 12832 3516 12844
rect 2915 12804 3516 12832
rect 2915 12801 2927 12804
rect 2869 12795 2927 12801
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 3878 12792 3884 12844
rect 3936 12832 3942 12844
rect 3973 12835 4031 12841
rect 3973 12832 3985 12835
rect 3936 12804 3985 12832
rect 3936 12792 3942 12804
rect 3973 12801 3985 12804
rect 4019 12801 4031 12835
rect 6914 12832 6920 12844
rect 3973 12795 4031 12801
rect 5736 12804 6920 12832
rect 4338 12724 4344 12776
rect 4396 12764 4402 12776
rect 5736 12773 5764 12804
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7300 12841 7328 12872
rect 7392 12872 7788 12900
rect 7009 12835 7067 12841
rect 7009 12801 7021 12835
rect 7055 12801 7067 12835
rect 7009 12795 7067 12801
rect 7285 12835 7343 12841
rect 7285 12801 7297 12835
rect 7331 12801 7343 12835
rect 7285 12795 7343 12801
rect 4801 12767 4859 12773
rect 4801 12764 4813 12767
rect 4396 12736 4813 12764
rect 4396 12724 4402 12736
rect 4801 12733 4813 12736
rect 4847 12733 4859 12767
rect 4801 12727 4859 12733
rect 5721 12767 5779 12773
rect 5721 12733 5733 12767
rect 5767 12733 5779 12767
rect 5902 12764 5908 12776
rect 5863 12736 5908 12764
rect 5721 12727 5779 12733
rect 5902 12724 5908 12736
rect 5960 12724 5966 12776
rect 7024 12764 7052 12795
rect 7392 12764 7420 12872
rect 7558 12841 7564 12844
rect 7552 12795 7564 12841
rect 7616 12832 7622 12844
rect 7760 12832 7788 12872
rect 7834 12860 7840 12912
rect 7892 12900 7898 12912
rect 11790 12909 11796 12912
rect 9186 12903 9244 12909
rect 9186 12900 9198 12903
rect 7892 12872 9198 12900
rect 7892 12860 7898 12872
rect 9186 12869 9198 12872
rect 9232 12869 9244 12903
rect 11784 12900 11796 12909
rect 11751 12872 11796 12900
rect 9186 12863 9244 12869
rect 11784 12863 11796 12872
rect 11790 12860 11796 12863
rect 11848 12860 11854 12912
rect 9766 12832 9772 12844
rect 7616 12804 7652 12832
rect 7760 12804 9772 12832
rect 7558 12792 7564 12795
rect 7616 12792 7622 12804
rect 9766 12792 9772 12804
rect 9824 12792 9830 12844
rect 12912 12832 12940 12928
rect 14553 12903 14611 12909
rect 14553 12869 14565 12903
rect 14599 12900 14611 12903
rect 15470 12900 15476 12912
rect 14599 12872 15476 12900
rect 14599 12869 14611 12872
rect 14553 12863 14611 12869
rect 13173 12835 13231 12841
rect 13173 12832 13185 12835
rect 12912 12804 13185 12832
rect 13173 12801 13185 12804
rect 13219 12801 13231 12835
rect 13173 12795 13231 12801
rect 7024 12736 7420 12764
rect 8294 12724 8300 12776
rect 8352 12764 8358 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8352 12736 8953 12764
rect 8352 12724 8358 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9950 12724 9956 12776
rect 10008 12764 10014 12776
rect 10965 12767 11023 12773
rect 10965 12764 10977 12767
rect 10008 12736 10977 12764
rect 10008 12724 10014 12736
rect 10965 12733 10977 12736
rect 11011 12733 11023 12767
rect 11514 12764 11520 12776
rect 11475 12736 11520 12764
rect 10965 12727 11023 12733
rect 11514 12724 11520 12736
rect 11572 12724 11578 12776
rect 3053 12699 3111 12705
rect 3053 12665 3065 12699
rect 3099 12696 3111 12699
rect 6638 12696 6644 12708
rect 3099 12668 6644 12696
rect 3099 12665 3111 12668
rect 3053 12659 3111 12665
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 14568 12696 14596 12863
rect 15470 12860 15476 12872
rect 15528 12860 15534 12912
rect 17954 12900 17960 12912
rect 17328 12872 17960 12900
rect 17328 12841 17356 12872
rect 17954 12860 17960 12872
rect 18012 12900 18018 12912
rect 19058 12900 19064 12912
rect 18012 12872 19064 12900
rect 18012 12860 18018 12872
rect 19058 12860 19064 12872
rect 19116 12900 19122 12912
rect 19116 12872 21404 12900
rect 19116 12860 19122 12872
rect 17586 12841 17592 12844
rect 15197 12835 15255 12841
rect 15197 12801 15209 12835
rect 15243 12832 15255 12835
rect 15841 12835 15899 12841
rect 15841 12832 15853 12835
rect 15243 12804 15853 12832
rect 15243 12801 15255 12804
rect 15197 12795 15255 12801
rect 15841 12801 15853 12804
rect 15887 12801 15899 12835
rect 15841 12795 15899 12801
rect 17313 12835 17371 12841
rect 17313 12801 17325 12835
rect 17359 12801 17371 12835
rect 17580 12832 17592 12841
rect 17547 12804 17592 12832
rect 17313 12795 17371 12801
rect 17580 12795 17592 12804
rect 17586 12792 17592 12795
rect 17644 12792 17650 12844
rect 21082 12832 21088 12844
rect 21140 12841 21146 12844
rect 21376 12841 21404 12872
rect 21052 12804 21088 12832
rect 21082 12792 21088 12804
rect 21140 12795 21152 12841
rect 21361 12835 21419 12841
rect 21361 12801 21373 12835
rect 21407 12801 21419 12835
rect 21361 12795 21419 12801
rect 21140 12792 21146 12795
rect 15013 12767 15071 12773
rect 15013 12733 15025 12767
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 15105 12767 15163 12773
rect 15105 12733 15117 12767
rect 15151 12764 15163 12767
rect 15286 12764 15292 12776
rect 15151 12736 15292 12764
rect 15151 12733 15163 12736
rect 15105 12727 15163 12733
rect 13648 12668 14596 12696
rect 15028 12696 15056 12727
rect 15286 12724 15292 12736
rect 15344 12724 15350 12776
rect 15378 12696 15384 12708
rect 15028 12668 15384 12696
rect 2130 12628 2136 12640
rect 2091 12600 2136 12628
rect 2130 12588 2136 12600
rect 2188 12588 2194 12640
rect 3326 12628 3332 12640
rect 3287 12600 3332 12628
rect 3326 12588 3332 12600
rect 3384 12588 3390 12640
rect 4614 12588 4620 12640
rect 4672 12628 4678 12640
rect 5261 12631 5319 12637
rect 5261 12628 5273 12631
rect 4672 12600 5273 12628
rect 4672 12588 4678 12600
rect 5261 12597 5273 12600
rect 5307 12597 5319 12631
rect 5261 12591 5319 12597
rect 6365 12631 6423 12637
rect 6365 12597 6377 12631
rect 6411 12628 6423 12631
rect 9582 12628 9588 12640
rect 6411 12600 9588 12628
rect 6411 12597 6423 12600
rect 6365 12591 6423 12597
rect 9582 12588 9588 12600
rect 9640 12588 9646 12640
rect 12158 12588 12164 12640
rect 12216 12628 12222 12640
rect 13648 12628 13676 12668
rect 15378 12656 15384 12668
rect 15436 12696 15442 12708
rect 16022 12696 16028 12708
rect 15436 12668 16028 12696
rect 15436 12656 15442 12668
rect 16022 12656 16028 12668
rect 16080 12656 16086 12708
rect 13814 12628 13820 12640
rect 12216 12600 13676 12628
rect 13775 12600 13820 12628
rect 12216 12588 12222 12600
rect 13814 12588 13820 12600
rect 13872 12588 13878 12640
rect 14274 12588 14280 12640
rect 14332 12628 14338 12640
rect 16669 12631 16727 12637
rect 16669 12628 16681 12631
rect 14332 12600 16681 12628
rect 14332 12588 14338 12600
rect 16669 12597 16681 12600
rect 16715 12628 16727 12631
rect 16942 12628 16948 12640
rect 16715 12600 16948 12628
rect 16715 12597 16727 12600
rect 16669 12591 16727 12597
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 18966 12588 18972 12640
rect 19024 12628 19030 12640
rect 19061 12631 19119 12637
rect 19061 12628 19073 12631
rect 19024 12600 19073 12628
rect 19024 12588 19030 12600
rect 19061 12597 19073 12600
rect 19107 12628 19119 12631
rect 19702 12628 19708 12640
rect 19107 12600 19708 12628
rect 19107 12597 19119 12600
rect 19061 12591 19119 12597
rect 19702 12588 19708 12600
rect 19760 12588 19766 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 1394 12424 1400 12436
rect 1355 12396 1400 12424
rect 1394 12384 1400 12396
rect 1452 12384 1458 12436
rect 2961 12427 3019 12433
rect 2961 12393 2973 12427
rect 3007 12424 3019 12427
rect 4062 12424 4068 12436
rect 3007 12396 4068 12424
rect 3007 12393 3019 12396
rect 2961 12387 3019 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 5074 12424 5080 12436
rect 4273 12396 5080 12424
rect 2498 12356 2504 12368
rect 2459 12328 2504 12356
rect 2498 12316 2504 12328
rect 2556 12316 2562 12368
rect 3510 12316 3516 12368
rect 3568 12356 3574 12368
rect 4273 12356 4301 12396
rect 5074 12384 5080 12396
rect 5132 12384 5138 12436
rect 5813 12427 5871 12433
rect 5813 12393 5825 12427
rect 5859 12424 5871 12427
rect 5902 12424 5908 12436
rect 5859 12396 5908 12424
rect 5859 12393 5871 12396
rect 5813 12387 5871 12393
rect 5902 12384 5908 12396
rect 5960 12424 5966 12436
rect 6546 12424 6552 12436
rect 5960 12396 6552 12424
rect 5960 12384 5966 12396
rect 6546 12384 6552 12396
rect 6604 12384 6610 12436
rect 14369 12427 14427 12433
rect 14369 12393 14381 12427
rect 14415 12424 14427 12427
rect 15378 12424 15384 12436
rect 14415 12396 15384 12424
rect 14415 12393 14427 12396
rect 14369 12387 14427 12393
rect 15378 12384 15384 12396
rect 15436 12384 15442 12436
rect 15746 12384 15752 12436
rect 15804 12424 15810 12436
rect 16669 12427 16727 12433
rect 16669 12424 16681 12427
rect 15804 12396 16681 12424
rect 15804 12384 15810 12396
rect 16669 12393 16681 12396
rect 16715 12393 16727 12427
rect 16669 12387 16727 12393
rect 17497 12427 17555 12433
rect 17497 12393 17509 12427
rect 17543 12424 17555 12427
rect 17678 12424 17684 12436
rect 17543 12396 17684 12424
rect 17543 12393 17555 12396
rect 17497 12387 17555 12393
rect 17678 12384 17684 12396
rect 17736 12384 17742 12436
rect 18046 12384 18052 12436
rect 18104 12424 18110 12436
rect 19245 12427 19303 12433
rect 19245 12424 19257 12427
rect 18104 12396 19257 12424
rect 18104 12384 18110 12396
rect 19245 12393 19257 12396
rect 19291 12393 19303 12427
rect 19245 12387 19303 12393
rect 3568 12328 4301 12356
rect 3568 12316 3574 12328
rect 7466 12316 7472 12368
rect 7524 12356 7530 12368
rect 8110 12356 8116 12368
rect 7524 12328 8116 12356
rect 7524 12316 7530 12328
rect 8110 12316 8116 12328
rect 8168 12316 8174 12368
rect 17586 12316 17592 12368
rect 17644 12356 17650 12368
rect 17644 12328 19840 12356
rect 17644 12316 17650 12328
rect 2958 12288 2964 12300
rect 2056 12260 2964 12288
rect 1394 12180 1400 12232
rect 1452 12220 1458 12232
rect 2056 12229 2084 12260
rect 2958 12248 2964 12260
rect 3016 12248 3022 12300
rect 8018 12248 8024 12300
rect 8076 12288 8082 12300
rect 8297 12291 8355 12297
rect 8297 12288 8309 12291
rect 8076 12260 8309 12288
rect 8076 12248 8082 12260
rect 8297 12257 8309 12260
rect 8343 12257 8355 12291
rect 8297 12251 8355 12257
rect 15749 12291 15807 12297
rect 15749 12257 15761 12291
rect 15795 12288 15807 12291
rect 16942 12288 16948 12300
rect 15795 12260 16948 12288
rect 15795 12257 15807 12260
rect 15749 12251 15807 12257
rect 16942 12248 16948 12260
rect 17000 12288 17006 12300
rect 17954 12288 17960 12300
rect 17000 12260 17960 12288
rect 17000 12248 17006 12260
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 18156 12297 18184 12328
rect 18141 12291 18199 12297
rect 18141 12257 18153 12291
rect 18187 12257 18199 12291
rect 19702 12288 19708 12300
rect 19663 12260 19708 12288
rect 18141 12251 18199 12257
rect 19702 12248 19708 12260
rect 19760 12248 19766 12300
rect 19812 12297 19840 12328
rect 19797 12291 19855 12297
rect 19797 12257 19809 12291
rect 19843 12257 19855 12291
rect 19797 12251 19855 12257
rect 1581 12223 1639 12229
rect 1581 12220 1593 12223
rect 1452 12192 1593 12220
rect 1452 12180 1458 12192
rect 1581 12189 1593 12192
rect 1627 12189 1639 12223
rect 1581 12183 1639 12189
rect 2041 12223 2099 12229
rect 2041 12189 2053 12223
rect 2087 12189 2099 12223
rect 2041 12183 2099 12189
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2332 12152 2360 12183
rect 2406 12180 2412 12232
rect 2464 12220 2470 12232
rect 2777 12223 2835 12229
rect 2777 12220 2789 12223
rect 2464 12192 2789 12220
rect 2464 12180 2470 12192
rect 2777 12189 2789 12192
rect 2823 12189 2835 12223
rect 2777 12183 2835 12189
rect 3418 12180 3424 12232
rect 3476 12220 3482 12232
rect 3973 12223 4031 12229
rect 3973 12220 3985 12223
rect 3476 12192 3985 12220
rect 3476 12180 3482 12192
rect 3973 12189 3985 12192
rect 4019 12189 4031 12223
rect 3973 12183 4031 12189
rect 4433 12223 4491 12229
rect 4433 12189 4445 12223
rect 4479 12220 4491 12223
rect 5718 12220 5724 12232
rect 4479 12192 5724 12220
rect 4479 12189 4491 12192
rect 4433 12183 4491 12189
rect 5718 12180 5724 12192
rect 5776 12180 5782 12232
rect 7190 12220 7196 12232
rect 7248 12229 7254 12232
rect 7160 12192 7196 12220
rect 7190 12180 7196 12192
rect 7248 12183 7260 12229
rect 7469 12223 7527 12229
rect 7469 12189 7481 12223
rect 7515 12220 7527 12223
rect 7515 12192 8340 12220
rect 7515 12189 7527 12192
rect 7469 12183 7527 12189
rect 7248 12180 7254 12183
rect 8312 12164 8340 12192
rect 8662 12180 8668 12232
rect 8720 12220 8726 12232
rect 11054 12220 11060 12232
rect 8720 12192 11060 12220
rect 8720 12180 8726 12192
rect 11054 12180 11060 12192
rect 11112 12180 11118 12232
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12220 11207 12223
rect 11514 12220 11520 12232
rect 11195 12192 11520 12220
rect 11195 12189 11207 12192
rect 11149 12183 11207 12189
rect 11514 12180 11520 12192
rect 11572 12220 11578 12232
rect 11882 12220 11888 12232
rect 11572 12192 11888 12220
rect 11572 12180 11578 12192
rect 11882 12180 11888 12192
rect 11940 12220 11946 12232
rect 12342 12220 12348 12232
rect 11940 12192 12348 12220
rect 11940 12180 11946 12192
rect 12342 12180 12348 12192
rect 12400 12220 12406 12232
rect 12897 12223 12955 12229
rect 12897 12220 12909 12223
rect 12400 12192 12909 12220
rect 12400 12180 12406 12192
rect 12897 12189 12909 12192
rect 12943 12189 12955 12223
rect 12897 12183 12955 12189
rect 12986 12180 12992 12232
rect 13044 12220 13050 12232
rect 16022 12220 16028 12232
rect 13044 12192 15608 12220
rect 15983 12192 16028 12220
rect 13044 12180 13050 12192
rect 2866 12152 2872 12164
rect 2332 12124 2872 12152
rect 2866 12112 2872 12124
rect 2924 12152 2930 12164
rect 3050 12152 3056 12164
rect 2924 12124 3056 12152
rect 2924 12112 2930 12124
rect 3050 12112 3056 12124
rect 3108 12112 3114 12164
rect 3326 12112 3332 12164
rect 3384 12152 3390 12164
rect 4678 12155 4736 12161
rect 4678 12152 4690 12155
rect 3384 12124 4690 12152
rect 3384 12112 3390 12124
rect 4678 12121 4690 12124
rect 4724 12121 4736 12155
rect 4678 12115 4736 12121
rect 4798 12112 4804 12164
rect 4856 12152 4862 12164
rect 4856 12124 7788 12152
rect 4856 12112 4862 12124
rect 1578 12044 1584 12096
rect 1636 12084 1642 12096
rect 1857 12087 1915 12093
rect 1857 12084 1869 12087
rect 1636 12056 1869 12084
rect 1636 12044 1642 12056
rect 1857 12053 1869 12056
rect 1903 12053 1915 12087
rect 1857 12047 1915 12053
rect 3421 12087 3479 12093
rect 3421 12053 3433 12087
rect 3467 12084 3479 12087
rect 3510 12084 3516 12096
rect 3467 12056 3516 12084
rect 3467 12053 3479 12056
rect 3421 12047 3479 12053
rect 3510 12044 3516 12056
rect 3568 12044 3574 12096
rect 3786 12084 3792 12096
rect 3747 12056 3792 12084
rect 3786 12044 3792 12056
rect 3844 12044 3850 12096
rect 5994 12044 6000 12096
rect 6052 12084 6058 12096
rect 7760 12093 7788 12124
rect 8294 12112 8300 12164
rect 8352 12112 8358 12164
rect 10870 12112 10876 12164
rect 10928 12161 10934 12164
rect 10928 12152 10940 12161
rect 12652 12155 12710 12161
rect 10928 12124 11560 12152
rect 10928 12115 10940 12124
rect 10928 12112 10934 12115
rect 6089 12087 6147 12093
rect 6089 12084 6101 12087
rect 6052 12056 6101 12084
rect 6052 12044 6058 12056
rect 6089 12053 6101 12056
rect 6135 12053 6147 12087
rect 6089 12047 6147 12053
rect 7745 12087 7803 12093
rect 7745 12053 7757 12087
rect 7791 12053 7803 12087
rect 8110 12084 8116 12096
rect 8071 12056 8116 12084
rect 7745 12047 7803 12053
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 8202 12044 8208 12096
rect 8260 12084 8266 12096
rect 8260 12056 8305 12084
rect 8260 12044 8266 12056
rect 8386 12044 8392 12096
rect 8444 12084 8450 12096
rect 9033 12087 9091 12093
rect 9033 12084 9045 12087
rect 8444 12056 9045 12084
rect 8444 12044 8450 12056
rect 9033 12053 9045 12056
rect 9079 12053 9091 12087
rect 9766 12084 9772 12096
rect 9679 12056 9772 12084
rect 9033 12047 9091 12053
rect 9766 12044 9772 12056
rect 9824 12084 9830 12096
rect 10502 12084 10508 12096
rect 9824 12056 10508 12084
rect 9824 12044 9830 12056
rect 10502 12044 10508 12056
rect 10560 12044 10566 12096
rect 11532 12093 11560 12124
rect 12652 12121 12664 12155
rect 12698 12152 12710 12155
rect 13814 12152 13820 12164
rect 12698 12124 13820 12152
rect 12698 12121 12710 12124
rect 12652 12115 12710 12121
rect 13814 12112 13820 12124
rect 13872 12112 13878 12164
rect 15378 12112 15384 12164
rect 15436 12152 15442 12164
rect 15482 12155 15540 12161
rect 15482 12152 15494 12155
rect 15436 12124 15494 12152
rect 15436 12112 15442 12124
rect 15482 12121 15494 12124
rect 15528 12121 15540 12155
rect 15580 12152 15608 12192
rect 16022 12180 16028 12192
rect 16080 12180 16086 12232
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 17034 12220 17040 12232
rect 16448 12192 17040 12220
rect 16448 12180 16454 12192
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 19610 12220 19616 12232
rect 19571 12192 19616 12220
rect 19610 12180 19616 12192
rect 19668 12180 19674 12232
rect 17957 12155 18015 12161
rect 17957 12152 17969 12155
rect 15580 12124 17969 12152
rect 15482 12115 15540 12121
rect 17957 12121 17969 12124
rect 18003 12152 18015 12155
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 18003 12124 18521 12152
rect 18003 12121 18015 12124
rect 17957 12115 18015 12121
rect 18509 12121 18521 12124
rect 18555 12121 18567 12155
rect 18509 12115 18567 12121
rect 11517 12087 11575 12093
rect 11517 12053 11529 12087
rect 11563 12053 11575 12087
rect 13170 12084 13176 12096
rect 13131 12056 13176 12084
rect 11517 12047 11575 12053
rect 13170 12044 13176 12056
rect 13228 12044 13234 12096
rect 13630 12084 13636 12096
rect 13591 12056 13636 12084
rect 13630 12044 13636 12056
rect 13688 12044 13694 12096
rect 13722 12044 13728 12096
rect 13780 12084 13786 12096
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 13780 12056 17877 12084
rect 13780 12044 13786 12056
rect 17865 12053 17877 12056
rect 17911 12084 17923 12087
rect 20714 12084 20720 12096
rect 17911 12056 20720 12084
rect 17911 12053 17923 12056
rect 17865 12047 17923 12053
rect 20714 12044 20720 12056
rect 20772 12044 20778 12096
rect 1104 11994 21896 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21896 11994
rect 1104 11920 21896 11942
rect 1397 11883 1455 11889
rect 1397 11849 1409 11883
rect 1443 11880 1455 11883
rect 1670 11880 1676 11892
rect 1443 11852 1676 11880
rect 1443 11849 1455 11852
rect 1397 11843 1455 11849
rect 1670 11840 1676 11852
rect 1728 11840 1734 11892
rect 3421 11883 3479 11889
rect 2332 11852 2774 11880
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1857 11747 1915 11753
rect 1857 11713 1869 11747
rect 1903 11744 1915 11747
rect 2222 11744 2228 11756
rect 1903 11716 2228 11744
rect 1903 11713 1915 11716
rect 1857 11707 1915 11713
rect 1596 11676 1624 11707
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2332 11753 2360 11852
rect 2746 11812 2774 11852
rect 3421 11849 3433 11883
rect 3467 11880 3479 11883
rect 5810 11880 5816 11892
rect 3467 11852 5816 11880
rect 3467 11849 3479 11852
rect 3421 11843 3479 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6104 11852 7972 11880
rect 4832 11815 4890 11821
rect 2746 11784 3924 11812
rect 2317 11747 2375 11753
rect 2317 11713 2329 11747
rect 2363 11713 2375 11747
rect 2958 11744 2964 11756
rect 2919 11716 2964 11744
rect 2317 11707 2375 11713
rect 2958 11704 2964 11716
rect 3016 11704 3022 11756
rect 3237 11747 3295 11753
rect 3237 11713 3249 11747
rect 3283 11744 3295 11747
rect 3786 11744 3792 11756
rect 3283 11716 3792 11744
rect 3283 11713 3295 11716
rect 3237 11707 3295 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 3896 11744 3924 11784
rect 4832 11781 4844 11815
rect 4878 11812 4890 11815
rect 5353 11815 5411 11821
rect 5353 11812 5365 11815
rect 4878 11784 5365 11812
rect 4878 11781 4890 11784
rect 4832 11775 4890 11781
rect 5353 11781 5365 11784
rect 5399 11781 5411 11815
rect 5353 11775 5411 11781
rect 5077 11747 5135 11753
rect 3896 11716 5028 11744
rect 3142 11676 3148 11688
rect 1596 11648 3148 11676
rect 3142 11636 3148 11648
rect 3200 11636 3206 11688
rect 5000 11676 5028 11716
rect 5077 11713 5089 11747
rect 5123 11744 5135 11747
rect 5718 11744 5724 11756
rect 5123 11716 5724 11744
rect 5123 11713 5135 11716
rect 5077 11707 5135 11713
rect 5718 11704 5724 11716
rect 5776 11704 5782 11756
rect 5994 11744 6000 11756
rect 5955 11716 6000 11744
rect 5994 11704 6000 11716
rect 6052 11704 6058 11756
rect 6104 11676 6132 11852
rect 6730 11812 6736 11824
rect 6691 11784 6736 11812
rect 6730 11772 6736 11784
rect 6788 11772 6794 11824
rect 7644 11815 7702 11821
rect 7644 11781 7656 11815
rect 7690 11812 7702 11815
rect 7834 11812 7840 11824
rect 7690 11784 7840 11812
rect 7690 11781 7702 11784
rect 7644 11775 7702 11781
rect 7834 11772 7840 11784
rect 7892 11772 7898 11824
rect 7944 11812 7972 11852
rect 8018 11840 8024 11892
rect 8076 11880 8082 11892
rect 8757 11883 8815 11889
rect 8757 11880 8769 11883
rect 8076 11852 8769 11880
rect 8076 11840 8082 11852
rect 8757 11849 8769 11852
rect 8803 11849 8815 11883
rect 8757 11843 8815 11849
rect 9769 11883 9827 11889
rect 9769 11849 9781 11883
rect 9815 11880 9827 11883
rect 9950 11880 9956 11892
rect 9815 11852 9956 11880
rect 9815 11849 9827 11852
rect 9769 11843 9827 11849
rect 9950 11840 9956 11852
rect 10008 11840 10014 11892
rect 10137 11883 10195 11889
rect 10137 11849 10149 11883
rect 10183 11849 10195 11883
rect 10137 11843 10195 11849
rect 10689 11883 10747 11889
rect 10689 11849 10701 11883
rect 10735 11880 10747 11883
rect 11793 11883 11851 11889
rect 11793 11880 11805 11883
rect 10735 11852 11805 11880
rect 10735 11849 10747 11852
rect 10689 11843 10747 11849
rect 11793 11849 11805 11852
rect 11839 11849 11851 11883
rect 11793 11843 11851 11849
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 12250 11880 12256 11892
rect 12207 11852 12256 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 10042 11812 10048 11824
rect 7944 11784 10048 11812
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 10152 11812 10180 11843
rect 12250 11840 12256 11852
rect 12308 11880 12314 11892
rect 13722 11880 13728 11892
rect 12308 11852 13728 11880
rect 12308 11840 12314 11852
rect 13722 11840 13728 11852
rect 13780 11840 13786 11892
rect 15286 11840 15292 11892
rect 15344 11880 15350 11892
rect 15381 11883 15439 11889
rect 15381 11880 15393 11883
rect 15344 11852 15393 11880
rect 15344 11840 15350 11852
rect 15381 11849 15393 11852
rect 15427 11849 15439 11883
rect 15381 11843 15439 11849
rect 15470 11840 15476 11892
rect 15528 11880 15534 11892
rect 15841 11883 15899 11889
rect 15841 11880 15853 11883
rect 15528 11852 15853 11880
rect 15528 11840 15534 11852
rect 15841 11849 15853 11852
rect 15887 11849 15899 11883
rect 15841 11843 15899 11849
rect 21082 11840 21088 11892
rect 21140 11880 21146 11892
rect 21177 11883 21235 11889
rect 21177 11880 21189 11883
rect 21140 11852 21189 11880
rect 21140 11840 21146 11852
rect 21177 11849 21189 11852
rect 21223 11849 21235 11883
rect 21177 11843 21235 11849
rect 10781 11815 10839 11821
rect 10781 11812 10793 11815
rect 10152 11784 10793 11812
rect 10781 11781 10793 11784
rect 10827 11781 10839 11815
rect 10781 11775 10839 11781
rect 11882 11772 11888 11824
rect 11940 11812 11946 11824
rect 18448 11815 18506 11821
rect 11940 11784 13768 11812
rect 11940 11772 11946 11784
rect 6825 11747 6883 11753
rect 6825 11713 6837 11747
rect 6871 11744 6883 11747
rect 10870 11744 10876 11756
rect 6871 11716 9444 11744
rect 6871 11713 6883 11716
rect 6825 11707 6883 11713
rect 5000 11648 6132 11676
rect 6917 11679 6975 11685
rect 6917 11645 6929 11679
rect 6963 11645 6975 11679
rect 6917 11639 6975 11645
rect 7377 11679 7435 11685
rect 7377 11645 7389 11679
rect 7423 11645 7435 11679
rect 7377 11639 7435 11645
rect 2041 11611 2099 11617
rect 2041 11577 2053 11611
rect 2087 11608 2099 11611
rect 2590 11608 2596 11620
rect 2087 11580 2596 11608
rect 2087 11577 2099 11580
rect 2041 11571 2099 11577
rect 2590 11568 2596 11580
rect 2648 11568 2654 11620
rect 3878 11608 3884 11620
rect 2700 11580 3884 11608
rect 2501 11543 2559 11549
rect 2501 11509 2513 11543
rect 2547 11540 2559 11543
rect 2700 11540 2728 11580
rect 3878 11568 3884 11580
rect 3936 11568 3942 11620
rect 5994 11568 6000 11620
rect 6052 11608 6058 11620
rect 6932 11608 6960 11639
rect 6052 11580 6960 11608
rect 6052 11568 6058 11580
rect 2547 11512 2728 11540
rect 2547 11509 2559 11512
rect 2501 11503 2559 11509
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 2832 11512 2877 11540
rect 2832 11500 2838 11512
rect 3050 11500 3056 11552
rect 3108 11540 3114 11552
rect 3418 11540 3424 11552
rect 3108 11512 3424 11540
rect 3108 11500 3114 11512
rect 3418 11500 3424 11512
rect 3476 11500 3482 11552
rect 3697 11543 3755 11549
rect 3697 11509 3709 11543
rect 3743 11540 3755 11543
rect 3970 11540 3976 11552
rect 3743 11512 3976 11540
rect 3743 11509 3755 11512
rect 3697 11503 3755 11509
rect 3970 11500 3976 11512
rect 4028 11500 4034 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 6365 11543 6423 11549
rect 6365 11540 6377 11543
rect 4856 11512 6377 11540
rect 4856 11500 4862 11512
rect 6365 11509 6377 11512
rect 6411 11509 6423 11543
rect 7392 11540 7420 11639
rect 8294 11540 8300 11552
rect 7392 11512 8300 11540
rect 6365 11503 6423 11509
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 8570 11500 8576 11552
rect 8628 11540 8634 11552
rect 9033 11543 9091 11549
rect 9033 11540 9045 11543
rect 8628 11512 9045 11540
rect 8628 11500 8634 11512
rect 9033 11509 9045 11512
rect 9079 11540 9091 11543
rect 9306 11540 9312 11552
rect 9079 11512 9312 11540
rect 9079 11509 9091 11512
rect 9033 11503 9091 11509
rect 9306 11500 9312 11512
rect 9364 11500 9370 11552
rect 9416 11540 9444 11716
rect 9600 11716 10876 11744
rect 9600 11685 9628 11716
rect 10870 11704 10876 11716
rect 10928 11704 10934 11756
rect 12253 11747 12311 11753
rect 12253 11713 12265 11747
rect 12299 11744 12311 11747
rect 12618 11744 12624 11756
rect 12299 11716 12624 11744
rect 12299 11713 12311 11716
rect 12253 11707 12311 11713
rect 12618 11704 12624 11716
rect 12676 11744 12682 11756
rect 12986 11744 12992 11756
rect 12676 11716 12992 11744
rect 12676 11704 12682 11716
rect 12986 11704 12992 11716
rect 13044 11704 13050 11756
rect 13446 11744 13452 11756
rect 13407 11716 13452 11744
rect 13446 11704 13452 11716
rect 13504 11704 13510 11756
rect 13740 11753 13768 11784
rect 18448 11781 18460 11815
rect 18494 11812 18506 11815
rect 19886 11812 19892 11824
rect 18494 11784 19892 11812
rect 18494 11781 18506 11784
rect 18448 11775 18506 11781
rect 19886 11772 19892 11784
rect 19944 11772 19950 11824
rect 13725 11747 13783 11753
rect 13725 11713 13737 11747
rect 13771 11713 13783 11747
rect 13725 11707 13783 11713
rect 13992 11747 14050 11753
rect 13992 11713 14004 11747
rect 14038 11744 14050 11747
rect 14274 11744 14280 11756
rect 14038 11716 14280 11744
rect 14038 11713 14050 11716
rect 13992 11707 14050 11713
rect 14274 11704 14280 11716
rect 14332 11704 14338 11756
rect 15746 11744 15752 11756
rect 15707 11716 15752 11744
rect 15746 11704 15752 11716
rect 15804 11744 15810 11756
rect 16669 11747 16727 11753
rect 16669 11744 16681 11747
rect 15804 11716 16681 11744
rect 15804 11704 15810 11716
rect 16669 11713 16681 11716
rect 16715 11713 16727 11747
rect 18969 11747 19027 11753
rect 18969 11744 18981 11747
rect 16669 11707 16727 11713
rect 17604 11716 18981 11744
rect 9585 11679 9643 11685
rect 9585 11645 9597 11679
rect 9631 11645 9643 11679
rect 9585 11639 9643 11645
rect 9677 11679 9735 11685
rect 9677 11645 9689 11679
rect 9723 11676 9735 11679
rect 9858 11676 9864 11688
rect 9723 11648 9864 11676
rect 9723 11645 9735 11648
rect 9677 11639 9735 11645
rect 9858 11636 9864 11648
rect 9916 11636 9922 11688
rect 10502 11676 10508 11688
rect 10463 11648 10508 11676
rect 10502 11636 10508 11648
rect 10560 11636 10566 11688
rect 10888 11676 10916 11704
rect 12345 11679 12403 11685
rect 12345 11676 12357 11679
rect 10888 11648 12357 11676
rect 12345 11645 12357 11648
rect 12391 11645 12403 11679
rect 12345 11639 12403 11645
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11645 15991 11679
rect 15933 11639 15991 11645
rect 11149 11611 11207 11617
rect 11149 11577 11161 11611
rect 11195 11608 11207 11611
rect 15948 11608 15976 11639
rect 17310 11608 17316 11620
rect 11195 11580 13400 11608
rect 11195 11577 11207 11580
rect 11149 11571 11207 11577
rect 11974 11540 11980 11552
rect 9416 11512 11980 11540
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12802 11540 12808 11552
rect 12763 11512 12808 11540
rect 12802 11500 12808 11512
rect 12860 11500 12866 11552
rect 13372 11540 13400 11580
rect 15120 11580 15976 11608
rect 17223 11580 17316 11608
rect 14458 11540 14464 11552
rect 13372 11512 14464 11540
rect 14458 11500 14464 11512
rect 14516 11500 14522 11552
rect 14734 11500 14740 11552
rect 14792 11540 14798 11552
rect 15120 11549 15148 11580
rect 17310 11568 17316 11580
rect 17368 11608 17374 11620
rect 17604 11608 17632 11716
rect 18969 11713 18981 11716
rect 19015 11713 19027 11747
rect 18969 11707 19027 11713
rect 20901 11747 20959 11753
rect 20901 11713 20913 11747
rect 20947 11744 20959 11747
rect 21358 11744 21364 11756
rect 20947 11716 21364 11744
rect 20947 11713 20959 11716
rect 20901 11707 20959 11713
rect 21358 11704 21364 11716
rect 21416 11704 21422 11756
rect 18693 11679 18751 11685
rect 18693 11645 18705 11679
rect 18739 11676 18751 11679
rect 19058 11676 19064 11688
rect 18739 11648 19064 11676
rect 18739 11645 18751 11648
rect 18693 11639 18751 11645
rect 19058 11636 19064 11648
rect 19116 11636 19122 11688
rect 17368 11580 17632 11608
rect 17368 11568 17374 11580
rect 15105 11543 15163 11549
rect 15105 11540 15117 11543
rect 14792 11512 15117 11540
rect 14792 11500 14798 11512
rect 15105 11509 15117 11512
rect 15151 11509 15163 11543
rect 15105 11503 15163 11509
rect 17494 11500 17500 11552
rect 17552 11540 17558 11552
rect 19613 11543 19671 11549
rect 19613 11540 19625 11543
rect 17552 11512 19625 11540
rect 17552 11500 17558 11512
rect 19613 11509 19625 11512
rect 19659 11509 19671 11543
rect 19613 11503 19671 11509
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2958 11296 2964 11348
rect 3016 11336 3022 11348
rect 4341 11339 4399 11345
rect 4341 11336 4353 11339
rect 3016 11308 4353 11336
rect 3016 11296 3022 11308
rect 4341 11305 4353 11308
rect 4387 11305 4399 11339
rect 4341 11299 4399 11305
rect 4430 11296 4436 11348
rect 4488 11336 4494 11348
rect 5810 11336 5816 11348
rect 4488 11308 5816 11336
rect 4488 11296 4494 11308
rect 5810 11296 5816 11308
rect 5868 11296 5874 11348
rect 6365 11339 6423 11345
rect 6365 11305 6377 11339
rect 6411 11336 6423 11339
rect 6411 11308 7880 11336
rect 6411 11305 6423 11308
rect 6365 11299 6423 11305
rect 7852 11280 7880 11308
rect 7926 11296 7932 11348
rect 7984 11336 7990 11348
rect 8021 11339 8079 11345
rect 8021 11336 8033 11339
rect 7984 11308 8033 11336
rect 7984 11296 7990 11308
rect 8021 11305 8033 11308
rect 8067 11305 8079 11339
rect 8021 11299 8079 11305
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8260 11308 8953 11336
rect 8260 11296 8266 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9398 11296 9404 11348
rect 9456 11336 9462 11348
rect 13630 11336 13636 11348
rect 9456 11308 13636 11336
rect 9456 11296 9462 11308
rect 13630 11296 13636 11308
rect 13688 11296 13694 11348
rect 15102 11336 15108 11348
rect 15063 11308 15108 11336
rect 15102 11296 15108 11308
rect 15160 11296 15166 11348
rect 18049 11339 18107 11345
rect 18049 11305 18061 11339
rect 18095 11336 18107 11339
rect 18230 11336 18236 11348
rect 18095 11308 18236 11336
rect 18095 11305 18107 11308
rect 18049 11299 18107 11305
rect 18230 11296 18236 11308
rect 18288 11296 18294 11348
rect 2685 11271 2743 11277
rect 2685 11268 2697 11271
rect 1964 11240 2697 11268
rect 1854 11200 1860 11212
rect 1815 11172 1860 11200
rect 1854 11160 1860 11172
rect 1912 11160 1918 11212
rect 1964 11209 1992 11240
rect 2685 11237 2697 11240
rect 2731 11237 2743 11271
rect 2685 11231 2743 11237
rect 3326 11228 3332 11280
rect 3384 11268 3390 11280
rect 3881 11271 3939 11277
rect 3881 11268 3893 11271
rect 3384 11240 3893 11268
rect 3384 11228 3390 11240
rect 3881 11237 3893 11240
rect 3927 11237 3939 11271
rect 5353 11271 5411 11277
rect 5353 11268 5365 11271
rect 3881 11231 3939 11237
rect 4724 11240 5365 11268
rect 1949 11203 2007 11209
rect 1949 11169 1961 11203
rect 1995 11169 2007 11203
rect 3234 11200 3240 11212
rect 3195 11172 3240 11200
rect 1949 11163 2007 11169
rect 3234 11160 3240 11172
rect 3292 11160 3298 11212
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4028 11172 4384 11200
rect 4028 11160 4034 11172
rect 2130 11092 2136 11144
rect 2188 11132 2194 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 2188 11104 4077 11132
rect 2188 11092 2194 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4065 11095 4123 11101
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11064 3203 11067
rect 4246 11064 4252 11076
rect 3191 11036 4252 11064
rect 3191 11033 3203 11036
rect 3145 11027 3203 11033
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4356 11064 4384 11172
rect 4724 11141 4752 11240
rect 5353 11237 5365 11240
rect 5399 11237 5411 11271
rect 5353 11231 5411 11237
rect 5442 11228 5448 11280
rect 5500 11268 5506 11280
rect 6730 11268 6736 11280
rect 5500 11240 6736 11268
rect 5500 11228 5506 11240
rect 6730 11228 6736 11240
rect 6788 11228 6794 11280
rect 7834 11228 7840 11280
rect 7892 11268 7898 11280
rect 13265 11271 13323 11277
rect 7892 11240 9536 11268
rect 7892 11228 7898 11240
rect 4798 11160 4804 11212
rect 4856 11200 4862 11212
rect 4985 11203 5043 11209
rect 4856 11172 4901 11200
rect 4856 11160 4862 11172
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 5994 11200 6000 11212
rect 5955 11172 6000 11200
rect 4985 11163 5043 11169
rect 4709 11135 4767 11141
rect 4709 11101 4721 11135
rect 4755 11101 4767 11135
rect 4709 11095 4767 11101
rect 5000 11064 5028 11163
rect 5994 11160 6000 11172
rect 6052 11160 6058 11212
rect 6748 11132 6776 11228
rect 7745 11203 7803 11209
rect 7745 11169 7757 11203
rect 7791 11200 7803 11203
rect 8294 11200 8300 11212
rect 7791 11172 8300 11200
rect 7791 11169 7803 11172
rect 7745 11163 7803 11169
rect 8294 11160 8300 11172
rect 8352 11200 8358 11212
rect 9398 11200 9404 11212
rect 8352 11172 9404 11200
rect 8352 11160 8358 11172
rect 9398 11160 9404 11172
rect 9456 11160 9462 11212
rect 9508 11209 9536 11240
rect 13265 11237 13277 11271
rect 13311 11237 13323 11271
rect 13265 11231 13323 11237
rect 9493 11203 9551 11209
rect 9493 11169 9505 11203
rect 9539 11169 9551 11203
rect 13280 11200 13308 11231
rect 13446 11200 13452 11212
rect 13280 11172 13452 11200
rect 9493 11163 9551 11169
rect 13446 11160 13452 11172
rect 13504 11200 13510 11212
rect 14185 11203 14243 11209
rect 14185 11200 14197 11203
rect 13504 11172 14197 11200
rect 13504 11160 13510 11172
rect 14185 11169 14197 11172
rect 14231 11169 14243 11203
rect 14185 11163 14243 11169
rect 14369 11203 14427 11209
rect 14369 11169 14381 11203
rect 14415 11200 14427 11203
rect 15120 11200 15148 11296
rect 17037 11271 17095 11277
rect 17037 11237 17049 11271
rect 17083 11237 17095 11271
rect 17037 11231 17095 11237
rect 14415 11172 15148 11200
rect 17052 11200 17080 11231
rect 17497 11203 17555 11209
rect 17497 11200 17509 11203
rect 17052 11172 17509 11200
rect 14415 11169 14427 11172
rect 14369 11163 14427 11169
rect 17497 11169 17509 11172
rect 17543 11200 17555 11203
rect 17678 11200 17684 11212
rect 17543 11172 17684 11200
rect 17543 11169 17555 11172
rect 17497 11163 17555 11169
rect 17678 11160 17684 11172
rect 17736 11160 17742 11212
rect 8205 11135 8263 11141
rect 6748 11104 8064 11132
rect 4356 11036 5028 11064
rect 5721 11067 5779 11073
rect 5721 11033 5733 11067
rect 5767 11064 5779 11067
rect 5994 11064 6000 11076
rect 5767 11036 6000 11064
rect 5767 11033 5779 11036
rect 5721 11027 5779 11033
rect 5994 11024 6000 11036
rect 6052 11024 6058 11076
rect 7374 11064 7380 11076
rect 6104 11036 7380 11064
rect 2038 10996 2044 11008
rect 1999 10968 2044 10996
rect 2038 10956 2044 10968
rect 2096 10956 2102 11008
rect 2406 10996 2412 11008
rect 2367 10968 2412 10996
rect 2406 10956 2412 10968
rect 2464 10956 2470 11008
rect 3050 10996 3056 11008
rect 3011 10968 3056 10996
rect 3050 10956 3056 10968
rect 3108 10956 3114 11008
rect 5813 10999 5871 11005
rect 5813 10965 5825 10999
rect 5859 10996 5871 10999
rect 6104 10996 6132 11036
rect 7374 11024 7380 11036
rect 7432 11024 7438 11076
rect 7500 11067 7558 11073
rect 7500 11033 7512 11067
rect 7546 11064 7558 11067
rect 7926 11064 7932 11076
rect 7546 11036 7932 11064
rect 7546 11033 7558 11036
rect 7500 11027 7558 11033
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 8036 11064 8064 11104
rect 8205 11101 8217 11135
rect 8251 11132 8263 11135
rect 9122 11132 9128 11144
rect 8251 11104 9128 11132
rect 8251 11101 8263 11104
rect 8205 11095 8263 11101
rect 9122 11092 9128 11104
rect 9180 11092 9186 11144
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9416 11132 9444 11160
rect 10137 11135 10195 11141
rect 10137 11132 10149 11135
rect 9416 11104 10149 11132
rect 9309 11095 9367 11101
rect 10137 11101 10149 11104
rect 10183 11101 10195 11135
rect 11882 11132 11888 11144
rect 11843 11104 11888 11132
rect 10137 11095 10195 11101
rect 8036 11036 8432 11064
rect 5859 10968 6132 10996
rect 8404 10996 8432 11036
rect 8478 11024 8484 11076
rect 8536 11064 8542 11076
rect 9324 11064 9352 11095
rect 11882 11092 11888 11104
rect 11940 11092 11946 11144
rect 12152 11135 12210 11141
rect 12152 11101 12164 11135
rect 12198 11132 12210 11135
rect 13814 11132 13820 11144
rect 12198 11104 13820 11132
rect 12198 11101 12210 11104
rect 12152 11095 12210 11101
rect 13814 11092 13820 11104
rect 13872 11092 13878 11144
rect 14458 11132 14464 11144
rect 14419 11104 14464 11132
rect 14458 11092 14464 11104
rect 14516 11092 14522 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 16942 11132 16948 11144
rect 15703 11104 16948 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 16942 11092 16948 11104
rect 17000 11092 17006 11144
rect 8536 11036 8581 11064
rect 8680 11036 9352 11064
rect 9401 11067 9459 11073
rect 8536 11024 8542 11036
rect 8680 10996 8708 11036
rect 9401 11033 9413 11067
rect 9447 11064 9459 11067
rect 9490 11064 9496 11076
rect 9447 11036 9496 11064
rect 9447 11033 9459 11036
rect 9401 11027 9459 11033
rect 9490 11024 9496 11036
rect 9548 11024 9554 11076
rect 9582 11024 9588 11076
rect 9640 11064 9646 11076
rect 10382 11067 10440 11073
rect 10382 11064 10394 11067
rect 9640 11036 10394 11064
rect 9640 11024 9646 11036
rect 10382 11033 10394 11036
rect 10428 11033 10440 11067
rect 10382 11027 10440 11033
rect 13725 11067 13783 11073
rect 13725 11033 13737 11067
rect 13771 11064 13783 11067
rect 14918 11064 14924 11076
rect 13771 11036 14924 11064
rect 13771 11033 13783 11036
rect 13725 11027 13783 11033
rect 14918 11024 14924 11036
rect 14976 11024 14982 11076
rect 15924 11067 15982 11073
rect 15924 11033 15936 11067
rect 15970 11064 15982 11067
rect 17494 11064 17500 11076
rect 15970 11036 17500 11064
rect 15970 11033 15982 11036
rect 15924 11027 15982 11033
rect 17494 11024 17500 11036
rect 17552 11024 17558 11076
rect 17681 11067 17739 11073
rect 17681 11033 17693 11067
rect 17727 11064 17739 11067
rect 18325 11067 18383 11073
rect 18325 11064 18337 11067
rect 17727 11036 18337 11064
rect 17727 11033 17739 11036
rect 17681 11027 17739 11033
rect 18325 11033 18337 11036
rect 18371 11033 18383 11067
rect 18325 11027 18383 11033
rect 8404 10968 8708 10996
rect 11517 10999 11575 11005
rect 5859 10965 5871 10968
rect 5813 10959 5871 10965
rect 11517 10965 11529 10999
rect 11563 10996 11575 10999
rect 11698 10996 11704 11008
rect 11563 10968 11704 10996
rect 11563 10965 11575 10968
rect 11517 10959 11575 10965
rect 11698 10956 11704 10968
rect 11756 10956 11762 11008
rect 14826 10996 14832 11008
rect 14787 10968 14832 10996
rect 14826 10956 14832 10968
rect 14884 10956 14890 11008
rect 17586 10996 17592 11008
rect 17547 10968 17592 10996
rect 17586 10956 17592 10968
rect 17644 10956 17650 11008
rect 1104 10906 21896 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21896 10906
rect 1104 10832 21896 10854
rect 1673 10795 1731 10801
rect 1673 10761 1685 10795
rect 1719 10792 1731 10795
rect 2038 10792 2044 10804
rect 1719 10764 2044 10792
rect 1719 10761 1731 10764
rect 1673 10755 1731 10761
rect 2038 10752 2044 10764
rect 2096 10752 2102 10804
rect 2685 10795 2743 10801
rect 2685 10761 2697 10795
rect 2731 10792 2743 10795
rect 3234 10792 3240 10804
rect 2731 10764 3240 10792
rect 2731 10761 2743 10764
rect 2685 10755 2743 10761
rect 2038 10656 2044 10668
rect 1999 10628 2044 10656
rect 2038 10616 2044 10628
rect 2096 10616 2102 10668
rect 2133 10659 2191 10665
rect 2133 10625 2145 10659
rect 2179 10656 2191 10659
rect 2958 10656 2964 10668
rect 2179 10628 2964 10656
rect 2179 10625 2191 10628
rect 2133 10619 2191 10625
rect 2958 10616 2964 10628
rect 3016 10616 3022 10668
rect 2317 10591 2375 10597
rect 2317 10557 2329 10591
rect 2363 10588 2375 10591
rect 2866 10588 2872 10600
rect 2363 10560 2872 10588
rect 2363 10557 2375 10560
rect 2317 10551 2375 10557
rect 2866 10548 2872 10560
rect 2924 10588 2930 10600
rect 3068 10588 3096 10764
rect 3234 10752 3240 10764
rect 3292 10752 3298 10804
rect 4246 10752 4252 10804
rect 4304 10792 4310 10804
rect 4341 10795 4399 10801
rect 4341 10792 4353 10795
rect 4304 10764 4353 10792
rect 4304 10752 4310 10764
rect 4341 10761 4353 10764
rect 4387 10761 4399 10795
rect 4341 10755 4399 10761
rect 4522 10752 4528 10804
rect 4580 10792 4586 10804
rect 4801 10795 4859 10801
rect 4801 10792 4813 10795
rect 4580 10764 4813 10792
rect 4580 10752 4586 10764
rect 4801 10761 4813 10764
rect 4847 10761 4859 10795
rect 5350 10792 5356 10804
rect 5311 10764 5356 10792
rect 4801 10755 4859 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 5994 10752 6000 10804
rect 6052 10792 6058 10804
rect 6365 10795 6423 10801
rect 6365 10792 6377 10795
rect 6052 10764 6377 10792
rect 6052 10752 6058 10764
rect 6365 10761 6377 10764
rect 6411 10761 6423 10795
rect 6365 10755 6423 10761
rect 7561 10795 7619 10801
rect 7561 10761 7573 10795
rect 7607 10792 7619 10795
rect 8110 10792 8116 10804
rect 7607 10764 8116 10792
rect 7607 10761 7619 10764
rect 7561 10755 7619 10761
rect 8110 10752 8116 10764
rect 8168 10752 8174 10804
rect 10229 10795 10287 10801
rect 10229 10761 10241 10795
rect 10275 10792 10287 10795
rect 10410 10792 10416 10804
rect 10275 10764 10416 10792
rect 10275 10761 10287 10764
rect 10229 10755 10287 10761
rect 10410 10752 10416 10764
rect 10468 10792 10474 10804
rect 11793 10795 11851 10801
rect 11793 10792 11805 10795
rect 10468 10764 11805 10792
rect 10468 10752 10474 10764
rect 11793 10761 11805 10764
rect 11839 10761 11851 10795
rect 11793 10755 11851 10761
rect 12066 10752 12072 10804
rect 12124 10792 12130 10804
rect 14826 10792 14832 10804
rect 12124 10764 13308 10792
rect 14787 10764 14832 10792
rect 12124 10752 12130 10764
rect 3820 10727 3878 10733
rect 3820 10693 3832 10727
rect 3866 10724 3878 10727
rect 3970 10724 3976 10736
rect 3866 10696 3976 10724
rect 3866 10693 3878 10696
rect 3820 10687 3878 10693
rect 3970 10684 3976 10696
rect 4028 10684 4034 10736
rect 5718 10724 5724 10736
rect 4080 10696 5724 10724
rect 4080 10668 4108 10696
rect 5718 10684 5724 10696
rect 5776 10684 5782 10736
rect 7006 10684 7012 10736
rect 7064 10724 7070 10736
rect 7837 10727 7895 10733
rect 7837 10724 7849 10727
rect 7064 10696 7849 10724
rect 7064 10684 7070 10696
rect 7837 10693 7849 10696
rect 7883 10724 7895 10727
rect 11238 10724 11244 10736
rect 7883 10696 11244 10724
rect 7883 10693 7895 10696
rect 7837 10687 7895 10693
rect 11238 10684 11244 10696
rect 11296 10684 11302 10736
rect 12618 10724 12624 10736
rect 12579 10696 12624 10724
rect 12618 10684 12624 10696
rect 12676 10684 12682 10736
rect 12802 10684 12808 10736
rect 12860 10724 12866 10736
rect 13142 10727 13200 10733
rect 13142 10724 13154 10727
rect 12860 10696 13154 10724
rect 12860 10684 12866 10696
rect 13142 10693 13154 10696
rect 13188 10693 13200 10727
rect 13280 10724 13308 10764
rect 14826 10752 14832 10764
rect 14884 10752 14890 10804
rect 14918 10752 14924 10804
rect 14976 10792 14982 10804
rect 14976 10764 15021 10792
rect 14976 10752 14982 10764
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15841 10795 15899 10801
rect 15841 10792 15853 10795
rect 15620 10764 15853 10792
rect 15620 10752 15626 10764
rect 15841 10761 15853 10764
rect 15887 10761 15899 10795
rect 15841 10755 15899 10761
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 17586 10792 17592 10804
rect 16347 10764 17592 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 17586 10752 17592 10764
rect 17644 10752 17650 10804
rect 13280 10696 15332 10724
rect 13142 10687 13200 10693
rect 4062 10656 4068 10668
rect 3975 10628 4068 10656
rect 4062 10616 4068 10628
rect 4120 10616 4126 10668
rect 4709 10659 4767 10665
rect 4709 10625 4721 10659
rect 4755 10656 4767 10659
rect 4798 10656 4804 10668
rect 4755 10628 4804 10656
rect 4755 10625 4767 10628
rect 4709 10619 4767 10625
rect 4798 10616 4804 10628
rect 4856 10656 4862 10668
rect 5442 10656 5448 10668
rect 4856 10628 5448 10656
rect 4856 10616 4862 10628
rect 5442 10616 5448 10628
rect 5500 10616 5506 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5960 10628 6009 10656
rect 5960 10616 5966 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10656 7251 10659
rect 8386 10656 8392 10668
rect 7239 10628 8392 10656
rect 7239 10625 7251 10628
rect 7193 10619 7251 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 11149 10659 11207 10665
rect 11149 10625 11161 10659
rect 11195 10625 11207 10659
rect 11149 10619 11207 10625
rect 11885 10659 11943 10665
rect 11885 10625 11897 10659
rect 11931 10625 11943 10659
rect 11885 10619 11943 10625
rect 2924 10560 3096 10588
rect 4985 10591 5043 10597
rect 2924 10548 2930 10560
rect 4985 10557 4997 10591
rect 5031 10588 5043 10591
rect 5074 10588 5080 10600
rect 5031 10560 5080 10588
rect 5031 10557 5043 10560
rect 4985 10551 5043 10557
rect 5074 10548 5080 10560
rect 5132 10548 5138 10600
rect 7009 10591 7067 10597
rect 7009 10557 7021 10591
rect 7055 10557 7067 10591
rect 7009 10551 7067 10557
rect 7101 10591 7159 10597
rect 7101 10557 7113 10591
rect 7147 10588 7159 10591
rect 7374 10588 7380 10600
rect 7147 10560 7380 10588
rect 7147 10557 7159 10560
rect 7101 10551 7159 10557
rect 7024 10520 7052 10551
rect 7374 10548 7380 10560
rect 7432 10548 7438 10600
rect 11164 10588 11192 10619
rect 11698 10588 11704 10600
rect 11164 10560 11704 10588
rect 11698 10548 11704 10560
rect 11756 10548 11762 10600
rect 7834 10520 7840 10532
rect 7024 10492 7840 10520
rect 7834 10480 7840 10492
rect 7892 10480 7898 10532
rect 11900 10520 11928 10619
rect 12897 10591 12955 10597
rect 12897 10557 12909 10591
rect 12943 10557 12955 10591
rect 12897 10551 12955 10557
rect 14737 10591 14795 10597
rect 14737 10557 14749 10591
rect 14783 10588 14795 10591
rect 14918 10588 14924 10600
rect 14783 10560 14924 10588
rect 14783 10557 14795 10560
rect 14737 10551 14795 10557
rect 12912 10520 12940 10551
rect 14918 10548 14924 10560
rect 14976 10548 14982 10600
rect 7944 10492 11928 10520
rect 11992 10492 12940 10520
rect 15304 10520 15332 10696
rect 15764 10696 16574 10724
rect 15764 10597 15792 10696
rect 15930 10656 15936 10668
rect 15891 10628 15936 10656
rect 15930 10616 15936 10628
rect 15988 10616 15994 10668
rect 16546 10656 16574 10696
rect 16942 10684 16948 10736
rect 17000 10724 17006 10736
rect 17000 10696 18092 10724
rect 17000 10684 17006 10696
rect 17310 10656 17316 10668
rect 16546 10628 17316 10656
rect 17310 10616 17316 10628
rect 17368 10616 17374 10668
rect 17793 10659 17851 10665
rect 17793 10625 17805 10659
rect 17839 10656 17851 10659
rect 17954 10656 17960 10668
rect 17839 10628 17960 10656
rect 17839 10625 17851 10628
rect 17793 10619 17851 10625
rect 17954 10616 17960 10628
rect 18012 10616 18018 10668
rect 18064 10665 18092 10696
rect 18049 10659 18107 10665
rect 18049 10625 18061 10659
rect 18095 10625 18107 10659
rect 18049 10619 18107 10625
rect 15749 10591 15807 10597
rect 15749 10557 15761 10591
rect 15795 10557 15807 10591
rect 15749 10551 15807 10557
rect 16669 10523 16727 10529
rect 16669 10520 16681 10523
rect 15304 10492 16681 10520
rect 2682 10412 2688 10464
rect 2740 10452 2746 10464
rect 5994 10452 6000 10464
rect 2740 10424 6000 10452
rect 2740 10412 2746 10424
rect 5994 10412 6000 10424
rect 6052 10412 6058 10464
rect 6914 10412 6920 10464
rect 6972 10452 6978 10464
rect 7944 10452 7972 10492
rect 6972 10424 7972 10452
rect 9309 10455 9367 10461
rect 6972 10412 6978 10424
rect 9309 10421 9321 10455
rect 9355 10452 9367 10455
rect 9398 10452 9404 10464
rect 9355 10424 9404 10452
rect 9355 10421 9367 10424
rect 9309 10415 9367 10421
rect 9398 10412 9404 10424
rect 9456 10412 9462 10464
rect 10505 10455 10563 10461
rect 10505 10421 10517 10455
rect 10551 10452 10563 10455
rect 11790 10452 11796 10464
rect 10551 10424 11796 10452
rect 10551 10421 10563 10424
rect 10505 10415 10563 10421
rect 11790 10412 11796 10424
rect 11848 10412 11854 10464
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 11992 10452 12020 10492
rect 16669 10489 16681 10492
rect 16715 10489 16727 10523
rect 16669 10483 16727 10489
rect 12250 10452 12256 10464
rect 11940 10424 12020 10452
rect 12211 10424 12256 10452
rect 11940 10412 11946 10424
rect 12250 10412 12256 10424
rect 12308 10412 12314 10464
rect 14277 10455 14335 10461
rect 14277 10421 14289 10455
rect 14323 10452 14335 10455
rect 14918 10452 14924 10464
rect 14323 10424 14924 10452
rect 14323 10421 14335 10424
rect 14277 10415 14335 10421
rect 14918 10412 14924 10424
rect 14976 10412 14982 10464
rect 15289 10455 15347 10461
rect 15289 10421 15301 10455
rect 15335 10452 15347 10455
rect 17770 10452 17776 10464
rect 15335 10424 17776 10452
rect 15335 10421 15347 10424
rect 15289 10415 15347 10421
rect 17770 10412 17776 10424
rect 17828 10412 17834 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1854 10248 1860 10260
rect 1815 10220 1860 10248
rect 1854 10208 1860 10220
rect 1912 10208 1918 10260
rect 3050 10208 3056 10260
rect 3108 10248 3114 10260
rect 3789 10251 3847 10257
rect 3789 10248 3801 10251
rect 3108 10220 3801 10248
rect 3108 10208 3114 10220
rect 3789 10217 3801 10220
rect 3835 10217 3847 10251
rect 3789 10211 3847 10217
rect 4154 10208 4160 10260
rect 4212 10248 4218 10260
rect 4801 10251 4859 10257
rect 4801 10248 4813 10251
rect 4212 10220 4813 10248
rect 4212 10208 4218 10220
rect 4801 10217 4813 10220
rect 4847 10217 4859 10251
rect 5718 10248 5724 10260
rect 5679 10220 5724 10248
rect 4801 10211 4859 10217
rect 5718 10208 5724 10220
rect 5776 10208 5782 10260
rect 7469 10251 7527 10257
rect 7469 10217 7481 10251
rect 7515 10248 7527 10251
rect 7558 10248 7564 10260
rect 7515 10220 7564 10248
rect 7515 10217 7527 10220
rect 7469 10211 7527 10217
rect 7558 10208 7564 10220
rect 7616 10208 7622 10260
rect 9122 10208 9128 10260
rect 9180 10248 9186 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9180 10220 9965 10248
rect 9180 10208 9186 10220
rect 9953 10217 9965 10220
rect 9999 10217 10011 10251
rect 9953 10211 10011 10217
rect 10873 10251 10931 10257
rect 10873 10217 10885 10251
rect 10919 10248 10931 10251
rect 11882 10248 11888 10260
rect 10919 10220 11888 10248
rect 10919 10217 10931 10220
rect 10873 10211 10931 10217
rect 11882 10208 11888 10220
rect 11940 10208 11946 10260
rect 13078 10208 13084 10260
rect 13136 10248 13142 10260
rect 13173 10251 13231 10257
rect 13173 10248 13185 10251
rect 13136 10220 13185 10248
rect 13136 10208 13142 10220
rect 13173 10217 13185 10220
rect 13219 10217 13231 10251
rect 15378 10248 15384 10260
rect 15339 10220 15384 10248
rect 13173 10211 13231 10217
rect 15378 10208 15384 10220
rect 15436 10208 15442 10260
rect 16942 10248 16948 10260
rect 16903 10220 16948 10248
rect 16942 10208 16948 10220
rect 17000 10208 17006 10260
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18325 10251 18383 10257
rect 18325 10248 18337 10251
rect 18012 10220 18337 10248
rect 18012 10208 18018 10220
rect 18325 10217 18337 10220
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 1397 10183 1455 10189
rect 1397 10149 1409 10183
rect 1443 10180 1455 10183
rect 1946 10180 1952 10192
rect 1443 10152 1952 10180
rect 1443 10149 1455 10152
rect 1397 10143 1455 10149
rect 1946 10140 1952 10152
rect 2004 10140 2010 10192
rect 3602 10140 3608 10192
rect 3660 10180 3666 10192
rect 3970 10180 3976 10192
rect 3660 10152 3976 10180
rect 3660 10140 3666 10152
rect 3970 10140 3976 10152
rect 4028 10180 4034 10192
rect 4028 10152 4476 10180
rect 4028 10140 4034 10152
rect 3234 10072 3240 10124
rect 3292 10112 3298 10124
rect 4062 10112 4068 10124
rect 3292 10084 4068 10112
rect 3292 10072 3298 10084
rect 4062 10072 4068 10084
rect 4120 10072 4126 10124
rect 4448 10121 4476 10152
rect 6730 10140 6736 10192
rect 6788 10180 6794 10192
rect 8941 10183 8999 10189
rect 8941 10180 8953 10183
rect 6788 10152 8953 10180
rect 6788 10140 6794 10152
rect 8941 10149 8953 10152
rect 8987 10149 8999 10183
rect 12066 10180 12072 10192
rect 8941 10143 8999 10149
rect 9048 10152 12072 10180
rect 4433 10115 4491 10121
rect 4433 10081 4445 10115
rect 4479 10112 4491 10115
rect 5074 10112 5080 10124
rect 4479 10084 5080 10112
rect 4479 10081 4491 10084
rect 4433 10075 4491 10081
rect 5074 10072 5080 10084
rect 5132 10112 5138 10124
rect 9048 10112 9076 10152
rect 12066 10140 12072 10152
rect 12124 10140 12130 10192
rect 12250 10140 12256 10192
rect 12308 10180 12314 10192
rect 12308 10152 12756 10180
rect 12308 10140 12314 10152
rect 9490 10112 9496 10124
rect 5132 10084 9076 10112
rect 9451 10084 9496 10112
rect 5132 10072 5138 10084
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 12618 10112 12624 10124
rect 12579 10084 12624 10112
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 12728 10121 12756 10152
rect 12713 10115 12771 10121
rect 12713 10081 12725 10115
rect 12759 10081 12771 10115
rect 12713 10075 12771 10081
rect 1578 10044 1584 10056
rect 1539 10016 1584 10044
rect 1578 10004 1584 10016
rect 1636 10004 1642 10056
rect 4982 10044 4988 10056
rect 4943 10016 4988 10044
rect 4982 10004 4988 10016
rect 5040 10004 5046 10056
rect 7006 10044 7012 10056
rect 6967 10016 7012 10044
rect 7006 10004 7012 10016
rect 7064 10004 7070 10056
rect 8018 10004 8024 10056
rect 8076 10044 8082 10056
rect 8113 10047 8171 10053
rect 8113 10044 8125 10047
rect 8076 10016 8125 10044
rect 8076 10004 8082 10016
rect 8113 10013 8125 10016
rect 8159 10013 8171 10047
rect 8113 10007 8171 10013
rect 8478 10004 8484 10056
rect 8536 10044 8542 10056
rect 9306 10044 9312 10056
rect 8536 10016 9312 10044
rect 8536 10004 8542 10016
rect 9306 10004 9312 10016
rect 9364 10004 9370 10056
rect 11238 10004 11244 10056
rect 11296 10044 11302 10056
rect 12161 10047 12219 10053
rect 12161 10044 12173 10047
rect 11296 10016 12173 10044
rect 11296 10004 11302 10016
rect 12161 10013 12173 10016
rect 12207 10013 12219 10047
rect 12161 10007 12219 10013
rect 12805 10047 12863 10053
rect 12805 10013 12817 10047
rect 12851 10044 12863 10047
rect 13170 10044 13176 10056
rect 12851 10016 13176 10044
rect 12851 10013 12863 10016
rect 12805 10007 12863 10013
rect 2866 9936 2872 9988
rect 2924 9976 2930 9988
rect 2970 9979 3028 9985
rect 2970 9976 2982 9979
rect 2924 9948 2982 9976
rect 2924 9936 2930 9948
rect 2970 9945 2982 9948
rect 3016 9945 3028 9979
rect 2970 9939 3028 9945
rect 4157 9979 4215 9985
rect 4157 9945 4169 9979
rect 4203 9976 4215 9979
rect 8496 9976 8524 10004
rect 4203 9948 8524 9976
rect 12176 9976 12204 10007
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 14734 10044 14740 10056
rect 14695 10016 14740 10044
rect 14734 10004 14740 10016
rect 14792 10004 14798 10056
rect 17678 10044 17684 10056
rect 17639 10016 17684 10044
rect 17678 10004 17684 10016
rect 17736 10004 17742 10056
rect 15657 9979 15715 9985
rect 15657 9976 15669 9979
rect 12176 9948 15669 9976
rect 4203 9945 4215 9948
rect 4157 9939 4215 9945
rect 15657 9945 15669 9948
rect 15703 9945 15715 9979
rect 15657 9939 15715 9945
rect 2590 9868 2596 9920
rect 2648 9908 2654 9920
rect 3786 9908 3792 9920
rect 2648 9880 3792 9908
rect 2648 9868 2654 9880
rect 3786 9868 3792 9880
rect 3844 9868 3850 9920
rect 4249 9911 4307 9917
rect 4249 9877 4261 9911
rect 4295 9908 4307 9911
rect 5258 9908 5264 9920
rect 4295 9880 5264 9908
rect 4295 9877 4307 9880
rect 4249 9871 4307 9877
rect 5258 9868 5264 9880
rect 5316 9868 5322 9920
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 8389 9911 8447 9917
rect 8389 9908 8401 9911
rect 5684 9880 8401 9908
rect 5684 9868 5690 9880
rect 8389 9877 8401 9880
rect 8435 9877 8447 9911
rect 9306 9908 9312 9920
rect 9267 9880 9312 9908
rect 8389 9871 8447 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 9401 9911 9459 9917
rect 9401 9877 9413 9911
rect 9447 9908 9459 9911
rect 9674 9908 9680 9920
rect 9447 9880 9680 9908
rect 9447 9877 9459 9880
rect 9401 9871 9459 9877
rect 9674 9868 9680 9880
rect 9732 9868 9738 9920
rect 1104 9818 21896 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21896 9818
rect 1104 9744 21896 9766
rect 2958 9704 2964 9716
rect 2919 9676 2964 9704
rect 2958 9664 2964 9676
rect 3016 9664 3022 9716
rect 4157 9707 4215 9713
rect 4157 9673 4169 9707
rect 4203 9673 4215 9707
rect 4157 9667 4215 9673
rect 4062 9596 4068 9648
rect 4120 9636 4126 9648
rect 4172 9636 4200 9667
rect 4246 9664 4252 9716
rect 4304 9704 4310 9716
rect 4706 9704 4712 9716
rect 4304 9676 4712 9704
rect 4304 9664 4310 9676
rect 4706 9664 4712 9676
rect 4764 9664 4770 9716
rect 5718 9664 5724 9716
rect 5776 9704 5782 9716
rect 5776 9676 7144 9704
rect 5776 9664 5782 9676
rect 4120 9608 4200 9636
rect 4120 9596 4126 9608
rect 1486 9568 1492 9580
rect 1447 9540 1492 9568
rect 1486 9528 1492 9540
rect 1544 9528 1550 9580
rect 1854 9528 1860 9580
rect 1912 9568 1918 9580
rect 1949 9571 2007 9577
rect 1949 9568 1961 9571
rect 1912 9540 1961 9568
rect 1912 9528 1918 9540
rect 1949 9537 1961 9540
rect 1995 9537 2007 9571
rect 3329 9571 3387 9577
rect 3329 9564 3341 9571
rect 3375 9564 3387 9571
rect 1949 9531 2007 9537
rect 3326 9512 3332 9564
rect 3384 9512 3390 9564
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 3973 9571 4031 9577
rect 3973 9568 3985 9571
rect 3844 9540 3985 9568
rect 3844 9528 3850 9540
rect 3973 9537 3985 9540
rect 4019 9537 4031 9571
rect 3973 9531 4031 9537
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 3421 9503 3479 9509
rect 3421 9469 3433 9503
rect 3467 9469 3479 9503
rect 3602 9500 3608 9512
rect 3563 9472 3608 9500
rect 3421 9463 3479 9469
rect 1670 9432 1676 9444
rect 1631 9404 1676 9432
rect 1670 9392 1676 9404
rect 1728 9392 1734 9444
rect 2866 9392 2872 9444
rect 2924 9432 2930 9444
rect 3050 9432 3056 9444
rect 2924 9404 3056 9432
rect 2924 9392 2930 9404
rect 3050 9392 3056 9404
rect 3108 9392 3114 9444
rect 3436 9432 3464 9463
rect 3602 9460 3608 9472
rect 3660 9460 3666 9512
rect 4154 9432 4160 9444
rect 3436 9404 4160 9432
rect 4154 9392 4160 9404
rect 4212 9392 4218 9444
rect 2590 9364 2596 9376
rect 2551 9336 2596 9364
rect 2590 9324 2596 9336
rect 2648 9324 2654 9376
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 4448 9364 4476 9531
rect 5074 9528 5080 9580
rect 5132 9568 5138 9580
rect 5261 9571 5319 9577
rect 5261 9568 5273 9571
rect 5132 9540 5273 9568
rect 5132 9528 5138 9540
rect 5261 9537 5273 9540
rect 5307 9537 5319 9571
rect 5261 9531 5319 9537
rect 4614 9432 4620 9444
rect 4575 9404 4620 9432
rect 4614 9392 4620 9404
rect 4672 9392 4678 9444
rect 5276 9432 5304 9531
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 6641 9571 6699 9577
rect 5408 9540 5453 9568
rect 5408 9528 5414 9540
rect 6641 9537 6653 9571
rect 6687 9568 6699 9571
rect 6822 9568 6828 9580
rect 6687 9540 6828 9568
rect 6687 9537 6699 9540
rect 6641 9531 6699 9537
rect 6822 9528 6828 9540
rect 6880 9528 6886 9580
rect 7116 9577 7144 9676
rect 8386 9664 8392 9716
rect 8444 9704 8450 9716
rect 8662 9704 8668 9716
rect 8444 9676 8668 9704
rect 8444 9664 8450 9676
rect 8662 9664 8668 9676
rect 8720 9664 8726 9716
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12897 9707 12955 9713
rect 12897 9704 12909 9707
rect 12676 9676 12909 9704
rect 12676 9664 12682 9676
rect 12897 9673 12909 9676
rect 12943 9673 12955 9707
rect 12897 9667 12955 9673
rect 15289 9707 15347 9713
rect 15289 9673 15301 9707
rect 15335 9704 15347 9707
rect 15562 9704 15568 9716
rect 15335 9676 15568 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 8294 9636 8300 9648
rect 7208 9608 8300 9636
rect 7101 9571 7159 9577
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7101 9531 7159 9537
rect 5442 9500 5448 9512
rect 5403 9472 5448 9500
rect 5442 9460 5448 9472
rect 5500 9460 5506 9512
rect 7208 9500 7236 9608
rect 8294 9596 8300 9608
rect 8352 9596 8358 9648
rect 9398 9636 9404 9648
rect 8956 9608 9404 9636
rect 7368 9571 7426 9577
rect 7368 9537 7380 9571
rect 7414 9568 7426 9571
rect 8662 9568 8668 9580
rect 7414 9540 8668 9568
rect 7414 9537 7426 9540
rect 7368 9531 7426 9537
rect 8662 9528 8668 9540
rect 8720 9528 8726 9580
rect 8956 9577 8984 9608
rect 9398 9596 9404 9608
rect 9456 9596 9462 9648
rect 9582 9596 9588 9648
rect 9640 9636 9646 9648
rect 11790 9645 11796 9648
rect 10597 9639 10655 9645
rect 10597 9636 10609 9639
rect 9640 9608 10609 9636
rect 9640 9596 9646 9608
rect 10597 9605 10609 9608
rect 10643 9605 10655 9639
rect 11784 9636 11796 9645
rect 11751 9608 11796 9636
rect 10597 9599 10655 9605
rect 11784 9599 11796 9608
rect 11790 9596 11796 9599
rect 11848 9596 11854 9648
rect 9214 9577 9220 9580
rect 8941 9571 8999 9577
rect 8941 9537 8953 9571
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9208 9531 9220 9577
rect 9272 9568 9278 9580
rect 9416 9568 9444 9596
rect 11517 9571 11575 9577
rect 11517 9568 11529 9571
rect 9272 9540 9308 9568
rect 9416 9540 11529 9568
rect 9214 9528 9220 9531
rect 9272 9528 9278 9540
rect 11517 9537 11529 9540
rect 11563 9537 11575 9571
rect 12912 9568 12940 9667
rect 15562 9664 15568 9676
rect 15620 9664 15626 9716
rect 13814 9636 13820 9648
rect 13775 9608 13820 9636
rect 13814 9596 13820 9608
rect 13872 9596 13878 9648
rect 14274 9636 14280 9648
rect 14235 9608 14280 9636
rect 14274 9596 14280 9608
rect 14332 9596 14338 9648
rect 13173 9571 13231 9577
rect 13173 9568 13185 9571
rect 12912 9540 13185 9568
rect 11517 9531 11575 9537
rect 13173 9537 13185 9540
rect 13219 9537 13231 9571
rect 14918 9568 14924 9580
rect 14879 9540 14924 9568
rect 13173 9531 13231 9537
rect 14918 9528 14924 9540
rect 14976 9528 14982 9580
rect 5920 9472 7236 9500
rect 5920 9441 5948 9472
rect 8294 9460 8300 9512
rect 8352 9500 8358 9512
rect 8478 9500 8484 9512
rect 8352 9472 8484 9500
rect 8352 9460 8358 9472
rect 8478 9460 8484 9472
rect 8536 9460 8542 9512
rect 5905 9435 5963 9441
rect 5905 9432 5917 9435
rect 5276 9404 5917 9432
rect 5905 9401 5917 9404
rect 5951 9401 5963 9435
rect 15565 9435 15623 9441
rect 15565 9432 15577 9435
rect 5905 9395 5963 9401
rect 14568 9404 15577 9432
rect 2832 9336 4476 9364
rect 2832 9324 2838 9336
rect 4706 9324 4712 9376
rect 4764 9364 4770 9376
rect 4893 9367 4951 9373
rect 4893 9364 4905 9367
rect 4764 9336 4905 9364
rect 4764 9324 4770 9336
rect 4893 9333 4905 9336
rect 4939 9333 4951 9367
rect 4893 9327 4951 9333
rect 6825 9367 6883 9373
rect 6825 9333 6837 9367
rect 6871 9364 6883 9367
rect 7742 9364 7748 9376
rect 6871 9336 7748 9364
rect 6871 9333 6883 9336
rect 6825 9327 6883 9333
rect 7742 9324 7748 9336
rect 7800 9324 7806 9376
rect 8478 9364 8484 9376
rect 8439 9336 8484 9364
rect 8478 9324 8484 9336
rect 8536 9324 8542 9376
rect 9582 9324 9588 9376
rect 9640 9364 9646 9376
rect 10321 9367 10379 9373
rect 10321 9364 10333 9367
rect 9640 9336 10333 9364
rect 9640 9324 9646 9336
rect 10321 9333 10333 9336
rect 10367 9333 10379 9367
rect 10962 9364 10968 9376
rect 10923 9336 10968 9364
rect 10321 9327 10379 9333
rect 10962 9324 10968 9336
rect 11020 9324 11026 9376
rect 11054 9324 11060 9376
rect 11112 9364 11118 9376
rect 14568 9364 14596 9404
rect 15565 9401 15577 9404
rect 15611 9432 15623 9435
rect 15930 9432 15936 9444
rect 15611 9404 15936 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 15930 9392 15936 9404
rect 15988 9392 15994 9444
rect 11112 9336 14596 9364
rect 11112 9324 11118 9336
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1302 9120 1308 9172
rect 1360 9160 1366 9172
rect 1360 9132 1440 9160
rect 1360 9120 1366 9132
rect 1412 8965 1440 9132
rect 1946 9120 1952 9172
rect 2004 9160 2010 9172
rect 4982 9160 4988 9172
rect 2004 9132 4988 9160
rect 2004 9120 2010 9132
rect 4982 9120 4988 9132
rect 5040 9120 5046 9172
rect 5442 9120 5448 9172
rect 5500 9120 5506 9172
rect 8021 9163 8079 9169
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 9306 9160 9312 9172
rect 8067 9132 9312 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 9306 9120 9312 9132
rect 9364 9120 9370 9172
rect 9674 9160 9680 9172
rect 9635 9132 9680 9160
rect 9674 9120 9680 9132
rect 9732 9120 9738 9172
rect 9766 9120 9772 9172
rect 9824 9160 9830 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 9824 9132 10609 9160
rect 9824 9120 9830 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 10965 9163 11023 9169
rect 10965 9129 10977 9163
rect 11011 9160 11023 9163
rect 17218 9160 17224 9172
rect 11011 9132 17224 9160
rect 11011 9129 11023 9132
rect 10965 9123 11023 9129
rect 3421 9095 3479 9101
rect 3421 9061 3433 9095
rect 3467 9061 3479 9095
rect 3421 9055 3479 9061
rect 3436 9024 3464 9055
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 4614 9092 4620 9104
rect 4212 9064 4620 9092
rect 4212 9052 4218 9064
rect 4614 9052 4620 9064
rect 4672 9092 4678 9104
rect 5166 9092 5172 9104
rect 4672 9064 5172 9092
rect 4672 9052 4678 9064
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5460 9092 5488 9120
rect 5276 9064 5488 9092
rect 3510 9024 3516 9036
rect 3423 8996 3516 9024
rect 3510 8984 3516 8996
rect 3568 9024 3574 9036
rect 4433 9027 4491 9033
rect 4433 9024 4445 9027
rect 3568 8996 4445 9024
rect 3568 8984 3574 8996
rect 4433 8993 4445 8996
rect 4479 9024 4491 9027
rect 5276 9024 5304 9064
rect 5810 9052 5816 9104
rect 5868 9092 5874 9104
rect 6273 9095 6331 9101
rect 6273 9092 6285 9095
rect 5868 9064 6285 9092
rect 5868 9052 5874 9064
rect 6273 9061 6285 9064
rect 6319 9061 6331 9095
rect 9490 9092 9496 9104
rect 6273 9055 6331 9061
rect 6564 9064 9496 9092
rect 4479 8996 5304 9024
rect 5445 9027 5503 9033
rect 4479 8993 4491 8996
rect 4433 8987 4491 8993
rect 5445 8993 5457 9027
rect 5491 9024 5503 9027
rect 6564 9024 6592 9064
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 6730 9024 6736 9036
rect 5491 8996 6592 9024
rect 6691 8996 6736 9024
rect 5491 8993 5503 8996
rect 5445 8987 5503 8993
rect 6730 8984 6736 8996
rect 6788 8984 6794 9036
rect 6825 9027 6883 9033
rect 6825 8993 6837 9027
rect 6871 8993 6883 9027
rect 6825 8987 6883 8993
rect 7469 9027 7527 9033
rect 7469 8993 7481 9027
rect 7515 9024 7527 9027
rect 8018 9024 8024 9036
rect 7515 8996 8024 9024
rect 7515 8993 7527 8996
rect 7469 8987 7527 8993
rect 1397 8959 1455 8965
rect 1397 8925 1409 8959
rect 1443 8956 1455 8959
rect 1854 8956 1860 8968
rect 1443 8928 1860 8956
rect 1443 8925 1455 8928
rect 1397 8919 1455 8925
rect 1854 8916 1860 8928
rect 1912 8916 1918 8968
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8956 2099 8959
rect 3234 8956 3240 8968
rect 2087 8928 3240 8956
rect 2087 8925 2099 8928
rect 2041 8919 2099 8925
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 4522 8916 4528 8968
rect 4580 8956 4586 8968
rect 4617 8959 4675 8965
rect 4617 8956 4629 8959
rect 4580 8928 4629 8956
rect 4580 8916 4586 8928
rect 4617 8925 4629 8928
rect 4663 8925 4675 8959
rect 5626 8956 5632 8968
rect 5587 8928 5632 8956
rect 4617 8919 4675 8925
rect 5626 8916 5632 8928
rect 5684 8916 5690 8968
rect 6840 8956 6868 8987
rect 8018 8984 8024 8996
rect 8076 9024 8082 9036
rect 9122 9024 9128 9036
rect 8076 8996 9128 9024
rect 8076 8984 8082 8996
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 9217 9027 9275 9033
rect 9217 8993 9229 9027
rect 9263 9024 9275 9027
rect 10980 9024 11008 9123
rect 17218 9120 17224 9132
rect 17276 9120 17282 9172
rect 9263 8996 11008 9024
rect 9263 8993 9275 8996
rect 9217 8987 9275 8993
rect 8478 8956 8484 8968
rect 6840 8928 8484 8956
rect 8478 8916 8484 8928
rect 8536 8956 8542 8968
rect 9953 8959 10011 8965
rect 9953 8956 9965 8959
rect 8536 8928 9965 8956
rect 8536 8916 8542 8928
rect 9953 8925 9965 8928
rect 9999 8925 10011 8959
rect 9953 8919 10011 8925
rect 2308 8891 2366 8897
rect 2308 8857 2320 8891
rect 2354 8888 2366 8891
rect 2590 8888 2596 8900
rect 2354 8860 2596 8888
rect 2354 8857 2366 8860
rect 2308 8851 2366 8857
rect 2590 8848 2596 8860
rect 2648 8848 2654 8900
rect 3789 8891 3847 8897
rect 3789 8888 3801 8891
rect 2746 8860 3801 8888
rect 1578 8820 1584 8832
rect 1539 8792 1584 8820
rect 1578 8780 1584 8792
rect 1636 8780 1642 8832
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 2746 8820 2774 8860
rect 3789 8857 3801 8860
rect 3835 8857 3847 8891
rect 6641 8891 6699 8897
rect 6641 8888 6653 8891
rect 3789 8851 3847 8857
rect 6012 8860 6653 8888
rect 2096 8792 2774 8820
rect 2096 8780 2102 8792
rect 2958 8780 2964 8832
rect 3016 8820 3022 8832
rect 4246 8820 4252 8832
rect 3016 8792 4252 8820
rect 3016 8780 3022 8792
rect 4246 8780 4252 8792
rect 4304 8780 4310 8832
rect 4430 8780 4436 8832
rect 4488 8820 4494 8832
rect 4525 8823 4583 8829
rect 4525 8820 4537 8823
rect 4488 8792 4537 8820
rect 4488 8780 4494 8792
rect 4525 8789 4537 8792
rect 4571 8789 4583 8823
rect 4982 8820 4988 8832
rect 4943 8792 4988 8820
rect 4525 8783 4583 8789
rect 4982 8780 4988 8792
rect 5040 8780 5046 8832
rect 5166 8780 5172 8832
rect 5224 8820 5230 8832
rect 5537 8823 5595 8829
rect 5537 8820 5549 8823
rect 5224 8792 5549 8820
rect 5224 8780 5230 8792
rect 5537 8789 5549 8792
rect 5583 8820 5595 8823
rect 5718 8820 5724 8832
rect 5583 8792 5724 8820
rect 5583 8789 5595 8792
rect 5537 8783 5595 8789
rect 5718 8780 5724 8792
rect 5776 8780 5782 8832
rect 6012 8829 6040 8860
rect 6641 8857 6653 8860
rect 6687 8857 6699 8891
rect 10962 8888 10968 8900
rect 6641 8851 6699 8857
rect 7668 8860 10968 8888
rect 7668 8832 7696 8860
rect 10962 8848 10968 8860
rect 11020 8848 11026 8900
rect 5997 8823 6055 8829
rect 5997 8789 6009 8823
rect 6043 8789 6055 8823
rect 5997 8783 6055 8789
rect 6546 8780 6552 8832
rect 6604 8820 6610 8832
rect 7561 8823 7619 8829
rect 7561 8820 7573 8823
rect 6604 8792 7573 8820
rect 6604 8780 6610 8792
rect 7561 8789 7573 8792
rect 7607 8789 7619 8823
rect 7561 8783 7619 8789
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8297 8823 8355 8829
rect 7708 8792 7753 8820
rect 7708 8780 7714 8792
rect 8297 8789 8309 8823
rect 8343 8820 8355 8823
rect 8754 8820 8760 8832
rect 8343 8792 8760 8820
rect 8343 8789 8355 8792
rect 8297 8783 8355 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9306 8820 9312 8832
rect 9267 8792 9312 8820
rect 9306 8780 9312 8792
rect 9364 8820 9370 8832
rect 11241 8823 11299 8829
rect 11241 8820 11253 8823
rect 9364 8792 11253 8820
rect 9364 8780 9370 8792
rect 11241 8789 11253 8792
rect 11287 8789 11299 8823
rect 11241 8783 11299 8789
rect 1104 8730 21896 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21896 8730
rect 1104 8656 21896 8678
rect 1397 8619 1455 8625
rect 1397 8585 1409 8619
rect 1443 8616 1455 8619
rect 1762 8616 1768 8628
rect 1443 8588 1768 8616
rect 1443 8585 1455 8588
rect 1397 8579 1455 8585
rect 1762 8576 1768 8588
rect 1820 8576 1826 8628
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 4890 8616 4896 8628
rect 4851 8588 4896 8616
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 7009 8619 7067 8625
rect 7009 8616 7021 8619
rect 5675 8588 7021 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 7009 8585 7021 8588
rect 7055 8585 7067 8619
rect 7009 8579 7067 8585
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 2682 8548 2688 8560
rect 1872 8520 2688 8548
rect 1578 8480 1584 8492
rect 1539 8452 1584 8480
rect 1578 8440 1584 8452
rect 1636 8440 1642 8492
rect 1872 8489 1900 8520
rect 2682 8508 2688 8520
rect 2740 8508 2746 8560
rect 4062 8548 4068 8560
rect 3252 8520 4068 8548
rect 3252 8492 3280 8520
rect 4062 8508 4068 8520
rect 4120 8508 4126 8560
rect 7392 8548 7420 8579
rect 8662 8576 8668 8628
rect 8720 8616 8726 8628
rect 9677 8619 9735 8625
rect 9677 8616 9689 8619
rect 8720 8588 9689 8616
rect 8720 8576 8726 8588
rect 9677 8585 9689 8588
rect 9723 8585 9735 8619
rect 9677 8579 9735 8585
rect 8754 8548 8760 8560
rect 7392 8520 8760 8548
rect 8754 8508 8760 8520
rect 8812 8508 8818 8560
rect 9490 8508 9496 8560
rect 9548 8548 9554 8560
rect 9548 8520 10364 8548
rect 9548 8508 9554 8520
rect 1857 8483 1915 8489
rect 1857 8449 1869 8483
rect 1903 8449 1915 8483
rect 2314 8480 2320 8492
rect 2275 8452 2320 8480
rect 1857 8443 1915 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2774 8440 2780 8492
rect 2832 8440 2838 8492
rect 2958 8440 2964 8492
rect 3016 8480 3022 8492
rect 3234 8480 3240 8492
rect 3016 8452 3061 8480
rect 3195 8452 3240 8480
rect 3016 8440 3022 8452
rect 3234 8440 3240 8452
rect 3292 8440 3298 8492
rect 3510 8489 3516 8492
rect 3504 8480 3516 8489
rect 3471 8452 3516 8480
rect 3504 8443 3516 8452
rect 3510 8440 3516 8443
rect 3568 8440 3574 8492
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 6454 8480 6460 8492
rect 4488 8452 6460 8480
rect 4488 8440 4494 8452
rect 6454 8440 6460 8452
rect 6512 8440 6518 8492
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8480 7527 8483
rect 8386 8480 8392 8492
rect 7515 8452 8392 8480
rect 7515 8449 7527 8452
rect 7469 8443 7527 8449
rect 2792 8412 2820 8440
rect 5718 8412 5724 8424
rect 2516 8384 2820 8412
rect 5679 8384 5724 8412
rect 2516 8353 2544 8384
rect 5718 8372 5724 8384
rect 5776 8372 5782 8424
rect 5902 8412 5908 8424
rect 5863 8384 5908 8412
rect 5902 8372 5908 8384
rect 5960 8372 5966 8424
rect 6086 8372 6092 8424
rect 6144 8412 6150 8424
rect 6564 8412 6592 8443
rect 8386 8440 8392 8452
rect 8444 8440 8450 8492
rect 9145 8483 9203 8489
rect 9145 8449 9157 8483
rect 9191 8480 9203 8483
rect 10226 8480 10232 8492
rect 9191 8452 10232 8480
rect 9191 8449 9203 8452
rect 9145 8443 9203 8449
rect 10226 8440 10232 8452
rect 10284 8440 10290 8492
rect 10336 8489 10364 8520
rect 10321 8483 10379 8489
rect 10321 8449 10333 8483
rect 10367 8449 10379 8483
rect 10321 8443 10379 8449
rect 6144 8384 6592 8412
rect 7653 8415 7711 8421
rect 6144 8372 6150 8384
rect 7653 8381 7665 8415
rect 7699 8412 7711 8415
rect 7742 8412 7748 8424
rect 7699 8384 7748 8412
rect 7699 8381 7711 8384
rect 7653 8375 7711 8381
rect 7742 8372 7748 8384
rect 7800 8372 7806 8424
rect 9398 8412 9404 8424
rect 9359 8384 9404 8412
rect 9398 8372 9404 8384
rect 9456 8372 9462 8424
rect 2501 8347 2559 8353
rect 2501 8313 2513 8347
rect 2547 8313 2559 8347
rect 2501 8307 2559 8313
rect 2777 8347 2835 8353
rect 2777 8313 2789 8347
rect 2823 8344 2835 8347
rect 3142 8344 3148 8356
rect 2823 8316 3148 8344
rect 2823 8313 2835 8316
rect 2777 8307 2835 8313
rect 3142 8304 3148 8316
rect 3200 8304 3206 8356
rect 5261 8347 5319 8353
rect 5261 8344 5273 8347
rect 4172 8316 5273 8344
rect 2866 8236 2872 8288
rect 2924 8276 2930 8288
rect 4172 8276 4200 8316
rect 5261 8313 5273 8316
rect 5307 8313 5319 8347
rect 5261 8307 5319 8313
rect 5534 8304 5540 8356
rect 5592 8344 5598 8356
rect 6365 8347 6423 8353
rect 6365 8344 6377 8347
rect 5592 8316 6377 8344
rect 5592 8304 5598 8316
rect 6365 8313 6377 8316
rect 6411 8313 6423 8347
rect 8018 8344 8024 8356
rect 7979 8316 8024 8344
rect 6365 8307 6423 8313
rect 8018 8304 8024 8316
rect 8076 8304 8082 8356
rect 18874 8304 18880 8356
rect 18932 8344 18938 8356
rect 20162 8344 20168 8356
rect 18932 8316 20168 8344
rect 18932 8304 18938 8316
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 2924 8248 4200 8276
rect 4617 8279 4675 8285
rect 2924 8236 2930 8248
rect 4617 8245 4629 8279
rect 4663 8276 4675 8279
rect 4798 8276 4804 8288
rect 4663 8248 4804 8276
rect 4663 8245 4675 8248
rect 4617 8239 4675 8245
rect 4798 8236 4804 8248
rect 4856 8236 4862 8288
rect 7098 8236 7104 8288
rect 7156 8276 7162 8288
rect 7650 8276 7656 8288
rect 7156 8248 7656 8276
rect 7156 8236 7162 8248
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 1486 8072 1492 8084
rect 1447 8044 1492 8072
rect 1486 8032 1492 8044
rect 1544 8032 1550 8084
rect 1578 8032 1584 8084
rect 1636 8072 1642 8084
rect 2225 8075 2283 8081
rect 2225 8072 2237 8075
rect 1636 8044 2237 8072
rect 1636 8032 1642 8044
rect 2225 8041 2237 8044
rect 2271 8041 2283 8075
rect 2225 8035 2283 8041
rect 2746 8044 3832 8072
rect 1946 8004 1952 8016
rect 1907 7976 1952 8004
rect 1946 7964 1952 7976
rect 2004 7964 2010 8016
rect 2130 7936 2136 7948
rect 1780 7908 2136 7936
rect 1780 7877 1808 7908
rect 2130 7896 2136 7908
rect 2188 7896 2194 7948
rect 1765 7871 1823 7877
rect 1765 7837 1777 7871
rect 1811 7837 1823 7871
rect 2406 7868 2412 7880
rect 2367 7840 2412 7868
rect 1765 7831 1823 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2130 7760 2136 7812
rect 2188 7800 2194 7812
rect 2746 7800 2774 8044
rect 3804 8013 3832 8044
rect 5902 8032 5908 8084
rect 5960 8072 5966 8084
rect 8573 8075 8631 8081
rect 8573 8072 8585 8075
rect 5960 8044 8585 8072
rect 5960 8032 5966 8044
rect 8573 8041 8585 8044
rect 8619 8041 8631 8075
rect 8573 8035 8631 8041
rect 3789 8007 3847 8013
rect 3789 7973 3801 8007
rect 3835 7973 3847 8007
rect 3789 7967 3847 7973
rect 4154 7964 4160 8016
rect 4212 8004 4218 8016
rect 8588 8004 8616 8035
rect 10226 8032 10232 8084
rect 10284 8072 10290 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10284 8044 10609 8072
rect 10284 8032 10290 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 18874 8072 18880 8084
rect 18835 8044 18880 8072
rect 10597 8035 10655 8041
rect 18874 8032 18880 8044
rect 18932 8032 18938 8084
rect 4212 7976 5304 8004
rect 8588 7976 9996 8004
rect 4212 7964 4218 7976
rect 3326 7936 3332 7948
rect 3287 7908 3332 7936
rect 3326 7896 3332 7908
rect 3384 7896 3390 7948
rect 4246 7936 4252 7948
rect 3896 7908 4252 7936
rect 3053 7871 3111 7877
rect 3053 7837 3065 7871
rect 3099 7868 3111 7871
rect 3896 7868 3924 7908
rect 4246 7896 4252 7908
rect 4304 7896 4310 7948
rect 4706 7936 4712 7948
rect 4667 7908 4712 7936
rect 4706 7896 4712 7908
rect 4764 7896 4770 7948
rect 4798 7896 4804 7948
rect 4856 7936 4862 7948
rect 5276 7945 5304 7976
rect 5261 7939 5319 7945
rect 4856 7908 4901 7936
rect 4856 7896 4862 7908
rect 5261 7905 5273 7939
rect 5307 7905 5319 7939
rect 5261 7899 5319 7905
rect 9306 7896 9312 7948
rect 9364 7936 9370 7948
rect 9493 7939 9551 7945
rect 9493 7936 9505 7939
rect 9364 7908 9505 7936
rect 9364 7896 9370 7908
rect 9493 7905 9505 7908
rect 9539 7905 9551 7939
rect 9493 7899 9551 7905
rect 3099 7840 3924 7868
rect 3099 7837 3111 7840
rect 3053 7831 3111 7837
rect 3970 7828 3976 7880
rect 4028 7868 4034 7880
rect 4617 7871 4675 7877
rect 4028 7840 4073 7868
rect 4028 7828 4034 7840
rect 4617 7837 4629 7871
rect 4663 7868 4675 7871
rect 4982 7868 4988 7880
rect 4663 7840 4988 7868
rect 4663 7837 4675 7840
rect 4617 7831 4675 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7868 7251 7871
rect 9398 7868 9404 7880
rect 7239 7840 9404 7868
rect 7239 7837 7251 7840
rect 7193 7831 7251 7837
rect 9398 7828 9404 7840
rect 9456 7828 9462 7880
rect 9968 7877 9996 7976
rect 9953 7871 10011 7877
rect 9953 7837 9965 7871
rect 9999 7837 10011 7871
rect 18690 7868 18696 7880
rect 18603 7840 18696 7868
rect 9953 7831 10011 7837
rect 18690 7828 18696 7840
rect 18748 7868 18754 7880
rect 19245 7871 19303 7877
rect 19245 7868 19257 7871
rect 18748 7840 19257 7868
rect 18748 7828 18754 7840
rect 19245 7837 19257 7840
rect 19291 7837 19303 7871
rect 19245 7831 19303 7837
rect 2188 7772 2774 7800
rect 5528 7803 5586 7809
rect 2188 7760 2194 7772
rect 5528 7769 5540 7803
rect 5574 7800 5586 7803
rect 5994 7800 6000 7812
rect 5574 7772 6000 7800
rect 5574 7769 5586 7772
rect 5528 7763 5586 7769
rect 5994 7760 6000 7772
rect 6052 7760 6058 7812
rect 7460 7803 7518 7809
rect 6472 7772 7052 7800
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2685 7735 2743 7741
rect 2685 7732 2697 7735
rect 2372 7704 2697 7732
rect 2372 7692 2378 7704
rect 2685 7701 2697 7704
rect 2731 7701 2743 7735
rect 2685 7695 2743 7701
rect 3145 7735 3203 7741
rect 3145 7701 3157 7735
rect 3191 7732 3203 7735
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 3191 7704 4261 7732
rect 3191 7701 3203 7704
rect 3145 7695 3203 7701
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 4890 7692 4896 7744
rect 4948 7732 4954 7744
rect 6472 7732 6500 7772
rect 6638 7732 6644 7744
rect 4948 7704 6500 7732
rect 6599 7704 6644 7732
rect 4948 7692 4954 7704
rect 6638 7692 6644 7704
rect 6696 7692 6702 7744
rect 7024 7732 7052 7772
rect 7460 7769 7472 7803
rect 7506 7800 7518 7803
rect 7742 7800 7748 7812
rect 7506 7772 7748 7800
rect 7506 7769 7518 7772
rect 7460 7763 7518 7769
rect 7742 7760 7748 7772
rect 7800 7760 7806 7812
rect 9309 7803 9367 7809
rect 9309 7800 9321 7803
rect 7852 7772 9321 7800
rect 7852 7732 7880 7772
rect 9309 7769 9321 7772
rect 9355 7769 9367 7803
rect 9309 7763 9367 7769
rect 7024 7704 7880 7732
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8720 7704 8953 7732
rect 8720 7692 8726 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 9401 7735 9459 7741
rect 9401 7701 9413 7735
rect 9447 7732 9459 7735
rect 10318 7732 10324 7744
rect 9447 7704 10324 7732
rect 9447 7701 9459 7704
rect 9401 7695 9459 7701
rect 10318 7692 10324 7704
rect 10376 7692 10382 7744
rect 1104 7642 21896 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21896 7642
rect 1104 7568 21896 7590
rect 1394 7488 1400 7540
rect 1452 7528 1458 7540
rect 2041 7531 2099 7537
rect 2041 7528 2053 7531
rect 1452 7500 2053 7528
rect 1452 7488 1458 7500
rect 2041 7497 2053 7500
rect 2087 7497 2099 7531
rect 2041 7491 2099 7497
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 2501 7531 2559 7537
rect 2501 7528 2513 7531
rect 2280 7500 2513 7528
rect 2280 7488 2286 7500
rect 2501 7497 2513 7500
rect 2547 7497 2559 7531
rect 2501 7491 2559 7497
rect 3326 7488 3332 7540
rect 3384 7528 3390 7540
rect 5534 7528 5540 7540
rect 3384 7500 5540 7528
rect 3384 7488 3390 7500
rect 5534 7488 5540 7500
rect 5592 7488 5598 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 6546 7528 6552 7540
rect 5951 7500 6552 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 6546 7488 6552 7500
rect 6604 7488 6610 7540
rect 8386 7488 8392 7540
rect 8444 7528 8450 7540
rect 9125 7531 9183 7537
rect 9125 7528 9137 7531
rect 8444 7500 9137 7528
rect 8444 7488 8450 7500
rect 9125 7497 9137 7500
rect 9171 7497 9183 7531
rect 9582 7528 9588 7540
rect 9543 7500 9588 7528
rect 9125 7491 9183 7497
rect 9582 7488 9588 7500
rect 9640 7488 9646 7540
rect 10229 7531 10287 7537
rect 10229 7497 10241 7531
rect 10275 7528 10287 7531
rect 10318 7528 10324 7540
rect 10275 7500 10324 7528
rect 10275 7497 10287 7500
rect 10229 7491 10287 7497
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 19429 7531 19487 7537
rect 19429 7497 19441 7531
rect 19475 7528 19487 7531
rect 19518 7528 19524 7540
rect 19475 7500 19524 7528
rect 19475 7497 19487 7500
rect 19429 7491 19487 7497
rect 19518 7488 19524 7500
rect 19576 7488 19582 7540
rect 2958 7460 2964 7472
rect 2148 7432 2964 7460
rect 2148 7404 2176 7432
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 3418 7460 3424 7472
rect 3379 7432 3424 7460
rect 3418 7420 3424 7432
rect 3476 7420 3482 7472
rect 6638 7469 6644 7472
rect 6632 7460 6644 7469
rect 4172 7432 6408 7460
rect 6599 7432 6644 7460
rect 4172 7404 4200 7432
rect 1397 7395 1455 7401
rect 1397 7361 1409 7395
rect 1443 7392 1455 7395
rect 2130 7392 2136 7404
rect 1443 7364 2136 7392
rect 1443 7361 1455 7364
rect 1397 7355 1455 7361
rect 2130 7352 2136 7364
rect 2188 7352 2194 7404
rect 2225 7395 2283 7401
rect 2225 7361 2237 7395
rect 2271 7361 2283 7395
rect 2682 7392 2688 7404
rect 2643 7364 2688 7392
rect 2225 7355 2283 7361
rect 934 7216 940 7268
rect 992 7256 998 7268
rect 1394 7256 1400 7268
rect 992 7228 1400 7256
rect 992 7216 998 7228
rect 1394 7216 1400 7228
rect 1452 7216 1458 7268
rect 1578 7256 1584 7268
rect 1539 7228 1584 7256
rect 1578 7216 1584 7228
rect 1636 7216 1642 7268
rect 2240 7188 2268 7355
rect 2682 7352 2688 7364
rect 2740 7352 2746 7404
rect 4154 7392 4160 7404
rect 4115 7364 4160 7392
rect 4154 7352 4160 7364
rect 4212 7352 4218 7404
rect 4424 7395 4482 7401
rect 4424 7361 4436 7395
rect 4470 7392 4482 7395
rect 4798 7392 4804 7404
rect 4470 7364 4804 7392
rect 4470 7361 4482 7364
rect 4424 7355 4482 7361
rect 4798 7352 4804 7364
rect 4856 7352 4862 7404
rect 6380 7401 6408 7432
rect 6632 7423 6644 7432
rect 6696 7460 6702 7472
rect 9306 7460 9312 7472
rect 6696 7432 9312 7460
rect 6638 7420 6644 7423
rect 6696 7420 6702 7432
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 8294 7352 8300 7404
rect 8352 7392 8358 7404
rect 8481 7395 8539 7401
rect 8481 7392 8493 7395
rect 8352 7364 8493 7392
rect 8352 7352 8358 7364
rect 8481 7361 8493 7364
rect 8527 7361 8539 7395
rect 8588 7392 8616 7432
rect 9306 7420 9312 7432
rect 9364 7460 9370 7472
rect 9364 7432 9628 7460
rect 9364 7420 9370 7432
rect 9493 7395 9551 7401
rect 8588 7364 8708 7392
rect 8481 7355 8539 7361
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7293 3939 7327
rect 8570 7324 8576 7336
rect 8531 7296 8576 7324
rect 3881 7287 3939 7293
rect 3896 7256 3924 7287
rect 8570 7284 8576 7296
rect 8628 7284 8634 7336
rect 8680 7333 8708 7364
rect 9493 7361 9505 7395
rect 9539 7361 9551 7395
rect 9493 7355 9551 7361
rect 8665 7327 8723 7333
rect 8665 7293 8677 7327
rect 8711 7293 8723 7327
rect 8665 7287 8723 7293
rect 4154 7256 4160 7268
rect 3896 7228 4160 7256
rect 4154 7216 4160 7228
rect 4212 7216 4218 7268
rect 7374 7216 7380 7268
rect 7432 7256 7438 7268
rect 9508 7256 9536 7355
rect 9600 7324 9628 7432
rect 17954 7352 17960 7404
rect 18012 7392 18018 7404
rect 19245 7395 19303 7401
rect 19245 7392 19257 7395
rect 18012 7364 19257 7392
rect 18012 7352 18018 7364
rect 19245 7361 19257 7364
rect 19291 7392 19303 7395
rect 19705 7395 19763 7401
rect 19705 7392 19717 7395
rect 19291 7364 19717 7392
rect 19291 7361 19303 7364
rect 19245 7355 19303 7361
rect 19705 7361 19717 7364
rect 19751 7361 19763 7395
rect 19705 7355 19763 7361
rect 9677 7327 9735 7333
rect 9677 7324 9689 7327
rect 9600 7296 9689 7324
rect 9677 7293 9689 7296
rect 9723 7293 9735 7327
rect 9677 7287 9735 7293
rect 7432 7228 9536 7256
rect 7432 7216 7438 7228
rect 5810 7188 5816 7200
rect 2240 7160 5816 7188
rect 5810 7148 5816 7160
rect 5868 7148 5874 7200
rect 7742 7188 7748 7200
rect 7703 7160 7748 7188
rect 7742 7148 7748 7160
rect 7800 7148 7806 7200
rect 8110 7188 8116 7200
rect 8071 7160 8116 7188
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 198 7080 204 7132
rect 256 7120 262 7132
rect 934 7120 940 7132
rect 256 7092 940 7120
rect 256 7080 262 7092
rect 934 7080 940 7092
rect 992 7080 998 7132
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 1578 6944 1584 6996
rect 1636 6984 1642 6996
rect 4157 6987 4215 6993
rect 1636 6956 3372 6984
rect 1636 6944 1642 6956
rect 3237 6919 3295 6925
rect 3237 6885 3249 6919
rect 3283 6885 3295 6919
rect 3344 6916 3372 6956
rect 4157 6953 4169 6987
rect 4203 6984 4215 6987
rect 4246 6984 4252 6996
rect 4203 6956 4252 6984
rect 4203 6953 4215 6956
rect 4157 6947 4215 6953
rect 4246 6944 4252 6956
rect 4304 6944 4310 6996
rect 5902 6984 5908 6996
rect 4356 6956 5908 6984
rect 4356 6916 4384 6956
rect 5902 6944 5908 6956
rect 5960 6944 5966 6996
rect 5994 6944 6000 6996
rect 6052 6984 6058 6996
rect 6181 6987 6239 6993
rect 6181 6984 6193 6987
rect 6052 6956 6193 6984
rect 6052 6944 6058 6956
rect 6181 6953 6193 6956
rect 6227 6953 6239 6987
rect 6181 6947 6239 6953
rect 3344 6888 4384 6916
rect 3237 6879 3295 6885
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 3252 6848 3280 6879
rect 4522 6876 4528 6928
rect 4580 6916 4586 6928
rect 5350 6916 5356 6928
rect 4580 6888 5356 6916
rect 4580 6876 4586 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 8941 6919 8999 6925
rect 8941 6916 8953 6919
rect 5460 6888 8953 6916
rect 3786 6848 3792 6860
rect 1268 6820 3280 6848
rect 3344 6820 3556 6848
rect 3747 6820 3792 6848
rect 1268 6808 1274 6820
rect 1394 6780 1400 6792
rect 1307 6752 1400 6780
rect 1394 6740 1400 6752
rect 1452 6780 1458 6792
rect 1670 6780 1676 6792
rect 1452 6752 1676 6780
rect 1452 6740 1458 6752
rect 1670 6740 1676 6752
rect 1728 6740 1734 6792
rect 1762 6740 1768 6792
rect 1820 6780 1826 6792
rect 1857 6783 1915 6789
rect 1857 6780 1869 6783
rect 1820 6752 1869 6780
rect 1820 6740 1826 6752
rect 1857 6749 1869 6752
rect 1903 6749 1915 6783
rect 1857 6743 1915 6749
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6780 2375 6783
rect 2777 6783 2835 6789
rect 2363 6752 2728 6780
rect 2363 6749 2375 6752
rect 2317 6743 2375 6749
rect 2700 6712 2728 6752
rect 2777 6749 2789 6783
rect 2823 6780 2835 6783
rect 2866 6780 2872 6792
rect 2823 6752 2872 6780
rect 2823 6749 2835 6752
rect 2777 6743 2835 6749
rect 2866 6740 2872 6752
rect 2924 6740 2930 6792
rect 3142 6712 3148 6724
rect 1596 6684 2636 6712
rect 2700 6684 3148 6712
rect 1596 6653 1624 6684
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6613 1639 6647
rect 2038 6644 2044 6656
rect 1999 6616 2044 6644
rect 1581 6607 1639 6613
rect 2038 6604 2044 6616
rect 2096 6604 2102 6656
rect 2498 6644 2504 6656
rect 2459 6616 2504 6644
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 2608 6644 2636 6684
rect 3142 6672 3148 6684
rect 3200 6712 3206 6724
rect 3344 6712 3372 6820
rect 3421 6783 3479 6789
rect 3421 6749 3433 6783
rect 3467 6749 3479 6783
rect 3528 6780 3556 6820
rect 3786 6808 3792 6820
rect 3844 6808 3850 6860
rect 4798 6848 4804 6860
rect 4759 6820 4804 6848
rect 4798 6808 4804 6820
rect 4856 6808 4862 6860
rect 5460 6848 5488 6888
rect 8941 6885 8953 6888
rect 8987 6916 8999 6919
rect 9582 6916 9588 6928
rect 8987 6888 9588 6916
rect 8987 6885 8999 6888
rect 8941 6879 8999 6885
rect 9582 6876 9588 6888
rect 9640 6876 9646 6928
rect 5276 6820 5488 6848
rect 3970 6780 3976 6792
rect 3528 6752 3976 6780
rect 3421 6743 3479 6749
rect 3200 6684 3372 6712
rect 3200 6672 3206 6684
rect 2682 6644 2688 6656
rect 2608 6616 2688 6644
rect 2682 6604 2688 6616
rect 2740 6604 2746 6656
rect 2961 6647 3019 6653
rect 2961 6613 2973 6647
rect 3007 6644 3019 6647
rect 3436 6644 3464 6743
rect 3970 6740 3976 6752
rect 4028 6740 4034 6792
rect 4154 6740 4160 6792
rect 4212 6780 4218 6792
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4212 6752 4537 6780
rect 4212 6740 4218 6752
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4614 6740 4620 6792
rect 4672 6780 4678 6792
rect 5276 6780 5304 6820
rect 7742 6808 7748 6860
rect 7800 6848 7806 6860
rect 8205 6851 8263 6857
rect 8205 6848 8217 6851
rect 7800 6820 8217 6848
rect 7800 6808 7806 6820
rect 8205 6817 8217 6820
rect 8251 6817 8263 6851
rect 8205 6811 8263 6817
rect 5534 6780 5540 6792
rect 4672 6752 5304 6780
rect 5495 6752 5540 6780
rect 4672 6740 4678 6752
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 8021 6783 8079 6789
rect 8021 6749 8033 6783
rect 8067 6780 8079 6783
rect 8110 6780 8116 6792
rect 8067 6752 8116 6780
rect 8067 6749 8079 6752
rect 8021 6743 8079 6749
rect 8110 6740 8116 6752
rect 8168 6740 8174 6792
rect 19610 6780 19616 6792
rect 19571 6752 19616 6780
rect 19610 6740 19616 6752
rect 19668 6740 19674 6792
rect 4246 6672 4252 6724
rect 4304 6712 4310 6724
rect 4430 6712 4436 6724
rect 4304 6684 4436 6712
rect 4304 6672 4310 6684
rect 4430 6672 4436 6684
rect 4488 6712 4494 6724
rect 5169 6715 5227 6721
rect 5169 6712 5181 6715
rect 4488 6684 5181 6712
rect 4488 6672 4494 6684
rect 5169 6681 5181 6684
rect 5215 6681 5227 6715
rect 5169 6675 5227 6681
rect 3007 6616 3464 6644
rect 3007 6613 3019 6616
rect 2961 6607 3019 6613
rect 4522 6604 4528 6656
rect 4580 6644 4586 6656
rect 4617 6647 4675 6653
rect 4617 6644 4629 6647
rect 4580 6616 4629 6644
rect 4580 6604 4586 6616
rect 4617 6613 4629 6616
rect 4663 6644 4675 6647
rect 5074 6644 5080 6656
rect 4663 6616 5080 6644
rect 4663 6613 4675 6616
rect 4617 6607 4675 6613
rect 5074 6604 5080 6616
rect 5132 6604 5138 6656
rect 5184 6644 5212 6675
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 5776 6684 7696 6712
rect 5776 6672 5782 6684
rect 6733 6647 6791 6653
rect 6733 6644 6745 6647
rect 5184 6616 6745 6644
rect 6733 6613 6745 6616
rect 6779 6613 6791 6647
rect 7098 6644 7104 6656
rect 7059 6616 7104 6644
rect 6733 6607 6791 6613
rect 7098 6604 7104 6616
rect 7156 6604 7162 6656
rect 7668 6653 7696 6684
rect 7653 6647 7711 6653
rect 7653 6613 7665 6647
rect 7699 6613 7711 6647
rect 7653 6607 7711 6613
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 8662 6644 8668 6656
rect 8159 6616 8668 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 8662 6604 8668 6616
rect 8720 6604 8726 6656
rect 19794 6644 19800 6656
rect 19755 6616 19800 6644
rect 19794 6604 19800 6616
rect 19852 6604 19858 6656
rect 1104 6554 21896 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21896 6554
rect 1104 6480 21896 6502
rect 1578 6440 1584 6452
rect 1539 6412 1584 6440
rect 1578 6400 1584 6412
rect 1636 6400 1642 6452
rect 2501 6443 2559 6449
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 2590 6440 2596 6452
rect 2547 6412 2596 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 2590 6400 2596 6412
rect 2648 6400 2654 6452
rect 2774 6400 2780 6452
rect 2832 6440 2838 6452
rect 2961 6443 3019 6449
rect 2961 6440 2973 6443
rect 2832 6412 2973 6440
rect 2832 6400 2838 6412
rect 2961 6409 2973 6412
rect 3007 6409 3019 6443
rect 3786 6440 3792 6452
rect 3747 6412 3792 6440
rect 2961 6403 3019 6409
rect 3786 6400 3792 6412
rect 3844 6400 3850 6452
rect 3970 6400 3976 6452
rect 4028 6440 4034 6452
rect 6365 6443 6423 6449
rect 6365 6440 6377 6443
rect 4028 6412 6377 6440
rect 4028 6400 4034 6412
rect 6365 6409 6377 6412
rect 6411 6409 6423 6443
rect 8294 6440 8300 6452
rect 8255 6412 8300 6440
rect 6365 6403 6423 6409
rect 8294 6400 8300 6412
rect 8352 6400 8358 6452
rect 20257 6443 20315 6449
rect 20257 6409 20269 6443
rect 20303 6440 20315 6443
rect 21634 6440 21640 6452
rect 20303 6412 21640 6440
rect 20303 6409 20315 6412
rect 20257 6403 20315 6409
rect 21634 6400 21640 6412
rect 21692 6400 21698 6452
rect 1670 6332 1676 6384
rect 1728 6372 1734 6384
rect 2682 6372 2688 6384
rect 1728 6344 2688 6372
rect 1728 6332 1734 6344
rect 2682 6332 2688 6344
rect 2740 6332 2746 6384
rect 4062 6372 4068 6384
rect 2792 6344 4068 6372
rect 1394 6304 1400 6316
rect 1355 6276 1400 6304
rect 1394 6264 1400 6276
rect 1452 6264 1458 6316
rect 1857 6307 1915 6313
rect 1857 6273 1869 6307
rect 1903 6273 1915 6307
rect 2314 6304 2320 6316
rect 2275 6276 2320 6304
rect 1857 6267 1915 6273
rect 1872 6236 1900 6267
rect 2314 6264 2320 6276
rect 2372 6264 2378 6316
rect 2792 6313 2820 6344
rect 4062 6332 4068 6344
rect 4120 6332 4126 6384
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 5721 6375 5779 6381
rect 5721 6372 5733 6375
rect 5684 6344 5733 6372
rect 5684 6332 5690 6344
rect 5721 6341 5733 6344
rect 5767 6341 5779 6375
rect 5721 6335 5779 6341
rect 2777 6307 2835 6313
rect 2777 6273 2789 6307
rect 2823 6273 2835 6307
rect 3234 6304 3240 6316
rect 3195 6276 3240 6304
rect 2777 6267 2835 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 20070 6304 20076 6316
rect 20031 6276 20076 6304
rect 20070 6264 20076 6276
rect 20128 6264 20134 6316
rect 2406 6236 2412 6248
rect 1872 6208 2412 6236
rect 2406 6196 2412 6208
rect 2464 6236 2470 6248
rect 6733 6239 6791 6245
rect 6733 6236 6745 6239
rect 2464 6208 6745 6236
rect 2464 6196 2470 6208
rect 6733 6205 6745 6208
rect 6779 6205 6791 6239
rect 6733 6199 6791 6205
rect 474 6128 480 6180
rect 532 6168 538 6180
rect 2041 6171 2099 6177
rect 2041 6168 2053 6171
rect 532 6140 2053 6168
rect 532 6128 538 6140
rect 2041 6137 2053 6140
rect 2087 6137 2099 6171
rect 3418 6168 3424 6180
rect 3379 6140 3424 6168
rect 2041 6131 2099 6137
rect 3418 6128 3424 6140
rect 3476 6128 3482 6180
rect 3970 6168 3976 6180
rect 3528 6140 3976 6168
rect 1762 6060 1768 6112
rect 1820 6100 1826 6112
rect 3528 6100 3556 6140
rect 3970 6128 3976 6140
rect 4028 6168 4034 6180
rect 4338 6168 4344 6180
rect 4028 6140 4344 6168
rect 4028 6128 4034 6140
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 4430 6128 4436 6180
rect 4488 6168 4494 6180
rect 5258 6168 5264 6180
rect 4488 6140 5264 6168
rect 4488 6128 4494 6140
rect 5258 6128 5264 6140
rect 5316 6168 5322 6180
rect 7929 6171 7987 6177
rect 7929 6168 7941 6171
rect 5316 6140 7941 6168
rect 5316 6128 5322 6140
rect 7929 6137 7941 6140
rect 7975 6168 7987 6171
rect 8570 6168 8576 6180
rect 7975 6140 8576 6168
rect 7975 6137 7987 6140
rect 7929 6131 7987 6137
rect 8570 6128 8576 6140
rect 8628 6128 8634 6180
rect 4154 6100 4160 6112
rect 1820 6072 3556 6100
rect 4115 6072 4160 6100
rect 1820 6060 1826 6072
rect 4154 6060 4160 6072
rect 4212 6100 4218 6112
rect 4614 6100 4620 6112
rect 4212 6072 4620 6100
rect 4212 6060 4218 6072
rect 4614 6060 4620 6072
rect 4672 6060 4678 6112
rect 4706 6060 4712 6112
rect 4764 6100 4770 6112
rect 4982 6100 4988 6112
rect 4764 6072 4988 6100
rect 4764 6060 4770 6072
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5074 6060 5080 6112
rect 5132 6100 5138 6112
rect 5350 6100 5356 6112
rect 5132 6072 5356 6100
rect 5132 6060 5138 6072
rect 5350 6060 5356 6072
rect 5408 6100 5414 6112
rect 7098 6100 7104 6112
rect 5408 6072 7104 6100
rect 5408 6060 5414 6072
rect 7098 6060 7104 6072
rect 7156 6060 7162 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 1780 5868 4568 5896
rect 1302 5652 1308 5704
rect 1360 5692 1366 5704
rect 1397 5695 1455 5701
rect 1397 5692 1409 5695
rect 1360 5664 1409 5692
rect 1360 5652 1366 5664
rect 1397 5661 1409 5664
rect 1443 5692 1455 5695
rect 1780 5692 1808 5868
rect 2498 5828 2504 5840
rect 2459 5800 2504 5828
rect 2498 5788 2504 5800
rect 2556 5788 2562 5840
rect 2866 5828 2872 5840
rect 2608 5800 2872 5828
rect 2608 5760 2636 5800
rect 2866 5788 2872 5800
rect 2924 5788 2930 5840
rect 2961 5831 3019 5837
rect 2961 5797 2973 5831
rect 3007 5828 3019 5831
rect 3050 5828 3056 5840
rect 3007 5800 3056 5828
rect 3007 5797 3019 5800
rect 2961 5791 3019 5797
rect 3050 5788 3056 5800
rect 3108 5788 3114 5840
rect 3326 5828 3332 5840
rect 3287 5800 3332 5828
rect 3326 5788 3332 5800
rect 3384 5788 3390 5840
rect 3786 5788 3792 5840
rect 3844 5828 3850 5840
rect 4430 5828 4436 5840
rect 3844 5800 4436 5828
rect 3844 5788 3850 5800
rect 4430 5788 4436 5800
rect 4488 5788 4494 5840
rect 4540 5828 4568 5868
rect 4614 5856 4620 5908
rect 4672 5896 4678 5908
rect 4982 5896 4988 5908
rect 4672 5868 4717 5896
rect 4943 5868 4988 5896
rect 4672 5856 4678 5868
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5350 5896 5356 5908
rect 5311 5868 5356 5896
rect 5350 5856 5356 5868
rect 5408 5856 5414 5908
rect 20717 5899 20775 5905
rect 20717 5865 20729 5899
rect 20763 5896 20775 5899
rect 21542 5896 21548 5908
rect 20763 5868 21548 5896
rect 20763 5865 20775 5868
rect 20717 5859 20775 5865
rect 21542 5856 21548 5868
rect 21600 5856 21606 5908
rect 6365 5831 6423 5837
rect 6365 5828 6377 5831
rect 4540 5800 6377 5828
rect 6365 5797 6377 5800
rect 6411 5797 6423 5831
rect 6365 5791 6423 5797
rect 20993 5831 21051 5837
rect 20993 5797 21005 5831
rect 21039 5828 21051 5831
rect 21818 5828 21824 5840
rect 21039 5800 21824 5828
rect 21039 5797 21051 5800
rect 20993 5791 21051 5797
rect 21818 5788 21824 5800
rect 21876 5788 21882 5840
rect 1872 5732 2636 5760
rect 1872 5701 1900 5732
rect 3234 5720 3240 5772
rect 3292 5760 3298 5772
rect 5629 5763 5687 5769
rect 5629 5760 5641 5763
rect 3292 5732 5641 5760
rect 3292 5720 3298 5732
rect 5629 5729 5641 5732
rect 5675 5729 5687 5763
rect 5629 5723 5687 5729
rect 1443 5664 1808 5692
rect 1857 5695 1915 5701
rect 1443 5661 1455 5664
rect 1397 5655 1455 5661
rect 1857 5661 1869 5695
rect 1903 5661 1915 5695
rect 1857 5655 1915 5661
rect 2222 5652 2228 5704
rect 2280 5692 2286 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2280 5664 2329 5692
rect 2280 5652 2286 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2038 5556 2044 5568
rect 1999 5528 2044 5556
rect 2038 5516 2044 5528
rect 2096 5516 2102 5568
rect 2332 5556 2360 5655
rect 2774 5652 2780 5704
rect 2832 5692 2838 5704
rect 5997 5695 6055 5701
rect 5997 5692 6009 5695
rect 2832 5664 6009 5692
rect 2832 5652 2838 5664
rect 5997 5661 6009 5664
rect 6043 5661 6055 5695
rect 20533 5695 20591 5701
rect 20533 5692 20545 5695
rect 5997 5655 6055 5661
rect 20180 5664 20545 5692
rect 5350 5624 5356 5636
rect 2746 5596 5356 5624
rect 2746 5556 2774 5596
rect 5350 5584 5356 5596
rect 5408 5584 5414 5636
rect 2332 5528 2774 5556
rect 3234 5516 3240 5568
rect 3292 5556 3298 5568
rect 3786 5556 3792 5568
rect 3292 5528 3792 5556
rect 3292 5516 3298 5528
rect 3786 5516 3792 5528
rect 3844 5516 3850 5568
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4338 5556 4344 5568
rect 4295 5528 4344 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4338 5516 4344 5528
rect 4396 5556 4402 5568
rect 5258 5556 5264 5568
rect 4396 5528 5264 5556
rect 4396 5516 4402 5528
rect 5258 5516 5264 5528
rect 5316 5516 5322 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 20180 5565 20208 5664
rect 20533 5661 20545 5664
rect 20579 5661 20591 5695
rect 20533 5655 20591 5661
rect 20806 5652 20812 5704
rect 20864 5692 20870 5704
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 20864 5664 21189 5692
rect 20864 5652 20870 5664
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 21177 5655 21235 5661
rect 20165 5559 20223 5565
rect 20165 5556 20177 5559
rect 8352 5528 20177 5556
rect 8352 5516 8358 5528
rect 20165 5525 20177 5528
rect 20211 5525 20223 5559
rect 20165 5519 20223 5525
rect 1104 5466 21896 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21896 5466
rect 1104 5392 21896 5414
rect 2038 5352 2044 5364
rect 1999 5324 2044 5352
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 2498 5352 2504 5364
rect 2459 5324 2504 5352
rect 2498 5312 2504 5324
rect 2556 5312 2562 5364
rect 2869 5355 2927 5361
rect 2869 5321 2881 5355
rect 2915 5352 2927 5355
rect 3050 5352 3056 5364
rect 2915 5324 3056 5352
rect 2915 5321 2927 5324
rect 2869 5315 2927 5321
rect 3050 5312 3056 5324
rect 3108 5312 3114 5364
rect 3970 5312 3976 5364
rect 4028 5312 4034 5364
rect 4614 5352 4620 5364
rect 4575 5324 4620 5352
rect 4614 5312 4620 5324
rect 4672 5312 4678 5364
rect 5350 5352 5356 5364
rect 5311 5324 5356 5352
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 5813 5355 5871 5361
rect 5813 5321 5825 5355
rect 5859 5352 5871 5355
rect 5902 5352 5908 5364
rect 5859 5324 5908 5352
rect 5859 5321 5871 5324
rect 5813 5315 5871 5321
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 934 5244 940 5296
rect 992 5284 998 5296
rect 3145 5287 3203 5293
rect 3145 5284 3157 5287
rect 992 5256 3157 5284
rect 992 5244 998 5256
rect 3145 5253 3157 5256
rect 3191 5253 3203 5287
rect 3988 5284 4016 5312
rect 4985 5287 5043 5293
rect 4985 5284 4997 5287
rect 3988 5256 4997 5284
rect 3145 5247 3203 5253
rect 4985 5253 4997 5256
rect 5031 5253 5043 5287
rect 4985 5247 5043 5253
rect 1302 5176 1308 5228
rect 1360 5216 1366 5228
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 1360 5188 1409 5216
rect 1360 5176 1366 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1854 5216 1860 5228
rect 1815 5188 1860 5216
rect 1397 5179 1455 5185
rect 1854 5176 1860 5188
rect 1912 5176 1918 5228
rect 2317 5219 2375 5225
rect 2317 5185 2329 5219
rect 2363 5216 2375 5219
rect 2774 5216 2780 5228
rect 2363 5188 2780 5216
rect 2363 5185 2375 5188
rect 2317 5179 2375 5185
rect 2774 5176 2780 5188
rect 2832 5216 2838 5228
rect 3970 5216 3976 5228
rect 2832 5188 3976 5216
rect 2832 5176 2838 5188
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 7466 5216 7472 5228
rect 4387 5188 7472 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 7466 5176 7472 5188
rect 7524 5176 7530 5228
rect 1872 5148 1900 5176
rect 3050 5148 3056 5160
rect 1872 5120 3056 5148
rect 3050 5108 3056 5120
rect 3108 5108 3114 5160
rect 20806 5148 20812 5160
rect 20767 5120 20812 5148
rect 20806 5108 20812 5120
rect 20864 5108 20870 5160
rect 5074 5080 5080 5092
rect 3528 5052 5080 5080
rect 1578 5012 1584 5024
rect 1539 4984 1584 5012
rect 1578 4972 1584 4984
rect 1636 4972 1642 5024
rect 2590 4972 2596 5024
rect 2648 5012 2654 5024
rect 3528 5021 3556 5052
rect 5074 5040 5080 5052
rect 5132 5040 5138 5092
rect 3513 5015 3571 5021
rect 3513 5012 3525 5015
rect 2648 4984 3525 5012
rect 2648 4972 2654 4984
rect 3513 4981 3525 4984
rect 3559 4981 3571 5015
rect 3513 4975 3571 4981
rect 3973 5015 4031 5021
rect 3973 4981 3985 5015
rect 4019 5012 4031 5015
rect 4246 5012 4252 5024
rect 4019 4984 4252 5012
rect 4019 4981 4031 4984
rect 3973 4975 4031 4981
rect 4246 4972 4252 4984
rect 4304 4972 4310 5024
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 658 4768 664 4820
rect 716 4808 722 4820
rect 2041 4811 2099 4817
rect 2041 4808 2053 4811
rect 716 4780 2053 4808
rect 716 4768 722 4780
rect 2041 4777 2053 4780
rect 2087 4777 2099 4811
rect 3878 4808 3884 4820
rect 3839 4780 3884 4808
rect 2041 4771 2099 4777
rect 3878 4768 3884 4780
rect 3936 4768 3942 4820
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 4157 4811 4215 4817
rect 4157 4808 4169 4811
rect 4120 4780 4169 4808
rect 4120 4768 4126 4780
rect 4157 4777 4169 4780
rect 4203 4777 4215 4811
rect 4157 4771 4215 4777
rect 750 4700 756 4752
rect 808 4740 814 4752
rect 2317 4743 2375 4749
rect 2317 4740 2329 4743
rect 808 4712 2329 4740
rect 808 4700 814 4712
rect 2317 4709 2329 4712
rect 2363 4709 2375 4743
rect 2317 4703 2375 4709
rect 2774 4700 2780 4752
rect 2832 4740 2838 4752
rect 4525 4743 4583 4749
rect 4525 4740 4537 4743
rect 2832 4712 4537 4740
rect 2832 4700 2838 4712
rect 4525 4709 4537 4712
rect 4571 4709 4583 4743
rect 4525 4703 4583 4709
rect 1118 4632 1124 4684
rect 1176 4672 1182 4684
rect 3145 4675 3203 4681
rect 3145 4672 3157 4675
rect 1176 4644 3157 4672
rect 1176 4632 1182 4644
rect 3145 4641 3157 4644
rect 3191 4641 3203 4675
rect 3145 4635 3203 4641
rect 1394 4604 1400 4616
rect 1307 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 1854 4604 1860 4616
rect 1767 4576 1860 4604
rect 1854 4564 1860 4576
rect 1912 4604 1918 4616
rect 4893 4607 4951 4613
rect 4893 4604 4905 4607
rect 1912 4576 4905 4604
rect 1912 4564 1918 4576
rect 4893 4573 4905 4576
rect 4939 4573 4951 4607
rect 4893 4567 4951 4573
rect 1412 4536 1440 4564
rect 3694 4536 3700 4548
rect 1412 4508 3700 4536
rect 3694 4496 3700 4508
rect 3752 4496 3758 4548
rect 1578 4468 1584 4480
rect 1539 4440 1584 4468
rect 1578 4428 1584 4440
rect 1636 4428 1642 4480
rect 2774 4468 2780 4480
rect 2735 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4468 2838 4480
rect 4154 4468 4160 4480
rect 2832 4440 4160 4468
rect 2832 4428 2838 4440
rect 4154 4428 4160 4440
rect 4212 4428 4218 4480
rect 1104 4378 21896 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21896 4378
rect 1104 4304 21896 4326
rect 2130 4224 2136 4276
rect 2188 4264 2194 4276
rect 3605 4267 3663 4273
rect 3605 4264 3617 4267
rect 2188 4236 3617 4264
rect 2188 4224 2194 4236
rect 3605 4233 3617 4236
rect 3651 4233 3663 4267
rect 3970 4264 3976 4276
rect 3931 4236 3976 4264
rect 3605 4227 3663 4233
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 7374 4196 7380 4208
rect 1964 4168 7380 4196
rect 1964 4137 1992 4168
rect 7374 4156 7380 4168
rect 7432 4156 7438 4208
rect 1949 4131 2007 4137
rect 1949 4097 1961 4131
rect 1995 4097 2007 4131
rect 1949 4091 2007 4097
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 4709 4131 4767 4137
rect 4709 4128 4721 4131
rect 3752 4100 4721 4128
rect 3752 4088 3758 4100
rect 4709 4097 4721 4100
rect 4755 4097 4767 4131
rect 4709 4091 4767 4097
rect 2222 4060 2228 4072
rect 2183 4032 2228 4060
rect 2222 4020 2228 4032
rect 2280 4020 2286 4072
rect 3050 4020 3056 4072
rect 3108 4060 3114 4072
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 3108 4032 4353 4060
rect 3108 4020 3114 4032
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 1946 3952 1952 4004
rect 2004 3992 2010 4004
rect 2869 3995 2927 4001
rect 2869 3992 2881 3995
rect 2004 3964 2881 3992
rect 2004 3952 2010 3964
rect 2869 3961 2881 3964
rect 2915 3961 2927 3995
rect 3234 3992 3240 4004
rect 3195 3964 3240 3992
rect 2869 3955 2927 3961
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 566 3884 572 3936
rect 624 3924 630 3936
rect 2501 3927 2559 3933
rect 2501 3924 2513 3927
rect 624 3896 2513 3924
rect 624 3884 630 3896
rect 2501 3893 2513 3896
rect 2547 3893 2559 3927
rect 2501 3887 2559 3893
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2222 3680 2228 3732
rect 2280 3720 2286 3732
rect 4157 3723 4215 3729
rect 4157 3720 4169 3723
rect 2280 3692 4169 3720
rect 2280 3680 2286 3692
rect 4157 3689 4169 3692
rect 4203 3689 4215 3723
rect 4157 3683 4215 3689
rect 2866 3612 2872 3664
rect 2924 3652 2930 3664
rect 3053 3655 3111 3661
rect 3053 3652 3065 3655
rect 2924 3624 3065 3652
rect 2924 3612 2930 3624
rect 3053 3621 3065 3624
rect 3099 3621 3111 3655
rect 3053 3615 3111 3621
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2777 3587 2835 3593
rect 2777 3553 2789 3587
rect 2823 3584 2835 3587
rect 4338 3584 4344 3596
rect 2823 3556 4344 3584
rect 2823 3553 2835 3556
rect 2777 3547 2835 3553
rect 4338 3544 4344 3556
rect 4396 3544 4402 3596
rect 2222 3516 2228 3528
rect 2183 3488 2228 3516
rect 2222 3476 2228 3488
rect 2280 3516 2286 3528
rect 4525 3519 4583 3525
rect 4525 3516 4537 3519
rect 2280 3488 4537 3516
rect 2280 3476 2286 3488
rect 4525 3485 4537 3488
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 2593 3451 2651 3457
rect 2593 3417 2605 3451
rect 2639 3448 2651 3451
rect 2866 3448 2872 3460
rect 2639 3420 2872 3448
rect 2639 3417 2651 3420
rect 2593 3411 2651 3417
rect 2866 3408 2872 3420
rect 2924 3408 2930 3460
rect 1302 3340 1308 3392
rect 1360 3380 1366 3392
rect 3789 3383 3847 3389
rect 3789 3380 3801 3383
rect 1360 3352 3801 3380
rect 1360 3340 1366 3352
rect 3789 3349 3801 3352
rect 3835 3349 3847 3383
rect 3789 3343 3847 3349
rect 1104 3290 21896 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21896 3290
rect 1104 3216 21896 3238
rect 2593 3179 2651 3185
rect 2593 3145 2605 3179
rect 2639 3176 2651 3179
rect 2774 3176 2780 3188
rect 2639 3148 2780 3176
rect 2639 3145 2651 3148
rect 2593 3139 2651 3145
rect 2774 3136 2780 3148
rect 2832 3136 2838 3188
rect 4706 3108 4712 3120
rect 1964 3080 4712 3108
rect 1964 3049 1992 3080
rect 4706 3068 4712 3080
rect 4764 3068 4770 3120
rect 1949 3043 2007 3049
rect 1949 3009 1961 3043
rect 1995 3009 2007 3043
rect 1949 3003 2007 3009
rect 2685 3043 2743 3049
rect 2685 3009 2697 3043
rect 2731 3040 2743 3043
rect 2774 3040 2780 3052
rect 2731 3012 2780 3040
rect 2731 3009 2743 3012
rect 2685 3003 2743 3009
rect 2774 3000 2780 3012
rect 2832 3040 2838 3052
rect 3789 3043 3847 3049
rect 3789 3040 3801 3043
rect 2832 3012 3801 3040
rect 2832 3000 2838 3012
rect 3789 3009 3801 3012
rect 3835 3009 3847 3043
rect 3789 3003 3847 3009
rect 2225 2975 2283 2981
rect 2225 2941 2237 2975
rect 2271 2972 2283 2975
rect 2866 2972 2872 2984
rect 2271 2944 2872 2972
rect 2271 2941 2283 2944
rect 2225 2935 2283 2941
rect 2866 2932 2872 2944
rect 2924 2972 2930 2984
rect 4157 2975 4215 2981
rect 4157 2972 4169 2975
rect 2924 2944 4169 2972
rect 2924 2932 2930 2944
rect 4157 2941 4169 2944
rect 4203 2941 4215 2975
rect 4157 2935 4215 2941
rect 2958 2864 2964 2916
rect 3016 2904 3022 2916
rect 4525 2907 4583 2913
rect 4525 2904 4537 2907
rect 3016 2876 4537 2904
rect 3016 2864 3022 2876
rect 4525 2873 4537 2876
rect 4571 2873 4583 2907
rect 4525 2867 4583 2873
rect 3050 2836 3056 2848
rect 3011 2808 3056 2836
rect 3050 2796 3056 2808
rect 3108 2796 3114 2848
rect 3234 2796 3240 2848
rect 3292 2836 3298 2848
rect 3421 2839 3479 2845
rect 3421 2836 3433 2839
rect 3292 2808 3433 2836
rect 3292 2796 3298 2808
rect 3421 2805 3433 2808
rect 3467 2805 3479 2839
rect 3421 2799 3479 2805
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2590 2592 2596 2644
rect 2648 2632 2654 2644
rect 2685 2635 2743 2641
rect 2685 2632 2697 2635
rect 2648 2604 2697 2632
rect 2648 2592 2654 2604
rect 2685 2601 2697 2604
rect 2731 2601 2743 2635
rect 2685 2595 2743 2601
rect 3145 2635 3203 2641
rect 3145 2601 3157 2635
rect 3191 2632 3203 2635
rect 3326 2632 3332 2644
rect 3191 2604 3332 2632
rect 3191 2601 3203 2604
rect 3145 2595 3203 2601
rect 3326 2592 3332 2604
rect 3384 2592 3390 2644
rect 4065 2635 4123 2641
rect 4065 2601 4077 2635
rect 4111 2632 4123 2635
rect 4246 2632 4252 2644
rect 4111 2604 4252 2632
rect 4111 2601 4123 2604
rect 4065 2595 4123 2601
rect 4246 2592 4252 2604
rect 4304 2592 4310 2644
rect 4890 2564 4896 2576
rect 1964 2536 4896 2564
rect 1964 2505 1992 2536
rect 4890 2524 4896 2536
rect 4948 2524 4954 2576
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 3418 2456 3424 2508
rect 3476 2496 3482 2508
rect 3476 2468 11928 2496
rect 3476 2456 3482 2468
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2397 2283 2431
rect 2225 2391 2283 2397
rect 2593 2431 2651 2437
rect 2593 2397 2605 2431
rect 2639 2428 2651 2431
rect 2774 2428 2780 2440
rect 2639 2400 2780 2428
rect 2639 2397 2651 2400
rect 2593 2391 2651 2397
rect 2240 2360 2268 2391
rect 2774 2388 2780 2400
rect 2832 2428 2838 2440
rect 11900 2437 11928 2468
rect 4893 2431 4951 2437
rect 4893 2428 4905 2431
rect 2832 2400 4905 2428
rect 2832 2388 2838 2400
rect 4893 2397 4905 2400
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2428 11943 2431
rect 12161 2431 12219 2437
rect 12161 2428 12173 2431
rect 11931 2400 12173 2428
rect 11931 2397 11943 2400
rect 11885 2391 11943 2397
rect 12161 2397 12173 2400
rect 12207 2397 12219 2431
rect 12161 2391 12219 2397
rect 2958 2360 2964 2372
rect 2240 2332 2964 2360
rect 2792 2304 2820 2332
rect 2958 2320 2964 2332
rect 3016 2320 3022 2372
rect 3234 2360 3240 2372
rect 3195 2332 3240 2360
rect 3234 2320 3240 2332
rect 3292 2320 3298 2372
rect 3970 2320 3976 2372
rect 4028 2360 4034 2372
rect 4157 2363 4215 2369
rect 4157 2360 4169 2363
rect 4028 2332 4169 2360
rect 4028 2320 4034 2332
rect 4157 2329 4169 2332
rect 4203 2360 4215 2363
rect 4525 2363 4583 2369
rect 4525 2360 4537 2363
rect 4203 2332 4537 2360
rect 4203 2329 4215 2332
rect 4157 2323 4215 2329
rect 4525 2329 4537 2332
rect 4571 2329 4583 2363
rect 4525 2323 4583 2329
rect 2774 2252 2780 2304
rect 2832 2252 2838 2304
rect 11698 2292 11704 2304
rect 11659 2264 11704 2292
rect 11698 2252 11704 2264
rect 11756 2252 11762 2304
rect 1104 2202 21896 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21896 2202
rect 1104 2128 21896 2150
<< via1 >>
rect 2780 21292 2832 21344
rect 9128 21292 9180 21344
rect 5632 20884 5684 20936
rect 6184 20884 6236 20936
rect 3976 20816 4028 20868
rect 6828 20816 6880 20868
rect 11244 20816 11296 20868
rect 16120 20816 16172 20868
rect 8392 20748 8444 20800
rect 8944 20748 8996 20800
rect 11704 20748 11756 20800
rect 12808 20748 12860 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 3424 20544 3476 20596
rect 3976 20544 4028 20596
rect 8484 20544 8536 20596
rect 9128 20587 9180 20596
rect 9128 20553 9137 20587
rect 9137 20553 9171 20587
rect 9171 20553 9180 20587
rect 9128 20544 9180 20553
rect 2044 20476 2096 20528
rect 848 20408 900 20460
rect 2964 20408 3016 20460
rect 6736 20451 6788 20460
rect 3332 20340 3384 20392
rect 3976 20340 4028 20392
rect 5540 20340 5592 20392
rect 5724 20383 5776 20392
rect 5724 20349 5733 20383
rect 5733 20349 5767 20383
rect 5767 20349 5776 20383
rect 5724 20340 5776 20349
rect 5816 20340 5868 20392
rect 6736 20417 6745 20451
rect 6745 20417 6779 20451
rect 6779 20417 6788 20451
rect 6736 20408 6788 20417
rect 8300 20408 8352 20460
rect 8668 20408 8720 20460
rect 8944 20451 8996 20460
rect 8944 20417 8953 20451
rect 8953 20417 8987 20451
rect 8987 20417 8996 20451
rect 8944 20408 8996 20417
rect 9496 20408 9548 20460
rect 12992 20544 13044 20596
rect 13084 20544 13136 20596
rect 13544 20544 13596 20596
rect 14464 20544 14516 20596
rect 15844 20544 15896 20596
rect 17224 20544 17276 20596
rect 18604 20544 18656 20596
rect 19432 20544 19484 20596
rect 12624 20476 12676 20528
rect 15936 20476 15988 20528
rect 11060 20408 11112 20460
rect 12716 20451 12768 20460
rect 12716 20417 12725 20451
rect 12725 20417 12759 20451
rect 12759 20417 12768 20451
rect 12716 20408 12768 20417
rect 13452 20451 13504 20460
rect 13452 20417 13461 20451
rect 13461 20417 13495 20451
rect 13495 20417 13504 20451
rect 13452 20408 13504 20417
rect 9404 20340 9456 20392
rect 9588 20340 9640 20392
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 6644 20204 6696 20256
rect 13636 20272 13688 20324
rect 14004 20272 14056 20324
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 12164 20247 12216 20256
rect 12164 20213 12173 20247
rect 12173 20213 12207 20247
rect 12207 20213 12216 20247
rect 12164 20204 12216 20213
rect 12256 20204 12308 20256
rect 15476 20451 15528 20460
rect 15476 20417 15485 20451
rect 15485 20417 15519 20451
rect 15519 20417 15528 20451
rect 15476 20408 15528 20417
rect 17592 20476 17644 20528
rect 17224 20340 17276 20392
rect 18052 20451 18104 20460
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 18604 20451 18656 20460
rect 18604 20417 18613 20451
rect 18613 20417 18647 20451
rect 18647 20417 18656 20451
rect 18604 20408 18656 20417
rect 17960 20340 18012 20392
rect 21088 20476 21140 20528
rect 20812 20408 20864 20460
rect 20536 20340 20588 20392
rect 20996 20340 21048 20392
rect 21456 20340 21508 20392
rect 22744 20340 22796 20392
rect 14924 20272 14976 20324
rect 16304 20272 16356 20324
rect 17684 20272 17736 20324
rect 18512 20204 18564 20256
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 8576 20000 8628 20052
rect 9680 20000 9732 20052
rect 8760 19932 8812 19984
rect 1216 19796 1268 19848
rect 1584 19796 1636 19848
rect 2504 19796 2556 19848
rect 5448 19864 5500 19916
rect 8668 19864 8720 19916
rect 10048 19864 10100 19916
rect 5172 19839 5224 19848
rect 5172 19805 5181 19839
rect 5181 19805 5215 19839
rect 5215 19805 5224 19839
rect 5172 19796 5224 19805
rect 5540 19796 5592 19848
rect 6644 19839 6696 19848
rect 6644 19805 6662 19839
rect 6662 19805 6696 19839
rect 6920 19839 6972 19848
rect 6644 19796 6696 19805
rect 6920 19805 6929 19839
rect 6929 19805 6963 19839
rect 6963 19805 6972 19839
rect 6920 19796 6972 19805
rect 9220 19796 9272 19848
rect 9588 19796 9640 19848
rect 10784 19796 10836 19848
rect 13452 20000 13504 20052
rect 15384 20000 15436 20052
rect 16948 20043 17000 20052
rect 16948 20009 16957 20043
rect 16957 20009 16991 20043
rect 16991 20009 17000 20043
rect 16948 20000 17000 20009
rect 17224 20000 17276 20052
rect 18144 20000 18196 20052
rect 19524 20000 19576 20052
rect 11796 19932 11848 19984
rect 19616 19932 19668 19984
rect 13912 19864 13964 19916
rect 11888 19796 11940 19848
rect 13176 19796 13228 19848
rect 14556 19839 14608 19848
rect 4160 19728 4212 19780
rect 3976 19660 4028 19712
rect 5540 19703 5592 19712
rect 5540 19669 5549 19703
rect 5549 19669 5583 19703
rect 5583 19669 5592 19703
rect 5540 19660 5592 19669
rect 6644 19660 6696 19712
rect 7196 19703 7248 19712
rect 7196 19669 7205 19703
rect 7205 19669 7239 19703
rect 7239 19669 7248 19703
rect 7196 19660 7248 19669
rect 8484 19660 8536 19712
rect 8852 19660 8904 19712
rect 9312 19703 9364 19712
rect 9312 19669 9321 19703
rect 9321 19669 9355 19703
rect 9355 19669 9364 19703
rect 9312 19660 9364 19669
rect 9588 19660 9640 19712
rect 9772 19703 9824 19712
rect 9772 19669 9781 19703
rect 9781 19669 9815 19703
rect 9815 19669 9824 19703
rect 9772 19660 9824 19669
rect 12164 19728 12216 19780
rect 13452 19728 13504 19780
rect 14556 19805 14565 19839
rect 14565 19805 14599 19839
rect 14599 19805 14608 19839
rect 14556 19796 14608 19805
rect 14280 19703 14332 19712
rect 14280 19669 14289 19703
rect 14289 19669 14323 19703
rect 14323 19669 14332 19703
rect 14280 19660 14332 19669
rect 15936 19796 15988 19848
rect 16396 19796 16448 19848
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 17132 19839 17184 19848
rect 16488 19796 16540 19805
rect 17132 19805 17141 19839
rect 17141 19805 17175 19839
rect 17175 19805 17184 19839
rect 17132 19796 17184 19805
rect 17868 19864 17920 19916
rect 19708 19864 19760 19916
rect 20720 19907 20772 19916
rect 20720 19873 20729 19907
rect 20729 19873 20763 19907
rect 20763 19873 20772 19907
rect 20720 19864 20772 19873
rect 19064 19796 19116 19848
rect 19340 19839 19392 19848
rect 19340 19805 19349 19839
rect 19349 19805 19383 19839
rect 19383 19805 19392 19839
rect 19340 19796 19392 19805
rect 20168 19796 20220 19848
rect 21364 19839 21416 19848
rect 21364 19805 21373 19839
rect 21373 19805 21407 19839
rect 21407 19805 21416 19839
rect 21364 19796 21416 19805
rect 22284 19796 22336 19848
rect 19432 19728 19484 19780
rect 16028 19703 16080 19712
rect 16028 19669 16037 19703
rect 16037 19669 16071 19703
rect 16071 19669 16080 19703
rect 16028 19660 16080 19669
rect 17132 19660 17184 19712
rect 17868 19660 17920 19712
rect 18144 19660 18196 19712
rect 18788 19703 18840 19712
rect 18788 19669 18797 19703
rect 18797 19669 18831 19703
rect 18831 19669 18840 19703
rect 18788 19660 18840 19669
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 2872 19456 2924 19508
rect 4068 19456 4120 19508
rect 5448 19456 5500 19508
rect 4988 19388 5040 19440
rect 5356 19388 5408 19440
rect 7012 19456 7064 19508
rect 7288 19456 7340 19508
rect 8668 19456 8720 19508
rect 2044 19320 2096 19372
rect 940 19252 992 19304
rect 1124 19252 1176 19304
rect 4436 19320 4488 19372
rect 5080 19320 5132 19372
rect 5172 19252 5224 19304
rect 7196 19388 7248 19440
rect 11888 19456 11940 19508
rect 5816 19320 5868 19372
rect 6092 19320 6144 19372
rect 6552 19363 6604 19372
rect 6552 19329 6561 19363
rect 6561 19329 6595 19363
rect 6595 19329 6604 19363
rect 6552 19320 6604 19329
rect 572 19184 624 19236
rect 2504 19184 2556 19236
rect 4528 19227 4580 19236
rect 4528 19193 4537 19227
rect 4537 19193 4571 19227
rect 4571 19193 4580 19227
rect 4528 19184 4580 19193
rect 5448 19184 5500 19236
rect 4620 19116 4672 19168
rect 7196 19252 7248 19304
rect 9956 19388 10008 19440
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 7380 19252 7432 19304
rect 8576 19363 8628 19372
rect 8576 19329 8585 19363
rect 8585 19329 8619 19363
rect 8619 19329 8628 19363
rect 8576 19320 8628 19329
rect 8852 19320 8904 19372
rect 9588 19320 9640 19372
rect 10508 19363 10560 19372
rect 10508 19329 10526 19363
rect 10526 19329 10560 19363
rect 10508 19320 10560 19329
rect 10784 19363 10836 19372
rect 10784 19329 10793 19363
rect 10793 19329 10827 19363
rect 10827 19329 10836 19363
rect 10784 19320 10836 19329
rect 11152 19320 11204 19372
rect 12348 19388 12400 19440
rect 13912 19499 13964 19508
rect 13912 19465 13921 19499
rect 13921 19465 13955 19499
rect 13955 19465 13964 19499
rect 13912 19456 13964 19465
rect 9680 19252 9732 19304
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 12992 19363 13044 19372
rect 12992 19329 13001 19363
rect 13001 19329 13035 19363
rect 13035 19329 13044 19363
rect 12992 19320 13044 19329
rect 12900 19252 12952 19304
rect 13728 19363 13780 19372
rect 13728 19329 13737 19363
rect 13737 19329 13771 19363
rect 13771 19329 13780 19363
rect 13728 19320 13780 19329
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 14740 19295 14792 19304
rect 12808 19184 12860 19236
rect 14464 19184 14516 19236
rect 14740 19261 14749 19295
rect 14749 19261 14783 19295
rect 14783 19261 14792 19295
rect 14740 19252 14792 19261
rect 15200 19252 15252 19304
rect 15292 19184 15344 19236
rect 15752 19456 15804 19508
rect 16948 19456 17000 19508
rect 17316 19456 17368 19508
rect 17592 19499 17644 19508
rect 17592 19465 17601 19499
rect 17601 19465 17635 19499
rect 17635 19465 17644 19499
rect 17592 19456 17644 19465
rect 18512 19499 18564 19508
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 16856 19363 16908 19372
rect 16856 19329 16865 19363
rect 16865 19329 16899 19363
rect 16899 19329 16908 19363
rect 16856 19320 16908 19329
rect 17408 19320 17460 19372
rect 18512 19465 18521 19499
rect 18521 19465 18555 19499
rect 18555 19465 18564 19499
rect 18512 19456 18564 19465
rect 19892 19456 19944 19508
rect 19984 19456 20036 19508
rect 20444 19456 20496 19508
rect 18328 19388 18380 19440
rect 19524 19388 19576 19440
rect 19432 19320 19484 19372
rect 19616 19363 19668 19372
rect 19616 19329 19625 19363
rect 19625 19329 19659 19363
rect 19659 19329 19668 19363
rect 19616 19320 19668 19329
rect 20628 19363 20680 19372
rect 20628 19329 20637 19363
rect 20637 19329 20671 19363
rect 20671 19329 20680 19363
rect 20628 19320 20680 19329
rect 21732 19320 21784 19372
rect 7840 19159 7892 19168
rect 7840 19125 7849 19159
rect 7849 19125 7883 19159
rect 7883 19125 7892 19159
rect 7840 19116 7892 19125
rect 10416 19116 10468 19168
rect 10876 19116 10928 19168
rect 14280 19116 14332 19168
rect 15844 19116 15896 19168
rect 21180 19159 21232 19168
rect 21180 19125 21189 19159
rect 21189 19125 21223 19159
rect 21223 19125 21232 19159
rect 21180 19116 21232 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 4160 18912 4212 18964
rect 3700 18844 3752 18896
rect 3884 18844 3936 18896
rect 5540 18912 5592 18964
rect 6736 18955 6788 18964
rect 6736 18921 6745 18955
rect 6745 18921 6779 18955
rect 6779 18921 6788 18955
rect 6736 18912 6788 18921
rect 8484 18912 8536 18964
rect 2872 18819 2924 18828
rect 2872 18785 2881 18819
rect 2881 18785 2915 18819
rect 2915 18785 2924 18819
rect 2872 18776 2924 18785
rect 4804 18844 4856 18896
rect 5264 18776 5316 18828
rect 7564 18844 7616 18896
rect 10232 18912 10284 18964
rect 10508 18912 10560 18964
rect 10968 18912 11020 18964
rect 15384 18912 15436 18964
rect 15476 18912 15528 18964
rect 18052 18912 18104 18964
rect 20904 18912 20956 18964
rect 3792 18751 3844 18760
rect 3792 18717 3801 18751
rect 3801 18717 3835 18751
rect 3835 18717 3844 18751
rect 3792 18708 3844 18717
rect 5172 18708 5224 18760
rect 8300 18776 8352 18828
rect 11060 18844 11112 18896
rect 6000 18708 6052 18760
rect 7012 18751 7064 18760
rect 7012 18717 7021 18751
rect 7021 18717 7055 18751
rect 7055 18717 7064 18751
rect 7012 18708 7064 18717
rect 8208 18708 8260 18760
rect 9772 18776 9824 18828
rect 13820 18844 13872 18896
rect 15752 18844 15804 18896
rect 12440 18776 12492 18828
rect 11244 18751 11296 18760
rect 11244 18717 11253 18751
rect 11253 18717 11287 18751
rect 11287 18717 11296 18751
rect 11244 18708 11296 18717
rect 12624 18708 12676 18760
rect 15108 18708 15160 18760
rect 2688 18640 2740 18692
rect 2964 18615 3016 18624
rect 2964 18581 2973 18615
rect 2973 18581 3007 18615
rect 3007 18581 3016 18615
rect 2964 18572 3016 18581
rect 3240 18572 3292 18624
rect 3424 18615 3476 18624
rect 3424 18581 3433 18615
rect 3433 18581 3467 18615
rect 3467 18581 3476 18615
rect 3424 18572 3476 18581
rect 3700 18572 3752 18624
rect 4436 18572 4488 18624
rect 4712 18615 4764 18624
rect 4712 18581 4721 18615
rect 4721 18581 4755 18615
rect 4755 18581 4764 18615
rect 4712 18572 4764 18581
rect 9496 18640 9548 18692
rect 11060 18640 11112 18692
rect 15844 18708 15896 18760
rect 16304 18708 16356 18760
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 7932 18615 7984 18624
rect 7932 18581 7941 18615
rect 7941 18581 7975 18615
rect 7975 18581 7984 18615
rect 7932 18572 7984 18581
rect 11704 18572 11756 18624
rect 12072 18615 12124 18624
rect 12072 18581 12081 18615
rect 12081 18581 12115 18615
rect 12115 18581 12124 18615
rect 12072 18572 12124 18581
rect 12164 18615 12216 18624
rect 12164 18581 12173 18615
rect 12173 18581 12207 18615
rect 12207 18581 12216 18615
rect 12532 18615 12584 18624
rect 12164 18572 12216 18581
rect 12532 18581 12541 18615
rect 12541 18581 12575 18615
rect 12575 18581 12584 18615
rect 12532 18572 12584 18581
rect 12808 18572 12860 18624
rect 14004 18572 14056 18624
rect 17132 18640 17184 18692
rect 17592 18640 17644 18692
rect 17960 18844 18012 18896
rect 21824 18844 21876 18896
rect 21180 18776 21232 18828
rect 18880 18708 18932 18760
rect 18420 18640 18472 18692
rect 18512 18640 18564 18692
rect 21640 18708 21692 18760
rect 21824 18640 21876 18692
rect 19800 18572 19852 18624
rect 20260 18572 20312 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 2044 18368 2096 18420
rect 2688 18411 2740 18420
rect 2688 18377 2697 18411
rect 2697 18377 2731 18411
rect 2731 18377 2740 18411
rect 2688 18368 2740 18377
rect 2964 18368 3016 18420
rect 4160 18368 4212 18420
rect 4620 18411 4672 18420
rect 4620 18377 4629 18411
rect 4629 18377 4663 18411
rect 4663 18377 4672 18411
rect 4620 18368 4672 18377
rect 5816 18368 5868 18420
rect 5172 18300 5224 18352
rect 3516 18232 3568 18284
rect 3884 18232 3936 18284
rect 4804 18232 4856 18284
rect 5724 18275 5776 18284
rect 5724 18241 5742 18275
rect 5742 18241 5776 18275
rect 5724 18232 5776 18241
rect 6828 18368 6880 18420
rect 7104 18368 7156 18420
rect 8300 18368 8352 18420
rect 8484 18368 8536 18420
rect 9588 18368 9640 18420
rect 10048 18411 10100 18420
rect 10048 18377 10057 18411
rect 10057 18377 10091 18411
rect 10091 18377 10100 18411
rect 10048 18368 10100 18377
rect 14740 18368 14792 18420
rect 15292 18368 15344 18420
rect 16304 18368 16356 18420
rect 18604 18368 18656 18420
rect 21272 18411 21324 18420
rect 21272 18377 21281 18411
rect 21281 18377 21315 18411
rect 21315 18377 21324 18411
rect 21272 18368 21324 18377
rect 11796 18300 11848 18352
rect 6460 18232 6512 18284
rect 2504 18096 2556 18148
rect 3792 18096 3844 18148
rect 3976 18096 4028 18148
rect 6920 18164 6972 18216
rect 9772 18232 9824 18284
rect 10416 18232 10468 18284
rect 12256 18300 12308 18352
rect 12716 18300 12768 18352
rect 13544 18300 13596 18352
rect 14004 18300 14056 18352
rect 14464 18300 14516 18352
rect 16396 18300 16448 18352
rect 17500 18300 17552 18352
rect 17592 18300 17644 18352
rect 13268 18232 13320 18284
rect 13636 18232 13688 18284
rect 13820 18275 13872 18284
rect 13820 18241 13829 18275
rect 13829 18241 13863 18275
rect 13863 18241 13872 18275
rect 13820 18232 13872 18241
rect 14096 18232 14148 18284
rect 14004 18207 14056 18216
rect 14004 18173 14013 18207
rect 14013 18173 14047 18207
rect 14047 18173 14056 18207
rect 14004 18164 14056 18173
rect 2872 18028 2924 18080
rect 3424 18028 3476 18080
rect 6828 18028 6880 18080
rect 7196 18028 7248 18080
rect 8208 18028 8260 18080
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 9680 18028 9732 18037
rect 10968 18071 11020 18080
rect 10968 18037 10977 18071
rect 10977 18037 11011 18071
rect 11011 18037 11020 18071
rect 10968 18028 11020 18037
rect 12440 18028 12492 18080
rect 13084 18028 13136 18080
rect 13360 18071 13412 18080
rect 13360 18037 13369 18071
rect 13369 18037 13403 18071
rect 13403 18037 13412 18071
rect 13360 18028 13412 18037
rect 14372 18071 14424 18080
rect 14372 18037 14381 18071
rect 14381 18037 14415 18071
rect 14415 18037 14424 18071
rect 14372 18028 14424 18037
rect 15752 18232 15804 18284
rect 16488 18232 16540 18284
rect 18328 18275 18380 18284
rect 18328 18241 18337 18275
rect 18337 18241 18371 18275
rect 18371 18241 18380 18275
rect 18328 18232 18380 18241
rect 18420 18232 18472 18284
rect 15384 18207 15436 18216
rect 15384 18173 15393 18207
rect 15393 18173 15427 18207
rect 15427 18173 15436 18207
rect 15384 18164 15436 18173
rect 19800 18232 19852 18284
rect 20352 18275 20404 18284
rect 20352 18241 20361 18275
rect 20361 18241 20395 18275
rect 20395 18241 20404 18275
rect 20352 18232 20404 18241
rect 20812 18275 20864 18284
rect 20812 18241 20821 18275
rect 20821 18241 20855 18275
rect 20855 18241 20864 18275
rect 20812 18232 20864 18241
rect 21548 18232 21600 18284
rect 21180 18164 21232 18216
rect 18052 18096 18104 18148
rect 19708 18139 19760 18148
rect 19708 18105 19717 18139
rect 19717 18105 19751 18139
rect 19751 18105 19760 18139
rect 19708 18096 19760 18105
rect 20628 18139 20680 18148
rect 20628 18105 20637 18139
rect 20637 18105 20671 18139
rect 20671 18105 20680 18139
rect 20628 18096 20680 18105
rect 18788 18028 18840 18080
rect 18972 18071 19024 18080
rect 18972 18037 18981 18071
rect 18981 18037 19015 18071
rect 19015 18037 19024 18071
rect 18972 18028 19024 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 5540 17824 5592 17876
rect 6000 17824 6052 17876
rect 10324 17824 10376 17876
rect 11244 17824 11296 17876
rect 12624 17824 12676 17876
rect 14832 17867 14884 17876
rect 14832 17833 14841 17867
rect 14841 17833 14875 17867
rect 14875 17833 14884 17867
rect 14832 17824 14884 17833
rect 16488 17867 16540 17876
rect 2872 17756 2924 17808
rect 4160 17756 4212 17808
rect 5448 17756 5500 17808
rect 7288 17756 7340 17808
rect 6000 17688 6052 17740
rect 7012 17688 7064 17740
rect 8944 17688 8996 17740
rect 9220 17731 9272 17740
rect 9220 17697 9229 17731
rect 9229 17697 9263 17731
rect 9263 17697 9272 17731
rect 9220 17688 9272 17697
rect 756 17620 808 17672
rect 1492 17620 1544 17672
rect 2688 17620 2740 17672
rect 5172 17663 5224 17672
rect 2872 17552 2924 17604
rect 2780 17527 2832 17536
rect 2780 17493 2789 17527
rect 2789 17493 2823 17527
rect 2823 17493 2832 17527
rect 5172 17629 5181 17663
rect 5181 17629 5215 17663
rect 5215 17629 5224 17663
rect 5172 17620 5224 17629
rect 3884 17552 3936 17604
rect 2780 17484 2832 17493
rect 4344 17484 4396 17536
rect 4436 17484 4488 17536
rect 6552 17620 6604 17672
rect 8484 17620 8536 17672
rect 11152 17663 11204 17672
rect 11152 17629 11186 17663
rect 11186 17629 11204 17663
rect 11152 17620 11204 17629
rect 5632 17552 5684 17604
rect 5908 17484 5960 17536
rect 6736 17484 6788 17536
rect 7288 17527 7340 17536
rect 7288 17493 7297 17527
rect 7297 17493 7331 17527
rect 7331 17493 7340 17527
rect 7288 17484 7340 17493
rect 7472 17484 7524 17536
rect 9680 17552 9732 17604
rect 9864 17552 9916 17604
rect 14740 17756 14792 17808
rect 13084 17731 13136 17740
rect 13084 17697 13093 17731
rect 13093 17697 13127 17731
rect 13127 17697 13136 17731
rect 13084 17688 13136 17697
rect 16488 17833 16497 17867
rect 16497 17833 16531 17867
rect 16531 17833 16540 17867
rect 16488 17824 16540 17833
rect 15108 17731 15160 17740
rect 15108 17697 15117 17731
rect 15117 17697 15151 17731
rect 15151 17697 15160 17731
rect 15108 17688 15160 17697
rect 13360 17620 13412 17672
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 12164 17552 12216 17604
rect 13636 17552 13688 17604
rect 15844 17620 15896 17672
rect 16948 17620 17000 17672
rect 14648 17552 14700 17604
rect 10508 17484 10560 17536
rect 12624 17484 12676 17536
rect 13084 17484 13136 17536
rect 15016 17484 15068 17536
rect 15108 17484 15160 17536
rect 17592 17688 17644 17740
rect 17960 17688 18012 17740
rect 18328 17688 18380 17740
rect 20352 17824 20404 17876
rect 20536 17824 20588 17876
rect 20904 17824 20956 17876
rect 19892 17688 19944 17740
rect 20352 17663 20404 17672
rect 20352 17629 20361 17663
rect 20361 17629 20395 17663
rect 20395 17629 20404 17663
rect 20352 17620 20404 17629
rect 20076 17552 20128 17604
rect 17408 17527 17460 17536
rect 17408 17493 17417 17527
rect 17417 17493 17451 17527
rect 17451 17493 17460 17527
rect 17408 17484 17460 17493
rect 18420 17527 18472 17536
rect 18420 17493 18429 17527
rect 18429 17493 18463 17527
rect 18463 17493 18472 17527
rect 18420 17484 18472 17493
rect 18604 17484 18656 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 1676 17323 1728 17332
rect 1676 17289 1685 17323
rect 1685 17289 1719 17323
rect 1719 17289 1728 17323
rect 1676 17280 1728 17289
rect 5264 17280 5316 17332
rect 5724 17280 5776 17332
rect 5908 17280 5960 17332
rect 6644 17280 6696 17332
rect 7012 17280 7064 17332
rect 2780 17212 2832 17264
rect 2228 17144 2280 17196
rect 3424 17144 3476 17196
rect 2688 17119 2740 17128
rect 2688 17085 2697 17119
rect 2697 17085 2731 17119
rect 2731 17085 2740 17119
rect 2688 17076 2740 17085
rect 3056 17076 3108 17128
rect 4804 17144 4856 17196
rect 7932 17212 7984 17264
rect 9312 17280 9364 17332
rect 9956 17280 10008 17332
rect 12072 17280 12124 17332
rect 13084 17280 13136 17332
rect 14648 17323 14700 17332
rect 14648 17289 14657 17323
rect 14657 17289 14691 17323
rect 14691 17289 14700 17323
rect 14648 17280 14700 17289
rect 15200 17280 15252 17332
rect 20720 17280 20772 17332
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 6276 17144 6328 17196
rect 6644 17187 6696 17196
rect 6644 17153 6653 17187
rect 6653 17153 6687 17187
rect 6687 17153 6696 17187
rect 6644 17144 6696 17153
rect 9312 17144 9364 17196
rect 9680 17187 9732 17196
rect 9680 17153 9689 17187
rect 9689 17153 9723 17187
rect 9723 17153 9732 17187
rect 9680 17144 9732 17153
rect 10048 17144 10100 17196
rect 4896 17076 4948 17128
rect 5172 17076 5224 17128
rect 8300 17119 8352 17128
rect 8300 17085 8309 17119
rect 8309 17085 8343 17119
rect 8343 17085 8352 17119
rect 8300 17076 8352 17085
rect 9220 17076 9272 17128
rect 1860 16940 1912 16992
rect 2412 16940 2464 16992
rect 9864 17076 9916 17128
rect 11244 17076 11296 17128
rect 11796 17144 11848 17196
rect 13360 17187 13412 17196
rect 13360 17153 13369 17187
rect 13369 17153 13403 17187
rect 13403 17153 13412 17187
rect 13360 17144 13412 17153
rect 13636 17144 13688 17196
rect 15292 17187 15344 17196
rect 12256 17076 12308 17128
rect 13544 17119 13596 17128
rect 13544 17085 13553 17119
rect 13553 17085 13587 17119
rect 13587 17085 13596 17119
rect 13544 17076 13596 17085
rect 15292 17153 15301 17187
rect 15301 17153 15335 17187
rect 15335 17153 15344 17187
rect 15292 17144 15344 17153
rect 15476 17144 15528 17196
rect 17132 17212 17184 17264
rect 18604 17144 18656 17196
rect 14280 17076 14332 17128
rect 4804 16940 4856 16992
rect 5172 16940 5224 16992
rect 9956 16940 10008 16992
rect 10692 16940 10744 16992
rect 13084 17008 13136 17060
rect 15568 17076 15620 17128
rect 16120 17119 16172 17128
rect 16120 17085 16129 17119
rect 16129 17085 16163 17119
rect 16163 17085 16172 17119
rect 16120 17076 16172 17085
rect 16212 17076 16264 17128
rect 19892 17187 19944 17196
rect 19892 17153 19901 17187
rect 19901 17153 19935 17187
rect 19935 17153 19944 17187
rect 19892 17144 19944 17153
rect 14372 16940 14424 16992
rect 15384 17008 15436 17060
rect 15844 17008 15896 17060
rect 16304 16940 16356 16992
rect 16580 16940 16632 16992
rect 20628 17076 20680 17128
rect 17960 17051 18012 17060
rect 17960 17017 17969 17051
rect 17969 17017 18003 17051
rect 18003 17017 18012 17051
rect 17960 17008 18012 17017
rect 20536 16983 20588 16992
rect 20536 16949 20545 16983
rect 20545 16949 20579 16983
rect 20579 16949 20588 16983
rect 20536 16940 20588 16949
rect 20812 16940 20864 16992
rect 20996 16983 21048 16992
rect 20996 16949 21005 16983
rect 21005 16949 21039 16983
rect 21039 16949 21048 16983
rect 20996 16940 21048 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 3424 16736 3476 16788
rect 2780 16668 2832 16720
rect 4436 16668 4488 16720
rect 4344 16643 4396 16652
rect 4344 16609 4353 16643
rect 4353 16609 4387 16643
rect 4387 16609 4396 16643
rect 4344 16600 4396 16609
rect 5172 16736 5224 16788
rect 6276 16779 6328 16788
rect 6276 16745 6285 16779
rect 6285 16745 6319 16779
rect 6319 16745 6328 16779
rect 6276 16736 6328 16745
rect 7288 16736 7340 16788
rect 7748 16736 7800 16788
rect 9220 16736 9272 16788
rect 9312 16668 9364 16720
rect 4896 16643 4948 16652
rect 1952 16532 2004 16584
rect 2964 16532 3016 16584
rect 3884 16532 3936 16584
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 4896 16609 4905 16643
rect 4905 16609 4939 16643
rect 4939 16609 4948 16643
rect 4896 16600 4948 16609
rect 7932 16643 7984 16652
rect 4528 16532 4580 16584
rect 6552 16575 6604 16584
rect 6552 16541 6561 16575
rect 6561 16541 6595 16575
rect 6595 16541 6604 16575
rect 6552 16532 6604 16541
rect 7932 16609 7941 16643
rect 7941 16609 7975 16643
rect 7975 16609 7984 16643
rect 7932 16600 7984 16609
rect 8116 16643 8168 16652
rect 8116 16609 8125 16643
rect 8125 16609 8159 16643
rect 8159 16609 8168 16643
rect 8116 16600 8168 16609
rect 11152 16600 11204 16652
rect 12716 16668 12768 16720
rect 13268 16736 13320 16788
rect 15752 16779 15804 16788
rect 14004 16668 14056 16720
rect 14280 16668 14332 16720
rect 11888 16643 11940 16652
rect 8392 16532 8444 16584
rect 8668 16532 8720 16584
rect 8760 16532 8812 16584
rect 9680 16532 9732 16584
rect 10968 16532 11020 16584
rect 11888 16609 11897 16643
rect 11897 16609 11931 16643
rect 11931 16609 11940 16643
rect 11888 16600 11940 16609
rect 13360 16600 13412 16652
rect 13544 16600 13596 16652
rect 15752 16745 15761 16779
rect 15761 16745 15795 16779
rect 15795 16745 15804 16779
rect 15752 16736 15804 16745
rect 17040 16736 17092 16788
rect 18420 16736 18472 16788
rect 16304 16643 16356 16652
rect 16304 16609 16313 16643
rect 16313 16609 16347 16643
rect 16347 16609 16356 16643
rect 16304 16600 16356 16609
rect 17132 16643 17184 16652
rect 17132 16609 17141 16643
rect 17141 16609 17175 16643
rect 17175 16609 17184 16643
rect 17132 16600 17184 16609
rect 18788 16643 18840 16652
rect 18788 16609 18797 16643
rect 18797 16609 18831 16643
rect 18831 16609 18840 16643
rect 18788 16600 18840 16609
rect 21272 16668 21324 16720
rect 12532 16532 12584 16584
rect 4344 16464 4396 16516
rect 940 16396 992 16448
rect 1584 16439 1636 16448
rect 1584 16405 1593 16439
rect 1593 16405 1627 16439
rect 1627 16405 1636 16439
rect 1584 16396 1636 16405
rect 2044 16439 2096 16448
rect 2044 16405 2053 16439
rect 2053 16405 2087 16439
rect 2087 16405 2096 16439
rect 2044 16396 2096 16405
rect 3424 16396 3476 16448
rect 4068 16396 4120 16448
rect 4436 16396 4488 16448
rect 10692 16464 10744 16516
rect 10784 16464 10836 16516
rect 12624 16507 12676 16516
rect 7196 16439 7248 16448
rect 7196 16405 7205 16439
rect 7205 16405 7239 16439
rect 7239 16405 7248 16439
rect 7196 16396 7248 16405
rect 7840 16439 7892 16448
rect 7840 16405 7849 16439
rect 7849 16405 7883 16439
rect 7883 16405 7892 16439
rect 7840 16396 7892 16405
rect 9864 16396 9916 16448
rect 10324 16396 10376 16448
rect 11244 16396 11296 16448
rect 12624 16473 12633 16507
rect 12633 16473 12667 16507
rect 12667 16473 12676 16507
rect 12624 16464 12676 16473
rect 13728 16464 13780 16516
rect 16580 16532 16632 16584
rect 17408 16575 17460 16584
rect 17408 16541 17442 16575
rect 17442 16541 17460 16575
rect 17408 16532 17460 16541
rect 17224 16464 17276 16516
rect 13360 16439 13412 16448
rect 13360 16405 13369 16439
rect 13369 16405 13403 16439
rect 13403 16405 13412 16439
rect 13360 16396 13412 16405
rect 14004 16396 14056 16448
rect 16396 16396 16448 16448
rect 20628 16532 20680 16584
rect 20996 16532 21048 16584
rect 19800 16464 19852 16516
rect 21088 16396 21140 16448
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 2136 16235 2188 16244
rect 2136 16201 2145 16235
rect 2145 16201 2179 16235
rect 2179 16201 2188 16235
rect 2136 16192 2188 16201
rect 3148 16235 3200 16244
rect 3148 16201 3157 16235
rect 3157 16201 3191 16235
rect 3191 16201 3200 16235
rect 3148 16192 3200 16201
rect 4528 16192 4580 16244
rect 8300 16235 8352 16244
rect 204 16124 256 16176
rect 6000 16167 6052 16176
rect 6000 16133 6009 16167
rect 6009 16133 6043 16167
rect 6043 16133 6052 16167
rect 8300 16201 8309 16235
rect 8309 16201 8343 16235
rect 8343 16201 8352 16235
rect 8300 16192 8352 16201
rect 10784 16192 10836 16244
rect 11060 16192 11112 16244
rect 13360 16192 13412 16244
rect 13728 16192 13780 16244
rect 14556 16192 14608 16244
rect 15844 16192 15896 16244
rect 16120 16192 16172 16244
rect 6000 16124 6052 16133
rect 1676 16056 1728 16108
rect 1768 16056 1820 16108
rect 3976 16099 4028 16108
rect 3976 16065 3985 16099
rect 3985 16065 4019 16099
rect 4019 16065 4028 16099
rect 3976 16056 4028 16065
rect 4068 16056 4120 16108
rect 4436 15988 4488 16040
rect 5448 16031 5500 16040
rect 5448 15997 5457 16031
rect 5457 15997 5491 16031
rect 5491 15997 5500 16031
rect 5448 15988 5500 15997
rect 5540 15988 5592 16040
rect 4804 15920 4856 15972
rect 1584 15895 1636 15904
rect 1584 15861 1593 15895
rect 1593 15861 1627 15895
rect 1627 15861 1636 15895
rect 1584 15852 1636 15861
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 6092 15920 6144 15972
rect 7104 16056 7156 16108
rect 8300 16056 8352 16108
rect 12440 16124 12492 16176
rect 12808 16056 12860 16108
rect 12992 16056 13044 16108
rect 13360 16056 13412 16108
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 10416 16031 10468 16040
rect 10416 15997 10425 16031
rect 10425 15997 10459 16031
rect 10459 15997 10468 16031
rect 10416 15988 10468 15997
rect 15476 16124 15528 16176
rect 13820 16056 13872 16108
rect 16948 16192 17000 16244
rect 19892 16235 19944 16244
rect 13912 15988 13964 16040
rect 14280 15988 14332 16040
rect 14740 16031 14792 16040
rect 14740 15997 14749 16031
rect 14749 15997 14783 16031
rect 14783 15997 14792 16031
rect 14740 15988 14792 15997
rect 7012 15920 7064 15972
rect 7104 15920 7156 15972
rect 7288 15852 7340 15904
rect 9588 15852 9640 15904
rect 10140 15852 10192 15904
rect 11152 15852 11204 15904
rect 13360 15920 13412 15972
rect 13636 15852 13688 15904
rect 16948 15988 17000 16040
rect 17132 16124 17184 16176
rect 19892 16201 19901 16235
rect 19901 16201 19935 16235
rect 19935 16201 19944 16235
rect 19892 16192 19944 16201
rect 18972 16124 19024 16176
rect 19064 16124 19116 16176
rect 20904 16192 20956 16244
rect 20260 16056 20312 16108
rect 17040 15852 17092 15904
rect 21732 15988 21784 16040
rect 20628 15920 20680 15972
rect 19984 15852 20036 15904
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 1492 15648 1544 15700
rect 2596 15648 2648 15700
rect 3240 15691 3292 15700
rect 3240 15657 3249 15691
rect 3249 15657 3283 15691
rect 3283 15657 3292 15691
rect 3240 15648 3292 15657
rect 4344 15691 4396 15700
rect 4344 15657 4353 15691
rect 4353 15657 4387 15691
rect 4387 15657 4396 15691
rect 4344 15648 4396 15657
rect 1400 15487 1452 15496
rect 1400 15453 1409 15487
rect 1409 15453 1443 15487
rect 1443 15453 1452 15487
rect 1400 15444 1452 15453
rect 3240 15512 3292 15564
rect 4896 15512 4948 15564
rect 5172 15512 5224 15564
rect 2136 15376 2188 15428
rect 2964 15444 3016 15496
rect 3884 15487 3936 15496
rect 3884 15453 3893 15487
rect 3893 15453 3927 15487
rect 3927 15453 3936 15487
rect 3884 15444 3936 15453
rect 4988 15487 5040 15496
rect 4988 15453 4997 15487
rect 4997 15453 5031 15487
rect 5031 15453 5040 15487
rect 4988 15444 5040 15453
rect 5448 15444 5500 15496
rect 5724 15444 5776 15496
rect 6092 15444 6144 15496
rect 8300 15648 8352 15700
rect 8576 15691 8628 15700
rect 8576 15657 8585 15691
rect 8585 15657 8619 15691
rect 8619 15657 8628 15691
rect 8576 15648 8628 15657
rect 9312 15648 9364 15700
rect 8392 15580 8444 15632
rect 10416 15648 10468 15700
rect 10784 15648 10836 15700
rect 12532 15648 12584 15700
rect 13728 15691 13780 15700
rect 13728 15657 13737 15691
rect 13737 15657 13771 15691
rect 13771 15657 13780 15691
rect 13728 15648 13780 15657
rect 17132 15691 17184 15700
rect 17132 15657 17141 15691
rect 17141 15657 17175 15691
rect 17175 15657 17184 15691
rect 17132 15648 17184 15657
rect 18512 15648 18564 15700
rect 20076 15648 20128 15700
rect 4160 15376 4212 15428
rect 4804 15376 4856 15428
rect 7840 15376 7892 15428
rect 10416 15512 10468 15564
rect 8668 15444 8720 15496
rect 8484 15376 8536 15428
rect 8576 15376 8628 15428
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 4528 15308 4580 15360
rect 6920 15308 6972 15360
rect 7380 15308 7432 15360
rect 7748 15351 7800 15360
rect 7748 15317 7757 15351
rect 7757 15317 7791 15351
rect 7791 15317 7800 15351
rect 7748 15308 7800 15317
rect 8300 15308 8352 15360
rect 10784 15444 10836 15496
rect 10876 15444 10928 15496
rect 11152 15512 11204 15564
rect 11888 15555 11940 15564
rect 11888 15521 11897 15555
rect 11897 15521 11931 15555
rect 11931 15521 11940 15555
rect 11888 15512 11940 15521
rect 15568 15580 15620 15632
rect 17224 15580 17276 15632
rect 14648 15512 14700 15564
rect 12532 15487 12584 15496
rect 12532 15453 12541 15487
rect 12541 15453 12575 15487
rect 12575 15453 12584 15487
rect 12532 15444 12584 15453
rect 13360 15487 13412 15496
rect 13360 15453 13369 15487
rect 13369 15453 13403 15487
rect 13403 15453 13412 15487
rect 13360 15444 13412 15453
rect 19432 15512 19484 15564
rect 19892 15555 19944 15564
rect 19892 15521 19901 15555
rect 19901 15521 19935 15555
rect 19935 15521 19944 15555
rect 19892 15512 19944 15521
rect 18236 15444 18288 15496
rect 9772 15376 9824 15428
rect 9680 15308 9732 15360
rect 11060 15308 11112 15360
rect 11980 15308 12032 15360
rect 12440 15376 12492 15428
rect 13268 15351 13320 15360
rect 13268 15317 13277 15351
rect 13277 15317 13311 15351
rect 13311 15317 13320 15351
rect 13268 15308 13320 15317
rect 14372 15351 14424 15360
rect 14372 15317 14381 15351
rect 14381 15317 14415 15351
rect 14415 15317 14424 15351
rect 14372 15308 14424 15317
rect 15108 15308 15160 15360
rect 18052 15351 18104 15360
rect 18052 15317 18061 15351
rect 18061 15317 18095 15351
rect 18095 15317 18104 15351
rect 18052 15308 18104 15317
rect 19616 15351 19668 15360
rect 19616 15317 19625 15351
rect 19625 15317 19659 15351
rect 19659 15317 19668 15351
rect 19616 15308 19668 15317
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 1492 15104 1544 15156
rect 3976 15104 4028 15156
rect 4988 15104 5040 15156
rect 5264 15104 5316 15156
rect 8484 15147 8536 15156
rect 8484 15113 8493 15147
rect 8493 15113 8527 15147
rect 8527 15113 8536 15147
rect 8484 15104 8536 15113
rect 9036 15104 9088 15156
rect 9312 15104 9364 15156
rect 10324 15104 10376 15156
rect 11060 15104 11112 15156
rect 11888 15147 11940 15156
rect 11888 15113 11897 15147
rect 11897 15113 11931 15147
rect 11931 15113 11940 15147
rect 11888 15104 11940 15113
rect 1216 14968 1268 15020
rect 5172 15036 5224 15088
rect 1492 14807 1544 14816
rect 1492 14773 1501 14807
rect 1501 14773 1535 14807
rect 1535 14773 1544 14807
rect 1492 14764 1544 14773
rect 2872 14968 2924 15020
rect 5448 14968 5500 15020
rect 7656 15036 7708 15088
rect 9680 15036 9732 15088
rect 10048 15079 10100 15088
rect 10048 15045 10057 15079
rect 10057 15045 10091 15079
rect 10091 15045 10100 15079
rect 10048 15036 10100 15045
rect 11244 15036 11296 15088
rect 11704 15036 11756 15088
rect 12900 15104 12952 15156
rect 13268 15104 13320 15156
rect 13544 15104 13596 15156
rect 15108 15104 15160 15156
rect 15476 15147 15528 15156
rect 15476 15113 15485 15147
rect 15485 15113 15519 15147
rect 15519 15113 15528 15147
rect 15476 15104 15528 15113
rect 16948 15104 17000 15156
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 9036 14943 9088 14952
rect 9036 14909 9045 14943
rect 9045 14909 9079 14943
rect 9079 14909 9088 14943
rect 9036 14900 9088 14909
rect 10600 14943 10652 14952
rect 10600 14909 10609 14943
rect 10609 14909 10643 14943
rect 10643 14909 10652 14943
rect 10600 14900 10652 14909
rect 12992 15036 13044 15088
rect 14372 15079 14424 15088
rect 13360 14968 13412 15020
rect 13636 14968 13688 15020
rect 14372 15045 14406 15079
rect 14406 15045 14424 15079
rect 14372 15036 14424 15045
rect 19432 15147 19484 15156
rect 12348 14900 12400 14952
rect 13728 14943 13780 14952
rect 13728 14909 13737 14943
rect 13737 14909 13771 14943
rect 13771 14909 13780 14943
rect 14740 14968 14792 15020
rect 13728 14900 13780 14909
rect 12900 14832 12952 14884
rect 16396 14900 16448 14952
rect 17132 15036 17184 15088
rect 19432 15113 19441 15147
rect 19441 15113 19475 15147
rect 19475 15113 19484 15147
rect 19432 15104 19484 15113
rect 21272 15104 21324 15156
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 17224 14943 17276 14952
rect 17224 14909 17233 14943
rect 17233 14909 17267 14943
rect 17267 14909 17276 14943
rect 17500 14968 17552 15020
rect 17960 14968 18012 15020
rect 20628 15036 20680 15088
rect 19432 14968 19484 15020
rect 17224 14900 17276 14909
rect 17776 14832 17828 14884
rect 4160 14764 4212 14816
rect 4344 14764 4396 14816
rect 7380 14764 7432 14816
rect 8392 14764 8444 14816
rect 17500 14764 17552 14816
rect 20536 14900 20588 14952
rect 19064 14764 19116 14816
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 2320 14560 2372 14612
rect 5448 14603 5500 14612
rect 5448 14569 5457 14603
rect 5457 14569 5491 14603
rect 5491 14569 5500 14603
rect 5448 14560 5500 14569
rect 5908 14560 5960 14612
rect 6552 14560 6604 14612
rect 8300 14560 8352 14612
rect 2872 14492 2924 14544
rect 3792 14424 3844 14476
rect 2412 14356 2464 14408
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 2320 14220 2372 14272
rect 3056 14263 3108 14272
rect 3056 14229 3065 14263
rect 3065 14229 3099 14263
rect 3099 14229 3108 14263
rect 3056 14220 3108 14229
rect 3148 14263 3200 14272
rect 3148 14229 3157 14263
rect 3157 14229 3191 14263
rect 3191 14229 3200 14263
rect 3792 14263 3844 14272
rect 3148 14220 3200 14229
rect 3792 14229 3801 14263
rect 3801 14229 3835 14263
rect 3835 14229 3844 14263
rect 3792 14220 3844 14229
rect 5172 14467 5224 14476
rect 5172 14433 5181 14467
rect 5181 14433 5215 14467
rect 5215 14433 5224 14467
rect 5172 14424 5224 14433
rect 4620 14356 4672 14408
rect 5724 14356 5776 14408
rect 6000 14356 6052 14408
rect 7104 14356 7156 14408
rect 10600 14560 10652 14612
rect 12072 14560 12124 14612
rect 12440 14560 12492 14612
rect 13820 14560 13872 14612
rect 16028 14560 16080 14612
rect 18880 14560 18932 14612
rect 21916 14560 21968 14612
rect 14648 14467 14700 14476
rect 14648 14433 14657 14467
rect 14657 14433 14691 14467
rect 14691 14433 14700 14467
rect 14648 14424 14700 14433
rect 17500 14467 17552 14476
rect 17500 14433 17509 14467
rect 17509 14433 17543 14467
rect 17543 14433 17552 14467
rect 17500 14424 17552 14433
rect 12992 14356 13044 14408
rect 15200 14356 15252 14408
rect 17132 14356 17184 14408
rect 17776 14399 17828 14408
rect 17776 14365 17785 14399
rect 17785 14365 17819 14399
rect 17819 14365 17828 14399
rect 17776 14356 17828 14365
rect 18052 14424 18104 14476
rect 18696 14424 18748 14476
rect 20536 14399 20588 14408
rect 20536 14365 20545 14399
rect 20545 14365 20579 14399
rect 20579 14365 20588 14399
rect 20536 14356 20588 14365
rect 6552 14288 6604 14340
rect 7472 14331 7524 14340
rect 7472 14297 7490 14331
rect 7490 14297 7524 14331
rect 7472 14288 7524 14297
rect 5448 14220 5500 14272
rect 8024 14263 8076 14272
rect 8024 14229 8033 14263
rect 8033 14229 8067 14263
rect 8067 14229 8076 14263
rect 8024 14220 8076 14229
rect 11152 14288 11204 14340
rect 11244 14331 11296 14340
rect 11244 14297 11262 14331
rect 11262 14297 11296 14331
rect 11244 14288 11296 14297
rect 11796 14220 11848 14272
rect 14556 14263 14608 14272
rect 14556 14229 14565 14263
rect 14565 14229 14599 14263
rect 14599 14229 14608 14263
rect 14556 14220 14608 14229
rect 17132 14263 17184 14272
rect 17132 14229 17141 14263
rect 17141 14229 17175 14263
rect 17175 14229 17184 14263
rect 17132 14220 17184 14229
rect 17408 14220 17460 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 3056 14016 3108 14068
rect 5540 14016 5592 14068
rect 6000 14059 6052 14068
rect 6000 14025 6009 14059
rect 6009 14025 6043 14059
rect 6043 14025 6052 14059
rect 6000 14016 6052 14025
rect 6552 14016 6604 14068
rect 8392 14059 8444 14068
rect 8392 14025 8401 14059
rect 8401 14025 8435 14059
rect 8435 14025 8444 14059
rect 8392 14016 8444 14025
rect 9128 14016 9180 14068
rect 10508 14016 10560 14068
rect 11888 14016 11940 14068
rect 11980 14016 12032 14068
rect 13084 14016 13136 14068
rect 13636 14016 13688 14068
rect 14648 14016 14700 14068
rect 17408 14059 17460 14068
rect 1768 13880 1820 13932
rect 2780 13880 2832 13932
rect 3056 13923 3108 13932
rect 3056 13889 3065 13923
rect 3065 13889 3099 13923
rect 3099 13889 3108 13923
rect 3056 13880 3108 13889
rect 1584 13787 1636 13796
rect 1584 13753 1593 13787
rect 1593 13753 1627 13787
rect 1627 13753 1636 13787
rect 1584 13744 1636 13753
rect 3148 13812 3200 13864
rect 4344 13880 4396 13932
rect 5724 13948 5776 14000
rect 8484 13948 8536 14000
rect 10232 13948 10284 14000
rect 4712 13880 4764 13932
rect 5172 13880 5224 13932
rect 7012 13880 7064 13932
rect 10048 13923 10100 13932
rect 10048 13889 10066 13923
rect 10066 13889 10100 13923
rect 10048 13880 10100 13889
rect 11152 13880 11204 13932
rect 12440 13880 12492 13932
rect 12992 13948 13044 14000
rect 13820 13880 13872 13932
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 17592 14016 17644 14068
rect 19984 14059 20036 14068
rect 16396 13880 16448 13932
rect 17500 13948 17552 14000
rect 19064 13948 19116 14000
rect 17132 13880 17184 13932
rect 19984 14025 19993 14059
rect 19993 14025 20027 14059
rect 20027 14025 20036 14059
rect 19984 14016 20036 14025
rect 21180 14016 21232 14068
rect 21364 14059 21416 14068
rect 21364 14025 21373 14059
rect 21373 14025 21407 14059
rect 21407 14025 21416 14059
rect 21364 14016 21416 14025
rect 3976 13812 4028 13864
rect 4252 13812 4304 13864
rect 7564 13855 7616 13864
rect 7564 13821 7573 13855
rect 7573 13821 7607 13855
rect 7607 13821 7616 13855
rect 7564 13812 7616 13821
rect 11060 13812 11112 13864
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 12348 13812 12400 13864
rect 16948 13812 17000 13864
rect 17040 13812 17092 13864
rect 19064 13855 19116 13864
rect 19064 13821 19073 13855
rect 19073 13821 19107 13855
rect 19107 13821 19116 13855
rect 19064 13812 19116 13821
rect 8668 13744 8720 13796
rect 16764 13744 16816 13796
rect 3884 13676 3936 13728
rect 6828 13676 6880 13728
rect 17592 13676 17644 13728
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 2964 13472 3016 13524
rect 4712 13472 4764 13524
rect 4344 13447 4396 13456
rect 1584 13311 1636 13320
rect 1584 13277 1593 13311
rect 1593 13277 1627 13311
rect 1627 13277 1636 13311
rect 1584 13268 1636 13277
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2596 13268 2648 13320
rect 4344 13413 4353 13447
rect 4353 13413 4387 13447
rect 4387 13413 4396 13447
rect 4344 13404 4396 13413
rect 6736 13472 6788 13524
rect 8576 13472 8628 13524
rect 10048 13472 10100 13524
rect 11152 13472 11204 13524
rect 14556 13472 14608 13524
rect 16396 13515 16448 13524
rect 16396 13481 16405 13515
rect 16405 13481 16439 13515
rect 16439 13481 16448 13515
rect 16396 13472 16448 13481
rect 20812 13472 20864 13524
rect 21456 13472 21508 13524
rect 3516 13336 3568 13388
rect 7564 13404 7616 13456
rect 5724 13379 5776 13388
rect 5724 13345 5733 13379
rect 5733 13345 5767 13379
rect 5767 13345 5776 13379
rect 5724 13336 5776 13345
rect 6552 13379 6604 13388
rect 6552 13345 6561 13379
rect 6561 13345 6595 13379
rect 6595 13345 6604 13379
rect 6552 13336 6604 13345
rect 3976 13268 4028 13320
rect 1492 13132 1544 13184
rect 2412 13132 2464 13184
rect 5632 13268 5684 13320
rect 7012 13268 7064 13320
rect 7472 13268 7524 13320
rect 8668 13336 8720 13388
rect 9128 13268 9180 13320
rect 12440 13379 12492 13388
rect 12440 13345 12449 13379
rect 12449 13345 12483 13379
rect 12483 13345 12492 13379
rect 12440 13336 12492 13345
rect 13820 13336 13872 13388
rect 10324 13268 10376 13320
rect 12348 13268 12400 13320
rect 20352 13404 20404 13456
rect 18696 13336 18748 13388
rect 5356 13200 5408 13252
rect 4712 13132 4764 13184
rect 7840 13132 7892 13184
rect 8484 13200 8536 13252
rect 11244 13200 11296 13252
rect 12532 13200 12584 13252
rect 13360 13243 13412 13252
rect 13360 13209 13369 13243
rect 13369 13209 13403 13243
rect 13403 13209 13412 13243
rect 13360 13200 13412 13209
rect 15752 13200 15804 13252
rect 16764 13268 16816 13320
rect 19984 13200 20036 13252
rect 9772 13132 9824 13184
rect 12256 13132 12308 13184
rect 17684 13175 17736 13184
rect 17684 13141 17693 13175
rect 17693 13141 17727 13175
rect 17727 13141 17736 13175
rect 17684 13132 17736 13141
rect 18052 13132 18104 13184
rect 19616 13132 19668 13184
rect 19892 13175 19944 13184
rect 19892 13141 19901 13175
rect 19901 13141 19935 13175
rect 19935 13141 19944 13175
rect 19892 13132 19944 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 1584 12928 1636 12980
rect 4712 12971 4764 12980
rect 4712 12937 4721 12971
rect 4721 12937 4755 12971
rect 4755 12937 4764 12971
rect 4712 12928 4764 12937
rect 8024 12928 8076 12980
rect 8668 12971 8720 12980
rect 8668 12937 8677 12971
rect 8677 12937 8711 12971
rect 8711 12937 8720 12971
rect 8668 12928 8720 12937
rect 10324 12971 10376 12980
rect 10324 12937 10333 12971
rect 10333 12937 10367 12971
rect 10367 12937 10376 12971
rect 10324 12928 10376 12937
rect 12164 12928 12216 12980
rect 12900 12971 12952 12980
rect 12900 12937 12909 12971
rect 12909 12937 12943 12971
rect 12943 12937 12952 12971
rect 12900 12928 12952 12937
rect 14280 12928 14332 12980
rect 18144 12928 18196 12980
rect 18696 12971 18748 12980
rect 18696 12937 18705 12971
rect 18705 12937 18739 12971
rect 18739 12937 18748 12971
rect 18696 12928 18748 12937
rect 19984 12971 20036 12980
rect 19984 12937 19993 12971
rect 19993 12937 20027 12971
rect 20027 12937 20036 12971
rect 19984 12928 20036 12937
rect 2228 12860 2280 12912
rect 4068 12860 4120 12912
rect 5172 12860 5224 12912
rect 5724 12860 5776 12912
rect 2688 12792 2740 12844
rect 3516 12792 3568 12844
rect 3884 12792 3936 12844
rect 4344 12724 4396 12776
rect 6920 12792 6972 12844
rect 5908 12767 5960 12776
rect 5908 12733 5917 12767
rect 5917 12733 5951 12767
rect 5951 12733 5960 12767
rect 5908 12724 5960 12733
rect 7564 12835 7616 12844
rect 7564 12801 7598 12835
rect 7598 12801 7616 12835
rect 7840 12860 7892 12912
rect 11796 12903 11848 12912
rect 11796 12869 11830 12903
rect 11830 12869 11848 12903
rect 11796 12860 11848 12869
rect 7564 12792 7616 12801
rect 9772 12792 9824 12844
rect 8300 12724 8352 12776
rect 9956 12724 10008 12776
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 6644 12656 6696 12708
rect 15476 12860 15528 12912
rect 17960 12860 18012 12912
rect 19064 12860 19116 12912
rect 17592 12835 17644 12844
rect 17592 12801 17626 12835
rect 17626 12801 17644 12835
rect 17592 12792 17644 12801
rect 21088 12835 21140 12844
rect 21088 12801 21106 12835
rect 21106 12801 21140 12835
rect 21088 12792 21140 12801
rect 15292 12724 15344 12776
rect 2136 12631 2188 12640
rect 2136 12597 2145 12631
rect 2145 12597 2179 12631
rect 2179 12597 2188 12631
rect 2136 12588 2188 12597
rect 3332 12631 3384 12640
rect 3332 12597 3341 12631
rect 3341 12597 3375 12631
rect 3375 12597 3384 12631
rect 3332 12588 3384 12597
rect 4620 12588 4672 12640
rect 9588 12588 9640 12640
rect 12164 12588 12216 12640
rect 15384 12656 15436 12708
rect 16028 12656 16080 12708
rect 13820 12631 13872 12640
rect 13820 12597 13829 12631
rect 13829 12597 13863 12631
rect 13863 12597 13872 12631
rect 13820 12588 13872 12597
rect 14280 12588 14332 12640
rect 16948 12588 17000 12640
rect 18972 12588 19024 12640
rect 19708 12588 19760 12640
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 1400 12427 1452 12436
rect 1400 12393 1409 12427
rect 1409 12393 1443 12427
rect 1443 12393 1452 12427
rect 1400 12384 1452 12393
rect 4068 12384 4120 12436
rect 2504 12359 2556 12368
rect 2504 12325 2513 12359
rect 2513 12325 2547 12359
rect 2547 12325 2556 12359
rect 2504 12316 2556 12325
rect 3516 12316 3568 12368
rect 5080 12384 5132 12436
rect 5908 12384 5960 12436
rect 6552 12384 6604 12436
rect 15384 12384 15436 12436
rect 15752 12384 15804 12436
rect 17684 12384 17736 12436
rect 18052 12384 18104 12436
rect 7472 12316 7524 12368
rect 8116 12316 8168 12368
rect 17592 12316 17644 12368
rect 1400 12180 1452 12232
rect 2964 12248 3016 12300
rect 8024 12248 8076 12300
rect 16948 12248 17000 12300
rect 17960 12248 18012 12300
rect 19708 12291 19760 12300
rect 19708 12257 19717 12291
rect 19717 12257 19751 12291
rect 19751 12257 19760 12291
rect 19708 12248 19760 12257
rect 2412 12180 2464 12232
rect 3424 12180 3476 12232
rect 5724 12180 5776 12232
rect 7196 12223 7248 12232
rect 7196 12189 7214 12223
rect 7214 12189 7248 12223
rect 7196 12180 7248 12189
rect 8668 12180 8720 12232
rect 11060 12180 11112 12232
rect 11520 12180 11572 12232
rect 11888 12180 11940 12232
rect 12348 12180 12400 12232
rect 12992 12180 13044 12232
rect 16028 12223 16080 12232
rect 2872 12112 2924 12164
rect 3056 12112 3108 12164
rect 3332 12112 3384 12164
rect 4804 12112 4856 12164
rect 1584 12044 1636 12096
rect 3516 12044 3568 12096
rect 3792 12087 3844 12096
rect 3792 12053 3801 12087
rect 3801 12053 3835 12087
rect 3835 12053 3844 12087
rect 3792 12044 3844 12053
rect 6000 12044 6052 12096
rect 8300 12112 8352 12164
rect 10876 12155 10928 12164
rect 10876 12121 10894 12155
rect 10894 12121 10928 12155
rect 10876 12112 10928 12121
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 8208 12087 8260 12096
rect 8208 12053 8217 12087
rect 8217 12053 8251 12087
rect 8251 12053 8260 12087
rect 8208 12044 8260 12053
rect 8392 12044 8444 12096
rect 9772 12087 9824 12096
rect 9772 12053 9781 12087
rect 9781 12053 9815 12087
rect 9815 12053 9824 12087
rect 9772 12044 9824 12053
rect 10508 12044 10560 12096
rect 13820 12112 13872 12164
rect 15384 12112 15436 12164
rect 16028 12189 16037 12223
rect 16037 12189 16071 12223
rect 16071 12189 16080 12223
rect 16028 12180 16080 12189
rect 16396 12180 16448 12232
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 19616 12223 19668 12232
rect 19616 12189 19625 12223
rect 19625 12189 19659 12223
rect 19659 12189 19668 12223
rect 19616 12180 19668 12189
rect 13176 12087 13228 12096
rect 13176 12053 13185 12087
rect 13185 12053 13219 12087
rect 13219 12053 13228 12087
rect 13176 12044 13228 12053
rect 13636 12087 13688 12096
rect 13636 12053 13645 12087
rect 13645 12053 13679 12087
rect 13679 12053 13688 12087
rect 13636 12044 13688 12053
rect 13728 12044 13780 12096
rect 20720 12044 20772 12096
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 1676 11840 1728 11892
rect 2228 11704 2280 11756
rect 5816 11840 5868 11892
rect 2964 11747 3016 11756
rect 2964 11713 2973 11747
rect 2973 11713 3007 11747
rect 3007 11713 3016 11747
rect 2964 11704 3016 11713
rect 3792 11704 3844 11756
rect 3148 11636 3200 11688
rect 5724 11704 5776 11756
rect 6000 11747 6052 11756
rect 6000 11713 6009 11747
rect 6009 11713 6043 11747
rect 6043 11713 6052 11747
rect 6000 11704 6052 11713
rect 6736 11815 6788 11824
rect 6736 11781 6745 11815
rect 6745 11781 6779 11815
rect 6779 11781 6788 11815
rect 6736 11772 6788 11781
rect 7840 11772 7892 11824
rect 8024 11840 8076 11892
rect 9956 11840 10008 11892
rect 10048 11772 10100 11824
rect 12256 11840 12308 11892
rect 13728 11840 13780 11892
rect 15292 11840 15344 11892
rect 15476 11840 15528 11892
rect 21088 11840 21140 11892
rect 11888 11772 11940 11824
rect 2596 11568 2648 11620
rect 3884 11568 3936 11620
rect 6000 11568 6052 11620
rect 2780 11543 2832 11552
rect 2780 11509 2789 11543
rect 2789 11509 2823 11543
rect 2823 11509 2832 11543
rect 2780 11500 2832 11509
rect 3056 11500 3108 11552
rect 3424 11500 3476 11552
rect 3976 11500 4028 11552
rect 4804 11500 4856 11552
rect 8300 11500 8352 11552
rect 8576 11500 8628 11552
rect 9312 11500 9364 11552
rect 10876 11704 10928 11756
rect 12624 11704 12676 11756
rect 12992 11704 13044 11756
rect 13452 11747 13504 11756
rect 13452 11713 13461 11747
rect 13461 11713 13495 11747
rect 13495 11713 13504 11747
rect 13452 11704 13504 11713
rect 19892 11772 19944 11824
rect 14280 11704 14332 11756
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 9864 11636 9916 11688
rect 10508 11679 10560 11688
rect 10508 11645 10517 11679
rect 10517 11645 10551 11679
rect 10551 11645 10560 11679
rect 10508 11636 10560 11645
rect 17316 11611 17368 11620
rect 11980 11500 12032 11552
rect 12808 11543 12860 11552
rect 12808 11509 12817 11543
rect 12817 11509 12851 11543
rect 12851 11509 12860 11543
rect 12808 11500 12860 11509
rect 14464 11500 14516 11552
rect 14740 11500 14792 11552
rect 17316 11577 17325 11611
rect 17325 11577 17359 11611
rect 17359 11577 17368 11611
rect 21364 11747 21416 11756
rect 21364 11713 21373 11747
rect 21373 11713 21407 11747
rect 21407 11713 21416 11747
rect 21364 11704 21416 11713
rect 19064 11636 19116 11688
rect 17316 11568 17368 11577
rect 17500 11500 17552 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2964 11296 3016 11348
rect 4436 11296 4488 11348
rect 5816 11296 5868 11348
rect 7932 11296 7984 11348
rect 8208 11296 8260 11348
rect 9404 11296 9456 11348
rect 13636 11296 13688 11348
rect 15108 11339 15160 11348
rect 15108 11305 15117 11339
rect 15117 11305 15151 11339
rect 15151 11305 15160 11339
rect 15108 11296 15160 11305
rect 18236 11296 18288 11348
rect 1860 11203 1912 11212
rect 1860 11169 1869 11203
rect 1869 11169 1903 11203
rect 1903 11169 1912 11203
rect 1860 11160 1912 11169
rect 3332 11228 3384 11280
rect 3240 11203 3292 11212
rect 3240 11169 3249 11203
rect 3249 11169 3283 11203
rect 3283 11169 3292 11203
rect 3240 11160 3292 11169
rect 3976 11160 4028 11212
rect 2136 11092 2188 11144
rect 4252 11024 4304 11076
rect 5448 11228 5500 11280
rect 6736 11228 6788 11280
rect 7840 11228 7892 11280
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 6000 11203 6052 11212
rect 6000 11169 6009 11203
rect 6009 11169 6043 11203
rect 6043 11169 6052 11203
rect 6000 11160 6052 11169
rect 8300 11160 8352 11212
rect 9404 11160 9456 11212
rect 13452 11160 13504 11212
rect 17684 11160 17736 11212
rect 6000 11024 6052 11076
rect 2044 10999 2096 11008
rect 2044 10965 2053 10999
rect 2053 10965 2087 10999
rect 2087 10965 2096 10999
rect 2044 10956 2096 10965
rect 2412 10999 2464 11008
rect 2412 10965 2421 10999
rect 2421 10965 2455 10999
rect 2455 10965 2464 10999
rect 2412 10956 2464 10965
rect 3056 10999 3108 11008
rect 3056 10965 3065 10999
rect 3065 10965 3099 10999
rect 3099 10965 3108 10999
rect 3056 10956 3108 10965
rect 7380 11024 7432 11076
rect 7932 11024 7984 11076
rect 9128 11092 9180 11144
rect 11888 11135 11940 11144
rect 8484 11067 8536 11076
rect 8484 11033 8493 11067
rect 8493 11033 8527 11067
rect 8527 11033 8536 11067
rect 11888 11101 11897 11135
rect 11897 11101 11931 11135
rect 11931 11101 11940 11135
rect 11888 11092 11940 11101
rect 13820 11092 13872 11144
rect 14464 11135 14516 11144
rect 14464 11101 14473 11135
rect 14473 11101 14507 11135
rect 14507 11101 14516 11135
rect 14464 11092 14516 11101
rect 16948 11092 17000 11144
rect 8484 11024 8536 11033
rect 9496 11024 9548 11076
rect 9588 11024 9640 11076
rect 14924 11024 14976 11076
rect 17500 11024 17552 11076
rect 11704 10956 11756 11008
rect 14832 10999 14884 11008
rect 14832 10965 14841 10999
rect 14841 10965 14875 10999
rect 14875 10965 14884 10999
rect 14832 10956 14884 10965
rect 17592 10999 17644 11008
rect 17592 10965 17601 10999
rect 17601 10965 17635 10999
rect 17635 10965 17644 10999
rect 17592 10956 17644 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 2044 10752 2096 10804
rect 2044 10659 2096 10668
rect 2044 10625 2053 10659
rect 2053 10625 2087 10659
rect 2087 10625 2096 10659
rect 2044 10616 2096 10625
rect 2964 10616 3016 10668
rect 2872 10548 2924 10600
rect 3240 10752 3292 10804
rect 4252 10752 4304 10804
rect 4528 10752 4580 10804
rect 5356 10795 5408 10804
rect 5356 10761 5365 10795
rect 5365 10761 5399 10795
rect 5399 10761 5408 10795
rect 5356 10752 5408 10761
rect 6000 10752 6052 10804
rect 8116 10752 8168 10804
rect 10416 10752 10468 10804
rect 12072 10752 12124 10804
rect 14832 10795 14884 10804
rect 3976 10684 4028 10736
rect 5724 10684 5776 10736
rect 7012 10684 7064 10736
rect 11244 10684 11296 10736
rect 12624 10727 12676 10736
rect 12624 10693 12633 10727
rect 12633 10693 12667 10727
rect 12667 10693 12676 10727
rect 12624 10684 12676 10693
rect 12808 10684 12860 10736
rect 14832 10761 14841 10795
rect 14841 10761 14875 10795
rect 14875 10761 14884 10795
rect 14832 10752 14884 10761
rect 14924 10795 14976 10804
rect 14924 10761 14933 10795
rect 14933 10761 14967 10795
rect 14967 10761 14976 10795
rect 14924 10752 14976 10761
rect 15568 10752 15620 10804
rect 17592 10752 17644 10804
rect 4068 10659 4120 10668
rect 4068 10625 4077 10659
rect 4077 10625 4111 10659
rect 4111 10625 4120 10659
rect 4068 10616 4120 10625
rect 4804 10616 4856 10668
rect 5448 10616 5500 10668
rect 5908 10616 5960 10668
rect 8392 10616 8444 10668
rect 5080 10548 5132 10600
rect 7380 10548 7432 10600
rect 11704 10591 11756 10600
rect 11704 10557 11713 10591
rect 11713 10557 11747 10591
rect 11747 10557 11756 10591
rect 11704 10548 11756 10557
rect 7840 10480 7892 10532
rect 14924 10548 14976 10600
rect 15936 10659 15988 10668
rect 15936 10625 15945 10659
rect 15945 10625 15979 10659
rect 15979 10625 15988 10659
rect 15936 10616 15988 10625
rect 16948 10684 17000 10736
rect 17316 10616 17368 10668
rect 17960 10616 18012 10668
rect 2688 10412 2740 10464
rect 6000 10412 6052 10464
rect 6920 10412 6972 10464
rect 9404 10412 9456 10464
rect 11796 10412 11848 10464
rect 11888 10412 11940 10464
rect 12256 10455 12308 10464
rect 12256 10421 12265 10455
rect 12265 10421 12299 10455
rect 12299 10421 12308 10455
rect 12256 10412 12308 10421
rect 14924 10412 14976 10464
rect 17776 10412 17828 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1860 10251 1912 10260
rect 1860 10217 1869 10251
rect 1869 10217 1903 10251
rect 1903 10217 1912 10251
rect 1860 10208 1912 10217
rect 3056 10208 3108 10260
rect 4160 10208 4212 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 7564 10208 7616 10260
rect 9128 10208 9180 10260
rect 11888 10208 11940 10260
rect 13084 10208 13136 10260
rect 15384 10251 15436 10260
rect 15384 10217 15393 10251
rect 15393 10217 15427 10251
rect 15427 10217 15436 10251
rect 15384 10208 15436 10217
rect 16948 10251 17000 10260
rect 16948 10217 16957 10251
rect 16957 10217 16991 10251
rect 16991 10217 17000 10251
rect 16948 10208 17000 10217
rect 17960 10208 18012 10260
rect 1952 10140 2004 10192
rect 3608 10140 3660 10192
rect 3976 10140 4028 10192
rect 3240 10115 3292 10124
rect 3240 10081 3249 10115
rect 3249 10081 3283 10115
rect 3283 10081 3292 10115
rect 3240 10072 3292 10081
rect 4068 10072 4120 10124
rect 6736 10140 6788 10192
rect 5080 10072 5132 10124
rect 12072 10140 12124 10192
rect 12256 10140 12308 10192
rect 9496 10115 9548 10124
rect 9496 10081 9505 10115
rect 9505 10081 9539 10115
rect 9539 10081 9548 10115
rect 9496 10072 9548 10081
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 1584 10047 1636 10056
rect 1584 10013 1593 10047
rect 1593 10013 1627 10047
rect 1627 10013 1636 10047
rect 1584 10004 1636 10013
rect 4988 10047 5040 10056
rect 4988 10013 4997 10047
rect 4997 10013 5031 10047
rect 5031 10013 5040 10047
rect 4988 10004 5040 10013
rect 7012 10047 7064 10056
rect 7012 10013 7021 10047
rect 7021 10013 7055 10047
rect 7055 10013 7064 10047
rect 7012 10004 7064 10013
rect 8024 10004 8076 10056
rect 8484 10004 8536 10056
rect 9312 10004 9364 10056
rect 11244 10004 11296 10056
rect 2872 9936 2924 9988
rect 13176 10004 13228 10056
rect 14740 10047 14792 10056
rect 14740 10013 14749 10047
rect 14749 10013 14783 10047
rect 14783 10013 14792 10047
rect 14740 10004 14792 10013
rect 17684 10047 17736 10056
rect 17684 10013 17693 10047
rect 17693 10013 17727 10047
rect 17727 10013 17736 10047
rect 17684 10004 17736 10013
rect 2596 9868 2648 9920
rect 3792 9868 3844 9920
rect 5264 9868 5316 9920
rect 5632 9868 5684 9920
rect 9312 9911 9364 9920
rect 9312 9877 9321 9911
rect 9321 9877 9355 9911
rect 9355 9877 9364 9911
rect 9312 9868 9364 9877
rect 9680 9868 9732 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 2964 9707 3016 9716
rect 2964 9673 2973 9707
rect 2973 9673 3007 9707
rect 3007 9673 3016 9707
rect 2964 9664 3016 9673
rect 4068 9596 4120 9648
rect 4252 9664 4304 9716
rect 4712 9664 4764 9716
rect 5724 9664 5776 9716
rect 1492 9571 1544 9580
rect 1492 9537 1501 9571
rect 1501 9537 1535 9571
rect 1535 9537 1544 9571
rect 1492 9528 1544 9537
rect 1860 9528 1912 9580
rect 3332 9537 3341 9564
rect 3341 9537 3375 9564
rect 3375 9537 3384 9564
rect 3332 9512 3384 9537
rect 3792 9528 3844 9580
rect 3608 9503 3660 9512
rect 1676 9435 1728 9444
rect 1676 9401 1685 9435
rect 1685 9401 1719 9435
rect 1719 9401 1728 9435
rect 1676 9392 1728 9401
rect 2872 9392 2924 9444
rect 3056 9392 3108 9444
rect 3608 9469 3617 9503
rect 3617 9469 3651 9503
rect 3651 9469 3660 9503
rect 3608 9460 3660 9469
rect 4160 9392 4212 9444
rect 2596 9367 2648 9376
rect 2596 9333 2605 9367
rect 2605 9333 2639 9367
rect 2639 9333 2648 9367
rect 2596 9324 2648 9333
rect 2780 9324 2832 9376
rect 5080 9528 5132 9580
rect 4620 9435 4672 9444
rect 4620 9401 4629 9435
rect 4629 9401 4663 9435
rect 4663 9401 4672 9435
rect 4620 9392 4672 9401
rect 5356 9571 5408 9580
rect 5356 9537 5365 9571
rect 5365 9537 5399 9571
rect 5399 9537 5408 9571
rect 5356 9528 5408 9537
rect 6828 9528 6880 9580
rect 8392 9664 8444 9716
rect 8668 9664 8720 9716
rect 12624 9664 12676 9716
rect 5448 9503 5500 9512
rect 5448 9469 5457 9503
rect 5457 9469 5491 9503
rect 5491 9469 5500 9503
rect 5448 9460 5500 9469
rect 8300 9596 8352 9648
rect 8668 9528 8720 9580
rect 9404 9596 9456 9648
rect 9588 9596 9640 9648
rect 11796 9639 11848 9648
rect 11796 9605 11830 9639
rect 11830 9605 11848 9639
rect 11796 9596 11848 9605
rect 9220 9571 9272 9580
rect 9220 9537 9254 9571
rect 9254 9537 9272 9571
rect 9220 9528 9272 9537
rect 15568 9664 15620 9716
rect 13820 9639 13872 9648
rect 13820 9605 13829 9639
rect 13829 9605 13863 9639
rect 13863 9605 13872 9639
rect 13820 9596 13872 9605
rect 14280 9639 14332 9648
rect 14280 9605 14289 9639
rect 14289 9605 14323 9639
rect 14323 9605 14332 9639
rect 14280 9596 14332 9605
rect 14924 9571 14976 9580
rect 14924 9537 14933 9571
rect 14933 9537 14967 9571
rect 14967 9537 14976 9571
rect 14924 9528 14976 9537
rect 8300 9460 8352 9512
rect 8484 9460 8536 9512
rect 4712 9324 4764 9376
rect 7748 9324 7800 9376
rect 8484 9367 8536 9376
rect 8484 9333 8493 9367
rect 8493 9333 8527 9367
rect 8527 9333 8536 9367
rect 8484 9324 8536 9333
rect 9588 9324 9640 9376
rect 10968 9367 11020 9376
rect 10968 9333 10977 9367
rect 10977 9333 11011 9367
rect 11011 9333 11020 9367
rect 10968 9324 11020 9333
rect 11060 9324 11112 9376
rect 15936 9392 15988 9444
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1308 9120 1360 9172
rect 1952 9120 2004 9172
rect 4988 9120 5040 9172
rect 5448 9120 5500 9172
rect 9312 9120 9364 9172
rect 9680 9163 9732 9172
rect 9680 9129 9689 9163
rect 9689 9129 9723 9163
rect 9723 9129 9732 9163
rect 9680 9120 9732 9129
rect 9772 9120 9824 9172
rect 4160 9052 4212 9104
rect 4620 9052 4672 9104
rect 5172 9052 5224 9104
rect 3516 8984 3568 9036
rect 5816 9052 5868 9104
rect 9496 9052 9548 9104
rect 6736 9027 6788 9036
rect 6736 8993 6745 9027
rect 6745 8993 6779 9027
rect 6779 8993 6788 9027
rect 6736 8984 6788 8993
rect 1860 8916 1912 8968
rect 3240 8916 3292 8968
rect 4528 8916 4580 8968
rect 5632 8959 5684 8968
rect 5632 8925 5641 8959
rect 5641 8925 5675 8959
rect 5675 8925 5684 8959
rect 5632 8916 5684 8925
rect 8024 8984 8076 9036
rect 9128 9027 9180 9036
rect 9128 8993 9137 9027
rect 9137 8993 9171 9027
rect 9171 8993 9180 9027
rect 9128 8984 9180 8993
rect 17224 9120 17276 9172
rect 8484 8916 8536 8968
rect 2596 8848 2648 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2044 8780 2096 8832
rect 2964 8780 3016 8832
rect 4252 8780 4304 8832
rect 4436 8780 4488 8832
rect 4988 8823 5040 8832
rect 4988 8789 4997 8823
rect 4997 8789 5031 8823
rect 5031 8789 5040 8823
rect 4988 8780 5040 8789
rect 5172 8780 5224 8832
rect 5724 8780 5776 8832
rect 10968 8848 11020 8900
rect 6552 8780 6604 8832
rect 7656 8823 7708 8832
rect 7656 8789 7665 8823
rect 7665 8789 7699 8823
rect 7699 8789 7708 8823
rect 7656 8780 7708 8789
rect 8760 8780 8812 8832
rect 9312 8823 9364 8832
rect 9312 8789 9321 8823
rect 9321 8789 9355 8823
rect 9355 8789 9364 8823
rect 9312 8780 9364 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 1768 8576 1820 8628
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 4896 8619 4948 8628
rect 4896 8585 4905 8619
rect 4905 8585 4939 8619
rect 4939 8585 4948 8619
rect 4896 8576 4948 8585
rect 1584 8483 1636 8492
rect 1584 8449 1593 8483
rect 1593 8449 1627 8483
rect 1627 8449 1636 8483
rect 1584 8440 1636 8449
rect 2688 8508 2740 8560
rect 4068 8508 4120 8560
rect 8668 8576 8720 8628
rect 8760 8508 8812 8560
rect 9496 8508 9548 8560
rect 2320 8483 2372 8492
rect 2320 8449 2329 8483
rect 2329 8449 2363 8483
rect 2363 8449 2372 8483
rect 2320 8440 2372 8449
rect 2780 8440 2832 8492
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 3240 8483 3292 8492
rect 2964 8440 3016 8449
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 3516 8483 3568 8492
rect 3516 8449 3550 8483
rect 3550 8449 3568 8483
rect 3516 8440 3568 8449
rect 4436 8440 4488 8492
rect 6460 8440 6512 8492
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 5908 8415 5960 8424
rect 5908 8381 5917 8415
rect 5917 8381 5951 8415
rect 5951 8381 5960 8415
rect 5908 8372 5960 8381
rect 6092 8372 6144 8424
rect 8392 8440 8444 8492
rect 10232 8440 10284 8492
rect 7748 8372 7800 8424
rect 9404 8415 9456 8424
rect 9404 8381 9413 8415
rect 9413 8381 9447 8415
rect 9447 8381 9456 8415
rect 9404 8372 9456 8381
rect 3148 8304 3200 8356
rect 2872 8236 2924 8288
rect 5540 8304 5592 8356
rect 8024 8347 8076 8356
rect 8024 8313 8033 8347
rect 8033 8313 8067 8347
rect 8067 8313 8076 8347
rect 8024 8304 8076 8313
rect 18880 8304 18932 8356
rect 20168 8304 20220 8356
rect 4804 8236 4856 8288
rect 7104 8236 7156 8288
rect 7656 8236 7708 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 1492 8075 1544 8084
rect 1492 8041 1501 8075
rect 1501 8041 1535 8075
rect 1535 8041 1544 8075
rect 1492 8032 1544 8041
rect 1584 8032 1636 8084
rect 1952 8007 2004 8016
rect 1952 7973 1961 8007
rect 1961 7973 1995 8007
rect 1995 7973 2004 8007
rect 1952 7964 2004 7973
rect 2136 7896 2188 7948
rect 2412 7871 2464 7880
rect 2412 7837 2421 7871
rect 2421 7837 2455 7871
rect 2455 7837 2464 7871
rect 2412 7828 2464 7837
rect 2136 7760 2188 7812
rect 5908 8032 5960 8084
rect 4160 7964 4212 8016
rect 10232 8032 10284 8084
rect 18880 8075 18932 8084
rect 18880 8041 18889 8075
rect 18889 8041 18923 8075
rect 18923 8041 18932 8075
rect 18880 8032 18932 8041
rect 3332 7939 3384 7948
rect 3332 7905 3341 7939
rect 3341 7905 3375 7939
rect 3375 7905 3384 7939
rect 3332 7896 3384 7905
rect 4252 7896 4304 7948
rect 4712 7939 4764 7948
rect 4712 7905 4721 7939
rect 4721 7905 4755 7939
rect 4755 7905 4764 7939
rect 4712 7896 4764 7905
rect 4804 7939 4856 7948
rect 4804 7905 4813 7939
rect 4813 7905 4847 7939
rect 4847 7905 4856 7939
rect 4804 7896 4856 7905
rect 9312 7896 9364 7948
rect 3976 7871 4028 7880
rect 3976 7837 3985 7871
rect 3985 7837 4019 7871
rect 4019 7837 4028 7871
rect 3976 7828 4028 7837
rect 4988 7828 5040 7880
rect 9404 7828 9456 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 6000 7760 6052 7812
rect 2320 7692 2372 7744
rect 4896 7692 4948 7744
rect 6644 7735 6696 7744
rect 6644 7701 6653 7735
rect 6653 7701 6687 7735
rect 6687 7701 6696 7735
rect 6644 7692 6696 7701
rect 7748 7760 7800 7812
rect 8668 7692 8720 7744
rect 10324 7692 10376 7744
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 1400 7488 1452 7540
rect 2228 7488 2280 7540
rect 3332 7488 3384 7540
rect 5540 7531 5592 7540
rect 5540 7497 5549 7531
rect 5549 7497 5583 7531
rect 5583 7497 5592 7531
rect 5540 7488 5592 7497
rect 6552 7488 6604 7540
rect 8392 7488 8444 7540
rect 9588 7531 9640 7540
rect 9588 7497 9597 7531
rect 9597 7497 9631 7531
rect 9631 7497 9640 7531
rect 9588 7488 9640 7497
rect 10324 7488 10376 7540
rect 19524 7488 19576 7540
rect 2964 7420 3016 7472
rect 3424 7463 3476 7472
rect 3424 7429 3433 7463
rect 3433 7429 3467 7463
rect 3467 7429 3476 7463
rect 3424 7420 3476 7429
rect 6644 7463 6696 7472
rect 2136 7352 2188 7404
rect 2688 7395 2740 7404
rect 940 7216 992 7268
rect 1400 7216 1452 7268
rect 1584 7259 1636 7268
rect 1584 7225 1593 7259
rect 1593 7225 1627 7259
rect 1627 7225 1636 7259
rect 1584 7216 1636 7225
rect 2688 7361 2697 7395
rect 2697 7361 2731 7395
rect 2731 7361 2740 7395
rect 2688 7352 2740 7361
rect 4160 7395 4212 7404
rect 4160 7361 4169 7395
rect 4169 7361 4203 7395
rect 4203 7361 4212 7395
rect 4160 7352 4212 7361
rect 4804 7352 4856 7404
rect 6644 7429 6678 7463
rect 6678 7429 6696 7463
rect 6644 7420 6696 7429
rect 8300 7352 8352 7404
rect 9312 7420 9364 7472
rect 8576 7327 8628 7336
rect 8576 7293 8585 7327
rect 8585 7293 8619 7327
rect 8619 7293 8628 7327
rect 8576 7284 8628 7293
rect 4160 7216 4212 7268
rect 7380 7216 7432 7268
rect 17960 7352 18012 7404
rect 5816 7148 5868 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 8116 7191 8168 7200
rect 8116 7157 8125 7191
rect 8125 7157 8159 7191
rect 8159 7157 8168 7191
rect 8116 7148 8168 7157
rect 204 7080 256 7132
rect 940 7080 992 7132
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 1584 6944 1636 6996
rect 4252 6944 4304 6996
rect 5908 6944 5960 6996
rect 6000 6944 6052 6996
rect 1216 6808 1268 6860
rect 4528 6876 4580 6928
rect 5356 6876 5408 6928
rect 3792 6851 3844 6860
rect 1400 6783 1452 6792
rect 1400 6749 1409 6783
rect 1409 6749 1443 6783
rect 1443 6749 1452 6783
rect 1400 6740 1452 6749
rect 1676 6740 1728 6792
rect 1768 6740 1820 6792
rect 2872 6740 2924 6792
rect 2044 6647 2096 6656
rect 2044 6613 2053 6647
rect 2053 6613 2087 6647
rect 2087 6613 2096 6647
rect 2044 6604 2096 6613
rect 2504 6647 2556 6656
rect 2504 6613 2513 6647
rect 2513 6613 2547 6647
rect 2547 6613 2556 6647
rect 2504 6604 2556 6613
rect 3148 6672 3200 6724
rect 3792 6817 3801 6851
rect 3801 6817 3835 6851
rect 3835 6817 3844 6851
rect 3792 6808 3844 6817
rect 4804 6851 4856 6860
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 9588 6876 9640 6928
rect 2688 6604 2740 6656
rect 3976 6740 4028 6792
rect 4160 6740 4212 6792
rect 4620 6740 4672 6792
rect 7748 6808 7800 6860
rect 5540 6783 5592 6792
rect 5540 6749 5549 6783
rect 5549 6749 5583 6783
rect 5583 6749 5592 6783
rect 5540 6740 5592 6749
rect 8116 6740 8168 6792
rect 19616 6783 19668 6792
rect 19616 6749 19625 6783
rect 19625 6749 19659 6783
rect 19659 6749 19668 6783
rect 19616 6740 19668 6749
rect 4252 6672 4304 6724
rect 4436 6672 4488 6724
rect 4528 6604 4580 6656
rect 5080 6604 5132 6656
rect 5724 6672 5776 6724
rect 7104 6647 7156 6656
rect 7104 6613 7113 6647
rect 7113 6613 7147 6647
rect 7147 6613 7156 6647
rect 7104 6604 7156 6613
rect 8668 6604 8720 6656
rect 19800 6647 19852 6656
rect 19800 6613 19809 6647
rect 19809 6613 19843 6647
rect 19843 6613 19852 6647
rect 19800 6604 19852 6613
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 1584 6443 1636 6452
rect 1584 6409 1593 6443
rect 1593 6409 1627 6443
rect 1627 6409 1636 6443
rect 1584 6400 1636 6409
rect 2596 6400 2648 6452
rect 2780 6400 2832 6452
rect 3792 6443 3844 6452
rect 3792 6409 3801 6443
rect 3801 6409 3835 6443
rect 3835 6409 3844 6443
rect 3792 6400 3844 6409
rect 3976 6400 4028 6452
rect 8300 6443 8352 6452
rect 8300 6409 8309 6443
rect 8309 6409 8343 6443
rect 8343 6409 8352 6443
rect 8300 6400 8352 6409
rect 21640 6400 21692 6452
rect 1676 6332 1728 6384
rect 2688 6332 2740 6384
rect 1400 6307 1452 6316
rect 1400 6273 1409 6307
rect 1409 6273 1443 6307
rect 1443 6273 1452 6307
rect 1400 6264 1452 6273
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 4068 6332 4120 6384
rect 5632 6332 5684 6384
rect 3240 6307 3292 6316
rect 3240 6273 3249 6307
rect 3249 6273 3283 6307
rect 3283 6273 3292 6307
rect 3240 6264 3292 6273
rect 20076 6307 20128 6316
rect 20076 6273 20085 6307
rect 20085 6273 20119 6307
rect 20119 6273 20128 6307
rect 20076 6264 20128 6273
rect 2412 6196 2464 6248
rect 480 6128 532 6180
rect 3424 6171 3476 6180
rect 3424 6137 3433 6171
rect 3433 6137 3467 6171
rect 3467 6137 3476 6171
rect 3424 6128 3476 6137
rect 1768 6060 1820 6112
rect 3976 6128 4028 6180
rect 4344 6128 4396 6180
rect 4436 6128 4488 6180
rect 5264 6128 5316 6180
rect 8576 6128 8628 6180
rect 4160 6103 4212 6112
rect 4160 6069 4169 6103
rect 4169 6069 4203 6103
rect 4203 6069 4212 6103
rect 4160 6060 4212 6069
rect 4620 6060 4672 6112
rect 4712 6103 4764 6112
rect 4712 6069 4721 6103
rect 4721 6069 4755 6103
rect 4755 6069 4764 6103
rect 4712 6060 4764 6069
rect 4988 6060 5040 6112
rect 5080 6103 5132 6112
rect 5080 6069 5089 6103
rect 5089 6069 5123 6103
rect 5123 6069 5132 6103
rect 5080 6060 5132 6069
rect 5356 6060 5408 6112
rect 7104 6060 7156 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 1308 5652 1360 5704
rect 2504 5831 2556 5840
rect 2504 5797 2513 5831
rect 2513 5797 2547 5831
rect 2547 5797 2556 5831
rect 2504 5788 2556 5797
rect 2872 5788 2924 5840
rect 3056 5788 3108 5840
rect 3332 5831 3384 5840
rect 3332 5797 3341 5831
rect 3341 5797 3375 5831
rect 3375 5797 3384 5831
rect 3332 5788 3384 5797
rect 3792 5788 3844 5840
rect 4436 5788 4488 5840
rect 4620 5899 4672 5908
rect 4620 5865 4629 5899
rect 4629 5865 4663 5899
rect 4663 5865 4672 5899
rect 4988 5899 5040 5908
rect 4620 5856 4672 5865
rect 4988 5865 4997 5899
rect 4997 5865 5031 5899
rect 5031 5865 5040 5899
rect 4988 5856 5040 5865
rect 5356 5899 5408 5908
rect 5356 5865 5365 5899
rect 5365 5865 5399 5899
rect 5399 5865 5408 5899
rect 5356 5856 5408 5865
rect 21548 5856 21600 5908
rect 21824 5788 21876 5840
rect 3240 5720 3292 5772
rect 2228 5652 2280 5704
rect 2044 5559 2096 5568
rect 2044 5525 2053 5559
rect 2053 5525 2087 5559
rect 2087 5525 2096 5559
rect 2044 5516 2096 5525
rect 2780 5695 2832 5704
rect 2780 5661 2789 5695
rect 2789 5661 2823 5695
rect 2823 5661 2832 5695
rect 2780 5652 2832 5661
rect 5356 5584 5408 5636
rect 3240 5516 3292 5568
rect 3792 5559 3844 5568
rect 3792 5525 3801 5559
rect 3801 5525 3835 5559
rect 3835 5525 3844 5559
rect 3792 5516 3844 5525
rect 4344 5516 4396 5568
rect 5264 5516 5316 5568
rect 8300 5516 8352 5568
rect 20812 5652 20864 5704
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 2044 5355 2096 5364
rect 2044 5321 2053 5355
rect 2053 5321 2087 5355
rect 2087 5321 2096 5355
rect 2044 5312 2096 5321
rect 2504 5355 2556 5364
rect 2504 5321 2513 5355
rect 2513 5321 2547 5355
rect 2547 5321 2556 5355
rect 2504 5312 2556 5321
rect 3056 5312 3108 5364
rect 3976 5312 4028 5364
rect 4620 5355 4672 5364
rect 4620 5321 4629 5355
rect 4629 5321 4663 5355
rect 4663 5321 4672 5355
rect 4620 5312 4672 5321
rect 5356 5355 5408 5364
rect 5356 5321 5365 5355
rect 5365 5321 5399 5355
rect 5399 5321 5408 5355
rect 5356 5312 5408 5321
rect 5908 5312 5960 5364
rect 940 5244 992 5296
rect 1308 5176 1360 5228
rect 1860 5219 1912 5228
rect 1860 5185 1869 5219
rect 1869 5185 1903 5219
rect 1903 5185 1912 5219
rect 1860 5176 1912 5185
rect 2780 5176 2832 5228
rect 3976 5176 4028 5228
rect 7472 5176 7524 5228
rect 3056 5108 3108 5160
rect 20812 5151 20864 5160
rect 20812 5117 20821 5151
rect 20821 5117 20855 5151
rect 20855 5117 20864 5151
rect 20812 5108 20864 5117
rect 1584 5015 1636 5024
rect 1584 4981 1593 5015
rect 1593 4981 1627 5015
rect 1627 4981 1636 5015
rect 1584 4972 1636 4981
rect 2596 4972 2648 5024
rect 5080 5040 5132 5092
rect 4252 4972 4304 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 664 4768 716 4820
rect 3884 4811 3936 4820
rect 3884 4777 3893 4811
rect 3893 4777 3927 4811
rect 3927 4777 3936 4811
rect 3884 4768 3936 4777
rect 4068 4768 4120 4820
rect 756 4700 808 4752
rect 2780 4700 2832 4752
rect 1124 4632 1176 4684
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 3700 4496 3752 4548
rect 1584 4471 1636 4480
rect 1584 4437 1593 4471
rect 1593 4437 1627 4471
rect 1627 4437 1636 4471
rect 1584 4428 1636 4437
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 4160 4428 4212 4480
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 2136 4224 2188 4276
rect 3976 4267 4028 4276
rect 3976 4233 3985 4267
rect 3985 4233 4019 4267
rect 4019 4233 4028 4267
rect 3976 4224 4028 4233
rect 7380 4156 7432 4208
rect 3700 4088 3752 4140
rect 2228 4063 2280 4072
rect 2228 4029 2237 4063
rect 2237 4029 2271 4063
rect 2271 4029 2280 4063
rect 2228 4020 2280 4029
rect 3056 4020 3108 4072
rect 1952 3952 2004 4004
rect 3240 3995 3292 4004
rect 3240 3961 3249 3995
rect 3249 3961 3283 3995
rect 3283 3961 3292 3995
rect 3240 3952 3292 3961
rect 572 3884 624 3936
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2228 3680 2280 3732
rect 2872 3612 2924 3664
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 4344 3544 4396 3596
rect 2228 3519 2280 3528
rect 2228 3485 2237 3519
rect 2237 3485 2271 3519
rect 2271 3485 2280 3519
rect 2228 3476 2280 3485
rect 2872 3408 2924 3460
rect 1308 3340 1360 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 2780 3136 2832 3188
rect 4712 3068 4764 3120
rect 2780 3000 2832 3052
rect 2872 2932 2924 2984
rect 2964 2864 3016 2916
rect 3056 2839 3108 2848
rect 3056 2805 3065 2839
rect 3065 2805 3099 2839
rect 3099 2805 3108 2839
rect 3056 2796 3108 2805
rect 3240 2796 3292 2848
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 2596 2592 2648 2644
rect 3332 2592 3384 2644
rect 4252 2592 4304 2644
rect 4896 2524 4948 2576
rect 3424 2456 3476 2508
rect 2780 2388 2832 2440
rect 2964 2320 3016 2372
rect 3240 2363 3292 2372
rect 3240 2329 3249 2363
rect 3249 2329 3283 2363
rect 3283 2329 3292 2363
rect 3240 2320 3292 2329
rect 3976 2320 4028 2372
rect 2780 2252 2832 2304
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
<< metal2 >>
rect 202 22200 258 23000
rect 662 22200 718 23000
rect 1122 22200 1178 23000
rect 1582 22200 1638 23000
rect 2042 22200 2098 23000
rect 2502 22200 2558 23000
rect 2594 22672 2650 22681
rect 2650 22630 2820 22658
rect 2594 22607 2650 22616
rect 216 16182 244 22200
rect 676 20097 704 22200
rect 848 20460 900 20466
rect 848 20402 900 20408
rect 662 20088 718 20097
rect 662 20023 718 20032
rect 572 19236 624 19242
rect 572 19178 624 19184
rect 204 16176 256 16182
rect 204 16118 256 16124
rect 216 7138 244 16118
rect 478 11656 534 11665
rect 478 11591 534 11600
rect 204 7132 256 7138
rect 204 7074 256 7080
rect 492 6186 520 11591
rect 480 6180 532 6186
rect 480 6122 532 6128
rect 584 3942 612 19178
rect 756 17672 808 17678
rect 756 17614 808 17620
rect 662 13560 718 13569
rect 662 13495 718 13504
rect 676 4826 704 13495
rect 664 4820 716 4826
rect 664 4762 716 4768
rect 768 4758 796 17614
rect 756 4752 808 4758
rect 756 4694 808 4700
rect 860 4026 888 20402
rect 1136 19310 1164 22200
rect 1596 19854 1624 22200
rect 1674 21312 1730 21321
rect 1674 21247 1730 21256
rect 1216 19848 1268 19854
rect 1216 19790 1268 19796
rect 1584 19848 1636 19854
rect 1584 19790 1636 19796
rect 940 19304 992 19310
rect 940 19246 992 19252
rect 1124 19304 1176 19310
rect 1124 19246 1176 19252
rect 952 16574 980 19246
rect 1228 16574 1256 19790
rect 1398 18864 1454 18873
rect 1398 18799 1454 18808
rect 952 16546 1072 16574
rect 940 16448 992 16454
rect 940 16390 992 16396
rect 952 12073 980 16390
rect 938 12064 994 12073
rect 938 11999 994 12008
rect 938 11928 994 11937
rect 938 11863 994 11872
rect 952 7274 980 11863
rect 940 7268 992 7274
rect 940 7210 992 7216
rect 940 7132 992 7138
rect 940 7074 992 7080
rect 952 5302 980 7074
rect 1044 5545 1072 16546
rect 1136 16546 1256 16574
rect 1030 5536 1086 5545
rect 1030 5471 1086 5480
rect 940 5296 992 5302
rect 940 5238 992 5244
rect 1136 4690 1164 16546
rect 1412 15586 1440 18799
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1504 17678 1532 17711
rect 1492 17672 1544 17678
rect 1492 17614 1544 17620
rect 1688 17338 1716 21247
rect 2056 20534 2084 22200
rect 2044 20528 2096 20534
rect 2044 20470 2096 20476
rect 2516 19854 2544 22200
rect 2792 21350 2820 22630
rect 2962 22200 3018 23000
rect 3422 22200 3478 23000
rect 3528 22222 3832 22250
rect 2780 21344 2832 21350
rect 2780 21286 2832 21292
rect 2976 20466 3004 22200
rect 3054 21720 3110 21729
rect 3054 21655 3110 21664
rect 2964 20460 3016 20466
rect 2964 20402 3016 20408
rect 2504 19848 2556 19854
rect 2134 19816 2190 19825
rect 2504 19790 2556 19796
rect 2134 19751 2190 19760
rect 2044 19372 2096 19378
rect 2044 19314 2096 19320
rect 2056 18426 2084 19314
rect 2044 18420 2096 18426
rect 2044 18362 2096 18368
rect 1676 17332 1728 17338
rect 1676 17274 1728 17280
rect 1490 17096 1546 17105
rect 1490 17031 1546 17040
rect 1504 15706 1532 17031
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1584 16448 1636 16454
rect 1584 16390 1636 16396
rect 1596 16153 1624 16390
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1676 16108 1728 16114
rect 1676 16050 1728 16056
rect 1768 16108 1820 16114
rect 1768 16050 1820 16056
rect 1584 15904 1636 15910
rect 1584 15846 1636 15852
rect 1492 15700 1544 15706
rect 1492 15642 1544 15648
rect 1596 15609 1624 15846
rect 1582 15600 1638 15609
rect 1412 15558 1532 15586
rect 1400 15496 1452 15502
rect 1400 15438 1452 15444
rect 1216 15020 1268 15026
rect 1216 14962 1268 14968
rect 1228 6866 1256 14962
rect 1306 13288 1362 13297
rect 1306 13223 1362 13232
rect 1320 9178 1348 13223
rect 1412 12442 1440 15438
rect 1504 15162 1532 15558
rect 1582 15535 1638 15544
rect 1584 15360 1636 15366
rect 1584 15302 1636 15308
rect 1596 15201 1624 15302
rect 1582 15192 1638 15201
rect 1492 15156 1544 15162
rect 1582 15127 1638 15136
rect 1492 15098 1544 15104
rect 1492 14816 1544 14822
rect 1492 14758 1544 14764
rect 1504 14657 1532 14758
rect 1490 14648 1546 14657
rect 1490 14583 1546 14592
rect 1492 14272 1544 14278
rect 1490 14240 1492 14249
rect 1544 14240 1546 14249
rect 1490 14175 1546 14184
rect 1582 13832 1638 13841
rect 1582 13767 1584 13776
rect 1636 13767 1638 13776
rect 1584 13738 1636 13744
rect 1584 13320 1636 13326
rect 1584 13262 1636 13268
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1400 12436 1452 12442
rect 1400 12378 1452 12384
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1308 9172 1360 9178
rect 1308 9114 1360 9120
rect 1306 9072 1362 9081
rect 1306 9007 1362 9016
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1320 5710 1348 9007
rect 1412 7546 1440 12174
rect 1504 9586 1532 13126
rect 1596 12986 1624 13262
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1584 12096 1636 12102
rect 1584 12038 1636 12044
rect 1596 10062 1624 12038
rect 1688 11898 1716 16050
rect 1780 15337 1808 16050
rect 1766 15328 1822 15337
rect 1766 15263 1822 15272
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1584 10056 1636 10062
rect 1584 9998 1636 10004
rect 1492 9580 1544 9586
rect 1492 9522 1544 9528
rect 1674 9480 1730 9489
rect 1674 9415 1676 9424
rect 1728 9415 1730 9424
rect 1676 9386 1728 9392
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1596 8838 1624 8871
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 1780 8634 1808 13874
rect 1872 13326 1900 16934
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 2042 16552 2098 16561
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 1860 11212 1912 11218
rect 1860 11154 1912 11160
rect 1872 10266 1900 11154
rect 1860 10260 1912 10266
rect 1860 10202 1912 10208
rect 1872 9586 1900 10202
rect 1964 10198 1992 16526
rect 2042 16487 2098 16496
rect 2056 16454 2084 16487
rect 2044 16448 2096 16454
rect 2044 16390 2096 16396
rect 2148 16250 2176 19751
rect 2516 19242 2544 19790
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2594 19408 2650 19417
rect 2594 19343 2650 19352
rect 2504 19236 2556 19242
rect 2504 19178 2556 19184
rect 2318 18456 2374 18465
rect 2318 18391 2374 18400
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2136 16244 2188 16250
rect 2136 16186 2188 16192
rect 2136 15428 2188 15434
rect 2136 15370 2188 15376
rect 2148 15337 2176 15370
rect 2134 15328 2190 15337
rect 2134 15263 2190 15272
rect 2240 12918 2268 17138
rect 2332 14618 2360 18391
rect 2504 18148 2556 18154
rect 2504 18090 2556 18096
rect 2412 16992 2464 16998
rect 2412 16934 2464 16940
rect 2320 14612 2372 14618
rect 2320 14554 2372 14560
rect 2424 14414 2452 16934
rect 2412 14408 2464 14414
rect 2412 14350 2464 14356
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 2136 12640 2188 12646
rect 2136 12582 2188 12588
rect 2148 11150 2176 12582
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2044 11008 2096 11014
rect 2044 10950 2096 10956
rect 2056 10810 2084 10950
rect 2044 10804 2096 10810
rect 2044 10746 2096 10752
rect 2044 10668 2096 10674
rect 2044 10610 2096 10616
rect 1952 10192 2004 10198
rect 1952 10134 2004 10140
rect 1860 9580 1912 9586
rect 1860 9522 1912 9528
rect 1952 9172 2004 9178
rect 1952 9114 2004 9120
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1504 8090 1532 8191
rect 1596 8090 1624 8434
rect 1492 8084 1544 8090
rect 1492 8026 1544 8032
rect 1584 8084 1636 8090
rect 1584 8026 1636 8032
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1582 7304 1638 7313
rect 1400 7268 1452 7274
rect 1582 7239 1584 7248
rect 1400 7210 1452 7216
rect 1636 7239 1638 7248
rect 1584 7210 1636 7216
rect 1412 6798 1440 7210
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1400 6792 1452 6798
rect 1400 6734 1452 6740
rect 1596 6644 1624 6938
rect 1872 6914 1900 8910
rect 1964 8022 1992 9114
rect 2056 8838 2084 10610
rect 2134 9616 2190 9625
rect 2134 9551 2190 9560
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 2042 8664 2098 8673
rect 2042 8599 2044 8608
rect 2096 8599 2098 8608
rect 2044 8570 2096 8576
rect 1952 8016 2004 8022
rect 1952 7958 2004 7964
rect 2148 7954 2176 9551
rect 2136 7948 2188 7954
rect 2136 7890 2188 7896
rect 2134 7848 2190 7857
rect 2134 7783 2136 7792
rect 2188 7783 2190 7792
rect 2136 7754 2188 7760
rect 2240 7546 2268 11698
rect 2332 8498 2360 14214
rect 2412 13184 2464 13190
rect 2412 13126 2464 13132
rect 2424 12238 2452 13126
rect 2516 12458 2544 18090
rect 2608 15706 2636 19343
rect 2884 18834 2912 19450
rect 2872 18828 2924 18834
rect 2872 18770 2924 18776
rect 2688 18692 2740 18698
rect 2688 18634 2740 18640
rect 2700 18426 2728 18634
rect 2688 18420 2740 18426
rect 2688 18362 2740 18368
rect 2884 18306 2912 18770
rect 2964 18624 3016 18630
rect 2964 18566 3016 18572
rect 2976 18426 3004 18566
rect 2964 18420 3016 18426
rect 2964 18362 3016 18368
rect 2884 18278 3004 18306
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2884 17814 2912 18022
rect 2872 17808 2924 17814
rect 2872 17750 2924 17756
rect 2688 17672 2740 17678
rect 2688 17614 2740 17620
rect 2700 17134 2728 17614
rect 2872 17604 2924 17610
rect 2872 17546 2924 17552
rect 2780 17536 2832 17542
rect 2780 17478 2832 17484
rect 2792 17270 2820 17478
rect 2780 17264 2832 17270
rect 2780 17206 2832 17212
rect 2688 17128 2740 17134
rect 2688 17070 2740 17076
rect 2780 16720 2832 16726
rect 2780 16662 2832 16668
rect 2596 15700 2648 15706
rect 2596 15642 2648 15648
rect 2792 13938 2820 16662
rect 2884 15026 2912 17546
rect 2976 16590 3004 18278
rect 3068 17134 3096 21655
rect 3436 20602 3464 22200
rect 3424 20596 3476 20602
rect 3424 20538 3476 20544
rect 3332 20392 3384 20398
rect 3528 20346 3556 22222
rect 3804 22114 3832 22222
rect 3882 22200 3938 23000
rect 4342 22200 4398 23000
rect 4802 22200 4858 23000
rect 5262 22200 5318 23000
rect 5722 22200 5778 23000
rect 6182 22200 6238 23000
rect 6642 22200 6698 23000
rect 7010 22264 7066 22273
rect 3896 22114 3924 22200
rect 3804 22086 3924 22114
rect 3976 20868 4028 20874
rect 3976 20810 4028 20816
rect 3988 20777 4016 20810
rect 3974 20768 4030 20777
rect 3974 20703 4030 20712
rect 3976 20596 4028 20602
rect 3976 20538 4028 20544
rect 3988 20398 4016 20538
rect 3976 20392 4028 20398
rect 3332 20334 3384 20340
rect 3240 18624 3292 18630
rect 3240 18566 3292 18572
rect 3252 18465 3280 18566
rect 3238 18456 3294 18465
rect 3238 18391 3294 18400
rect 3238 18048 3294 18057
rect 3238 17983 3294 17992
rect 3146 17504 3202 17513
rect 3146 17439 3202 17448
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 2964 16584 3016 16590
rect 2964 16526 3016 16532
rect 3160 16250 3188 17439
rect 3148 16244 3200 16250
rect 3148 16186 3200 16192
rect 3252 15706 3280 17983
rect 3240 15700 3292 15706
rect 3240 15642 3292 15648
rect 3240 15564 3292 15570
rect 3240 15506 3292 15512
rect 2964 15496 3016 15502
rect 2964 15438 3016 15444
rect 2872 15020 2924 15026
rect 2872 14962 2924 14968
rect 2872 14544 2924 14550
rect 2872 14486 2924 14492
rect 2780 13932 2832 13938
rect 2780 13874 2832 13880
rect 2792 13705 2820 13874
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2686 13424 2742 13433
rect 2686 13359 2742 13368
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2608 12594 2636 13262
rect 2700 12850 2728 13359
rect 2884 13138 2912 14486
rect 2976 13530 3004 15438
rect 3056 14272 3108 14278
rect 3056 14214 3108 14220
rect 3148 14272 3200 14278
rect 3148 14214 3200 14220
rect 3068 14074 3096 14214
rect 3056 14068 3108 14074
rect 3056 14010 3108 14016
rect 3056 13932 3108 13938
rect 3056 13874 3108 13880
rect 2964 13524 3016 13530
rect 2964 13466 3016 13472
rect 2884 13110 3004 13138
rect 2870 12880 2926 12889
rect 2688 12844 2740 12850
rect 2870 12815 2926 12824
rect 2688 12786 2740 12792
rect 2608 12566 2728 12594
rect 2516 12430 2636 12458
rect 2504 12368 2556 12374
rect 2502 12336 2504 12345
rect 2556 12336 2558 12345
rect 2502 12271 2558 12280
rect 2412 12232 2464 12238
rect 2412 12174 2464 12180
rect 2608 11626 2636 12430
rect 2700 11665 2728 12566
rect 2884 12170 2912 12815
rect 2976 12306 3004 13110
rect 3068 12345 3096 13874
rect 3160 13870 3188 14214
rect 3148 13864 3200 13870
rect 3148 13806 3200 13812
rect 3054 12336 3110 12345
rect 2964 12300 3016 12306
rect 3054 12271 3110 12280
rect 2964 12242 3016 12248
rect 2872 12164 2924 12170
rect 2872 12106 2924 12112
rect 3056 12164 3108 12170
rect 3056 12106 3108 12112
rect 2870 12064 2926 12073
rect 2870 11999 2926 12008
rect 2686 11656 2742 11665
rect 2596 11620 2648 11626
rect 2686 11591 2742 11600
rect 2596 11562 2648 11568
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2594 11384 2650 11393
rect 2594 11319 2650 11328
rect 2412 11008 2464 11014
rect 2412 10950 2464 10956
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 2424 7886 2452 10950
rect 2502 10024 2558 10033
rect 2502 9959 2558 9968
rect 2412 7880 2464 7886
rect 2412 7822 2464 7828
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1872 6886 1992 6914
rect 1676 6792 1728 6798
rect 1676 6734 1728 6740
rect 1768 6792 1820 6798
rect 1768 6734 1820 6740
rect 1412 6616 1624 6644
rect 1412 6322 1440 6616
rect 1584 6452 1636 6458
rect 1584 6394 1636 6400
rect 1596 6361 1624 6394
rect 1688 6390 1716 6734
rect 1676 6384 1728 6390
rect 1582 6352 1638 6361
rect 1400 6316 1452 6322
rect 1676 6326 1728 6332
rect 1582 6287 1638 6296
rect 1400 6258 1452 6264
rect 1780 6118 1808 6734
rect 1858 6624 1914 6633
rect 1858 6559 1914 6568
rect 1768 6112 1820 6118
rect 1768 6054 1820 6060
rect 1582 5944 1638 5953
rect 1582 5879 1584 5888
rect 1636 5879 1638 5888
rect 1584 5850 1636 5856
rect 1308 5704 1360 5710
rect 1308 5646 1360 5652
rect 1306 5400 1362 5409
rect 1306 5335 1362 5344
rect 1320 5234 1348 5335
rect 1398 5264 1454 5273
rect 1308 5228 1360 5234
rect 1872 5234 1900 6559
rect 1398 5199 1454 5208
rect 1860 5228 1912 5234
rect 1308 5170 1360 5176
rect 1124 4684 1176 4690
rect 1124 4626 1176 4632
rect 938 4040 994 4049
rect 860 3998 938 4026
rect 938 3975 994 3984
rect 572 3936 624 3942
rect 572 3878 624 3884
rect 1320 3398 1348 5170
rect 1412 4622 1440 5199
rect 1860 5170 1912 5176
rect 1584 5024 1636 5030
rect 1584 4966 1636 4972
rect 1596 4729 1624 4966
rect 1582 4720 1638 4729
rect 1582 4655 1638 4664
rect 1400 4616 1452 4622
rect 1860 4616 1912 4622
rect 1400 4558 1452 4564
rect 1582 4584 1638 4593
rect 1860 4558 1912 4564
rect 1582 4519 1638 4528
rect 1596 4486 1624 4519
rect 1584 4480 1636 4486
rect 1872 4457 1900 4558
rect 1584 4422 1636 4428
rect 1858 4448 1914 4457
rect 1858 4383 1914 4392
rect 1964 4010 1992 6886
rect 2044 6656 2096 6662
rect 2042 6624 2044 6633
rect 2096 6624 2098 6633
rect 2042 6559 2098 6568
rect 2042 5672 2098 5681
rect 2042 5607 2098 5616
rect 2056 5574 2084 5607
rect 2044 5568 2096 5574
rect 2044 5510 2096 5516
rect 2042 5400 2098 5409
rect 2042 5335 2044 5344
rect 2096 5335 2098 5344
rect 2044 5306 2096 5312
rect 2148 4282 2176 7346
rect 2226 7168 2282 7177
rect 2226 7103 2282 7112
rect 2240 5710 2268 7103
rect 2332 6322 2360 7686
rect 2516 6914 2544 9959
rect 2608 9926 2636 11319
rect 2688 10464 2740 10470
rect 2686 10432 2688 10441
rect 2740 10432 2742 10441
rect 2686 10367 2742 10376
rect 2596 9920 2648 9926
rect 2596 9862 2648 9868
rect 2792 9738 2820 11494
rect 2884 10713 2912 11999
rect 2964 11756 3016 11762
rect 2964 11698 3016 11704
rect 2976 11354 3004 11698
rect 3068 11558 3096 12106
rect 3148 11688 3200 11694
rect 3148 11630 3200 11636
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 2964 11348 3016 11354
rect 2964 11290 3016 11296
rect 3056 11008 3108 11014
rect 3056 10950 3108 10956
rect 2870 10704 2926 10713
rect 2870 10639 2926 10648
rect 2964 10668 3016 10674
rect 2964 10610 3016 10616
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2884 9994 2912 10542
rect 2872 9988 2924 9994
rect 2872 9930 2924 9936
rect 2700 9710 2820 9738
rect 2976 9722 3004 10610
rect 3068 10266 3096 10950
rect 3056 10260 3108 10266
rect 3056 10202 3108 10208
rect 3054 10160 3110 10169
rect 3054 10095 3110 10104
rect 2964 9716 3016 9722
rect 2596 9376 2648 9382
rect 2596 9318 2648 9324
rect 2608 8906 2636 9318
rect 2596 8900 2648 8906
rect 2596 8842 2648 8848
rect 2700 8566 2728 9710
rect 2964 9658 3016 9664
rect 3068 9450 3096 10095
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2688 8560 2740 8566
rect 2688 8502 2740 8508
rect 2792 8498 2820 9318
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2686 8392 2742 8401
rect 2884 8378 2912 9386
rect 3054 9344 3110 9353
rect 3054 9279 3110 9288
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8498 3004 8774
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 2884 8350 3004 8378
rect 2686 8327 2742 8336
rect 2594 7984 2650 7993
rect 2594 7919 2650 7928
rect 2424 6886 2544 6914
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2424 6254 2452 6886
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 2516 6662 2544 6695
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2608 6458 2636 7919
rect 2700 7410 2728 8327
rect 2872 8288 2924 8294
rect 2872 8230 2924 8236
rect 2778 8120 2834 8129
rect 2778 8055 2834 8064
rect 2688 7404 2740 7410
rect 2688 7346 2740 7352
rect 2686 6760 2742 6769
rect 2686 6695 2742 6704
rect 2700 6662 2728 6695
rect 2688 6656 2740 6662
rect 2792 6644 2820 8055
rect 2884 6798 2912 8230
rect 2976 7478 3004 8350
rect 3068 8242 3096 9279
rect 3160 8362 3188 11630
rect 3252 11370 3280 15506
rect 3344 13433 3372 20334
rect 3436 20318 3556 20346
rect 3882 20360 3938 20369
rect 3436 18714 3464 20318
rect 3976 20334 4028 20340
rect 3882 20295 3938 20304
rect 3549 20156 3857 20176
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20080 3857 20100
rect 3549 19068 3857 19088
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 18992 3857 19012
rect 3896 18902 3924 20295
rect 3988 20233 4016 20334
rect 3974 20224 4030 20233
rect 3974 20159 4030 20168
rect 4160 19780 4212 19786
rect 4160 19722 4212 19728
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3700 18896 3752 18902
rect 3700 18838 3752 18844
rect 3884 18896 3936 18902
rect 3884 18838 3936 18844
rect 3436 18686 3556 18714
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3436 18086 3464 18566
rect 3528 18290 3556 18686
rect 3712 18630 3740 18838
rect 3792 18760 3844 18766
rect 3792 18702 3844 18708
rect 3700 18624 3752 18630
rect 3700 18566 3752 18572
rect 3516 18284 3568 18290
rect 3516 18226 3568 18232
rect 3804 18154 3832 18702
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 3792 18148 3844 18154
rect 3792 18090 3844 18096
rect 3424 18080 3476 18086
rect 3424 18022 3476 18028
rect 3549 17980 3857 18000
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17904 3857 17924
rect 3896 17762 3924 18226
rect 3988 18154 4016 19654
rect 4068 19508 4120 19514
rect 4068 19450 4120 19456
rect 3976 18148 4028 18154
rect 3976 18090 4028 18096
rect 3896 17734 4016 17762
rect 3884 17604 3936 17610
rect 3884 17546 3936 17552
rect 3424 17196 3476 17202
rect 3424 17138 3476 17144
rect 3436 16794 3464 17138
rect 3549 16892 3857 16912
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3549 16816 3857 16836
rect 3424 16788 3476 16794
rect 3424 16730 3476 16736
rect 3896 16590 3924 17546
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3424 16448 3476 16454
rect 3988 16402 4016 17734
rect 4080 16454 4108 19450
rect 4172 18970 4200 19722
rect 4160 18964 4212 18970
rect 4160 18906 4212 18912
rect 4160 18420 4212 18426
rect 4160 18362 4212 18368
rect 4172 18193 4200 18362
rect 4158 18184 4214 18193
rect 4158 18119 4214 18128
rect 4160 17808 4212 17814
rect 4160 17750 4212 17756
rect 4172 16590 4200 17750
rect 4356 17626 4384 22200
rect 4434 19952 4490 19961
rect 4434 19887 4490 19896
rect 4448 19417 4476 19887
rect 4434 19408 4490 19417
rect 4434 19343 4436 19352
rect 4488 19343 4490 19352
rect 4436 19314 4488 19320
rect 4528 19236 4580 19242
rect 4528 19178 4580 19184
rect 4540 18737 4568 19178
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4526 18728 4582 18737
rect 4526 18663 4582 18672
rect 4436 18624 4488 18630
rect 4436 18566 4488 18572
rect 4264 17598 4384 17626
rect 4448 17626 4476 18566
rect 4632 18426 4660 19110
rect 4816 18986 4844 22200
rect 5276 20346 5304 22200
rect 5632 20936 5684 20942
rect 5632 20878 5684 20884
rect 5540 20392 5592 20398
rect 5276 20318 5396 20346
rect 5540 20334 5592 20340
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 4986 19952 5042 19961
rect 4986 19887 5042 19896
rect 5000 19446 5028 19887
rect 5172 19848 5224 19854
rect 5172 19790 5224 19796
rect 4988 19440 5040 19446
rect 4988 19382 5040 19388
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4816 18958 4936 18986
rect 4804 18896 4856 18902
rect 4804 18838 4856 18844
rect 4712 18624 4764 18630
rect 4712 18566 4764 18572
rect 4620 18420 4672 18426
rect 4620 18362 4672 18368
rect 4724 18057 4752 18566
rect 4816 18290 4844 18838
rect 4908 18329 4936 18958
rect 4894 18320 4950 18329
rect 4804 18284 4856 18290
rect 4894 18255 4950 18264
rect 4804 18226 4856 18232
rect 4710 18048 4766 18057
rect 4710 17983 4766 17992
rect 4448 17598 4660 17626
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 3424 16390 3476 16396
rect 3330 13424 3386 13433
rect 3330 13359 3386 13368
rect 3332 12640 3384 12646
rect 3332 12582 3384 12588
rect 3344 12170 3372 12582
rect 3436 12238 3464 16390
rect 3896 16374 4016 16402
rect 4068 16448 4120 16454
rect 4068 16390 4120 16396
rect 3549 15804 3857 15824
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15728 3857 15748
rect 3896 15502 3924 16374
rect 3976 16108 4028 16114
rect 3976 16050 4028 16056
rect 4068 16108 4120 16114
rect 4068 16050 4120 16056
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3549 14716 3857 14736
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14640 3857 14660
rect 3792 14476 3844 14482
rect 3792 14418 3844 14424
rect 3804 14278 3832 14418
rect 3792 14272 3844 14278
rect 3790 14240 3792 14249
rect 3844 14240 3846 14249
rect 3790 14175 3846 14184
rect 3896 13734 3924 15438
rect 3988 15162 4016 16050
rect 3976 15156 4028 15162
rect 3976 15098 4028 15104
rect 3988 13870 4016 15098
rect 3976 13864 4028 13870
rect 3976 13806 4028 13812
rect 3884 13728 3936 13734
rect 3884 13670 3936 13676
rect 3549 13628 3857 13648
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13552 3857 13572
rect 3974 13560 4030 13569
rect 3974 13495 4030 13504
rect 3516 13388 3568 13394
rect 3516 13330 3568 13336
rect 3528 12850 3556 13330
rect 3988 13326 4016 13495
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 4080 12918 4108 16050
rect 4172 15434 4200 16526
rect 4160 15428 4212 15434
rect 4160 15370 4212 15376
rect 4160 14816 4212 14822
rect 4160 14758 4212 14764
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 3549 12540 3857 12560
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12464 3857 12484
rect 3896 12434 3924 12786
rect 4068 12436 4120 12442
rect 3896 12406 4016 12434
rect 3516 12368 3568 12374
rect 3516 12310 3568 12316
rect 3424 12232 3476 12238
rect 3424 12174 3476 12180
rect 3332 12164 3384 12170
rect 3332 12106 3384 12112
rect 3528 12102 3556 12310
rect 3516 12096 3568 12102
rect 3516 12038 3568 12044
rect 3792 12096 3844 12102
rect 3792 12038 3844 12044
rect 3804 11762 3832 12038
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3884 11620 3936 11626
rect 3884 11562 3936 11568
rect 3424 11552 3476 11558
rect 3424 11494 3476 11500
rect 3252 11342 3372 11370
rect 3344 11286 3372 11342
rect 3332 11280 3384 11286
rect 3332 11222 3384 11228
rect 3240 11212 3292 11218
rect 3240 11154 3292 11160
rect 3252 10810 3280 11154
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3240 10124 3292 10130
rect 3240 10066 3292 10072
rect 3252 8974 3280 10066
rect 3332 9564 3384 9570
rect 3332 9506 3384 9512
rect 3344 9081 3372 9506
rect 3330 9072 3386 9081
rect 3330 9007 3386 9016
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8498 3280 8910
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3148 8356 3200 8362
rect 3148 8298 3200 8304
rect 3068 8214 3188 8242
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2872 6792 2924 6798
rect 2872 6734 2924 6740
rect 3054 6760 3110 6769
rect 3160 6730 3188 8214
rect 3436 8072 3464 11494
rect 3549 11452 3857 11472
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11376 3857 11396
rect 3549 10364 3857 10384
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10288 3857 10308
rect 3608 10192 3660 10198
rect 3608 10134 3660 10140
rect 3620 9518 3648 10134
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9586 3832 9862
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 3608 9512 3660 9518
rect 3804 9489 3832 9522
rect 3608 9454 3660 9460
rect 3790 9480 3846 9489
rect 3790 9415 3846 9424
rect 3549 9276 3857 9296
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9200 3857 9220
rect 3516 9036 3568 9042
rect 3516 8978 3568 8984
rect 3528 8498 3556 8978
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3549 8188 3857 8208
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8112 3857 8132
rect 3252 8044 3464 8072
rect 3054 6695 3110 6704
rect 3148 6724 3200 6730
rect 2792 6616 2912 6644
rect 2688 6598 2740 6604
rect 2778 6488 2834 6497
rect 2596 6452 2648 6458
rect 2778 6423 2780 6432
rect 2596 6394 2648 6400
rect 2832 6423 2834 6432
rect 2780 6394 2832 6400
rect 2688 6384 2740 6390
rect 2688 6326 2740 6332
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 2504 5840 2556 5846
rect 2502 5808 2504 5817
rect 2556 5808 2558 5817
rect 2502 5743 2558 5752
rect 2228 5704 2280 5710
rect 2228 5646 2280 5652
rect 2504 5364 2556 5370
rect 2504 5306 2556 5312
rect 2516 5273 2544 5306
rect 2502 5264 2558 5273
rect 2502 5199 2558 5208
rect 2596 5024 2648 5030
rect 2596 4966 2648 4972
rect 2136 4276 2188 4282
rect 2136 4218 2188 4224
rect 2228 4072 2280 4078
rect 2228 4014 2280 4020
rect 1952 4004 2004 4010
rect 1952 3946 2004 3952
rect 2240 3913 2268 4014
rect 2226 3904 2282 3913
rect 2226 3839 2282 3848
rect 2240 3738 2268 3839
rect 2228 3732 2280 3738
rect 2228 3674 2280 3680
rect 1950 3632 2006 3641
rect 1950 3567 1952 3576
rect 2004 3567 2006 3576
rect 1952 3538 2004 3544
rect 2228 3528 2280 3534
rect 2226 3496 2228 3505
rect 2280 3496 2282 3505
rect 2226 3431 2282 3440
rect 1308 3392 1360 3398
rect 1308 3334 1360 3340
rect 2608 2650 2636 4966
rect 2700 4706 2728 6326
rect 2778 6216 2834 6225
rect 2778 6151 2834 6160
rect 2792 5710 2820 6151
rect 2884 5846 2912 6616
rect 3068 5846 3096 6695
rect 3148 6666 3200 6672
rect 3252 6440 3280 8044
rect 3332 7948 3384 7954
rect 3332 7890 3384 7896
rect 3344 7546 3372 7890
rect 3896 7868 3924 11562
rect 3988 11558 4016 12406
rect 4068 12378 4120 12384
rect 4080 12345 4108 12378
rect 4066 12336 4122 12345
rect 4066 12271 4122 12280
rect 3976 11552 4028 11558
rect 3976 11494 4028 11500
rect 3988 11218 4016 11494
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3976 10736 4028 10742
rect 3976 10678 4028 10684
rect 3988 10198 4016 10678
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 3976 10192 4028 10198
rect 3976 10134 4028 10140
rect 4080 10130 4108 10610
rect 4172 10266 4200 14758
rect 4264 13870 4292 17598
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4436 17536 4488 17542
rect 4436 17478 4488 17484
rect 4356 16658 4384 17478
rect 4448 16726 4476 17478
rect 4436 16720 4488 16726
rect 4436 16662 4488 16668
rect 4344 16652 4396 16658
rect 4344 16594 4396 16600
rect 4528 16584 4580 16590
rect 4528 16526 4580 16532
rect 4344 16516 4396 16522
rect 4344 16458 4396 16464
rect 4356 15706 4384 16458
rect 4436 16448 4488 16454
rect 4436 16390 4488 16396
rect 4448 16046 4476 16390
rect 4540 16250 4568 16526
rect 4528 16244 4580 16250
rect 4528 16186 4580 16192
rect 4436 16040 4488 16046
rect 4632 16017 4660 17598
rect 4804 17196 4856 17202
rect 4804 17138 4856 17144
rect 4816 16998 4844 17138
rect 4896 17128 4948 17134
rect 4896 17070 4948 17076
rect 4804 16992 4856 16998
rect 4804 16934 4856 16940
rect 4908 16658 4936 17070
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4436 15982 4488 15988
rect 4618 16008 4674 16017
rect 4618 15943 4674 15952
rect 4804 15972 4856 15978
rect 4804 15914 4856 15920
rect 4620 15904 4672 15910
rect 4816 15881 4844 15914
rect 4620 15846 4672 15852
rect 4802 15872 4858 15881
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4528 15360 4580 15366
rect 4528 15302 4580 15308
rect 4344 14816 4396 14822
rect 4344 14758 4396 14764
rect 4356 13938 4384 14758
rect 4344 13932 4396 13938
rect 4396 13892 4476 13920
rect 4344 13874 4396 13880
rect 4252 13864 4304 13870
rect 4252 13806 4304 13812
rect 4344 13456 4396 13462
rect 4344 13398 4396 13404
rect 4356 12782 4384 13398
rect 4344 12776 4396 12782
rect 4344 12718 4396 12724
rect 4448 11354 4476 13892
rect 4436 11348 4488 11354
rect 4436 11290 4488 11296
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4264 10810 4292 11018
rect 4342 10976 4398 10985
rect 4342 10911 4398 10920
rect 4252 10804 4304 10810
rect 4252 10746 4304 10752
rect 4160 10260 4212 10266
rect 4160 10202 4212 10208
rect 4068 10124 4120 10130
rect 4068 10066 4120 10072
rect 4252 9716 4304 9722
rect 4252 9658 4304 9664
rect 4068 9648 4120 9654
rect 4068 9590 4120 9596
rect 4080 9353 4108 9590
rect 4160 9444 4212 9450
rect 4160 9386 4212 9392
rect 4066 9344 4122 9353
rect 4066 9279 4122 9288
rect 4172 9110 4200 9386
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4264 8838 4292 9658
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4068 8560 4120 8566
rect 3974 8528 4030 8537
rect 4068 8502 4120 8508
rect 3974 8463 4030 8472
rect 3988 8276 4016 8463
rect 4080 8378 4108 8502
rect 4080 8350 4200 8378
rect 3988 8248 4108 8276
rect 3976 7880 4028 7886
rect 3896 7840 3976 7868
rect 3976 7822 4028 7828
rect 3422 7576 3478 7585
rect 3332 7540 3384 7546
rect 3422 7511 3478 7520
rect 3332 7482 3384 7488
rect 3436 7478 3464 7511
rect 3424 7472 3476 7478
rect 3424 7414 3476 7420
rect 3549 7100 3857 7120
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7024 3857 7044
rect 3790 6896 3846 6905
rect 3790 6831 3792 6840
rect 3844 6831 3846 6840
rect 3792 6802 3844 6808
rect 3976 6792 4028 6798
rect 3976 6734 4028 6740
rect 3160 6412 3280 6440
rect 3790 6488 3846 6497
rect 3988 6458 4016 6734
rect 3790 6423 3792 6432
rect 2872 5840 2924 5846
rect 2872 5782 2924 5788
rect 3056 5840 3108 5846
rect 3056 5782 3108 5788
rect 2780 5704 2832 5710
rect 2780 5646 2832 5652
rect 2780 5228 2832 5234
rect 2780 5170 2832 5176
rect 2792 4865 2820 5170
rect 2778 4856 2834 4865
rect 2778 4791 2834 4800
rect 2780 4752 2832 4758
rect 2700 4700 2780 4706
rect 2700 4694 2832 4700
rect 2700 4678 2820 4694
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 3194 2820 4422
rect 2884 3670 2912 5782
rect 3056 5364 3108 5370
rect 3160 5352 3188 6412
rect 3844 6423 3846 6432
rect 3976 6452 4028 6458
rect 3792 6394 3844 6400
rect 3976 6394 4028 6400
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 3252 5953 3280 6258
rect 3422 6216 3478 6225
rect 3804 6202 3832 6394
rect 4080 6390 4108 8248
rect 4172 8022 4200 8350
rect 4160 8016 4212 8022
rect 4160 7958 4212 7964
rect 4172 7410 4200 7958
rect 4252 7948 4304 7954
rect 4252 7890 4304 7896
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4160 7268 4212 7274
rect 4160 7210 4212 7216
rect 4172 6798 4200 7210
rect 4264 7002 4292 7890
rect 4252 6996 4304 7002
rect 4252 6938 4304 6944
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4252 6724 4304 6730
rect 4252 6666 4304 6672
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3804 6174 3924 6202
rect 3422 6151 3424 6160
rect 3476 6151 3478 6160
rect 3424 6122 3476 6128
rect 3330 6080 3386 6089
rect 3330 6015 3386 6024
rect 3238 5944 3294 5953
rect 3238 5879 3294 5888
rect 3252 5778 3280 5879
rect 3344 5846 3372 6015
rect 3549 6012 3857 6032
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5936 3857 5956
rect 3332 5840 3384 5846
rect 3332 5782 3384 5788
rect 3792 5840 3844 5846
rect 3792 5782 3844 5788
rect 3240 5772 3292 5778
rect 3240 5714 3292 5720
rect 3804 5574 3832 5782
rect 3240 5568 3292 5574
rect 3240 5510 3292 5516
rect 3792 5568 3844 5574
rect 3792 5510 3844 5516
rect 3108 5324 3188 5352
rect 3056 5306 3108 5312
rect 3252 5250 3280 5510
rect 3896 5352 3924 6174
rect 3976 6180 4028 6186
rect 3976 6122 4028 6128
rect 3988 5370 4016 6122
rect 3160 5222 3280 5250
rect 3620 5324 3924 5352
rect 3976 5364 4028 5370
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 3068 4078 3096 5102
rect 3056 4072 3108 4078
rect 3056 4014 3108 4020
rect 3160 3754 3188 5222
rect 3620 5012 3648 5324
rect 3976 5306 4028 5312
rect 3882 5264 3938 5273
rect 3882 5199 3938 5208
rect 3976 5228 4028 5234
rect 3344 4984 3648 5012
rect 3238 4040 3294 4049
rect 3238 3975 3240 3984
rect 3292 3975 3294 3984
rect 3240 3946 3292 3952
rect 3344 3890 3372 4984
rect 3549 4924 3857 4944
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4848 3857 4868
rect 3896 4826 3924 5199
rect 3976 5170 4028 5176
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3700 4548 3752 4554
rect 3700 4490 3752 4496
rect 3712 4146 3740 4490
rect 3988 4282 4016 5170
rect 4080 4826 4108 6326
rect 4160 6112 4212 6118
rect 4160 6054 4212 6060
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4172 4486 4200 6054
rect 4264 5030 4292 6666
rect 4356 6186 4384 10911
rect 4540 10810 4568 15302
rect 4632 14414 4660 15846
rect 4802 15807 4858 15816
rect 4908 15570 4936 16594
rect 4896 15564 4948 15570
rect 4896 15506 4948 15512
rect 4988 15496 5040 15502
rect 4988 15438 5040 15444
rect 4804 15428 4856 15434
rect 4804 15370 4856 15376
rect 4816 14906 4844 15370
rect 5000 15162 5028 15438
rect 4988 15156 5040 15162
rect 4988 15098 5040 15104
rect 4816 14878 5028 14906
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4724 13530 4752 13874
rect 4894 13560 4950 13569
rect 4712 13524 4764 13530
rect 4894 13495 4950 13504
rect 4712 13466 4764 13472
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4724 12986 4752 13126
rect 4712 12980 4764 12986
rect 4712 12922 4764 12928
rect 4620 12640 4672 12646
rect 4620 12582 4672 12588
rect 4528 10804 4580 10810
rect 4528 10746 4580 10752
rect 4526 10704 4582 10713
rect 4526 10639 4582 10648
rect 4540 8974 4568 10639
rect 4632 9625 4660 12582
rect 4804 12164 4856 12170
rect 4804 12106 4856 12112
rect 4816 11642 4844 12106
rect 4724 11614 4844 11642
rect 4724 9722 4752 11614
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4816 11218 4844 11494
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 4804 10668 4856 10674
rect 4804 10610 4856 10616
rect 4712 9716 4764 9722
rect 4712 9658 4764 9664
rect 4618 9616 4674 9625
rect 4618 9551 4674 9560
rect 4618 9480 4674 9489
rect 4618 9415 4620 9424
rect 4672 9415 4674 9424
rect 4620 9386 4672 9392
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 9104 4672 9110
rect 4620 9046 4672 9052
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4448 8498 4476 8774
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4448 6730 4476 8434
rect 4540 6934 4568 8910
rect 4528 6928 4580 6934
rect 4528 6870 4580 6876
rect 4632 6798 4660 9046
rect 4724 7954 4752 9318
rect 4816 8514 4844 10610
rect 4908 8634 4936 13495
rect 5000 10690 5028 14878
rect 5092 12442 5120 19314
rect 5184 19310 5212 19790
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 18766 5212 19246
rect 5276 18834 5304 20198
rect 5368 19446 5396 20318
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 5460 19514 5488 19858
rect 5552 19854 5580 20334
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5540 19712 5592 19718
rect 5540 19654 5592 19660
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5448 19236 5500 19242
rect 5448 19178 5500 19184
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5172 18760 5224 18766
rect 5172 18702 5224 18708
rect 5184 18358 5212 18702
rect 5172 18352 5224 18358
rect 5172 18294 5224 18300
rect 5184 17678 5212 18294
rect 5460 17814 5488 19178
rect 5552 18970 5580 19654
rect 5540 18964 5592 18970
rect 5540 18906 5592 18912
rect 5644 18873 5672 20878
rect 5736 20482 5764 22200
rect 6196 20942 6224 22200
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6148 20700 6456 20720
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20624 6456 20644
rect 6656 20584 6684 22200
rect 7010 22199 7066 22208
rect 7102 22200 7158 23000
rect 7562 22200 7618 23000
rect 7668 22222 7972 22250
rect 6828 20868 6880 20874
rect 6828 20810 6880 20816
rect 6472 20556 6684 20584
rect 5736 20454 5948 20482
rect 5724 20392 5776 20398
rect 5724 20334 5776 20340
rect 5816 20392 5868 20398
rect 5816 20334 5868 20340
rect 5630 18864 5686 18873
rect 5630 18799 5686 18808
rect 5736 18408 5764 20334
rect 5828 19378 5856 20334
rect 5816 19372 5868 19378
rect 5816 19314 5868 19320
rect 5552 18380 5764 18408
rect 5816 18420 5868 18426
rect 5552 17882 5580 18380
rect 5816 18362 5868 18368
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5540 17876 5592 17882
rect 5540 17818 5592 17824
rect 5448 17808 5500 17814
rect 5448 17750 5500 17756
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 17134 5212 17614
rect 5632 17604 5684 17610
rect 5632 17546 5684 17552
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5172 17128 5224 17134
rect 5172 17070 5224 17076
rect 5172 16992 5224 16998
rect 5172 16934 5224 16940
rect 5184 16794 5212 16934
rect 5172 16788 5224 16794
rect 5172 16730 5224 16736
rect 5172 15564 5224 15570
rect 5172 15506 5224 15512
rect 5184 15094 5212 15506
rect 5276 15162 5304 17274
rect 5448 16040 5500 16046
rect 5448 15982 5500 15988
rect 5540 16040 5592 16046
rect 5540 15982 5592 15988
rect 5460 15502 5488 15982
rect 5448 15496 5500 15502
rect 5448 15438 5500 15444
rect 5264 15156 5316 15162
rect 5264 15098 5316 15104
rect 5172 15088 5224 15094
rect 5172 15030 5224 15036
rect 5184 14482 5212 15030
rect 5448 15020 5500 15026
rect 5448 14962 5500 14968
rect 5460 14618 5488 14962
rect 5448 14612 5500 14618
rect 5448 14554 5500 14560
rect 5172 14476 5224 14482
rect 5172 14418 5224 14424
rect 5448 14272 5500 14278
rect 5448 14214 5500 14220
rect 5460 13954 5488 14214
rect 5552 14074 5580 15982
rect 5540 14068 5592 14074
rect 5540 14010 5592 14016
rect 5172 13932 5224 13938
rect 5460 13926 5580 13954
rect 5172 13874 5224 13880
rect 5184 12918 5212 13874
rect 5356 13252 5408 13258
rect 5356 13194 5408 13200
rect 5172 12912 5224 12918
rect 5172 12854 5224 12860
rect 5080 12436 5132 12442
rect 5080 12378 5132 12384
rect 5368 10810 5396 13194
rect 5448 11280 5500 11286
rect 5448 11222 5500 11228
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5000 10662 5212 10690
rect 5460 10674 5488 11222
rect 5080 10600 5132 10606
rect 5080 10542 5132 10548
rect 5092 10130 5120 10542
rect 5080 10124 5132 10130
rect 5080 10066 5132 10072
rect 4988 10056 5040 10062
rect 4988 9998 5040 10004
rect 5000 9178 5028 9998
rect 5080 9580 5132 9586
rect 5080 9522 5132 9528
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 4988 8832 5040 8838
rect 4988 8774 5040 8780
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 4816 8486 4936 8514
rect 4804 8288 4856 8294
rect 4804 8230 4856 8236
rect 4816 7954 4844 8230
rect 4712 7948 4764 7954
rect 4712 7890 4764 7896
rect 4804 7948 4856 7954
rect 4804 7890 4856 7896
rect 4816 7410 4844 7890
rect 4908 7750 4936 8486
rect 5000 7886 5028 8774
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 4896 7744 4948 7750
rect 5092 7732 5120 9522
rect 5184 9110 5212 10662
rect 5448 10668 5500 10674
rect 5448 10610 5500 10616
rect 5354 10568 5410 10577
rect 5354 10503 5410 10512
rect 5264 9920 5316 9926
rect 5264 9862 5316 9868
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5172 8832 5224 8838
rect 5172 8774 5224 8780
rect 4896 7686 4948 7692
rect 5000 7704 5120 7732
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 4816 6866 4844 7346
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4620 6792 4672 6798
rect 4620 6734 4672 6740
rect 4436 6724 4488 6730
rect 4436 6666 4488 6672
rect 4528 6656 4580 6662
rect 4528 6598 4580 6604
rect 4344 6180 4396 6186
rect 4344 6122 4396 6128
rect 4436 6180 4488 6186
rect 4436 6122 4488 6128
rect 4448 5846 4476 6122
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4344 5568 4396 5574
rect 4344 5510 4396 5516
rect 4252 5024 4304 5030
rect 4252 4966 4304 4972
rect 4160 4480 4212 4486
rect 4160 4422 4212 4428
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3344 3862 3464 3890
rect 3160 3726 3372 3754
rect 2872 3664 2924 3670
rect 2872 3606 2924 3612
rect 2872 3460 2924 3466
rect 2872 3402 2924 3408
rect 2884 3346 2912 3402
rect 2884 3318 3096 3346
rect 2780 3188 2832 3194
rect 2780 3130 2832 3136
rect 2780 3052 2832 3058
rect 2780 2994 2832 3000
rect 2792 2961 2820 2994
rect 2872 2984 2924 2990
rect 2778 2952 2834 2961
rect 2872 2926 2924 2932
rect 2778 2887 2834 2896
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 2778 2544 2834 2553
rect 2778 2479 2834 2488
rect 2792 2446 2820 2479
rect 2780 2440 2832 2446
rect 2780 2382 2832 2388
rect 2780 2304 2832 2310
rect 2780 2246 2832 2252
rect 2792 241 2820 2246
rect 2884 649 2912 2926
rect 2964 2916 3016 2922
rect 2964 2858 3016 2864
rect 2976 2378 3004 2858
rect 3068 2854 3096 3318
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3240 2848 3292 2854
rect 3240 2790 3292 2796
rect 2964 2372 3016 2378
rect 2964 2314 3016 2320
rect 3068 2009 3096 2790
rect 3252 2378 3280 2790
rect 3344 2650 3372 3726
rect 3332 2644 3384 2650
rect 3332 2586 3384 2592
rect 3436 2514 3464 3862
rect 3549 3836 3857 3856
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3760 3857 3780
rect 3549 2748 3857 2768
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2672 3857 2692
rect 4264 2650 4292 4966
rect 4356 3602 4384 5510
rect 4540 3641 4568 6598
rect 4632 6118 4660 6734
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4712 6112 4764 6118
rect 4712 6054 4764 6060
rect 4618 5944 4674 5953
rect 4618 5879 4620 5888
rect 4672 5879 4674 5888
rect 4620 5850 4672 5856
rect 4618 5536 4674 5545
rect 4618 5471 4674 5480
rect 4632 5370 4660 5471
rect 4620 5364 4672 5370
rect 4620 5306 4672 5312
rect 4526 3632 4582 3641
rect 4344 3596 4396 3602
rect 4526 3567 4582 3576
rect 4344 3538 4396 3544
rect 4724 3126 4752 6054
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4908 2582 4936 7686
rect 5000 6118 5028 7704
rect 5080 6656 5132 6662
rect 5184 6644 5212 8774
rect 5132 6616 5212 6644
rect 5080 6598 5132 6604
rect 5276 6186 5304 9862
rect 5368 9586 5396 10503
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5368 8378 5396 9522
rect 5448 9512 5500 9518
rect 5448 9454 5500 9460
rect 5460 9178 5488 9454
rect 5448 9172 5500 9178
rect 5448 9114 5500 9120
rect 5368 8350 5488 8378
rect 5552 8362 5580 13926
rect 5644 13326 5672 17546
rect 5736 17338 5764 18226
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5736 14414 5764 15438
rect 5724 14408 5776 14414
rect 5724 14350 5776 14356
rect 5724 14000 5776 14006
rect 5724 13942 5776 13948
rect 5736 13394 5764 13942
rect 5724 13388 5776 13394
rect 5724 13330 5776 13336
rect 5632 13320 5684 13326
rect 5632 13262 5684 13268
rect 5736 12918 5764 13330
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 5736 12238 5764 12854
rect 5724 12232 5776 12238
rect 5724 12174 5776 12180
rect 5736 11762 5764 12174
rect 5828 11898 5856 18362
rect 5920 17785 5948 20454
rect 5998 19816 6054 19825
rect 5998 19751 6054 19760
rect 6012 18766 6040 19751
rect 6472 19700 6500 20556
rect 6736 20460 6788 20466
rect 6736 20402 6788 20408
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 19854 6684 20198
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6644 19712 6696 19718
rect 6472 19672 6592 19700
rect 6148 19612 6456 19632
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19536 6456 19556
rect 6564 19496 6592 19672
rect 6644 19654 6696 19660
rect 6472 19468 6592 19496
rect 6092 19372 6144 19378
rect 6092 19314 6144 19320
rect 6104 18873 6132 19314
rect 6090 18864 6146 18873
rect 6090 18799 6146 18808
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 6472 18612 6500 19468
rect 6550 19408 6606 19417
rect 6550 19343 6552 19352
rect 6604 19343 6606 19352
rect 6552 19314 6604 19320
rect 6472 18584 6592 18612
rect 6148 18524 6456 18544
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 5998 18456 6054 18465
rect 6148 18448 6456 18468
rect 5998 18391 6054 18400
rect 6012 17882 6040 18391
rect 6458 18320 6514 18329
rect 6458 18255 6460 18264
rect 6512 18255 6514 18264
rect 6460 18226 6512 18232
rect 6000 17876 6052 17882
rect 6000 17818 6052 17824
rect 5906 17776 5962 17785
rect 5906 17711 5962 17720
rect 6000 17740 6052 17746
rect 6000 17682 6052 17688
rect 5908 17536 5960 17542
rect 5906 17504 5908 17513
rect 5960 17504 5962 17513
rect 5906 17439 5962 17448
rect 5908 17332 5960 17338
rect 5908 17274 5960 17280
rect 5920 17082 5948 17274
rect 6012 17202 6040 17682
rect 6564 17678 6592 18584
rect 6552 17672 6604 17678
rect 6552 17614 6604 17620
rect 6148 17436 6456 17456
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17360 6456 17380
rect 6656 17338 6684 19654
rect 6748 18970 6776 20402
rect 6736 18964 6788 18970
rect 6736 18906 6788 18912
rect 6840 18426 6868 20810
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 6828 18420 6880 18426
rect 6828 18362 6880 18368
rect 6932 18222 6960 19790
rect 7024 19514 7052 22199
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 7012 18760 7064 18766
rect 7012 18702 7064 18708
rect 6920 18216 6972 18222
rect 6920 18158 6972 18164
rect 6828 18080 6880 18086
rect 6828 18022 6880 18028
rect 6736 17536 6788 17542
rect 6736 17478 6788 17484
rect 6644 17332 6696 17338
rect 6644 17274 6696 17280
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 6276 17196 6328 17202
rect 6276 17138 6328 17144
rect 6644 17196 6696 17202
rect 6644 17138 6696 17144
rect 5920 17054 6040 17082
rect 6012 16182 6040 17054
rect 6288 16794 6316 17138
rect 6276 16788 6328 16794
rect 6276 16730 6328 16736
rect 6552 16584 6604 16590
rect 6552 16526 6604 16532
rect 6148 16348 6456 16368
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16272 6456 16292
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 6092 15972 6144 15978
rect 6092 15914 6144 15920
rect 6104 15502 6132 15914
rect 6092 15496 6144 15502
rect 6092 15438 6144 15444
rect 6148 15260 6456 15280
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15184 6456 15204
rect 6564 14618 6592 16526
rect 5908 14612 5960 14618
rect 5908 14554 5960 14560
rect 6552 14612 6604 14618
rect 6552 14554 6604 14560
rect 5920 12782 5948 14554
rect 6000 14408 6052 14414
rect 6000 14350 6052 14356
rect 6012 14074 6040 14350
rect 6552 14340 6604 14346
rect 6552 14282 6604 14288
rect 6148 14172 6456 14192
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14096 6456 14116
rect 6564 14074 6592 14282
rect 6000 14068 6052 14074
rect 6000 14010 6052 14016
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6552 13388 6604 13394
rect 6552 13330 6604 13336
rect 6148 13084 6456 13104
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13008 6456 13028
rect 5908 12776 5960 12782
rect 5908 12718 5960 12724
rect 6564 12442 6592 13330
rect 6656 12714 6684 17138
rect 6748 13530 6776 17478
rect 6840 16096 6868 18022
rect 7024 17746 7052 18702
rect 7116 18426 7144 22200
rect 7196 19712 7248 19718
rect 7196 19654 7248 19660
rect 7208 19446 7236 19654
rect 7288 19508 7340 19514
rect 7288 19450 7340 19456
rect 7196 19440 7248 19446
rect 7196 19382 7248 19388
rect 7196 19304 7248 19310
rect 7196 19246 7248 19252
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7208 18086 7236 19246
rect 7196 18080 7248 18086
rect 7196 18022 7248 18028
rect 7300 17814 7328 19450
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7380 19304 7432 19310
rect 7380 19246 7432 19252
rect 7392 18329 7420 19246
rect 7378 18320 7434 18329
rect 7378 18255 7434 18264
rect 7484 18193 7512 19314
rect 7576 18902 7604 22200
rect 7564 18896 7616 18902
rect 7564 18838 7616 18844
rect 7668 18714 7696 22222
rect 7944 22114 7972 22222
rect 8022 22200 8078 23000
rect 8482 22200 8538 23000
rect 8588 22222 8892 22250
rect 8036 22114 8064 22200
rect 7944 22086 8064 22114
rect 8496 22114 8524 22200
rect 8588 22114 8616 22222
rect 8496 22086 8616 22114
rect 8392 20800 8444 20806
rect 8392 20742 8444 20748
rect 8300 20460 8352 20466
rect 8300 20402 8352 20408
rect 8022 20224 8078 20233
rect 8022 20159 8078 20168
rect 7840 19168 7892 19174
rect 7840 19110 7892 19116
rect 7576 18686 7696 18714
rect 7746 18728 7802 18737
rect 7470 18184 7526 18193
rect 7470 18119 7526 18128
rect 7288 17808 7340 17814
rect 7288 17750 7340 17756
rect 7012 17740 7064 17746
rect 7012 17682 7064 17688
rect 7024 17338 7052 17682
rect 7288 17536 7340 17542
rect 7288 17478 7340 17484
rect 7472 17536 7524 17542
rect 7472 17478 7524 17484
rect 7012 17332 7064 17338
rect 7012 17274 7064 17280
rect 7300 16794 7328 17478
rect 7288 16788 7340 16794
rect 7288 16730 7340 16736
rect 7196 16448 7248 16454
rect 7196 16390 7248 16396
rect 7104 16108 7156 16114
rect 6840 16068 7104 16096
rect 7104 16050 7156 16056
rect 6826 16008 6882 16017
rect 6882 15978 7052 15994
rect 6882 15972 7064 15978
rect 6882 15966 7012 15972
rect 6826 15943 6882 15952
rect 7012 15914 7064 15920
rect 7104 15972 7156 15978
rect 7104 15914 7156 15920
rect 7116 15881 7144 15914
rect 7102 15872 7158 15881
rect 7102 15807 7158 15816
rect 6920 15360 6972 15366
rect 6920 15302 6972 15308
rect 6828 13728 6880 13734
rect 6828 13670 6880 13676
rect 6736 13524 6788 13530
rect 6736 13466 6788 13472
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6840 12594 6868 13670
rect 6932 12850 6960 15302
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7116 14414 7144 14962
rect 7104 14408 7156 14414
rect 7104 14350 7156 14356
rect 7012 13932 7064 13938
rect 7012 13874 7064 13880
rect 7024 13326 7052 13874
rect 7012 13320 7064 13326
rect 7012 13262 7064 13268
rect 6920 12844 6972 12850
rect 6920 12786 6972 12792
rect 6656 12566 6868 12594
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6552 12436 6604 12442
rect 6552 12378 6604 12384
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5724 11756 5776 11762
rect 5724 11698 5776 11704
rect 5736 10742 5764 11698
rect 5816 11348 5868 11354
rect 5816 11290 5868 11296
rect 5724 10736 5776 10742
rect 5724 10678 5776 10684
rect 5736 10266 5764 10678
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 8974 5672 9862
rect 5736 9722 5764 10202
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5828 9466 5856 11290
rect 5920 10674 5948 12378
rect 6000 12096 6052 12102
rect 6000 12038 6052 12044
rect 6012 11762 6040 12038
rect 6148 11996 6456 12016
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11920 6456 11940
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6012 11626 6040 11698
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 6012 11218 6040 11562
rect 6550 11520 6606 11529
rect 6550 11455 6606 11464
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6012 10810 6040 11018
rect 6148 10908 6456 10928
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10832 6456 10852
rect 6000 10804 6052 10810
rect 6000 10746 6052 10752
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 6000 10464 6052 10470
rect 6000 10406 6052 10412
rect 5736 9438 5856 9466
rect 5632 8968 5684 8974
rect 5632 8910 5684 8916
rect 5736 8838 5764 9438
rect 5816 9104 5868 9110
rect 5816 9046 5868 9052
rect 5724 8832 5776 8838
rect 5724 8774 5776 8780
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5460 8242 5488 8350
rect 5540 8356 5592 8362
rect 5540 8298 5592 8304
rect 5460 8214 5672 8242
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5264 6180 5316 6186
rect 5264 6122 5316 6128
rect 5368 6118 5396 6870
rect 5552 6798 5580 7482
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5644 6390 5672 8214
rect 5736 6730 5764 8366
rect 5828 7206 5856 9046
rect 5908 8424 5960 8430
rect 5908 8366 5960 8372
rect 5920 8090 5948 8366
rect 5908 8084 5960 8090
rect 5908 8026 5960 8032
rect 6012 7936 6040 10406
rect 6148 9820 6456 9840
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9744 6456 9764
rect 6564 8838 6592 11455
rect 6552 8832 6604 8838
rect 6552 8774 6604 8780
rect 6148 8732 6456 8752
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8656 6456 8676
rect 6460 8492 6512 8498
rect 6564 8480 6592 8774
rect 6512 8452 6592 8480
rect 6460 8434 6512 8440
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 6104 7993 6132 8366
rect 5920 7908 6040 7936
rect 6090 7984 6146 7993
rect 6090 7919 6146 7928
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5920 7002 5948 7908
rect 6656 7868 6684 12566
rect 7208 12238 7236 16390
rect 7288 15904 7340 15910
rect 7288 15846 7340 15852
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 6736 11824 6788 11830
rect 6736 11766 6788 11772
rect 6748 11286 6776 11766
rect 6736 11280 6788 11286
rect 6736 11222 6788 11228
rect 7012 10736 7064 10742
rect 7012 10678 7064 10684
rect 6920 10464 6972 10470
rect 6920 10406 6972 10412
rect 6736 10192 6788 10198
rect 6736 10134 6788 10140
rect 6748 9042 6776 10134
rect 6826 9616 6882 9625
rect 6826 9551 6828 9560
rect 6880 9551 6882 9560
rect 6828 9522 6880 9528
rect 6932 9353 6960 10406
rect 7024 10062 7052 10678
rect 7012 10056 7064 10062
rect 7012 9998 7064 10004
rect 6918 9344 6974 9353
rect 6918 9279 6974 9288
rect 6736 9036 6788 9042
rect 6736 8978 6788 8984
rect 7300 8401 7328 15846
rect 7380 15360 7432 15366
rect 7380 15302 7432 15308
rect 7392 14822 7420 15302
rect 7380 14816 7432 14822
rect 7380 14758 7432 14764
rect 7484 14346 7512 17478
rect 7576 14906 7604 18686
rect 7746 18663 7802 18672
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7668 15094 7696 18566
rect 7760 16794 7788 18663
rect 7852 18329 7880 19110
rect 7932 18624 7984 18630
rect 7932 18566 7984 18572
rect 7838 18320 7894 18329
rect 7838 18255 7894 18264
rect 7944 17270 7972 18566
rect 7932 17264 7984 17270
rect 7932 17206 7984 17212
rect 7748 16788 7800 16794
rect 7748 16730 7800 16736
rect 7932 16652 7984 16658
rect 7932 16594 7984 16600
rect 7840 16448 7892 16454
rect 7840 16390 7892 16396
rect 7852 15434 7880 16390
rect 7840 15428 7892 15434
rect 7840 15370 7892 15376
rect 7748 15360 7800 15366
rect 7748 15302 7800 15308
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7576 14878 7696 14906
rect 7472 14340 7524 14346
rect 7472 14282 7524 14288
rect 7564 13864 7616 13870
rect 7564 13806 7616 13812
rect 7576 13462 7604 13806
rect 7564 13456 7616 13462
rect 7564 13398 7616 13404
rect 7472 13320 7524 13326
rect 7472 13262 7524 13268
rect 7484 12434 7512 13262
rect 7564 12844 7616 12850
rect 7564 12786 7616 12792
rect 7392 12406 7512 12434
rect 7392 12345 7420 12406
rect 7472 12368 7524 12374
rect 7378 12336 7434 12345
rect 7472 12310 7524 12316
rect 7378 12271 7434 12280
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7392 10606 7420 11018
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7392 9081 7420 10542
rect 7378 9072 7434 9081
rect 7378 9007 7434 9016
rect 7286 8392 7342 8401
rect 7286 8327 7342 8336
rect 7104 8288 7156 8294
rect 7104 8230 7156 8236
rect 6564 7840 6684 7868
rect 6000 7812 6052 7818
rect 6000 7754 6052 7760
rect 6012 7002 6040 7754
rect 6148 7644 6456 7664
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7568 6456 7588
rect 6564 7546 6592 7840
rect 6644 7744 6696 7750
rect 6644 7686 6696 7692
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6656 7478 6684 7686
rect 6644 7472 6696 7478
rect 6644 7414 6696 7420
rect 5908 6996 5960 7002
rect 5908 6938 5960 6944
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5080 6112 5132 6118
rect 5080 6054 5132 6060
rect 5356 6112 5408 6118
rect 5356 6054 5408 6060
rect 4986 5944 5042 5953
rect 4986 5879 4988 5888
rect 5040 5879 5042 5888
rect 4988 5850 5040 5856
rect 5092 5098 5120 6054
rect 5354 5944 5410 5953
rect 5354 5879 5356 5888
rect 5408 5879 5410 5888
rect 5356 5850 5408 5856
rect 5368 5794 5396 5850
rect 5276 5766 5396 5794
rect 5276 5574 5304 5766
rect 5356 5636 5408 5642
rect 5356 5578 5408 5584
rect 5264 5568 5316 5574
rect 5264 5510 5316 5516
rect 5368 5370 5396 5578
rect 5920 5370 5948 6938
rect 7116 6662 7144 8230
rect 7392 7274 7420 9007
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 6148 6556 6456 6576
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6480 6456 6500
rect 7116 6118 7144 6598
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 6148 5468 6456 5488
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5392 6456 5412
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5080 5092 5132 5098
rect 5080 5034 5132 5040
rect 6148 4380 6456 4400
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4304 6456 4324
rect 7392 4214 7420 7210
rect 7484 5234 7512 12310
rect 7576 10266 7604 12786
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7668 9625 7696 14878
rect 7654 9616 7710 9625
rect 7654 9551 7710 9560
rect 7760 9382 7788 15302
rect 7840 13184 7892 13190
rect 7840 13126 7892 13132
rect 7852 12918 7880 13126
rect 7840 12912 7892 12918
rect 7840 12854 7892 12860
rect 7840 11824 7892 11830
rect 7840 11766 7892 11772
rect 7852 11286 7880 11766
rect 7944 11354 7972 16594
rect 8036 16538 8064 20159
rect 8312 18834 8340 20402
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8208 18760 8260 18766
rect 8208 18702 8260 18708
rect 8220 18086 8248 18702
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8208 18080 8260 18086
rect 8128 18040 8208 18068
rect 8128 16658 8156 18040
rect 8208 18022 8260 18028
rect 8312 17218 8340 18362
rect 8220 17190 8340 17218
rect 8116 16652 8168 16658
rect 8116 16594 8168 16600
rect 8036 16510 8156 16538
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 8036 12986 8064 14214
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 8128 12374 8156 16510
rect 8220 15586 8248 17190
rect 8300 17128 8352 17134
rect 8300 17070 8352 17076
rect 8312 16266 8340 17070
rect 8404 16590 8432 20742
rect 8864 20618 8892 22222
rect 8942 22200 8998 23000
rect 9402 22200 9458 23000
rect 9862 22200 9918 23000
rect 10322 22200 10378 23000
rect 10782 22200 10838 23000
rect 11242 22200 11298 23000
rect 11702 22200 11758 23000
rect 12162 22200 12218 23000
rect 12622 22200 12678 23000
rect 13082 22200 13138 23000
rect 13542 22200 13598 23000
rect 14002 22200 14058 23000
rect 14462 22200 14518 23000
rect 14922 22200 14978 23000
rect 15382 22200 15438 23000
rect 15842 22200 15898 23000
rect 16302 22200 16358 23000
rect 16762 22200 16818 23000
rect 17222 22200 17278 23000
rect 17682 22200 17738 23000
rect 18142 22200 18198 23000
rect 18602 22200 18658 23000
rect 19062 22200 19118 23000
rect 19522 22200 19578 23000
rect 19982 22200 20038 23000
rect 20442 22200 20498 23000
rect 20902 22200 20958 23000
rect 21362 22200 21418 23000
rect 21822 22200 21878 23000
rect 22282 22200 22338 23000
rect 22742 22200 22798 23000
rect 8956 20806 8984 22200
rect 9128 21344 9180 21350
rect 9128 21286 9180 21292
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8484 20596 8536 20602
rect 8864 20590 9076 20618
rect 9140 20602 9168 21286
rect 8484 20538 8536 20544
rect 8496 19718 8524 20538
rect 8668 20460 8720 20466
rect 8668 20402 8720 20408
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8484 19712 8536 19718
rect 8484 19654 8536 19660
rect 8588 19530 8616 19994
rect 8680 19922 8708 20402
rect 8956 20369 8984 20402
rect 8942 20360 8998 20369
rect 9048 20346 9076 20590
rect 9128 20596 9180 20602
rect 9128 20538 9180 20544
rect 9416 20398 9444 22200
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9404 20392 9456 20398
rect 9048 20318 9168 20346
rect 9404 20334 9456 20340
rect 8942 20295 8998 20304
rect 8747 20156 9055 20176
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20080 9055 20100
rect 8760 19984 8812 19990
rect 8758 19952 8760 19961
rect 8812 19952 8814 19961
rect 8668 19916 8720 19922
rect 8758 19887 8814 19896
rect 8668 19858 8720 19864
rect 8496 19502 8616 19530
rect 8680 19514 8708 19858
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8668 19508 8720 19514
rect 8496 18970 8524 19502
rect 8668 19450 8720 19456
rect 8864 19378 8892 19654
rect 8576 19372 8628 19378
rect 8576 19314 8628 19320
rect 8852 19372 8904 19378
rect 8852 19314 8904 19320
rect 8484 18964 8536 18970
rect 8484 18906 8536 18912
rect 8496 18426 8524 18906
rect 8484 18420 8536 18426
rect 8484 18362 8536 18368
rect 8484 17672 8536 17678
rect 8484 17614 8536 17620
rect 8392 16584 8444 16590
rect 8392 16526 8444 16532
rect 8312 16250 8432 16266
rect 8300 16244 8432 16250
rect 8352 16238 8432 16244
rect 8300 16186 8352 16192
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8312 15706 8340 16050
rect 8300 15700 8352 15706
rect 8300 15642 8352 15648
rect 8404 15638 8432 16238
rect 8392 15632 8444 15638
rect 8220 15558 8340 15586
rect 8392 15574 8444 15580
rect 8312 15366 8340 15558
rect 8496 15434 8524 17614
rect 8588 15706 8616 19314
rect 8747 19068 9055 19088
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 18992 9055 19012
rect 8747 17980 9055 18000
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17904 9055 17924
rect 8944 17740 8996 17746
rect 8944 17682 8996 17688
rect 8956 17649 8984 17682
rect 8942 17640 8998 17649
rect 8942 17575 8998 17584
rect 8747 16892 9055 16912
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16816 9055 16836
rect 9140 16674 9168 20318
rect 9220 19848 9272 19854
rect 9220 19790 9272 19796
rect 9232 17746 9260 19790
rect 9312 19712 9364 19718
rect 9312 19654 9364 19660
rect 9220 17740 9272 17746
rect 9220 17682 9272 17688
rect 9232 17134 9260 17682
rect 9324 17338 9352 19654
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9416 17218 9444 20334
rect 9508 18698 9536 20402
rect 9588 20392 9640 20398
rect 9588 20334 9640 20340
rect 9600 19854 9628 20334
rect 9680 20052 9732 20058
rect 9680 19994 9732 20000
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19378 9628 19654
rect 9588 19372 9640 19378
rect 9588 19314 9640 19320
rect 9496 18692 9548 18698
rect 9496 18634 9548 18640
rect 9600 18578 9628 19314
rect 9692 19310 9720 19994
rect 9772 19712 9824 19718
rect 9772 19654 9824 19660
rect 9680 19304 9732 19310
rect 9680 19246 9732 19252
rect 9784 18834 9812 19654
rect 9772 18828 9824 18834
rect 9772 18770 9824 18776
rect 9324 17202 9444 17218
rect 9312 17196 9444 17202
rect 9364 17190 9444 17196
rect 9508 18550 9628 18578
rect 9312 17138 9364 17144
rect 9220 17128 9272 17134
rect 9508 17082 9536 18550
rect 9588 18420 9640 18426
rect 9588 18362 9640 18368
rect 9600 17354 9628 18362
rect 9772 18284 9824 18290
rect 9772 18226 9824 18232
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17610 9720 18022
rect 9680 17604 9732 17610
rect 9680 17546 9732 17552
rect 9784 17490 9812 18226
rect 9876 17610 9904 22200
rect 10048 19916 10100 19922
rect 10048 19858 10100 19864
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9864 17604 9916 17610
rect 9864 17546 9916 17552
rect 9784 17462 9904 17490
rect 9678 17368 9734 17377
rect 9600 17326 9678 17354
rect 9678 17303 9734 17312
rect 9680 17196 9732 17202
rect 9680 17138 9732 17144
rect 9220 17070 9272 17076
rect 9232 16794 9260 17070
rect 9416 17054 9536 17082
rect 9586 17096 9642 17105
rect 9220 16788 9272 16794
rect 9220 16730 9272 16736
rect 9312 16720 9364 16726
rect 9140 16646 9260 16674
rect 9312 16662 9364 16668
rect 8668 16584 8720 16590
rect 8760 16584 8812 16590
rect 8668 16526 8720 16532
rect 8758 16552 8760 16561
rect 8812 16552 8814 16561
rect 8576 15700 8628 15706
rect 8576 15642 8628 15648
rect 8680 15502 8708 16526
rect 8758 16487 8814 16496
rect 9126 16008 9182 16017
rect 9126 15943 9182 15952
rect 8747 15804 9055 15824
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15728 9055 15748
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 8484 15428 8536 15434
rect 8484 15370 8536 15376
rect 8576 15428 8628 15434
rect 8576 15370 8628 15376
rect 8300 15360 8352 15366
rect 8300 15302 8352 15308
rect 8312 14618 8340 15302
rect 8496 15162 8524 15370
rect 8484 15156 8536 15162
rect 8484 15098 8536 15104
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8300 14612 8352 14618
rect 8300 14554 8352 14560
rect 8404 14074 8432 14758
rect 8392 14068 8444 14074
rect 8392 14010 8444 14016
rect 8484 14000 8536 14006
rect 8484 13942 8536 13948
rect 8496 13258 8524 13942
rect 8588 13530 8616 15370
rect 9140 15178 9168 15943
rect 9048 15162 9168 15178
rect 9036 15156 9168 15162
rect 9088 15150 9168 15156
rect 9036 15098 9088 15104
rect 9036 14952 9088 14958
rect 9088 14900 9168 14906
rect 9036 14894 9168 14900
rect 9048 14878 9168 14894
rect 8747 14716 9055 14736
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14640 9055 14660
rect 9140 14074 9168 14878
rect 9128 14068 9180 14074
rect 9128 14010 9180 14016
rect 8668 13796 8720 13802
rect 8668 13738 8720 13744
rect 8576 13524 8628 13530
rect 8576 13466 8628 13472
rect 8680 13394 8708 13738
rect 8747 13628 9055 13648
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13552 9055 13572
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8484 13252 8536 13258
rect 8484 13194 8536 13200
rect 8680 12986 8708 13330
rect 9140 13326 9168 14010
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8668 12980 8720 12986
rect 8668 12922 8720 12928
rect 8300 12776 8352 12782
rect 8300 12718 8352 12724
rect 8116 12368 8168 12374
rect 8116 12310 8168 12316
rect 8024 12300 8076 12306
rect 8024 12242 8076 12248
rect 8036 11898 8064 12242
rect 8312 12170 8340 12718
rect 8747 12540 9055 12560
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12464 9055 12484
rect 9232 12434 9260 16646
rect 9324 15706 9352 16662
rect 9312 15700 9364 15706
rect 9312 15642 9364 15648
rect 9312 15156 9364 15162
rect 9312 15098 9364 15104
rect 9140 12406 9260 12434
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 8300 12164 8352 12170
rect 8300 12106 8352 12112
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8208 12096 8260 12102
rect 8208 12038 8260 12044
rect 8024 11892 8076 11898
rect 8024 11834 8076 11840
rect 7932 11348 7984 11354
rect 7932 11290 7984 11296
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 7852 10538 7880 11222
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7944 10985 7972 11018
rect 7930 10976 7986 10985
rect 7930 10911 7986 10920
rect 7840 10532 7892 10538
rect 7840 10474 7892 10480
rect 8036 10062 8064 11834
rect 8128 10810 8156 12038
rect 8220 11354 8248 12038
rect 8312 11558 8340 12106
rect 8392 12096 8444 12102
rect 8392 12038 8444 12044
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 8312 11218 8340 11494
rect 8300 11212 8352 11218
rect 8300 11154 8352 11160
rect 8116 10804 8168 10810
rect 8116 10746 8168 10752
rect 8404 10674 8432 12038
rect 8496 11082 8524 12271
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 11552 8628 11558
rect 8576 11494 8628 11500
rect 8484 11076 8536 11082
rect 8484 11018 8536 11024
rect 8392 10668 8444 10674
rect 8392 10610 8444 10616
rect 8496 10282 8524 11018
rect 8312 10254 8524 10282
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8312 9654 8340 10254
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8392 9716 8444 9722
rect 8392 9658 8444 9664
rect 8300 9648 8352 9654
rect 8220 9608 8300 9636
rect 7748 9376 7800 9382
rect 7748 9318 7800 9324
rect 8220 9081 8248 9608
rect 8300 9590 8352 9596
rect 8300 9512 8352 9518
rect 8300 9454 8352 9460
rect 8206 9072 8262 9081
rect 8024 9036 8076 9042
rect 8206 9007 8262 9016
rect 8024 8978 8076 8984
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 8294 7696 8774
rect 7748 8424 7800 8430
rect 7748 8366 7800 8372
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7760 7818 7788 8366
rect 8036 8362 8064 8978
rect 8024 8356 8076 8362
rect 8024 8298 8076 8304
rect 7748 7812 7800 7818
rect 7748 7754 7800 7760
rect 7760 7206 7788 7754
rect 8312 7410 8340 9454
rect 8404 8650 8432 9658
rect 8496 9518 8524 9998
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8484 9376 8536 9382
rect 8484 9318 8536 9324
rect 8496 8974 8524 9318
rect 8484 8968 8536 8974
rect 8484 8910 8536 8916
rect 8404 8622 8524 8650
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8404 7546 8432 8434
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8496 7449 8524 8622
rect 8482 7440 8538 7449
rect 8300 7404 8352 7410
rect 8482 7375 8538 7384
rect 8300 7346 8352 7352
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 7562 6896 7618 6905
rect 7760 6866 7788 7142
rect 7562 6831 7618 6840
rect 7748 6860 7800 6866
rect 7576 5681 7604 6831
rect 7748 6802 7800 6808
rect 8128 6798 8156 7142
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8312 6458 8340 7346
rect 8588 7342 8616 11494
rect 8680 9722 8708 12174
rect 8747 11452 9055 11472
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11376 9055 11396
rect 9140 11150 9168 12406
rect 9324 11558 9352 15098
rect 9312 11552 9364 11558
rect 9312 11494 9364 11500
rect 9416 11370 9444 17054
rect 9586 17031 9642 17040
rect 9600 15910 9628 17031
rect 9692 16590 9720 17138
rect 9876 17134 9904 17462
rect 9968 17338 9996 19382
rect 10060 18426 10088 19858
rect 10336 19360 10364 22200
rect 10796 20516 10824 22200
rect 11256 20874 11284 22200
rect 11244 20868 11296 20874
rect 11244 20810 11296 20816
rect 11716 20806 11744 22200
rect 11704 20800 11756 20806
rect 11704 20742 11756 20748
rect 11346 20700 11654 20720
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20624 11654 20644
rect 10796 20488 11008 20516
rect 10784 19848 10836 19854
rect 10784 19790 10836 19796
rect 10796 19378 10824 19790
rect 10508 19372 10560 19378
rect 10336 19332 10456 19360
rect 10428 19174 10456 19332
rect 10508 19314 10560 19320
rect 10784 19372 10836 19378
rect 10784 19314 10836 19320
rect 10416 19168 10468 19174
rect 10416 19110 10468 19116
rect 10520 18970 10548 19314
rect 10876 19168 10928 19174
rect 10876 19110 10928 19116
rect 10232 18964 10284 18970
rect 10232 18906 10284 18912
rect 10508 18964 10560 18970
rect 10508 18906 10560 18912
rect 10048 18420 10100 18426
rect 10048 18362 10100 18368
rect 9956 17332 10008 17338
rect 10060 17320 10088 18362
rect 10060 17292 10180 17320
rect 9956 17274 10008 17280
rect 10152 17241 10180 17292
rect 10138 17232 10194 17241
rect 10048 17196 10100 17202
rect 10138 17167 10194 17176
rect 10048 17138 10100 17144
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9876 16454 9904 17070
rect 9956 16992 10008 16998
rect 9956 16934 10008 16940
rect 9864 16448 9916 16454
rect 9864 16390 9916 16396
rect 9588 15904 9640 15910
rect 9588 15846 9640 15852
rect 9772 15428 9824 15434
rect 9772 15370 9824 15376
rect 9680 15360 9732 15366
rect 9680 15302 9732 15308
rect 9692 15094 9720 15302
rect 9680 15088 9732 15094
rect 9680 15030 9732 15036
rect 9784 13190 9812 15370
rect 9968 13841 9996 16934
rect 10060 15094 10088 17138
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 9954 13832 10010 13841
rect 9954 13767 10010 13776
rect 10060 13530 10088 13874
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9772 12844 9824 12850
rect 9772 12786 9824 12792
rect 9494 12744 9550 12753
rect 9494 12679 9550 12688
rect 9324 11354 9444 11370
rect 9324 11348 9456 11354
rect 9324 11342 9404 11348
rect 9128 11144 9180 11150
rect 9128 11086 9180 11092
rect 8747 10364 9055 10384
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10288 9055 10308
rect 9140 10266 9168 11086
rect 9128 10260 9180 10266
rect 9128 10202 9180 10208
rect 9324 10062 9352 11342
rect 9404 11290 9456 11296
rect 9404 11212 9456 11218
rect 9404 11154 9456 11160
rect 9416 10470 9444 11154
rect 9508 11082 9536 12679
rect 9588 12640 9640 12646
rect 9588 12582 9640 12588
rect 9600 11082 9628 12582
rect 9784 12102 9812 12786
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9772 12096 9824 12102
rect 9772 12038 9824 12044
rect 9968 11898 9996 12718
rect 10152 12434 10180 15846
rect 10244 14006 10272 18906
rect 10416 18284 10468 18290
rect 10416 18226 10468 18232
rect 10324 17876 10376 17882
rect 10324 17818 10376 17824
rect 10336 16454 10364 17818
rect 10324 16448 10376 16454
rect 10324 16390 10376 16396
rect 10428 16046 10456 18226
rect 10508 17536 10560 17542
rect 10508 17478 10560 17484
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10336 15162 10364 15982
rect 10428 15706 10456 15982
rect 10416 15700 10468 15706
rect 10416 15642 10468 15648
rect 10416 15564 10468 15570
rect 10416 15506 10468 15512
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10232 14000 10284 14006
rect 10232 13942 10284 13948
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12986 10364 13262
rect 10324 12980 10376 12986
rect 10324 12922 10376 12928
rect 10060 12406 10180 12434
rect 9956 11892 10008 11898
rect 9956 11834 10008 11840
rect 10060 11830 10088 12406
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9864 11688 9916 11694
rect 9864 11630 9916 11636
rect 9496 11076 9548 11082
rect 9496 11018 9548 11024
rect 9588 11076 9640 11082
rect 9588 11018 9640 11024
rect 9770 10976 9826 10985
rect 9770 10911 9826 10920
rect 9404 10464 9456 10470
rect 9404 10406 9456 10412
rect 9312 10056 9364 10062
rect 9312 9998 9364 10004
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8668 9716 8720 9722
rect 8668 9658 8720 9664
rect 8668 9580 8720 9586
rect 8668 9522 8720 9528
rect 9220 9580 9272 9586
rect 9220 9522 9272 9528
rect 8680 8634 8708 9522
rect 8747 9276 9055 9296
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9200 9055 9220
rect 9232 9194 9260 9522
rect 9140 9166 9260 9194
rect 9324 9178 9352 9862
rect 9416 9654 9444 10406
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9312 9172 9364 9178
rect 9140 9042 9168 9166
rect 9312 9114 9364 9120
rect 9310 9072 9366 9081
rect 9128 9036 9180 9042
rect 9310 9007 9366 9016
rect 9128 8978 9180 8984
rect 9324 8838 9352 9007
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 9312 8832 9364 8838
rect 9312 8774 9364 8780
rect 8668 8628 8720 8634
rect 8668 8570 8720 8576
rect 8772 8566 8800 8774
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 9416 8430 9444 9590
rect 9508 9364 9536 10066
rect 9680 9920 9732 9926
rect 9680 9862 9732 9868
rect 9588 9648 9640 9654
rect 9586 9616 9588 9625
rect 9640 9616 9642 9625
rect 9586 9551 9642 9560
rect 9588 9376 9640 9382
rect 9508 9336 9588 9364
rect 9508 9110 9536 9336
rect 9588 9318 9640 9324
rect 9692 9178 9720 9862
rect 9784 9178 9812 10911
rect 9680 9172 9732 9178
rect 9680 9114 9732 9120
rect 9772 9172 9824 9178
rect 9772 9114 9824 9120
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9508 8566 9536 9046
rect 9496 8560 9548 8566
rect 9496 8502 9548 8508
rect 9404 8424 9456 8430
rect 9404 8366 9456 8372
rect 8747 8188 9055 8208
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8112 9055 8132
rect 9312 7948 9364 7954
rect 9312 7890 9364 7896
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8576 7336 8628 7342
rect 8576 7278 8628 7284
rect 8300 6452 8352 6458
rect 8300 6394 8352 6400
rect 8312 5953 8340 6394
rect 8588 6186 8616 7278
rect 8680 6662 8708 7686
rect 9324 7478 9352 7890
rect 9416 7886 9444 8366
rect 9404 7880 9456 7886
rect 9404 7822 9456 7828
rect 9588 7540 9640 7546
rect 9588 7482 9640 7488
rect 9312 7472 9364 7478
rect 9312 7414 9364 7420
rect 8747 7100 9055 7120
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7024 9055 7044
rect 9600 6934 9628 7482
rect 9876 7313 9904 11630
rect 10428 10810 10456 15506
rect 10520 14074 10548 17478
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16522 10732 16934
rect 10692 16516 10744 16522
rect 10692 16458 10744 16464
rect 10784 16516 10836 16522
rect 10784 16458 10836 16464
rect 10796 16250 10824 16458
rect 10784 16244 10836 16250
rect 10784 16186 10836 16192
rect 10784 15700 10836 15706
rect 10784 15642 10836 15648
rect 10796 15502 10824 15642
rect 10888 15502 10916 19110
rect 10980 18970 11008 20488
rect 11060 20460 11112 20466
rect 11060 20402 11112 20408
rect 11072 20262 11100 20402
rect 12176 20369 12204 22200
rect 12636 20534 12664 22200
rect 12808 20800 12860 20806
rect 12808 20742 12860 20748
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12716 20460 12768 20466
rect 12716 20402 12768 20408
rect 12162 20360 12218 20369
rect 12162 20295 12218 20304
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 12256 20256 12308 20262
rect 12256 20198 12308 20204
rect 10968 18964 11020 18970
rect 10968 18906 11020 18912
rect 11072 18902 11100 20198
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11346 19612 11654 19632
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19536 11654 19556
rect 11152 19372 11204 19378
rect 11152 19314 11204 19320
rect 11060 18896 11112 18902
rect 11060 18838 11112 18844
rect 11060 18692 11112 18698
rect 11060 18634 11112 18640
rect 10968 18080 11020 18086
rect 10968 18022 11020 18028
rect 10980 16590 11008 18022
rect 10968 16584 11020 16590
rect 10968 16526 11020 16532
rect 11072 16250 11100 18634
rect 11164 17678 11192 19314
rect 11244 18760 11296 18766
rect 11244 18702 11296 18708
rect 11256 17882 11284 18702
rect 11704 18624 11756 18630
rect 11704 18566 11756 18572
rect 11346 18524 11654 18544
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18448 11654 18468
rect 11244 17876 11296 17882
rect 11244 17818 11296 17824
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11150 17368 11206 17377
rect 11150 17303 11206 17312
rect 11164 16658 11192 17303
rect 11256 17134 11284 17818
rect 11346 17436 11654 17456
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11346 17360 11654 17380
rect 11244 17128 11296 17134
rect 11244 17070 11296 17076
rect 11152 16652 11204 16658
rect 11152 16594 11204 16600
rect 11244 16448 11296 16454
rect 11244 16390 11296 16396
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11152 15904 11204 15910
rect 11152 15846 11204 15852
rect 11164 15570 11192 15846
rect 11152 15564 11204 15570
rect 11152 15506 11204 15512
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 11060 15360 11112 15366
rect 11060 15302 11112 15308
rect 11072 15162 11100 15302
rect 11060 15156 11112 15162
rect 11060 15098 11112 15104
rect 10600 14952 10652 14958
rect 10600 14894 10652 14900
rect 11164 14906 11192 15506
rect 11256 15094 11284 16390
rect 11346 16348 11654 16368
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16272 11654 16292
rect 11346 15260 11654 15280
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15184 11654 15204
rect 11716 15094 11744 18566
rect 11808 18358 11836 19926
rect 11888 19848 11940 19854
rect 11888 19790 11940 19796
rect 11900 19514 11928 19790
rect 12176 19786 12204 20198
rect 12268 19825 12296 20198
rect 12728 19961 12756 20402
rect 12714 19952 12770 19961
rect 12714 19887 12770 19896
rect 12254 19816 12310 19825
rect 12164 19780 12216 19786
rect 12254 19751 12310 19760
rect 12164 19722 12216 19728
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 12348 19440 12400 19446
rect 12348 19382 12400 19388
rect 12072 18624 12124 18630
rect 12072 18566 12124 18572
rect 12164 18624 12216 18630
rect 12164 18566 12216 18572
rect 11796 18352 11848 18358
rect 11796 18294 11848 18300
rect 11978 17640 12034 17649
rect 11978 17575 12034 17584
rect 11796 17196 11848 17202
rect 11796 17138 11848 17144
rect 11244 15088 11296 15094
rect 11244 15030 11296 15036
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 10612 14618 10640 14894
rect 11164 14878 11284 14906
rect 10600 14612 10652 14618
rect 10600 14554 10652 14560
rect 11256 14346 11284 14878
rect 11808 14396 11836 17138
rect 11888 16652 11940 16658
rect 11888 16594 11940 16600
rect 11900 15570 11928 16594
rect 11888 15564 11940 15570
rect 11888 15506 11940 15512
rect 11992 15366 12020 17575
rect 12084 17338 12112 18566
rect 12176 17610 12204 18566
rect 12254 18456 12310 18465
rect 12254 18391 12310 18400
rect 12268 18358 12296 18391
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12072 17332 12124 17338
rect 12072 17274 12124 17280
rect 12256 17128 12308 17134
rect 12256 17070 12308 17076
rect 11980 15360 12032 15366
rect 11980 15302 12032 15308
rect 11888 15156 11940 15162
rect 11888 15098 11940 15104
rect 11716 14368 11836 14396
rect 11152 14340 11204 14346
rect 11152 14282 11204 14288
rect 11244 14340 11296 14346
rect 11244 14282 11296 14288
rect 10508 14068 10560 14074
rect 10508 14010 10560 14016
rect 11164 13938 11192 14282
rect 11346 14172 11654 14192
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14096 11654 14116
rect 11152 13932 11204 13938
rect 11152 13874 11204 13880
rect 11060 13864 11112 13870
rect 11060 13806 11112 13812
rect 11072 12238 11100 13806
rect 11164 13530 11192 13874
rect 11152 13524 11204 13530
rect 11152 13466 11204 13472
rect 11244 13252 11296 13258
rect 11244 13194 11296 13200
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10876 12164 10928 12170
rect 10876 12106 10928 12112
rect 10508 12096 10560 12102
rect 10508 12038 10560 12044
rect 10520 11694 10548 12038
rect 10888 11762 10916 12106
rect 10876 11756 10928 11762
rect 10876 11698 10928 11704
rect 10508 11688 10560 11694
rect 10508 11630 10560 11636
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 11256 10742 11284 13194
rect 11346 13084 11654 13104
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13008 11654 13028
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11532 12238 11560 12718
rect 11520 12232 11572 12238
rect 11716 12209 11744 14368
rect 11796 14272 11848 14278
rect 11796 14214 11848 14220
rect 11808 12918 11836 14214
rect 11900 14074 11928 15098
rect 11992 14770 12020 15302
rect 11992 14742 12204 14770
rect 12072 14612 12124 14618
rect 12072 14554 12124 14560
rect 11888 14068 11940 14074
rect 11888 14010 11940 14016
rect 11980 14068 12032 14074
rect 11980 14010 12032 14016
rect 11796 12912 11848 12918
rect 11796 12854 11848 12860
rect 11888 12232 11940 12238
rect 11520 12174 11572 12180
rect 11702 12200 11758 12209
rect 11888 12174 11940 12180
rect 11702 12135 11758 12144
rect 11346 11996 11654 12016
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11920 11654 11940
rect 11900 11830 11928 12174
rect 11888 11824 11940 11830
rect 11888 11766 11940 11772
rect 11900 11150 11928 11766
rect 11992 11558 12020 14010
rect 12084 13870 12112 14554
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12176 12986 12204 14742
rect 12268 13190 12296 17070
rect 12360 14958 12388 19382
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12452 18834 12480 19314
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12452 18086 12480 18770
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 12532 18624 12584 18630
rect 12532 18566 12584 18572
rect 12440 18080 12492 18086
rect 12440 18022 12492 18028
rect 12544 16590 12572 18566
rect 12636 17882 12664 18702
rect 12728 18358 12756 19887
rect 12820 19242 12848 20742
rect 13096 20602 13124 22200
rect 13556 20602 13584 22200
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 13084 20596 13136 20602
rect 13084 20538 13136 20544
rect 13544 20596 13596 20602
rect 13544 20538 13596 20544
rect 13004 19378 13032 20538
rect 13452 20460 13504 20466
rect 13452 20402 13504 20408
rect 13464 20058 13492 20402
rect 13818 20360 13874 20369
rect 13636 20324 13688 20330
rect 14016 20330 14044 22200
rect 14476 20602 14504 22200
rect 14464 20596 14516 20602
rect 14464 20538 14516 20544
rect 14936 20330 14964 22200
rect 13818 20295 13874 20304
rect 14004 20324 14056 20330
rect 13636 20266 13688 20272
rect 13452 20052 13504 20058
rect 13452 19994 13504 20000
rect 13176 19848 13228 19854
rect 13648 19825 13676 20266
rect 13176 19790 13228 19796
rect 13634 19816 13690 19825
rect 12992 19372 13044 19378
rect 12992 19314 13044 19320
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 12808 19236 12860 19242
rect 12808 19178 12860 19184
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12716 18352 12768 18358
rect 12716 18294 12768 18300
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12636 17626 12664 17818
rect 12636 17598 12756 17626
rect 12624 17536 12676 17542
rect 12624 17478 12676 17484
rect 12532 16584 12584 16590
rect 12532 16526 12584 16532
rect 12636 16522 12664 17478
rect 12728 16726 12756 17598
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12452 15434 12480 16118
rect 12820 16114 12848 18566
rect 12912 17105 12940 19246
rect 13084 18080 13136 18086
rect 13084 18022 13136 18028
rect 13096 17746 13124 18022
rect 13084 17740 13136 17746
rect 13084 17682 13136 17688
rect 13084 17536 13136 17542
rect 13084 17478 13136 17484
rect 13096 17338 13124 17478
rect 13084 17332 13136 17338
rect 13084 17274 13136 17280
rect 12898 17096 12954 17105
rect 12898 17031 12954 17040
rect 13084 17060 13136 17066
rect 13084 17002 13136 17008
rect 13096 16266 13124 17002
rect 12912 16238 13124 16266
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12544 15502 12572 15642
rect 12532 15496 12584 15502
rect 12532 15438 12584 15444
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12348 14952 12400 14958
rect 12348 14894 12400 14900
rect 12452 14618 12480 15370
rect 12912 15162 12940 16238
rect 12992 16108 13044 16114
rect 12992 16050 13044 16056
rect 12900 15156 12952 15162
rect 12900 15098 12952 15104
rect 13004 15094 13032 16050
rect 12992 15088 13044 15094
rect 12992 15030 13044 15036
rect 12900 14884 12952 14890
rect 12900 14826 12952 14832
rect 12440 14612 12492 14618
rect 12492 14572 12572 14600
rect 12440 14554 12492 14560
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12348 13864 12400 13870
rect 12348 13806 12400 13812
rect 12360 13326 12388 13806
rect 12452 13394 12480 13874
rect 12440 13388 12492 13394
rect 12440 13330 12492 13336
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12256 13184 12308 13190
rect 12256 13126 12308 13132
rect 12164 12980 12216 12986
rect 12164 12922 12216 12928
rect 12176 12646 12204 12922
rect 12164 12640 12216 12646
rect 12164 12582 12216 12588
rect 12268 11898 12296 13126
rect 12360 12238 12388 13262
rect 12544 13258 12572 14572
rect 12532 13252 12584 13258
rect 12532 13194 12584 13200
rect 12912 12986 12940 14826
rect 13004 14414 13032 15030
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14006 13032 14350
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 13096 13852 13124 14010
rect 13004 13824 13124 13852
rect 12900 12980 12952 12986
rect 12900 12922 12952 12928
rect 13004 12238 13032 13824
rect 13188 12434 13216 19790
rect 13452 19780 13504 19786
rect 13634 19751 13690 19760
rect 13452 19722 13504 19728
rect 13268 18284 13320 18290
rect 13268 18226 13320 18232
rect 13280 16794 13308 18226
rect 13360 18080 13412 18086
rect 13360 18022 13412 18028
rect 13372 17678 13400 18022
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13358 17232 13414 17241
rect 13358 17167 13360 17176
rect 13412 17167 13414 17176
rect 13360 17138 13412 17144
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13280 16130 13308 16730
rect 13372 16658 13400 17138
rect 13360 16652 13412 16658
rect 13360 16594 13412 16600
rect 13360 16448 13412 16454
rect 13360 16390 13412 16396
rect 13372 16250 13400 16390
rect 13360 16244 13412 16250
rect 13360 16186 13412 16192
rect 13280 16114 13400 16130
rect 13280 16108 13412 16114
rect 13280 16102 13360 16108
rect 13360 16050 13412 16056
rect 13360 15972 13412 15978
rect 13360 15914 13412 15920
rect 13372 15502 13400 15914
rect 13360 15496 13412 15502
rect 13360 15438 13412 15444
rect 13268 15360 13320 15366
rect 13268 15302 13320 15308
rect 13280 15162 13308 15302
rect 13268 15156 13320 15162
rect 13268 15098 13320 15104
rect 13464 15042 13492 19722
rect 13544 18352 13596 18358
rect 13544 18294 13596 18300
rect 13556 17134 13584 18294
rect 13648 18290 13676 19751
rect 13728 19372 13780 19378
rect 13728 19314 13780 19320
rect 13636 18284 13688 18290
rect 13636 18226 13688 18232
rect 13636 17604 13688 17610
rect 13636 17546 13688 17552
rect 13648 17202 13676 17546
rect 13636 17196 13688 17202
rect 13636 17138 13688 17144
rect 13544 17128 13596 17134
rect 13544 17070 13596 17076
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13556 15162 13584 16594
rect 13648 15910 13676 17138
rect 13740 16522 13768 19314
rect 13832 19281 13860 20295
rect 14004 20266 14056 20272
rect 14924 20324 14976 20330
rect 14924 20266 14976 20272
rect 13945 20156 14253 20176
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20080 14253 20100
rect 15396 20058 15424 22200
rect 15856 20602 15884 22200
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 15844 20596 15896 20602
rect 15844 20538 15896 20544
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 15476 20460 15528 20466
rect 15476 20402 15528 20408
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 13912 19916 13964 19922
rect 13912 19858 13964 19864
rect 13924 19514 13952 19858
rect 14556 19848 14608 19854
rect 14556 19790 14608 19796
rect 14280 19712 14332 19718
rect 14280 19654 14332 19660
rect 13912 19508 13964 19514
rect 13912 19450 13964 19456
rect 13818 19272 13874 19281
rect 13818 19207 13874 19216
rect 14292 19174 14320 19654
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14280 19168 14332 19174
rect 14476 19145 14504 19178
rect 14280 19110 14332 19116
rect 14462 19136 14518 19145
rect 13945 19068 14253 19088
rect 14462 19071 14518 19080
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 18992 14253 19012
rect 13820 18896 13872 18902
rect 13818 18864 13820 18873
rect 13872 18864 13874 18873
rect 13818 18799 13874 18808
rect 13832 18290 13860 18799
rect 14004 18624 14056 18630
rect 14004 18566 14056 18572
rect 14016 18358 14044 18566
rect 14094 18456 14150 18465
rect 14094 18391 14150 18400
rect 14004 18352 14056 18358
rect 14004 18294 14056 18300
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13832 16266 13860 18226
rect 14016 18222 14044 18294
rect 14108 18290 14136 18391
rect 14464 18352 14516 18358
rect 14464 18294 14516 18300
rect 14096 18284 14148 18290
rect 14096 18226 14148 18232
rect 14004 18216 14056 18222
rect 14004 18158 14056 18164
rect 14372 18080 14424 18086
rect 14372 18022 14424 18028
rect 13945 17980 14253 18000
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17904 14253 17924
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 13945 16892 14253 16912
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16816 14253 16836
rect 14292 16726 14320 17070
rect 14384 16998 14412 18022
rect 14476 17678 14504 18294
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14462 17504 14518 17513
rect 14462 17439 14518 17448
rect 14372 16992 14424 16998
rect 14372 16934 14424 16940
rect 14004 16720 14056 16726
rect 14004 16662 14056 16668
rect 14280 16720 14332 16726
rect 14280 16662 14332 16668
rect 14016 16454 14044 16662
rect 14004 16448 14056 16454
rect 14004 16390 14056 16396
rect 13728 16244 13780 16250
rect 13832 16238 13952 16266
rect 13728 16186 13780 16192
rect 13636 15904 13688 15910
rect 13636 15846 13688 15852
rect 13544 15156 13596 15162
rect 13544 15098 13596 15104
rect 13372 15026 13492 15042
rect 13648 15026 13676 15846
rect 13740 15706 13768 16186
rect 13820 16108 13872 16114
rect 13820 16050 13872 16056
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13360 15020 13492 15026
rect 13412 15014 13492 15020
rect 13636 15020 13688 15026
rect 13360 14962 13412 14968
rect 13636 14962 13688 14968
rect 13648 14074 13676 14962
rect 13728 14952 13780 14958
rect 13728 14894 13780 14900
rect 13740 14498 13768 14894
rect 13832 14618 13860 16050
rect 13924 16046 13952 16238
rect 13912 16040 13964 16046
rect 13912 15982 13964 15988
rect 14280 16040 14332 16046
rect 14280 15982 14332 15988
rect 13945 15804 14253 15824
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15728 14253 15748
rect 13945 14716 14253 14736
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14640 14253 14660
rect 13820 14612 13872 14618
rect 13820 14554 13872 14560
rect 13740 14470 13860 14498
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 13832 13938 13860 14470
rect 13820 13932 13872 13938
rect 13820 13874 13872 13880
rect 13832 13394 13860 13874
rect 13945 13628 14253 13648
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13552 14253 13572
rect 13820 13388 13872 13394
rect 13820 13330 13872 13336
rect 13358 13288 13414 13297
rect 13358 13223 13360 13232
rect 13412 13223 13414 13232
rect 13360 13194 13412 13200
rect 14292 12986 14320 15982
rect 14372 15360 14424 15366
rect 14372 15302 14424 15308
rect 14384 15094 14412 15302
rect 14372 15088 14424 15094
rect 14372 15030 14424 15036
rect 14280 12980 14332 12986
rect 14280 12922 14332 12928
rect 14292 12646 14320 12922
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 14280 12640 14332 12646
rect 14280 12582 14332 12588
rect 13096 12406 13216 12434
rect 12348 12232 12400 12238
rect 12348 12174 12400 12180
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 12256 11892 12308 11898
rect 12256 11834 12308 11840
rect 13004 11762 13032 12174
rect 12624 11756 12676 11762
rect 12624 11698 12676 11704
rect 12992 11756 13044 11762
rect 12992 11698 13044 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 11888 11144 11940 11150
rect 11888 11086 11940 11092
rect 11704 11008 11756 11014
rect 11704 10950 11756 10956
rect 11346 10908 11654 10928
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10832 11654 10852
rect 11244 10736 11296 10742
rect 11244 10678 11296 10684
rect 11256 10062 11284 10678
rect 11716 10606 11744 10950
rect 11704 10600 11756 10606
rect 11704 10542 11756 10548
rect 11900 10470 11928 11086
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11796 10464 11848 10470
rect 11796 10406 11848 10412
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11244 10056 11296 10062
rect 11244 9998 11296 10004
rect 11346 9820 11654 9840
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9744 11654 9764
rect 11808 9654 11836 10406
rect 11900 10266 11928 10406
rect 11888 10260 11940 10266
rect 11888 10202 11940 10208
rect 12084 10198 12112 10746
rect 12636 10742 12664 11698
rect 12808 11552 12860 11558
rect 12808 11494 12860 11500
rect 12820 10742 12848 11494
rect 12624 10736 12676 10742
rect 12624 10678 12676 10684
rect 12808 10736 12860 10742
rect 12808 10678 12860 10684
rect 12256 10464 12308 10470
rect 12256 10406 12308 10412
rect 12268 10198 12296 10406
rect 13096 10266 13124 12406
rect 13832 12170 13860 12582
rect 13945 12540 14253 12560
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12464 14253 12484
rect 13820 12164 13872 12170
rect 13820 12106 13872 12112
rect 13176 12096 13228 12102
rect 13176 12038 13228 12044
rect 13636 12096 13688 12102
rect 13636 12038 13688 12044
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 12256 10192 12308 10198
rect 12256 10134 12308 10140
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12636 9722 12664 10066
rect 13188 10062 13216 12038
rect 13452 11756 13504 11762
rect 13452 11698 13504 11704
rect 13464 11218 13492 11698
rect 13648 11354 13676 12038
rect 13740 11898 13768 12038
rect 13728 11892 13780 11898
rect 13728 11834 13780 11840
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 13945 11452 14253 11472
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11376 14253 11396
rect 13636 11348 13688 11354
rect 13636 11290 13688 11296
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 13832 9654 13860 11086
rect 13945 10364 14253 10384
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10288 14253 10308
rect 14292 9654 14320 11698
rect 14476 11558 14504 17439
rect 14568 16250 14596 19790
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14752 18426 14780 19246
rect 14740 18420 14792 18426
rect 14740 18362 14792 18368
rect 14844 17882 14872 19314
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15108 18760 15160 18766
rect 15108 18702 15160 18708
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14740 17808 14792 17814
rect 14792 17756 14872 17762
rect 14740 17750 14872 17756
rect 14752 17734 14872 17750
rect 15120 17746 15148 18702
rect 14844 17626 14872 17734
rect 15108 17740 15160 17746
rect 15108 17682 15160 17688
rect 14648 17604 14700 17610
rect 14844 17598 15148 17626
rect 14648 17546 14700 17552
rect 14660 17338 14688 17546
rect 15120 17542 15148 17598
rect 15016 17536 15068 17542
rect 15016 17478 15068 17484
rect 15108 17536 15160 17542
rect 15212 17513 15240 19246
rect 15292 19236 15344 19242
rect 15292 19178 15344 19184
rect 15304 18426 15332 19178
rect 15488 18970 15516 20402
rect 15948 19854 15976 20470
rect 15936 19848 15988 19854
rect 15936 19790 15988 19796
rect 16028 19712 16080 19718
rect 16028 19654 16080 19660
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15764 19417 15792 19450
rect 16040 19417 16068 19654
rect 15750 19408 15806 19417
rect 15750 19343 15806 19352
rect 16026 19408 16082 19417
rect 16132 19378 16160 20810
rect 16316 20330 16344 22200
rect 16776 21026 16804 22200
rect 16776 20998 16988 21026
rect 16544 20700 16852 20720
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20624 16852 20644
rect 16304 20324 16356 20330
rect 16304 20266 16356 20272
rect 16960 20058 16988 20998
rect 17236 20602 17264 22200
rect 17224 20596 17276 20602
rect 17224 20538 17276 20544
rect 17592 20528 17644 20534
rect 17592 20470 17644 20476
rect 17224 20392 17276 20398
rect 17224 20334 17276 20340
rect 17236 20058 17264 20334
rect 16948 20052 17000 20058
rect 16948 19994 17000 20000
rect 17224 20052 17276 20058
rect 17224 19994 17276 20000
rect 16396 19848 16448 19854
rect 16488 19848 16540 19854
rect 16396 19790 16448 19796
rect 16486 19816 16488 19825
rect 17132 19848 17184 19854
rect 16540 19816 16542 19825
rect 16026 19343 16082 19352
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 15844 19168 15896 19174
rect 15844 19110 15896 19116
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15396 18850 15424 18906
rect 15752 18896 15804 18902
rect 15396 18844 15752 18850
rect 15396 18838 15804 18844
rect 15396 18822 15792 18838
rect 15856 18766 15884 19110
rect 15844 18760 15896 18766
rect 15844 18702 15896 18708
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15752 18284 15804 18290
rect 15752 18226 15804 18232
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15108 17478 15160 17484
rect 15198 17504 15254 17513
rect 14648 17332 14700 17338
rect 14648 17274 14700 17280
rect 15028 16697 15056 17478
rect 15198 17439 15254 17448
rect 15200 17332 15252 17338
rect 15200 17274 15252 17280
rect 15014 16688 15070 16697
rect 15014 16623 15070 16632
rect 14556 16244 14608 16250
rect 14556 16186 14608 16192
rect 14740 16040 14792 16046
rect 14740 15982 14792 15988
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14660 14482 14688 15506
rect 14752 15026 14780 15982
rect 14740 15020 14792 15026
rect 14740 14962 14792 14968
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14556 14272 14608 14278
rect 14556 14214 14608 14220
rect 14568 13530 14596 14214
rect 14660 14074 14688 14418
rect 14648 14068 14700 14074
rect 14648 14010 14700 14016
rect 14556 13524 14608 13530
rect 14556 13466 14608 13472
rect 14464 11552 14516 11558
rect 14464 11494 14516 11500
rect 14740 11552 14792 11558
rect 14740 11494 14792 11500
rect 14464 11144 14516 11150
rect 14464 11086 14516 11092
rect 11796 9648 11848 9654
rect 11796 9590 11848 9596
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 10968 9376 11020 9382
rect 10968 9318 11020 9324
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10980 8906 11008 9318
rect 10968 8900 11020 8906
rect 10968 8842 11020 8848
rect 10232 8492 10284 8498
rect 10232 8434 10284 8440
rect 10244 8090 10272 8434
rect 10322 8392 10378 8401
rect 10322 8327 10378 8336
rect 10232 8084 10284 8090
rect 10232 8026 10284 8032
rect 10336 7750 10364 8327
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7546 10364 7686
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9862 7304 9918 7313
rect 9862 7239 9918 7248
rect 9588 6928 9640 6934
rect 9588 6870 9640 6876
rect 8668 6656 8720 6662
rect 8668 6598 8720 6604
rect 8576 6180 8628 6186
rect 8576 6122 8628 6128
rect 8747 6012 9055 6032
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8298 5944 8354 5953
rect 8747 5936 9055 5956
rect 8298 5879 8354 5888
rect 7562 5672 7618 5681
rect 7562 5607 7618 5616
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 8312 4593 8340 5510
rect 8747 4924 9055 4944
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4848 9055 4868
rect 11072 4729 11100 9318
rect 13945 9276 14253 9296
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9200 14253 9220
rect 11346 8732 11654 8752
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8656 11654 8676
rect 13945 8188 14253 8208
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8112 14253 8132
rect 14476 7857 14504 11086
rect 14752 10062 14780 11494
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 14832 11008 14884 11014
rect 14832 10950 14884 10956
rect 14844 10810 14872 10950
rect 14936 10810 14964 11018
rect 14832 10804 14884 10810
rect 14832 10746 14884 10752
rect 14924 10804 14976 10810
rect 14924 10746 14976 10752
rect 14924 10600 14976 10606
rect 14924 10542 14976 10548
rect 14936 10470 14964 10542
rect 14924 10464 14976 10470
rect 14924 10406 14976 10412
rect 14740 10056 14792 10062
rect 14740 9998 14792 10004
rect 14936 9586 14964 10406
rect 14924 9580 14976 9586
rect 14924 9522 14976 9528
rect 15028 8945 15056 16623
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15120 15162 15148 15302
rect 15108 15156 15160 15162
rect 15108 15098 15160 15104
rect 15120 11354 15148 15098
rect 15212 14414 15240 17274
rect 15290 17232 15346 17241
rect 15290 17167 15292 17176
rect 15344 17167 15346 17176
rect 15292 17138 15344 17144
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 15304 14362 15332 17138
rect 15396 17066 15424 18158
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15384 17060 15436 17066
rect 15384 17002 15436 17008
rect 15488 16182 15516 17138
rect 15568 17128 15620 17134
rect 15568 17070 15620 17076
rect 15580 16561 15608 17070
rect 15764 16794 15792 18226
rect 16132 17954 16160 19314
rect 16304 18760 16356 18766
rect 16304 18702 16356 18708
rect 16316 18426 16344 18702
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16408 18358 16436 19790
rect 16486 19751 16542 19760
rect 17038 19816 17094 19825
rect 17132 19790 17184 19796
rect 17038 19751 17094 19760
rect 16544 19612 16852 19632
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19536 16852 19556
rect 16948 19508 17000 19514
rect 16948 19450 17000 19456
rect 16960 19417 16988 19450
rect 16946 19408 17002 19417
rect 16856 19372 16908 19378
rect 16946 19343 17002 19352
rect 16856 19314 16908 19320
rect 16868 19281 16896 19314
rect 16854 19272 16910 19281
rect 16854 19207 16910 19216
rect 16544 18524 16852 18544
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18448 16852 18468
rect 16396 18352 16448 18358
rect 16396 18294 16448 18300
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16040 17926 16160 17954
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15856 17066 15884 17614
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15752 16788 15804 16794
rect 15752 16730 15804 16736
rect 15566 16552 15622 16561
rect 15566 16487 15622 16496
rect 15476 16176 15528 16182
rect 15476 16118 15528 16124
rect 15488 15162 15516 16118
rect 15580 15638 15608 16487
rect 15856 16250 15884 17002
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 15568 15632 15620 15638
rect 15568 15574 15620 15580
rect 15476 15156 15528 15162
rect 15476 15098 15528 15104
rect 15304 14334 15516 14362
rect 15488 12918 15516 14334
rect 15476 12912 15528 12918
rect 15476 12854 15528 12860
rect 15292 12776 15344 12782
rect 15292 12718 15344 12724
rect 15304 11898 15332 12718
rect 15384 12708 15436 12714
rect 15384 12650 15436 12656
rect 15396 12442 15424 12650
rect 15384 12436 15436 12442
rect 15384 12378 15436 12384
rect 15384 12164 15436 12170
rect 15384 12106 15436 12112
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15108 11348 15160 11354
rect 15108 11290 15160 11296
rect 15396 10266 15424 12106
rect 15488 11898 15516 12854
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15580 10810 15608 15574
rect 16040 14618 16068 17926
rect 16500 17882 16528 18226
rect 16488 17876 16540 17882
rect 16488 17818 16540 17824
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16544 17436 16852 17456
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17360 16852 17380
rect 16210 17232 16266 17241
rect 16210 17167 16266 17176
rect 16224 17134 16252 17167
rect 16120 17128 16172 17134
rect 16120 17070 16172 17076
rect 16212 17128 16264 17134
rect 16212 17070 16264 17076
rect 16132 16250 16160 17070
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16580 16992 16632 16998
rect 16580 16934 16632 16940
rect 16316 16658 16344 16934
rect 16304 16652 16356 16658
rect 16304 16594 16356 16600
rect 16592 16590 16620 16934
rect 16580 16584 16632 16590
rect 16580 16526 16632 16532
rect 16396 16448 16448 16454
rect 16396 16390 16448 16396
rect 16120 16244 16172 16250
rect 16120 16186 16172 16192
rect 16408 14958 16436 16390
rect 16544 16348 16852 16368
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16272 16852 16292
rect 16960 16250 16988 17614
rect 17052 16794 17080 19751
rect 17144 19718 17172 19790
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17604 19514 17632 20470
rect 17696 20330 17724 22200
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17960 20392 18012 20398
rect 17960 20334 18012 20340
rect 17684 20324 17736 20330
rect 17684 20266 17736 20272
rect 17868 19916 17920 19922
rect 17868 19858 17920 19864
rect 17880 19718 17908 19858
rect 17868 19712 17920 19718
rect 17868 19654 17920 19660
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17592 19508 17644 19514
rect 17592 19450 17644 19456
rect 17132 18692 17184 18698
rect 17132 18634 17184 18640
rect 17144 17270 17172 18634
rect 17132 17264 17184 17270
rect 17132 17206 17184 17212
rect 17040 16788 17092 16794
rect 17040 16730 17092 16736
rect 16948 16244 17000 16250
rect 16948 16186 17000 16192
rect 16948 16040 17000 16046
rect 16948 15982 17000 15988
rect 16544 15260 16852 15280
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15184 16852 15204
rect 16960 15162 16988 15982
rect 17052 15910 17080 16730
rect 17144 16658 17172 17206
rect 17132 16652 17184 16658
rect 17132 16594 17184 16600
rect 17144 16182 17172 16594
rect 17224 16516 17276 16522
rect 17224 16458 17276 16464
rect 17132 16176 17184 16182
rect 17132 16118 17184 16124
rect 17040 15904 17092 15910
rect 17040 15846 17092 15852
rect 17144 15706 17172 16118
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17144 15094 17172 15642
rect 17236 15638 17264 16458
rect 17224 15632 17276 15638
rect 17224 15574 17276 15580
rect 17132 15088 17184 15094
rect 17038 15056 17094 15065
rect 17132 15030 17184 15036
rect 17038 14991 17040 15000
rect 17092 14991 17094 15000
rect 17040 14962 17092 14968
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 16028 14612 16080 14618
rect 16028 14554 16080 14560
rect 17144 14414 17172 15030
rect 17224 14952 17276 14958
rect 17224 14894 17276 14900
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 17132 14272 17184 14278
rect 17236 14260 17264 14894
rect 17184 14232 17264 14260
rect 17132 14214 17184 14220
rect 16544 14172 16852 14192
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14096 16852 14116
rect 17144 13938 17172 14214
rect 16396 13932 16448 13938
rect 16396 13874 16448 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16408 13530 16436 13874
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 17040 13864 17092 13870
rect 17040 13806 17092 13812
rect 16764 13796 16816 13802
rect 16764 13738 16816 13744
rect 16396 13524 16448 13530
rect 16396 13466 16448 13472
rect 16776 13326 16804 13738
rect 16764 13320 16816 13326
rect 16764 13262 16816 13268
rect 15752 13252 15804 13258
rect 15752 13194 15804 13200
rect 15764 12442 15792 13194
rect 16544 13084 16852 13104
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13008 16852 13028
rect 16028 12708 16080 12714
rect 16028 12650 16080 12656
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 16040 12238 16068 12650
rect 16960 12646 16988 13806
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16408 11801 16436 12174
rect 16544 11996 16852 12016
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11920 16852 11940
rect 16394 11792 16450 11801
rect 15752 11756 15804 11762
rect 16394 11727 16450 11736
rect 15752 11698 15804 11704
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15384 10260 15436 10266
rect 15384 10202 15436 10208
rect 15580 9722 15608 10746
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15014 8936 15070 8945
rect 15014 8871 15070 8880
rect 14462 7848 14518 7857
rect 14462 7783 14518 7792
rect 11346 7644 11654 7664
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7568 11654 7588
rect 13945 7100 14253 7120
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7024 14253 7044
rect 11346 6556 11654 6576
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6480 11654 6500
rect 15764 6361 15792 11698
rect 16960 11150 16988 12242
rect 17052 12238 17080 13806
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17328 11778 17356 19450
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17420 19145 17448 19314
rect 17406 19136 17462 19145
rect 17406 19071 17462 19080
rect 17972 18902 18000 20334
rect 18064 18970 18092 20402
rect 18156 20058 18184 22200
rect 18616 20602 18644 22200
rect 19076 20618 19104 22200
rect 19076 20602 19472 20618
rect 18604 20596 18656 20602
rect 19076 20596 19484 20602
rect 19076 20590 19432 20596
rect 18604 20538 18656 20544
rect 19432 20538 19484 20544
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18144 20052 18196 20058
rect 18144 19994 18196 20000
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17960 18896 18012 18902
rect 18156 18873 18184 19654
rect 18524 19514 18552 20198
rect 18512 19508 18564 19514
rect 18512 19450 18564 19456
rect 18328 19440 18380 19446
rect 18328 19382 18380 19388
rect 17960 18838 18012 18844
rect 18142 18864 18198 18873
rect 18142 18799 18198 18808
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17592 18692 17644 18698
rect 17592 18634 17644 18640
rect 17604 18358 17632 18634
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17512 17626 17540 18294
rect 17590 17776 17646 17785
rect 17590 17711 17592 17720
rect 17644 17711 17646 17720
rect 17592 17682 17644 17688
rect 17512 17598 17632 17626
rect 17408 17536 17460 17542
rect 17408 17478 17460 17484
rect 17420 16590 17448 17478
rect 17408 16584 17460 16590
rect 17408 16526 17460 16532
rect 17500 15020 17552 15026
rect 17500 14962 17552 14968
rect 17512 14822 17540 14962
rect 17500 14816 17552 14822
rect 17500 14758 17552 14764
rect 17500 14476 17552 14482
rect 17500 14418 17552 14424
rect 17408 14272 17460 14278
rect 17408 14214 17460 14220
rect 17420 14074 17448 14214
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17512 14006 17540 14418
rect 17604 14074 17632 17598
rect 17696 14260 17724 18702
rect 18340 18408 18368 19382
rect 18420 18692 18472 18698
rect 18420 18634 18472 18640
rect 18512 18692 18564 18698
rect 18512 18634 18564 18640
rect 18156 18380 18368 18408
rect 18052 18148 18104 18154
rect 18052 18090 18104 18096
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17972 17066 18000 17682
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 18064 15586 18092 18090
rect 17972 15558 18092 15586
rect 17972 15026 18000 15558
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17776 14884 17828 14890
rect 17776 14826 17828 14832
rect 17788 14414 17816 14826
rect 18064 14482 18092 15302
rect 18052 14476 18104 14482
rect 18052 14418 18104 14424
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17696 14232 17816 14260
rect 17592 14068 17644 14074
rect 17592 14010 17644 14016
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17592 13728 17644 13734
rect 17592 13670 17644 13676
rect 17604 12850 17632 13670
rect 17684 13184 17736 13190
rect 17684 13126 17736 13132
rect 17592 12844 17644 12850
rect 17592 12786 17644 12792
rect 17604 12374 17632 12786
rect 17696 12442 17724 13126
rect 17684 12436 17736 12442
rect 17684 12378 17736 12384
rect 17592 12368 17644 12374
rect 17592 12310 17644 12316
rect 17236 11750 17356 11778
rect 16948 11144 17000 11150
rect 16948 11086 17000 11092
rect 16544 10908 16852 10928
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10832 16852 10852
rect 16960 10742 16988 11086
rect 16948 10736 17000 10742
rect 16948 10678 17000 10684
rect 15936 10668 15988 10674
rect 15936 10610 15988 10616
rect 15948 9450 15976 10610
rect 16960 10266 16988 10678
rect 16948 10260 17000 10266
rect 16948 10202 17000 10208
rect 16544 9820 16852 9840
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9744 16852 9764
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 17236 9178 17264 11750
rect 17316 11620 17368 11626
rect 17316 11562 17368 11568
rect 17328 10674 17356 11562
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17512 11082 17540 11494
rect 17684 11212 17736 11218
rect 17684 11154 17736 11160
rect 17500 11076 17552 11082
rect 17500 11018 17552 11024
rect 17592 11008 17644 11014
rect 17592 10950 17644 10956
rect 17604 10810 17632 10950
rect 17592 10804 17644 10810
rect 17592 10746 17644 10752
rect 17316 10668 17368 10674
rect 17316 10610 17368 10616
rect 17696 10062 17724 11154
rect 17788 10470 17816 14232
rect 18052 13184 18104 13190
rect 18052 13126 18104 13132
rect 17960 12912 18012 12918
rect 17960 12854 18012 12860
rect 17972 12306 18000 12854
rect 18064 12442 18092 13126
rect 18156 12986 18184 18380
rect 18432 18290 18460 18634
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18420 18284 18472 18290
rect 18420 18226 18472 18232
rect 18340 17746 18368 18226
rect 18328 17740 18380 17746
rect 18328 17682 18380 17688
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18432 16794 18460 17478
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18524 15706 18552 18634
rect 18616 18426 18644 20402
rect 19143 20156 19451 20176
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20080 19451 20100
rect 19536 20058 19564 22200
rect 19524 20052 19576 20058
rect 19524 19994 19576 20000
rect 19616 19984 19668 19990
rect 19338 19952 19394 19961
rect 19616 19926 19668 19932
rect 19338 19887 19394 19896
rect 19352 19854 19380 19887
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 19340 19848 19392 19854
rect 19340 19790 19392 19796
rect 18788 19712 18840 19718
rect 18788 19654 18840 19660
rect 18694 19136 18750 19145
rect 18694 19071 18750 19080
rect 18604 18420 18656 18426
rect 18604 18362 18656 18368
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18616 17202 18644 17478
rect 18604 17196 18656 17202
rect 18604 17138 18656 17144
rect 18512 15700 18564 15706
rect 18512 15642 18564 15648
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18144 12980 18196 12986
rect 18144 12922 18196 12928
rect 18052 12436 18104 12442
rect 18052 12378 18104 12384
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 18248 11354 18276 15438
rect 18708 14482 18736 19071
rect 18800 18086 18828 19654
rect 18880 18760 18932 18766
rect 18880 18702 18932 18708
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18786 16688 18842 16697
rect 18786 16623 18788 16632
rect 18840 16623 18842 16632
rect 18788 16594 18840 16600
rect 18892 14618 18920 18702
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 16182 19012 18022
rect 19076 16182 19104 19790
rect 19432 19780 19484 19786
rect 19432 19722 19484 19728
rect 19444 19378 19472 19722
rect 19524 19440 19576 19446
rect 19524 19382 19576 19388
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19143 19068 19451 19088
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 18992 19451 19012
rect 19143 17980 19451 18000
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17904 19451 17924
rect 19143 16892 19451 16912
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16816 19451 16836
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 19064 16176 19116 16182
rect 19064 16118 19116 16124
rect 19143 15804 19451 15824
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15728 19451 15748
rect 19432 15564 19484 15570
rect 19432 15506 19484 15512
rect 19444 15162 19472 15506
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19444 15026 19472 15098
rect 19432 15020 19484 15026
rect 19432 14962 19484 14968
rect 19064 14816 19116 14822
rect 19064 14758 19116 14764
rect 18880 14612 18932 14618
rect 18880 14554 18932 14560
rect 18696 14476 18748 14482
rect 18696 14418 18748 14424
rect 19076 14006 19104 14758
rect 19143 14716 19451 14736
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14640 19451 14660
rect 19064 14000 19116 14006
rect 19064 13942 19116 13948
rect 19064 13864 19116 13870
rect 19064 13806 19116 13812
rect 18696 13388 18748 13394
rect 18696 13330 18748 13336
rect 18708 12986 18736 13330
rect 18696 12980 18748 12986
rect 18696 12922 18748 12928
rect 19076 12918 19104 13806
rect 19143 13628 19451 13648
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13552 19451 13572
rect 19064 12912 19116 12918
rect 19064 12854 19116 12860
rect 18972 12640 19024 12646
rect 18972 12582 19024 12588
rect 18236 11348 18288 11354
rect 18236 11290 18288 11296
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17776 10464 17828 10470
rect 17776 10406 17828 10412
rect 17972 10266 18000 10610
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17684 10056 17736 10062
rect 17684 9998 17736 10004
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 16544 8732 16852 8752
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8656 16852 8676
rect 18880 8356 18932 8362
rect 18880 8298 18932 8304
rect 18892 8090 18920 8298
rect 18880 8084 18932 8090
rect 18880 8026 18932 8032
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 16544 7644 16852 7664
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16544 7568 16852 7588
rect 17960 7404 18012 7410
rect 17960 7346 18012 7352
rect 16544 6556 16852 6576
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6480 16852 6500
rect 15750 6352 15806 6361
rect 15750 6287 15806 6296
rect 13945 6012 14253 6032
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5936 14253 5956
rect 11346 5468 11654 5488
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5392 11654 5412
rect 16544 5468 16852 5488
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5392 16852 5412
rect 17972 5273 18000 7346
rect 18708 5817 18736 7822
rect 18984 6914 19012 12582
rect 19076 11694 19104 12854
rect 19143 12540 19451 12560
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12464 19451 12484
rect 19064 11688 19116 11694
rect 19064 11630 19116 11636
rect 19143 11452 19451 11472
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11376 19451 11396
rect 19143 10364 19451 10384
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10288 19451 10308
rect 19143 9276 19451 9296
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9200 19451 9220
rect 19143 8188 19451 8208
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 19143 8112 19451 8132
rect 19536 7546 19564 19382
rect 19628 19378 19656 19926
rect 19708 19916 19760 19922
rect 19708 19858 19760 19864
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19720 18154 19748 19858
rect 19996 19514 20024 22200
rect 20168 19848 20220 19854
rect 20168 19790 20220 19796
rect 19892 19508 19944 19514
rect 19892 19450 19944 19456
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19800 18624 19852 18630
rect 19800 18566 19852 18572
rect 19812 18290 19840 18566
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19708 18148 19760 18154
rect 19708 18090 19760 18096
rect 19904 17746 19932 19450
rect 19892 17740 19944 17746
rect 19892 17682 19944 17688
rect 20076 17604 20128 17610
rect 20076 17546 20128 17552
rect 19892 17196 19944 17202
rect 19892 17138 19944 17144
rect 19800 16516 19852 16522
rect 19800 16458 19852 16464
rect 19616 15360 19668 15366
rect 19614 15328 19616 15337
rect 19668 15328 19670 15337
rect 19614 15263 19670 15272
rect 19812 14385 19840 16458
rect 19904 16250 19932 17138
rect 19892 16244 19944 16250
rect 19892 16186 19944 16192
rect 19904 15570 19932 16186
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19892 15564 19944 15570
rect 19892 15506 19944 15512
rect 19798 14376 19854 14385
rect 19798 14311 19854 14320
rect 19996 14074 20024 15846
rect 20088 15706 20116 17546
rect 20076 15700 20128 15706
rect 20076 15642 20128 15648
rect 19984 14068 20036 14074
rect 19984 14010 20036 14016
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19616 13184 19668 13190
rect 19616 13126 19668 13132
rect 19892 13184 19944 13190
rect 19892 13126 19944 13132
rect 19628 12238 19656 13126
rect 19708 12640 19760 12646
rect 19708 12582 19760 12588
rect 19720 12306 19748 12582
rect 19708 12300 19760 12306
rect 19708 12242 19760 12248
rect 19616 12232 19668 12238
rect 19616 12174 19668 12180
rect 19904 11830 19932 13126
rect 19996 12986 20024 13194
rect 19984 12980 20036 12986
rect 19984 12922 20036 12928
rect 19892 11824 19944 11830
rect 19892 11766 19944 11772
rect 20180 8362 20208 19790
rect 20456 19514 20484 22200
rect 20812 20460 20864 20466
rect 20812 20402 20864 20408
rect 20536 20392 20588 20398
rect 20536 20334 20588 20340
rect 20444 19508 20496 19514
rect 20444 19450 20496 19456
rect 20260 18624 20312 18630
rect 20260 18566 20312 18572
rect 20272 16114 20300 18566
rect 20352 18284 20404 18290
rect 20352 18226 20404 18232
rect 20364 17882 20392 18226
rect 20548 17882 20576 20334
rect 20720 19916 20772 19922
rect 20720 19858 20772 19864
rect 20626 19408 20682 19417
rect 20626 19343 20628 19352
rect 20680 19343 20682 19352
rect 20628 19314 20680 19320
rect 20626 18184 20682 18193
rect 20626 18119 20628 18128
rect 20680 18119 20682 18128
rect 20628 18090 20680 18096
rect 20352 17876 20404 17882
rect 20352 17818 20404 17824
rect 20536 17876 20588 17882
rect 20536 17818 20588 17824
rect 20352 17672 20404 17678
rect 20352 17614 20404 17620
rect 20260 16108 20312 16114
rect 20260 16050 20312 16056
rect 20364 13462 20392 17614
rect 20732 17338 20760 19858
rect 20824 18408 20852 20402
rect 20916 18970 20944 22200
rect 21088 20528 21140 20534
rect 21088 20470 21140 20476
rect 20996 20392 21048 20398
rect 20996 20334 21048 20340
rect 20904 18964 20956 18970
rect 20904 18906 20956 18912
rect 20824 18380 20944 18408
rect 20810 18320 20866 18329
rect 20810 18255 20812 18264
rect 20864 18255 20866 18264
rect 20812 18226 20864 18232
rect 20916 17882 20944 18380
rect 20904 17876 20956 17882
rect 20904 17818 20956 17824
rect 20720 17332 20772 17338
rect 20720 17274 20772 17280
rect 20628 17128 20680 17134
rect 21008 17082 21036 20334
rect 20628 17070 20680 17076
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20548 14958 20576 16934
rect 20640 16590 20668 17070
rect 20732 17054 21036 17082
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20640 15094 20668 15914
rect 20628 15088 20680 15094
rect 20628 15030 20680 15036
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20536 14408 20588 14414
rect 20534 14376 20536 14385
rect 20588 14376 20590 14385
rect 20534 14311 20590 14320
rect 20352 13456 20404 13462
rect 20352 13398 20404 13404
rect 20732 12102 20760 17054
rect 20812 16992 20864 16998
rect 20812 16934 20864 16940
rect 20996 16992 21048 16998
rect 20996 16934 21048 16940
rect 20824 13530 20852 16934
rect 21008 16590 21036 16934
rect 20996 16584 21048 16590
rect 20902 16552 20958 16561
rect 20996 16526 21048 16532
rect 20902 16487 20958 16496
rect 20916 16250 20944 16487
rect 21100 16454 21128 20470
rect 21376 19972 21404 22200
rect 21456 20392 21508 20398
rect 21456 20334 21508 20340
rect 21284 19944 21404 19972
rect 21180 19168 21232 19174
rect 21180 19110 21232 19116
rect 21192 18834 21220 19110
rect 21180 18828 21232 18834
rect 21180 18770 21232 18776
rect 21284 18426 21312 19944
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21272 18420 21324 18426
rect 21272 18362 21324 18368
rect 21180 18216 21232 18222
rect 21180 18158 21232 18164
rect 21088 16448 21140 16454
rect 21088 16390 21140 16396
rect 20904 16244 20956 16250
rect 20904 16186 20956 16192
rect 21192 14074 21220 18158
rect 21272 16720 21324 16726
rect 21272 16662 21324 16668
rect 21284 15162 21312 16662
rect 21272 15156 21324 15162
rect 21272 15098 21324 15104
rect 21376 14074 21404 19790
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 21364 14068 21416 14074
rect 21364 14010 21416 14016
rect 21468 13530 21496 20334
rect 21732 19372 21784 19378
rect 21732 19314 21784 19320
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21548 18284 21600 18290
rect 21548 18226 21600 18232
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 21456 13524 21508 13530
rect 21456 13466 21508 13472
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20720 12096 20772 12102
rect 20720 12038 20772 12044
rect 21100 11898 21128 12786
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21364 11756 21416 11762
rect 21364 11698 21416 11704
rect 21376 11529 21404 11698
rect 21362 11520 21418 11529
rect 21362 11455 21418 11464
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19143 7100 19451 7120
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7024 19451 7044
rect 18984 6905 19104 6914
rect 18984 6896 19118 6905
rect 18984 6886 19062 6896
rect 19062 6831 19118 6840
rect 19616 6792 19668 6798
rect 19614 6760 19616 6769
rect 19668 6760 19670 6769
rect 19614 6695 19670 6704
rect 19798 6760 19854 6769
rect 19798 6695 19854 6704
rect 19812 6662 19840 6695
rect 19800 6656 19852 6662
rect 19800 6598 19852 6604
rect 20076 6316 20128 6322
rect 20076 6258 20128 6264
rect 20088 6225 20116 6258
rect 20074 6216 20130 6225
rect 20074 6151 20130 6160
rect 19143 6012 19451 6032
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5936 19451 5956
rect 21560 5914 21588 18226
rect 21652 6458 21680 18702
rect 21744 16046 21772 19314
rect 21836 18902 21864 22200
rect 22296 19854 22324 22200
rect 22756 20398 22784 22200
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 22284 19848 22336 19854
rect 22284 19790 22336 19796
rect 21914 19272 21970 19281
rect 21914 19207 21970 19216
rect 21824 18896 21876 18902
rect 21824 18838 21876 18844
rect 21824 18692 21876 18698
rect 21824 18634 21876 18640
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21640 6452 21692 6458
rect 21640 6394 21692 6400
rect 21548 5908 21600 5914
rect 21548 5850 21600 5856
rect 21836 5846 21864 18634
rect 21928 14618 21956 19207
rect 21916 14612 21968 14618
rect 21916 14554 21968 14560
rect 21824 5840 21876 5846
rect 18694 5808 18750 5817
rect 21824 5782 21876 5788
rect 18694 5743 18750 5752
rect 20812 5704 20864 5710
rect 20812 5646 20864 5652
rect 17958 5264 18014 5273
rect 17958 5199 18014 5208
rect 20824 5166 20852 5646
rect 20812 5160 20864 5166
rect 20810 5128 20812 5137
rect 20864 5128 20866 5137
rect 20810 5063 20866 5072
rect 13945 4924 14253 4944
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4848 14253 4868
rect 19143 4924 19451 4944
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4848 19451 4868
rect 11058 4720 11114 4729
rect 11058 4655 11114 4664
rect 8298 4584 8354 4593
rect 8298 4519 8354 4528
rect 11346 4380 11654 4400
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4304 11654 4324
rect 16544 4380 16852 4400
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4304 16852 4324
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 8747 3836 9055 3856
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3760 9055 3780
rect 13945 3836 14253 3856
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3760 14253 3780
rect 19143 3836 19451 3856
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3760 19451 3780
rect 6148 3292 6456 3312
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3216 6456 3236
rect 11346 3292 11654 3312
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3216 11654 3236
rect 16544 3292 16852 3312
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3216 16852 3236
rect 8747 2748 9055 2768
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2672 9055 2692
rect 13945 2748 14253 2768
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2672 14253 2692
rect 19143 2748 19451 2768
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2672 19451 2692
rect 4896 2576 4948 2582
rect 4896 2518 4948 2524
rect 3424 2508 3476 2514
rect 3424 2450 3476 2456
rect 3240 2372 3292 2378
rect 3240 2314 3292 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 3054 2000 3110 2009
rect 3054 1935 3110 1944
rect 3252 1057 3280 2314
rect 3988 1601 4016 2314
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 6148 2204 6456 2224
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2128 6456 2148
rect 11346 2204 11654 2224
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2128 11654 2148
rect 3974 1592 4030 1601
rect 3974 1527 4030 1536
rect 11716 1170 11744 2246
rect 16544 2204 16852 2224
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2128 16852 2148
rect 11532 1142 11744 1170
rect 3238 1048 3294 1057
rect 3238 983 3294 992
rect 11532 800 11560 1142
rect 2870 640 2926 649
rect 2870 575 2926 584
rect 2778 232 2834 241
rect 2778 167 2834 176
rect 11518 0 11574 800
<< via2 >>
rect 2594 22616 2650 22672
rect 662 20032 718 20088
rect 478 11600 534 11656
rect 662 13504 718 13560
rect 1674 21256 1730 21312
rect 1398 18808 1454 18864
rect 938 12008 994 12064
rect 938 11872 994 11928
rect 1030 5480 1086 5536
rect 1490 17720 1546 17776
rect 3054 21664 3110 21720
rect 2134 19760 2190 19816
rect 1490 17040 1546 17096
rect 1582 16088 1638 16144
rect 1306 13232 1362 13288
rect 1582 15544 1638 15600
rect 1582 15136 1638 15192
rect 1490 14592 1546 14648
rect 1490 14220 1492 14240
rect 1492 14220 1544 14240
rect 1544 14220 1546 14240
rect 1490 14184 1546 14220
rect 1582 13796 1638 13832
rect 1582 13776 1584 13796
rect 1584 13776 1636 13796
rect 1636 13776 1638 13796
rect 1306 9016 1362 9072
rect 1766 15272 1822 15328
rect 1674 9444 1730 9480
rect 1674 9424 1676 9444
rect 1676 9424 1728 9444
rect 1728 9424 1730 9444
rect 1582 8880 1638 8936
rect 2042 16496 2098 16552
rect 2594 19352 2650 19408
rect 2318 18400 2374 18456
rect 2134 15272 2190 15328
rect 1490 8200 1546 8256
rect 1582 7268 1638 7304
rect 1582 7248 1584 7268
rect 1584 7248 1636 7268
rect 1636 7248 1638 7268
rect 2134 9560 2190 9616
rect 2042 8628 2098 8664
rect 2042 8608 2044 8628
rect 2044 8608 2096 8628
rect 2096 8608 2098 8628
rect 2134 7812 2190 7848
rect 2134 7792 2136 7812
rect 2136 7792 2188 7812
rect 2188 7792 2190 7812
rect 7010 22208 7066 22264
rect 3974 20712 4030 20768
rect 3238 18400 3294 18456
rect 3238 17992 3294 18048
rect 3146 17448 3202 17504
rect 2778 13640 2834 13696
rect 2686 13368 2742 13424
rect 2870 12824 2926 12880
rect 2502 12316 2504 12336
rect 2504 12316 2556 12336
rect 2556 12316 2558 12336
rect 2502 12280 2558 12316
rect 3054 12280 3110 12336
rect 2870 12008 2926 12064
rect 2686 11600 2742 11656
rect 2594 11328 2650 11384
rect 2502 9968 2558 10024
rect 1582 6296 1638 6352
rect 1858 6568 1914 6624
rect 1582 5908 1638 5944
rect 1582 5888 1584 5908
rect 1584 5888 1636 5908
rect 1636 5888 1638 5908
rect 1306 5344 1362 5400
rect 1398 5208 1454 5264
rect 938 3984 994 4040
rect 1582 4664 1638 4720
rect 1582 4528 1638 4584
rect 1858 4392 1914 4448
rect 2042 6604 2044 6624
rect 2044 6604 2096 6624
rect 2096 6604 2098 6624
rect 2042 6568 2098 6604
rect 2042 5616 2098 5672
rect 2042 5364 2098 5400
rect 2042 5344 2044 5364
rect 2044 5344 2096 5364
rect 2096 5344 2098 5364
rect 2226 7112 2282 7168
rect 2686 10412 2688 10432
rect 2688 10412 2740 10432
rect 2740 10412 2742 10432
rect 2686 10376 2742 10412
rect 2870 10648 2926 10704
rect 3054 10104 3110 10160
rect 2686 8336 2742 8392
rect 3054 9288 3110 9344
rect 2594 7928 2650 7984
rect 2502 6704 2558 6760
rect 2778 8064 2834 8120
rect 2686 6704 2742 6760
rect 3882 20304 3938 20360
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 3974 20168 4030 20224
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 4158 18128 4214 18184
rect 4434 19896 4490 19952
rect 4434 19372 4490 19408
rect 4434 19352 4436 19372
rect 4436 19352 4488 19372
rect 4488 19352 4490 19372
rect 4526 18672 4582 18728
rect 4986 19896 5042 19952
rect 4894 18264 4950 18320
rect 4710 17992 4766 18048
rect 3330 13368 3386 13424
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3790 14220 3792 14240
rect 3792 14220 3844 14240
rect 3844 14220 3846 14240
rect 3790 14184 3846 14220
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3974 13504 4030 13560
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3330 9016 3386 9072
rect 3054 6704 3110 6760
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3790 9424 3846 9480
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 2778 6452 2834 6488
rect 2778 6432 2780 6452
rect 2780 6432 2832 6452
rect 2832 6432 2834 6452
rect 2502 5788 2504 5808
rect 2504 5788 2556 5808
rect 2556 5788 2558 5808
rect 2502 5752 2558 5788
rect 2502 5208 2558 5264
rect 2226 3848 2282 3904
rect 1950 3596 2006 3632
rect 1950 3576 1952 3596
rect 1952 3576 2004 3596
rect 2004 3576 2006 3596
rect 2226 3476 2228 3496
rect 2228 3476 2280 3496
rect 2280 3476 2282 3496
rect 2226 3440 2282 3476
rect 2778 6160 2834 6216
rect 4066 12280 4122 12336
rect 4618 15952 4674 16008
rect 4342 10920 4398 10976
rect 4066 9288 4122 9344
rect 3974 8472 4030 8528
rect 3422 7520 3478 7576
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3790 6860 3846 6896
rect 3790 6840 3792 6860
rect 3792 6840 3844 6860
rect 3844 6840 3846 6860
rect 3790 6452 3846 6488
rect 3790 6432 3792 6452
rect 3792 6432 3844 6452
rect 3844 6432 3846 6452
rect 2778 4800 2834 4856
rect 3422 6180 3478 6216
rect 3422 6160 3424 6180
rect 3424 6160 3476 6180
rect 3476 6160 3478 6180
rect 3330 6024 3386 6080
rect 3238 5888 3294 5944
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 3882 5208 3938 5264
rect 3238 4004 3294 4040
rect 3238 3984 3240 4004
rect 3240 3984 3292 4004
rect 3292 3984 3294 4004
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 4802 15816 4858 15872
rect 4894 13504 4950 13560
rect 4526 10648 4582 10704
rect 4618 9560 4674 9616
rect 4618 9444 4674 9480
rect 4618 9424 4620 9444
rect 4620 9424 4672 9444
rect 4672 9424 4674 9444
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 5630 18808 5686 18864
rect 5354 10512 5410 10568
rect 2778 2896 2834 2952
rect 2778 2488 2834 2544
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 4618 5908 4674 5944
rect 4618 5888 4620 5908
rect 4620 5888 4672 5908
rect 4672 5888 4674 5908
rect 4618 5480 4674 5536
rect 4526 3576 4582 3632
rect 5998 19760 6054 19816
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6090 18808 6146 18864
rect 6550 19372 6606 19408
rect 6550 19352 6552 19372
rect 6552 19352 6604 19372
rect 6604 19352 6606 19372
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 5998 18400 6054 18456
rect 6458 18284 6514 18320
rect 6458 18264 6460 18284
rect 6460 18264 6512 18284
rect 6512 18264 6514 18284
rect 5906 17720 5962 17776
rect 5906 17484 5908 17504
rect 5908 17484 5960 17504
rect 5960 17484 5962 17504
rect 5906 17448 5962 17484
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 7378 18264 7434 18320
rect 8022 20168 8078 20224
rect 7470 18128 7526 18184
rect 6826 15952 6882 16008
rect 7102 15816 7158 15872
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 6550 11464 6606 11520
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6090 7928 6146 7984
rect 6826 9580 6882 9616
rect 6826 9560 6828 9580
rect 6828 9560 6880 9580
rect 6880 9560 6882 9580
rect 6918 9288 6974 9344
rect 7746 18672 7802 18728
rect 7838 18264 7894 18320
rect 7378 12280 7434 12336
rect 7378 9016 7434 9072
rect 7286 8336 7342 8392
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 4986 5908 5042 5944
rect 4986 5888 4988 5908
rect 4988 5888 5040 5908
rect 5040 5888 5042 5908
rect 5354 5908 5410 5944
rect 5354 5888 5356 5908
rect 5356 5888 5408 5908
rect 5408 5888 5410 5908
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 7654 9560 7710 9616
rect 8942 20304 8998 20360
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8758 19932 8760 19952
rect 8760 19932 8812 19952
rect 8812 19932 8814 19952
rect 8758 19896 8814 19932
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8942 17584 8998 17640
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9678 17312 9734 17368
rect 8758 16532 8760 16552
rect 8760 16532 8812 16552
rect 8812 16532 8814 16552
rect 8758 16496 8814 16532
rect 9126 15952 9182 16008
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8482 12280 8538 12336
rect 7930 10920 7986 10976
rect 8206 9016 8262 9072
rect 8482 7384 8538 7440
rect 7562 6840 7618 6896
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 9586 17040 9642 17096
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 10138 17176 10194 17232
rect 9954 13776 10010 13832
rect 9494 12688 9550 12744
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 9770 10920 9826 10976
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 9310 9016 9366 9072
rect 9586 9596 9588 9616
rect 9588 9596 9640 9616
rect 9640 9596 9642 9616
rect 9586 9560 9642 9596
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 12162 20304 12218 20360
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11150 17312 11206 17368
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 12714 19896 12770 19952
rect 12254 19760 12310 19816
rect 11978 17584 12034 17640
rect 12254 18400 12310 18456
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11702 12144 11758 12200
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 13818 20304 13874 20360
rect 12898 17040 12954 17096
rect 13634 19760 13690 19816
rect 13358 17196 13414 17232
rect 13358 17176 13360 17196
rect 13360 17176 13412 17196
rect 13412 17176 13414 17196
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 13818 19216 13874 19272
rect 14462 19080 14518 19136
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13818 18844 13820 18864
rect 13820 18844 13872 18864
rect 13872 18844 13874 18864
rect 13818 18808 13874 18844
rect 14094 18400 14150 18456
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 14462 17448 14518 17504
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13358 13252 13414 13288
rect 13358 13232 13360 13252
rect 13360 13232 13412 13252
rect 13412 13232 13414 13252
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 15750 19352 15806 19408
rect 16026 19352 16082 19408
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16486 19796 16488 19816
rect 16488 19796 16540 19816
rect 16540 19796 16542 19816
rect 15198 17448 15254 17504
rect 15014 16632 15070 16688
rect 10322 8336 10378 8392
rect 9862 7248 9918 7304
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8298 5888 8354 5944
rect 7562 5616 7618 5672
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 15290 17196 15346 17232
rect 15290 17176 15292 17196
rect 15292 17176 15344 17196
rect 15344 17176 15346 17196
rect 16486 19760 16542 19796
rect 17038 19760 17094 19816
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 16946 19352 17002 19408
rect 16854 19216 16910 19272
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 15566 16496 15622 16552
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16210 17176 16266 17232
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 17038 15020 17094 15056
rect 17038 15000 17040 15020
rect 17040 15000 17092 15020
rect 17092 15000 17094 15020
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16394 11736 16450 11792
rect 15014 8880 15070 8936
rect 14462 7792 14518 7848
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 17406 19080 17462 19136
rect 18142 18808 18198 18864
rect 17590 17740 17646 17776
rect 17590 17720 17592 17740
rect 17592 17720 17644 17740
rect 17644 17720 17646 17740
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19338 19896 19394 19952
rect 18694 19080 18750 19136
rect 18786 16652 18842 16688
rect 18786 16632 18788 16652
rect 18788 16632 18840 16652
rect 18840 16632 18842 16652
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 15750 6296 15806 6352
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 19614 15308 19616 15328
rect 19616 15308 19668 15328
rect 19668 15308 19670 15328
rect 19614 15272 19670 15308
rect 19798 14320 19854 14376
rect 20626 19372 20682 19408
rect 20626 19352 20628 19372
rect 20628 19352 20680 19372
rect 20680 19352 20682 19372
rect 20626 18148 20682 18184
rect 20626 18128 20628 18148
rect 20628 18128 20680 18148
rect 20680 18128 20682 18148
rect 20810 18284 20866 18320
rect 20810 18264 20812 18284
rect 20812 18264 20864 18284
rect 20864 18264 20866 18284
rect 20534 14356 20536 14376
rect 20536 14356 20588 14376
rect 20588 14356 20590 14376
rect 20534 14320 20590 14356
rect 20902 16496 20958 16552
rect 21362 11464 21418 11520
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 19062 6840 19118 6896
rect 19614 6740 19616 6760
rect 19616 6740 19668 6760
rect 19668 6740 19670 6760
rect 19614 6704 19670 6740
rect 19798 6704 19854 6760
rect 20074 6160 20130 6216
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 21914 19216 21970 19272
rect 18694 5752 18750 5808
rect 17958 5208 18014 5264
rect 20810 5108 20812 5128
rect 20812 5108 20864 5128
rect 20864 5108 20866 5128
rect 20810 5072 20866 5108
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 11058 4664 11114 4720
rect 8298 4528 8354 4584
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 3054 1944 3110 2000
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 3974 1536 4030 1592
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 3238 992 3294 1048
rect 2870 584 2926 640
rect 2778 176 2834 232
<< metal3 >>
rect 0 22674 800 22704
rect 2589 22674 2655 22677
rect 0 22672 2655 22674
rect 0 22616 2594 22672
rect 2650 22616 2655 22672
rect 0 22614 2655 22616
rect 0 22584 800 22614
rect 2589 22611 2655 22614
rect 0 22266 800 22296
rect 7005 22266 7071 22269
rect 0 22264 7071 22266
rect 0 22208 7010 22264
rect 7066 22208 7071 22264
rect 0 22206 7071 22208
rect 0 22176 800 22206
rect 7005 22203 7071 22206
rect 0 21722 800 21752
rect 3049 21722 3115 21725
rect 0 21720 3115 21722
rect 0 21664 3054 21720
rect 3110 21664 3115 21720
rect 0 21662 3115 21664
rect 0 21632 800 21662
rect 3049 21659 3115 21662
rect 0 21314 800 21344
rect 1669 21314 1735 21317
rect 0 21312 1735 21314
rect 0 21256 1674 21312
rect 1730 21256 1735 21312
rect 0 21254 1735 21256
rect 0 21224 800 21254
rect 1669 21251 1735 21254
rect 0 20770 800 20800
rect 3969 20770 4035 20773
rect 0 20768 4035 20770
rect 0 20712 3974 20768
rect 4030 20712 4035 20768
rect 0 20710 4035 20712
rect 0 20680 800 20710
rect 3969 20707 4035 20710
rect 6142 20704 6462 20705
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 20639 6462 20640
rect 11340 20704 11660 20705
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 20639 11660 20640
rect 16538 20704 16858 20705
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 20639 16858 20640
rect 0 20362 800 20392
rect 3877 20362 3943 20365
rect 0 20360 3943 20362
rect 0 20304 3882 20360
rect 3938 20304 3943 20360
rect 0 20302 3943 20304
rect 0 20272 800 20302
rect 3877 20299 3943 20302
rect 8518 20300 8524 20364
rect 8588 20362 8594 20364
rect 8937 20362 9003 20365
rect 8588 20360 9003 20362
rect 8588 20304 8942 20360
rect 8998 20304 9003 20360
rect 8588 20302 9003 20304
rect 8588 20300 8594 20302
rect 8937 20299 9003 20302
rect 12157 20362 12223 20365
rect 13813 20362 13879 20365
rect 12157 20360 13879 20362
rect 12157 20304 12162 20360
rect 12218 20304 13818 20360
rect 13874 20304 13879 20360
rect 12157 20302 13879 20304
rect 12157 20299 12223 20302
rect 13813 20299 13879 20302
rect 3969 20226 4035 20229
rect 8017 20226 8083 20229
rect 3969 20224 8083 20226
rect 3969 20168 3974 20224
rect 4030 20168 8022 20224
rect 8078 20168 8083 20224
rect 3969 20166 8083 20168
rect 3969 20163 4035 20166
rect 8017 20163 8083 20166
rect 3543 20160 3863 20161
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 20095 3863 20096
rect 8741 20160 9061 20161
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 20095 9061 20096
rect 13939 20160 14259 20161
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 20095 14259 20096
rect 19137 20160 19457 20161
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 20095 19457 20096
rect 657 20090 723 20093
rect 657 20088 2790 20090
rect 657 20032 662 20088
rect 718 20032 2790 20088
rect 657 20030 2790 20032
rect 657 20027 723 20030
rect 2730 19954 2790 20030
rect 4429 19954 4495 19957
rect 2730 19952 4495 19954
rect 2730 19896 4434 19952
rect 4490 19896 4495 19952
rect 2730 19894 4495 19896
rect 4429 19891 4495 19894
rect 4981 19954 5047 19957
rect 8753 19954 8819 19957
rect 4981 19952 8819 19954
rect 4981 19896 4986 19952
rect 5042 19896 8758 19952
rect 8814 19896 8819 19952
rect 4981 19894 8819 19896
rect 4981 19891 5047 19894
rect 8753 19891 8819 19894
rect 12709 19954 12775 19957
rect 19333 19954 19399 19957
rect 12709 19952 19399 19954
rect 12709 19896 12714 19952
rect 12770 19896 19338 19952
rect 19394 19896 19399 19952
rect 12709 19894 19399 19896
rect 12709 19891 12775 19894
rect 19333 19891 19399 19894
rect 0 19818 800 19848
rect 2129 19818 2195 19821
rect 0 19816 2195 19818
rect 0 19760 2134 19816
rect 2190 19760 2195 19816
rect 0 19758 2195 19760
rect 0 19728 800 19758
rect 2129 19755 2195 19758
rect 5993 19818 6059 19821
rect 12249 19818 12315 19821
rect 5993 19816 12315 19818
rect 5993 19760 5998 19816
rect 6054 19760 12254 19816
rect 12310 19760 12315 19816
rect 5993 19758 12315 19760
rect 5993 19755 6059 19758
rect 12249 19755 12315 19758
rect 13629 19818 13695 19821
rect 16481 19818 16547 19821
rect 17033 19818 17099 19821
rect 13629 19816 17099 19818
rect 13629 19760 13634 19816
rect 13690 19760 16486 19816
rect 16542 19760 17038 19816
rect 17094 19760 17099 19816
rect 13629 19758 17099 19760
rect 13629 19755 13695 19758
rect 16481 19755 16547 19758
rect 17033 19755 17099 19758
rect 6142 19616 6462 19617
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 6142 19551 6462 19552
rect 11340 19616 11660 19617
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 19551 11660 19552
rect 16538 19616 16858 19617
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 19551 16858 19552
rect 0 19410 800 19440
rect 2589 19410 2655 19413
rect 0 19408 2655 19410
rect 0 19352 2594 19408
rect 2650 19352 2655 19408
rect 0 19350 2655 19352
rect 0 19320 800 19350
rect 2589 19347 2655 19350
rect 4429 19410 4495 19413
rect 5022 19410 5028 19412
rect 4429 19408 5028 19410
rect 4429 19352 4434 19408
rect 4490 19352 5028 19408
rect 4429 19350 5028 19352
rect 4429 19347 4495 19350
rect 5022 19348 5028 19350
rect 5092 19348 5098 19412
rect 6545 19410 6611 19413
rect 6678 19410 6684 19412
rect 6545 19408 6684 19410
rect 6545 19352 6550 19408
rect 6606 19352 6684 19408
rect 6545 19350 6684 19352
rect 6545 19347 6611 19350
rect 6678 19348 6684 19350
rect 6748 19348 6754 19412
rect 15142 19348 15148 19412
rect 15212 19410 15218 19412
rect 15745 19410 15811 19413
rect 15212 19408 15811 19410
rect 15212 19352 15750 19408
rect 15806 19352 15811 19408
rect 15212 19350 15811 19352
rect 15212 19348 15218 19350
rect 15745 19347 15811 19350
rect 16021 19412 16087 19413
rect 16941 19412 17007 19413
rect 16021 19408 16068 19412
rect 16132 19410 16138 19412
rect 16021 19352 16026 19408
rect 16021 19348 16068 19352
rect 16132 19350 16178 19410
rect 16941 19408 16988 19412
rect 17052 19410 17058 19412
rect 16941 19352 16946 19408
rect 16132 19348 16138 19350
rect 16941 19348 16988 19352
rect 17052 19350 17098 19410
rect 17052 19348 17058 19350
rect 19926 19348 19932 19412
rect 19996 19410 20002 19412
rect 20621 19410 20687 19413
rect 19996 19408 20687 19410
rect 19996 19352 20626 19408
rect 20682 19352 20687 19408
rect 19996 19350 20687 19352
rect 19996 19348 20002 19350
rect 16021 19347 16087 19348
rect 16941 19347 17007 19348
rect 20621 19347 20687 19350
rect 13813 19274 13879 19277
rect 16849 19274 16915 19277
rect 21909 19274 21975 19277
rect 13813 19272 21975 19274
rect 13813 19216 13818 19272
rect 13874 19216 16854 19272
rect 16910 19216 21914 19272
rect 21970 19216 21975 19272
rect 13813 19214 21975 19216
rect 13813 19211 13879 19214
rect 16849 19211 16915 19214
rect 21909 19211 21975 19214
rect 14457 19138 14523 19141
rect 17401 19138 17467 19141
rect 18689 19138 18755 19141
rect 14457 19136 18755 19138
rect 14457 19080 14462 19136
rect 14518 19080 17406 19136
rect 17462 19080 18694 19136
rect 18750 19080 18755 19136
rect 14457 19078 18755 19080
rect 14457 19075 14523 19078
rect 17401 19075 17467 19078
rect 18689 19075 18755 19078
rect 3543 19072 3863 19073
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 19007 3863 19008
rect 8741 19072 9061 19073
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 19007 9061 19008
rect 13939 19072 14259 19073
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 19007 14259 19008
rect 19137 19072 19457 19073
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 19007 19457 19008
rect 0 18866 800 18896
rect 1393 18866 1459 18869
rect 0 18864 1459 18866
rect 0 18808 1398 18864
rect 1454 18808 1459 18864
rect 0 18806 1459 18808
rect 0 18776 800 18806
rect 1393 18803 1459 18806
rect 4470 18804 4476 18868
rect 4540 18866 4546 18868
rect 5625 18866 5691 18869
rect 4540 18864 5691 18866
rect 4540 18808 5630 18864
rect 5686 18808 5691 18864
rect 4540 18806 5691 18808
rect 4540 18804 4546 18806
rect 5625 18803 5691 18806
rect 5942 18804 5948 18868
rect 6012 18866 6018 18868
rect 6085 18866 6151 18869
rect 6012 18864 6151 18866
rect 6012 18808 6090 18864
rect 6146 18808 6151 18864
rect 6012 18806 6151 18808
rect 6012 18804 6018 18806
rect 6085 18803 6151 18806
rect 13813 18866 13879 18869
rect 18137 18866 18203 18869
rect 13813 18864 18203 18866
rect 13813 18808 13818 18864
rect 13874 18808 18142 18864
rect 18198 18808 18203 18864
rect 13813 18806 18203 18808
rect 13813 18803 13879 18806
rect 18137 18803 18203 18806
rect 4521 18730 4587 18733
rect 7741 18730 7807 18733
rect 4521 18728 7807 18730
rect 4521 18672 4526 18728
rect 4582 18672 7746 18728
rect 7802 18672 7807 18728
rect 4521 18670 7807 18672
rect 4521 18667 4587 18670
rect 7741 18667 7807 18670
rect 6142 18528 6462 18529
rect 0 18458 800 18488
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 18463 6462 18464
rect 11340 18528 11660 18529
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 18463 11660 18464
rect 16538 18528 16858 18529
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 18463 16858 18464
rect 2313 18458 2379 18461
rect 0 18456 2379 18458
rect 0 18400 2318 18456
rect 2374 18400 2379 18456
rect 0 18398 2379 18400
rect 0 18368 800 18398
rect 2313 18395 2379 18398
rect 3233 18458 3299 18461
rect 5993 18458 6059 18461
rect 3233 18456 6059 18458
rect 3233 18400 3238 18456
rect 3294 18400 5998 18456
rect 6054 18400 6059 18456
rect 3233 18398 6059 18400
rect 3233 18395 3299 18398
rect 5993 18395 6059 18398
rect 12249 18458 12315 18461
rect 14089 18458 14155 18461
rect 12249 18456 14155 18458
rect 12249 18400 12254 18456
rect 12310 18400 14094 18456
rect 14150 18400 14155 18456
rect 12249 18398 14155 18400
rect 12249 18395 12315 18398
rect 14089 18395 14155 18398
rect 4889 18322 4955 18325
rect 6453 18322 6519 18325
rect 7373 18322 7439 18325
rect 4889 18320 6519 18322
rect 4889 18264 4894 18320
rect 4950 18264 6458 18320
rect 6514 18264 6519 18320
rect 4889 18262 6519 18264
rect 4889 18259 4955 18262
rect 6453 18259 6519 18262
rect 7238 18320 7439 18322
rect 7238 18264 7378 18320
rect 7434 18264 7439 18320
rect 7238 18262 7439 18264
rect 4153 18186 4219 18189
rect 4286 18186 4292 18188
rect 4153 18184 4292 18186
rect 4153 18128 4158 18184
rect 4214 18128 4292 18184
rect 4153 18126 4292 18128
rect 4153 18123 4219 18126
rect 4286 18124 4292 18126
rect 4356 18186 4362 18188
rect 7238 18186 7298 18262
rect 7373 18259 7439 18262
rect 7833 18322 7899 18325
rect 20805 18322 20871 18325
rect 7833 18320 20871 18322
rect 7833 18264 7838 18320
rect 7894 18264 20810 18320
rect 20866 18264 20871 18320
rect 7833 18262 20871 18264
rect 7833 18259 7899 18262
rect 20805 18259 20871 18262
rect 4356 18126 7298 18186
rect 7465 18186 7531 18189
rect 7465 18184 12450 18186
rect 7465 18128 7470 18184
rect 7526 18128 12450 18184
rect 7465 18126 12450 18128
rect 4356 18124 4362 18126
rect 7465 18123 7531 18126
rect 0 18050 800 18080
rect 3233 18050 3299 18053
rect 0 18048 3299 18050
rect 0 17992 3238 18048
rect 3294 17992 3299 18048
rect 0 17990 3299 17992
rect 0 17960 800 17990
rect 3233 17987 3299 17990
rect 4705 18050 4771 18053
rect 4838 18050 4844 18052
rect 4705 18048 4844 18050
rect 4705 17992 4710 18048
rect 4766 17992 4844 18048
rect 4705 17990 4844 17992
rect 4705 17987 4771 17990
rect 4838 17988 4844 17990
rect 4908 17988 4914 18052
rect 3543 17984 3863 17985
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 17919 3863 17920
rect 8741 17984 9061 17985
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 17919 9061 17920
rect 1485 17778 1551 17781
rect 5901 17778 5967 17781
rect 1485 17776 5967 17778
rect 1485 17720 1490 17776
rect 1546 17720 5906 17776
rect 5962 17720 5967 17776
rect 1485 17718 5967 17720
rect 12390 17778 12450 18126
rect 17166 18124 17172 18188
rect 17236 18186 17242 18188
rect 20621 18186 20687 18189
rect 17236 18184 20687 18186
rect 17236 18128 20626 18184
rect 20682 18128 20687 18184
rect 17236 18126 20687 18128
rect 17236 18124 17242 18126
rect 20621 18123 20687 18126
rect 13939 17984 14259 17985
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 17919 14259 17920
rect 19137 17984 19457 17985
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 17919 19457 17920
rect 17585 17778 17651 17781
rect 12390 17776 17651 17778
rect 12390 17720 17590 17776
rect 17646 17720 17651 17776
rect 12390 17718 17651 17720
rect 1485 17715 1551 17718
rect 5901 17715 5967 17718
rect 17585 17715 17651 17718
rect 8937 17642 9003 17645
rect 11973 17642 12039 17645
rect 8937 17640 12039 17642
rect 8937 17584 8942 17640
rect 8998 17584 11978 17640
rect 12034 17584 12039 17640
rect 8937 17582 12039 17584
rect 8937 17579 9003 17582
rect 11973 17579 12039 17582
rect 0 17506 800 17536
rect 3141 17506 3207 17509
rect 5901 17508 5967 17509
rect 5901 17506 5948 17508
rect 0 17504 3207 17506
rect 0 17448 3146 17504
rect 3202 17448 3207 17504
rect 0 17446 3207 17448
rect 5856 17504 5948 17506
rect 5856 17448 5906 17504
rect 5856 17446 5948 17448
rect 0 17416 800 17446
rect 3141 17443 3207 17446
rect 5901 17444 5948 17446
rect 6012 17444 6018 17508
rect 14457 17506 14523 17509
rect 15193 17506 15259 17509
rect 14457 17504 15259 17506
rect 14457 17448 14462 17504
rect 14518 17448 15198 17504
rect 15254 17448 15259 17504
rect 14457 17446 15259 17448
rect 5901 17443 5967 17444
rect 14457 17443 14523 17446
rect 15193 17443 15259 17446
rect 6142 17440 6462 17441
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 17375 6462 17376
rect 11340 17440 11660 17441
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 17375 11660 17376
rect 16538 17440 16858 17441
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 17375 16858 17376
rect 9673 17370 9739 17373
rect 11145 17370 11211 17373
rect 9673 17368 11211 17370
rect 9673 17312 9678 17368
rect 9734 17312 11150 17368
rect 11206 17312 11211 17368
rect 9673 17310 11211 17312
rect 9673 17307 9739 17310
rect 11145 17307 11211 17310
rect 10133 17234 10199 17237
rect 13353 17234 13419 17237
rect 10133 17232 13419 17234
rect 10133 17176 10138 17232
rect 10194 17176 13358 17232
rect 13414 17176 13419 17232
rect 10133 17174 13419 17176
rect 10133 17171 10199 17174
rect 13353 17171 13419 17174
rect 15285 17234 15351 17237
rect 16205 17234 16271 17237
rect 15285 17232 16271 17234
rect 15285 17176 15290 17232
rect 15346 17176 16210 17232
rect 16266 17176 16271 17232
rect 15285 17174 16271 17176
rect 15285 17171 15351 17174
rect 16205 17171 16271 17174
rect 0 17098 800 17128
rect 1485 17098 1551 17101
rect 0 17096 1551 17098
rect 0 17040 1490 17096
rect 1546 17040 1551 17096
rect 0 17038 1551 17040
rect 0 17008 800 17038
rect 1485 17035 1551 17038
rect 9581 17098 9647 17101
rect 12893 17098 12959 17101
rect 9581 17096 12959 17098
rect 9581 17040 9586 17096
rect 9642 17040 12898 17096
rect 12954 17040 12959 17096
rect 9581 17038 12959 17040
rect 9581 17035 9647 17038
rect 12893 17035 12959 17038
rect 3543 16896 3863 16897
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 16831 3863 16832
rect 8741 16896 9061 16897
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 16831 9061 16832
rect 13939 16896 14259 16897
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 16831 14259 16832
rect 19137 16896 19457 16897
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 16831 19457 16832
rect 15009 16690 15075 16693
rect 18781 16690 18847 16693
rect 15009 16688 18847 16690
rect 15009 16632 15014 16688
rect 15070 16632 18786 16688
rect 18842 16632 18847 16688
rect 15009 16630 18847 16632
rect 15009 16627 15075 16630
rect 18781 16627 18847 16630
rect 0 16554 800 16584
rect 2037 16554 2103 16557
rect 0 16552 2103 16554
rect 0 16496 2042 16552
rect 2098 16496 2103 16552
rect 0 16494 2103 16496
rect 0 16464 800 16494
rect 2037 16491 2103 16494
rect 5942 16492 5948 16556
rect 6012 16554 6018 16556
rect 8753 16554 8819 16557
rect 6012 16552 8819 16554
rect 6012 16496 8758 16552
rect 8814 16496 8819 16552
rect 6012 16494 8819 16496
rect 6012 16492 6018 16494
rect 8753 16491 8819 16494
rect 15561 16554 15627 16557
rect 20897 16554 20963 16557
rect 15561 16552 20963 16554
rect 15561 16496 15566 16552
rect 15622 16496 20902 16552
rect 20958 16496 20963 16552
rect 15561 16494 20963 16496
rect 15561 16491 15627 16494
rect 20897 16491 20963 16494
rect 6142 16352 6462 16353
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 16287 6462 16288
rect 11340 16352 11660 16353
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 16287 11660 16288
rect 16538 16352 16858 16353
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 16287 16858 16288
rect 0 16146 800 16176
rect 1577 16146 1643 16149
rect 0 16144 1643 16146
rect 0 16088 1582 16144
rect 1638 16088 1643 16144
rect 0 16086 1643 16088
rect 0 16056 800 16086
rect 1577 16083 1643 16086
rect 4613 16010 4679 16013
rect 6821 16010 6887 16013
rect 9121 16010 9187 16013
rect 4613 16008 9187 16010
rect 4613 15952 4618 16008
rect 4674 15952 6826 16008
rect 6882 15952 9126 16008
rect 9182 15952 9187 16008
rect 4613 15950 9187 15952
rect 4613 15947 4679 15950
rect 6821 15947 6887 15950
rect 9121 15947 9187 15950
rect 4797 15874 4863 15877
rect 7097 15874 7163 15877
rect 4797 15872 7163 15874
rect 4797 15816 4802 15872
rect 4858 15816 7102 15872
rect 7158 15816 7163 15872
rect 4797 15814 7163 15816
rect 4797 15811 4863 15814
rect 7097 15811 7163 15814
rect 3543 15808 3863 15809
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3543 15743 3863 15744
rect 8741 15808 9061 15809
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 15743 9061 15744
rect 13939 15808 14259 15809
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 15743 14259 15744
rect 19137 15808 19457 15809
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 15743 19457 15744
rect 0 15602 800 15632
rect 1577 15602 1643 15605
rect 0 15600 1643 15602
rect 0 15544 1582 15600
rect 1638 15544 1643 15600
rect 0 15542 1643 15544
rect 0 15512 800 15542
rect 1577 15539 1643 15542
rect 1761 15332 1827 15333
rect 2129 15332 2195 15333
rect 1710 15330 1716 15332
rect 1670 15270 1716 15330
rect 1780 15328 1827 15332
rect 2078 15330 2084 15332
rect 1822 15272 1827 15328
rect 1710 15268 1716 15270
rect 1780 15268 1827 15272
rect 2038 15270 2084 15330
rect 2148 15328 2195 15332
rect 2190 15272 2195 15328
rect 2078 15268 2084 15270
rect 2148 15268 2195 15272
rect 1761 15267 1827 15268
rect 2129 15267 2195 15268
rect 19609 15330 19675 15333
rect 19742 15330 19748 15332
rect 19609 15328 19748 15330
rect 19609 15272 19614 15328
rect 19670 15272 19748 15328
rect 19609 15270 19748 15272
rect 19609 15267 19675 15270
rect 19742 15268 19748 15270
rect 19812 15268 19818 15332
rect 6142 15264 6462 15265
rect 0 15194 800 15224
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 15199 6462 15200
rect 11340 15264 11660 15265
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 15199 11660 15200
rect 16538 15264 16858 15265
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 15199 16858 15200
rect 1577 15194 1643 15197
rect 0 15192 1643 15194
rect 0 15136 1582 15192
rect 1638 15136 1643 15192
rect 0 15134 1643 15136
rect 0 15104 800 15134
rect 1577 15131 1643 15134
rect 1158 14996 1164 15060
rect 1228 15058 1234 15060
rect 17033 15058 17099 15061
rect 1228 15056 17099 15058
rect 1228 15000 17038 15056
rect 17094 15000 17099 15056
rect 1228 14998 17099 15000
rect 1228 14996 1234 14998
rect 17033 14995 17099 14998
rect 3543 14720 3863 14721
rect 0 14650 800 14680
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3543 14655 3863 14656
rect 8741 14720 9061 14721
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 14655 9061 14656
rect 13939 14720 14259 14721
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 14655 14259 14656
rect 19137 14720 19457 14721
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 14655 19457 14656
rect 1485 14650 1551 14653
rect 0 14648 1551 14650
rect 0 14592 1490 14648
rect 1546 14592 1551 14648
rect 0 14590 1551 14592
rect 0 14560 800 14590
rect 1485 14587 1551 14590
rect 974 14316 980 14380
rect 1044 14378 1050 14380
rect 19793 14378 19859 14381
rect 20529 14378 20595 14381
rect 1044 14376 20595 14378
rect 1044 14320 19798 14376
rect 19854 14320 20534 14376
rect 20590 14320 20595 14376
rect 1044 14318 20595 14320
rect 1044 14316 1050 14318
rect 19793 14315 19859 14318
rect 20529 14315 20595 14318
rect 0 14242 800 14272
rect 1485 14242 1551 14245
rect 0 14240 1551 14242
rect 0 14184 1490 14240
rect 1546 14184 1551 14240
rect 0 14182 1551 14184
rect 0 14152 800 14182
rect 1485 14179 1551 14182
rect 3785 14242 3851 14245
rect 3918 14242 3924 14244
rect 3785 14240 3924 14242
rect 3785 14184 3790 14240
rect 3846 14184 3924 14240
rect 3785 14182 3924 14184
rect 3785 14179 3851 14182
rect 3918 14180 3924 14182
rect 3988 14180 3994 14244
rect 6142 14176 6462 14177
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 14111 6462 14112
rect 11340 14176 11660 14177
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 14111 11660 14112
rect 16538 14176 16858 14177
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 14111 16858 14112
rect 0 13834 800 13864
rect 1577 13834 1643 13837
rect 9949 13834 10015 13837
rect 0 13832 1643 13834
rect 0 13776 1582 13832
rect 1638 13776 1643 13832
rect 0 13774 1643 13776
rect 0 13744 800 13774
rect 1577 13771 1643 13774
rect 3374 13832 10015 13834
rect 3374 13776 9954 13832
rect 10010 13776 10015 13832
rect 3374 13774 10015 13776
rect 2630 13636 2636 13700
rect 2700 13698 2706 13700
rect 2773 13698 2839 13701
rect 2700 13696 2839 13698
rect 2700 13640 2778 13696
rect 2834 13640 2839 13696
rect 2700 13638 2839 13640
rect 2700 13636 2706 13638
rect 2773 13635 2839 13638
rect 657 13562 723 13565
rect 3374 13562 3434 13774
rect 9949 13771 10015 13774
rect 3543 13632 3863 13633
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 13567 3863 13568
rect 8741 13632 9061 13633
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 13567 9061 13568
rect 13939 13632 14259 13633
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 13567 14259 13568
rect 19137 13632 19457 13633
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 13567 19457 13568
rect 657 13560 1594 13562
rect 657 13504 662 13560
rect 718 13504 1594 13560
rect 657 13502 1594 13504
rect 657 13499 723 13502
rect 0 13290 800 13320
rect 1301 13290 1367 13293
rect 0 13288 1367 13290
rect 0 13232 1306 13288
rect 1362 13232 1367 13288
rect 0 13230 1367 13232
rect 1534 13290 1594 13502
rect 2730 13502 3434 13562
rect 3969 13562 4035 13565
rect 4470 13562 4476 13564
rect 3969 13560 4476 13562
rect 3969 13504 3974 13560
rect 4030 13504 4476 13560
rect 3969 13502 4476 13504
rect 2730 13429 2790 13502
rect 3969 13499 4035 13502
rect 4470 13500 4476 13502
rect 4540 13562 4546 13564
rect 4889 13562 4955 13565
rect 4540 13560 4955 13562
rect 4540 13504 4894 13560
rect 4950 13504 4955 13560
rect 4540 13502 4955 13504
rect 4540 13500 4546 13502
rect 4889 13499 4955 13502
rect 2681 13424 2790 13429
rect 2681 13368 2686 13424
rect 2742 13368 2790 13424
rect 2681 13366 2790 13368
rect 3325 13426 3391 13429
rect 4102 13426 4108 13428
rect 3325 13424 4108 13426
rect 3325 13368 3330 13424
rect 3386 13368 4108 13424
rect 3325 13366 4108 13368
rect 2681 13363 2747 13366
rect 3325 13363 3391 13366
rect 4102 13364 4108 13366
rect 4172 13364 4178 13428
rect 13353 13290 13419 13293
rect 1534 13288 13419 13290
rect 1534 13232 13358 13288
rect 13414 13232 13419 13288
rect 1534 13230 13419 13232
rect 0 13200 800 13230
rect 1301 13227 1367 13230
rect 13353 13227 13419 13230
rect 6142 13088 6462 13089
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 13023 6462 13024
rect 11340 13088 11660 13089
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 13023 11660 13024
rect 16538 13088 16858 13089
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 13023 16858 13024
rect 0 12882 800 12912
rect 2865 12882 2931 12885
rect 0 12880 2931 12882
rect 0 12824 2870 12880
rect 2926 12824 2931 12880
rect 0 12822 2931 12824
rect 0 12792 800 12822
rect 2865 12819 2931 12822
rect 9489 12746 9555 12749
rect 15142 12746 15148 12748
rect 9489 12744 15148 12746
rect 9489 12688 9494 12744
rect 9550 12688 15148 12744
rect 9489 12686 15148 12688
rect 9489 12683 9555 12686
rect 15142 12684 15148 12686
rect 15212 12684 15218 12748
rect 3543 12544 3863 12545
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 12479 3863 12480
rect 8741 12544 9061 12545
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 12479 9061 12480
rect 13939 12544 14259 12545
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 12479 14259 12480
rect 19137 12544 19457 12545
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19137 12479 19457 12480
rect 0 12338 800 12368
rect 2497 12338 2563 12341
rect 3049 12338 3115 12341
rect 3182 12338 3188 12340
rect 0 12278 2146 12338
rect 0 12248 800 12278
rect 933 12066 999 12069
rect 1342 12066 1348 12068
rect 933 12064 1348 12066
rect 933 12008 938 12064
rect 994 12008 1348 12064
rect 933 12006 1348 12008
rect 933 12003 999 12006
rect 1342 12004 1348 12006
rect 1412 12004 1418 12068
rect 2086 12066 2146 12278
rect 2497 12336 2790 12338
rect 2497 12280 2502 12336
rect 2558 12280 2790 12336
rect 2497 12278 2790 12280
rect 2497 12275 2563 12278
rect 2730 12202 2790 12278
rect 3049 12336 3188 12338
rect 3049 12280 3054 12336
rect 3110 12280 3188 12336
rect 3049 12278 3188 12280
rect 3049 12275 3115 12278
rect 3182 12276 3188 12278
rect 3252 12276 3258 12340
rect 4061 12338 4127 12341
rect 6678 12338 6684 12340
rect 4061 12336 6684 12338
rect 4061 12280 4066 12336
rect 4122 12280 6684 12336
rect 4061 12278 6684 12280
rect 4061 12275 4127 12278
rect 6678 12276 6684 12278
rect 6748 12276 6754 12340
rect 7373 12338 7439 12341
rect 8477 12338 8543 12341
rect 7373 12336 8543 12338
rect 7373 12280 7378 12336
rect 7434 12280 8482 12336
rect 8538 12280 8543 12336
rect 7373 12278 8543 12280
rect 7373 12275 7439 12278
rect 8477 12275 8543 12278
rect 11697 12202 11763 12205
rect 2730 12200 11763 12202
rect 2730 12144 11702 12200
rect 11758 12144 11763 12200
rect 2730 12142 11763 12144
rect 11697 12139 11763 12142
rect 2865 12066 2931 12069
rect 2086 12064 2931 12066
rect 2086 12008 2870 12064
rect 2926 12008 2931 12064
rect 2086 12006 2931 12008
rect 2865 12003 2931 12006
rect 6142 12000 6462 12001
rect 0 11930 800 11960
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 11935 6462 11936
rect 11340 12000 11660 12001
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 11935 11660 11936
rect 16538 12000 16858 12001
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 11935 16858 11936
rect 933 11930 999 11933
rect 0 11928 999 11930
rect 0 11872 938 11928
rect 994 11872 999 11928
rect 0 11870 999 11872
rect 0 11840 800 11870
rect 933 11867 999 11870
rect 16389 11794 16455 11797
rect 17166 11794 17172 11796
rect 982 11792 16455 11794
rect 982 11736 16394 11792
rect 16450 11736 16455 11792
rect 982 11734 16455 11736
rect 473 11658 539 11661
rect 982 11658 1042 11734
rect 16389 11731 16455 11734
rect 16530 11734 17172 11794
rect 473 11656 1042 11658
rect 473 11600 478 11656
rect 534 11600 1042 11656
rect 473 11598 1042 11600
rect 2681 11658 2747 11661
rect 3366 11658 3372 11660
rect 2681 11656 3372 11658
rect 2681 11600 2686 11656
rect 2742 11600 3372 11656
rect 2681 11598 3372 11600
rect 473 11595 539 11598
rect 2681 11595 2747 11598
rect 3366 11596 3372 11598
rect 3436 11658 3442 11660
rect 16530 11658 16590 11734
rect 17166 11732 17172 11734
rect 17236 11732 17242 11796
rect 3436 11598 16590 11658
rect 3436 11596 3442 11598
rect 5942 11460 5948 11524
rect 6012 11522 6018 11524
rect 6545 11522 6611 11525
rect 6012 11520 6611 11522
rect 6012 11464 6550 11520
rect 6606 11464 6611 11520
rect 6012 11462 6611 11464
rect 6012 11460 6018 11462
rect 6545 11459 6611 11462
rect 21357 11522 21423 11525
rect 22200 11522 23000 11552
rect 21357 11520 23000 11522
rect 21357 11464 21362 11520
rect 21418 11464 23000 11520
rect 21357 11462 23000 11464
rect 21357 11459 21423 11462
rect 3543 11456 3863 11457
rect 0 11386 800 11416
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 11391 3863 11392
rect 8741 11456 9061 11457
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 11391 9061 11392
rect 13939 11456 14259 11457
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 11391 14259 11392
rect 19137 11456 19457 11457
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 22200 11432 23000 11462
rect 19137 11391 19457 11392
rect 2589 11386 2655 11389
rect 0 11384 2655 11386
rect 0 11328 2594 11384
rect 2650 11328 2655 11384
rect 0 11326 2655 11328
rect 0 11296 800 11326
rect 2589 11323 2655 11326
rect 0 10978 800 11008
rect 4337 10978 4403 10981
rect 0 10976 4403 10978
rect 0 10920 4342 10976
rect 4398 10920 4403 10976
rect 0 10918 4403 10920
rect 0 10888 800 10918
rect 4337 10915 4403 10918
rect 7925 10978 7991 10981
rect 9765 10978 9831 10981
rect 7925 10976 9831 10978
rect 7925 10920 7930 10976
rect 7986 10920 9770 10976
rect 9826 10920 9831 10976
rect 7925 10918 9831 10920
rect 7925 10915 7991 10918
rect 9765 10915 9831 10918
rect 6142 10912 6462 10913
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 10847 6462 10848
rect 11340 10912 11660 10913
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 10847 11660 10848
rect 16538 10912 16858 10913
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 10847 16858 10848
rect 2865 10706 2931 10709
rect 2865 10704 3066 10706
rect 2865 10648 2870 10704
rect 2926 10648 3066 10704
rect 2865 10646 3066 10648
rect 2865 10643 2931 10646
rect 0 10434 800 10464
rect 2681 10434 2747 10437
rect 0 10432 2747 10434
rect 0 10376 2686 10432
rect 2742 10376 2747 10432
rect 0 10374 2747 10376
rect 0 10344 800 10374
rect 2681 10371 2747 10374
rect 3006 10165 3066 10646
rect 4286 10644 4292 10708
rect 4356 10706 4362 10708
rect 4521 10706 4587 10709
rect 4356 10704 4587 10706
rect 4356 10648 4526 10704
rect 4582 10648 4587 10704
rect 4356 10646 4587 10648
rect 4356 10644 4362 10646
rect 4521 10643 4587 10646
rect 5349 10570 5415 10573
rect 16062 10570 16068 10572
rect 5349 10568 16068 10570
rect 5349 10512 5354 10568
rect 5410 10512 16068 10568
rect 5349 10510 16068 10512
rect 5349 10507 5415 10510
rect 16062 10508 16068 10510
rect 16132 10508 16138 10572
rect 3543 10368 3863 10369
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 10303 3863 10304
rect 8741 10368 9061 10369
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8741 10303 9061 10304
rect 13939 10368 14259 10369
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 10303 14259 10304
rect 19137 10368 19457 10369
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 10303 19457 10304
rect 3006 10160 3115 10165
rect 3006 10104 3054 10160
rect 3110 10104 3115 10160
rect 3006 10102 3115 10104
rect 3049 10099 3115 10102
rect 0 10026 800 10056
rect 2497 10026 2563 10029
rect 0 10024 2563 10026
rect 0 9968 2502 10024
rect 2558 9968 2563 10024
rect 0 9966 2563 9968
rect 0 9936 800 9966
rect 2497 9963 2563 9966
rect 6142 9824 6462 9825
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 9759 6462 9760
rect 11340 9824 11660 9825
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 9759 11660 9760
rect 16538 9824 16858 9825
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 9759 16858 9760
rect 2129 9618 2195 9621
rect 4613 9618 4679 9621
rect 2129 9616 4679 9618
rect 2129 9560 2134 9616
rect 2190 9560 4618 9616
rect 4674 9560 4679 9616
rect 2129 9558 4679 9560
rect 2129 9555 2195 9558
rect 4613 9555 4679 9558
rect 6821 9618 6887 9621
rect 7649 9618 7715 9621
rect 9581 9618 9647 9621
rect 6821 9616 9647 9618
rect 6821 9560 6826 9616
rect 6882 9560 7654 9616
rect 7710 9560 9586 9616
rect 9642 9560 9647 9616
rect 6821 9558 9647 9560
rect 6821 9555 6887 9558
rect 7649 9555 7715 9558
rect 9581 9555 9647 9558
rect 0 9482 800 9512
rect 1669 9484 1735 9485
rect 1669 9482 1716 9484
rect 0 9422 1410 9482
rect 1624 9480 1716 9482
rect 1624 9424 1674 9480
rect 1624 9422 1716 9424
rect 0 9392 800 9422
rect 1350 9346 1410 9422
rect 1669 9420 1716 9422
rect 1780 9420 1786 9484
rect 3785 9482 3851 9485
rect 4286 9482 4292 9484
rect 3785 9480 4292 9482
rect 3785 9424 3790 9480
rect 3846 9424 4292 9480
rect 3785 9422 4292 9424
rect 1669 9419 1735 9420
rect 3785 9419 3851 9422
rect 4286 9420 4292 9422
rect 4356 9420 4362 9484
rect 4613 9482 4679 9485
rect 8518 9482 8524 9484
rect 4613 9480 8524 9482
rect 4613 9424 4618 9480
rect 4674 9424 8524 9480
rect 4613 9422 8524 9424
rect 4613 9419 4679 9422
rect 8518 9420 8524 9422
rect 8588 9420 8594 9484
rect 3049 9346 3115 9349
rect 1350 9344 3115 9346
rect 1350 9288 3054 9344
rect 3110 9288 3115 9344
rect 1350 9286 3115 9288
rect 3049 9283 3115 9286
rect 4061 9346 4127 9349
rect 6913 9346 6979 9349
rect 4061 9344 6979 9346
rect 4061 9288 4066 9344
rect 4122 9288 6918 9344
rect 6974 9288 6979 9344
rect 4061 9286 6979 9288
rect 4061 9283 4127 9286
rect 6913 9283 6979 9286
rect 3543 9280 3863 9281
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 9215 3863 9216
rect 8741 9280 9061 9281
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 9215 9061 9216
rect 13939 9280 14259 9281
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 9215 14259 9216
rect 19137 9280 19457 9281
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 9215 19457 9216
rect 0 9074 800 9104
rect 1301 9074 1367 9077
rect 0 9072 1367 9074
rect 0 9016 1306 9072
rect 1362 9016 1367 9072
rect 0 9014 1367 9016
rect 0 8984 800 9014
rect 1301 9011 1367 9014
rect 3325 9074 3391 9077
rect 7373 9074 7439 9077
rect 3325 9072 7439 9074
rect 3325 9016 3330 9072
rect 3386 9016 7378 9072
rect 7434 9016 7439 9072
rect 3325 9014 7439 9016
rect 3325 9011 3391 9014
rect 7373 9011 7439 9014
rect 8201 9074 8267 9077
rect 9305 9074 9371 9077
rect 8201 9072 9371 9074
rect 8201 9016 8206 9072
rect 8262 9016 9310 9072
rect 9366 9016 9371 9072
rect 8201 9014 9371 9016
rect 8201 9011 8267 9014
rect 9305 9011 9371 9014
rect 1577 8938 1643 8941
rect 15009 8938 15075 8941
rect 1577 8936 15075 8938
rect 1577 8880 1582 8936
rect 1638 8880 15014 8936
rect 15070 8880 15075 8936
rect 1577 8878 15075 8880
rect 1577 8875 1643 8878
rect 15009 8875 15075 8878
rect 6142 8736 6462 8737
rect 0 8666 800 8696
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 8671 6462 8672
rect 11340 8736 11660 8737
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 8671 11660 8672
rect 16538 8736 16858 8737
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 8671 16858 8672
rect 2037 8668 2103 8669
rect 2037 8666 2084 8668
rect 0 8606 1594 8666
rect 1992 8664 2084 8666
rect 1992 8608 2042 8664
rect 1992 8606 2084 8608
rect 0 8576 800 8606
rect 1534 8530 1594 8606
rect 2037 8604 2084 8606
rect 2148 8604 2154 8668
rect 2037 8603 2103 8604
rect 3969 8530 4035 8533
rect 1534 8528 4035 8530
rect 1534 8472 3974 8528
rect 4030 8472 4035 8528
rect 1534 8470 4035 8472
rect 3969 8467 4035 8470
rect 2681 8394 2747 8397
rect 7281 8394 7347 8397
rect 2681 8392 7347 8394
rect 2681 8336 2686 8392
rect 2742 8336 7286 8392
rect 7342 8336 7347 8392
rect 2681 8334 7347 8336
rect 2681 8331 2747 8334
rect 7281 8331 7347 8334
rect 10317 8394 10383 8397
rect 16982 8394 16988 8396
rect 10317 8392 16988 8394
rect 10317 8336 10322 8392
rect 10378 8336 16988 8392
rect 10317 8334 16988 8336
rect 10317 8331 10383 8334
rect 16982 8332 16988 8334
rect 17052 8332 17058 8396
rect 1485 8258 1551 8261
rect 2630 8258 2636 8260
rect 1485 8256 2636 8258
rect 1485 8200 1490 8256
rect 1546 8200 2636 8256
rect 1485 8198 2636 8200
rect 1485 8195 1551 8198
rect 2630 8196 2636 8198
rect 2700 8196 2706 8260
rect 3543 8192 3863 8193
rect 0 8122 800 8152
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 8127 3863 8128
rect 8741 8192 9061 8193
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 8127 9061 8128
rect 13939 8192 14259 8193
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 8127 14259 8128
rect 19137 8192 19457 8193
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 8127 19457 8128
rect 2773 8122 2839 8125
rect 0 8120 2839 8122
rect 0 8064 2778 8120
rect 2834 8064 2839 8120
rect 0 8062 2839 8064
rect 0 8032 800 8062
rect 2773 8059 2839 8062
rect 2589 7986 2655 7989
rect 6085 7986 6151 7989
rect 2589 7984 6151 7986
rect 2589 7928 2594 7984
rect 2650 7928 6090 7984
rect 6146 7928 6151 7984
rect 2589 7926 6151 7928
rect 2589 7923 2655 7926
rect 6085 7923 6151 7926
rect 1342 7788 1348 7852
rect 1412 7850 1418 7852
rect 2129 7850 2195 7853
rect 1412 7848 2195 7850
rect 1412 7792 2134 7848
rect 2190 7792 2195 7848
rect 1412 7790 2195 7792
rect 1412 7788 1418 7790
rect 2129 7787 2195 7790
rect 5390 7788 5396 7852
rect 5460 7850 5466 7852
rect 14457 7850 14523 7853
rect 5460 7848 14523 7850
rect 5460 7792 14462 7848
rect 14518 7792 14523 7848
rect 5460 7790 14523 7792
rect 5460 7788 5466 7790
rect 14457 7787 14523 7790
rect 0 7714 800 7744
rect 1342 7714 1348 7716
rect 0 7654 1348 7714
rect 0 7624 800 7654
rect 1342 7652 1348 7654
rect 1412 7652 1418 7716
rect 6142 7648 6462 7649
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 7583 6462 7584
rect 11340 7648 11660 7649
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 7583 11660 7584
rect 16538 7648 16858 7649
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 7583 16858 7584
rect 3417 7578 3483 7581
rect 4838 7578 4844 7580
rect 3417 7576 4844 7578
rect 3417 7520 3422 7576
rect 3478 7520 4844 7576
rect 3417 7518 4844 7520
rect 3417 7515 3483 7518
rect 4838 7516 4844 7518
rect 4908 7516 4914 7580
rect 8477 7442 8543 7445
rect 2730 7440 8543 7442
rect 2730 7384 8482 7440
rect 8538 7384 8543 7440
rect 2730 7382 8543 7384
rect 1577 7306 1643 7309
rect 2730 7306 2790 7382
rect 8477 7379 8543 7382
rect 9857 7306 9923 7309
rect 1577 7304 2790 7306
rect 1577 7248 1582 7304
rect 1638 7248 2790 7304
rect 1577 7246 2790 7248
rect 3374 7304 9923 7306
rect 3374 7248 9862 7304
rect 9918 7248 9923 7304
rect 3374 7246 9923 7248
rect 1577 7243 1643 7246
rect 0 7170 800 7200
rect 2221 7170 2287 7173
rect 0 7168 2287 7170
rect 0 7112 2226 7168
rect 2282 7112 2287 7168
rect 0 7110 2287 7112
rect 0 7080 800 7110
rect 2221 7107 2287 7110
rect 3374 7034 3434 7246
rect 9857 7243 9923 7246
rect 3543 7104 3863 7105
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 7039 3863 7040
rect 8741 7104 9061 7105
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 7039 9061 7040
rect 13939 7104 14259 7105
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 7039 14259 7040
rect 19137 7104 19457 7105
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 7039 19457 7040
rect 3006 6974 3434 7034
rect 3006 6898 3066 6974
rect 2730 6838 3066 6898
rect 0 6762 800 6792
rect 2730 6765 2790 6838
rect 3182 6836 3188 6900
rect 3252 6898 3258 6900
rect 3785 6898 3851 6901
rect 3252 6896 3851 6898
rect 3252 6840 3790 6896
rect 3846 6840 3851 6896
rect 3252 6838 3851 6840
rect 3252 6836 3258 6838
rect 3785 6835 3851 6838
rect 7557 6898 7623 6901
rect 19057 6898 19123 6901
rect 7557 6896 19123 6898
rect 7557 6840 7562 6896
rect 7618 6840 19062 6896
rect 19118 6840 19123 6896
rect 7557 6838 19123 6840
rect 7557 6835 7623 6838
rect 19057 6835 19123 6838
rect 0 6702 1042 6762
rect 0 6672 800 6702
rect 982 6626 1042 6702
rect 1158 6700 1164 6764
rect 1228 6762 1234 6764
rect 2497 6762 2563 6765
rect 1228 6760 2563 6762
rect 1228 6704 2502 6760
rect 2558 6704 2563 6760
rect 1228 6702 2563 6704
rect 1228 6700 1234 6702
rect 2497 6699 2563 6702
rect 2681 6760 2790 6765
rect 2681 6704 2686 6760
rect 2742 6704 2790 6760
rect 2681 6702 2790 6704
rect 3049 6762 3115 6765
rect 19609 6762 19675 6765
rect 3049 6760 19675 6762
rect 3049 6704 3054 6760
rect 3110 6704 19614 6760
rect 19670 6704 19675 6760
rect 3049 6702 19675 6704
rect 2681 6699 2747 6702
rect 3049 6699 3115 6702
rect 19609 6699 19675 6702
rect 19793 6762 19859 6765
rect 19926 6762 19932 6764
rect 19793 6760 19932 6762
rect 19793 6704 19798 6760
rect 19854 6704 19932 6760
rect 19793 6702 19932 6704
rect 19793 6699 19859 6702
rect 19926 6700 19932 6702
rect 19996 6700 20002 6764
rect 1853 6626 1919 6629
rect 982 6624 1919 6626
rect 982 6568 1858 6624
rect 1914 6568 1919 6624
rect 982 6566 1919 6568
rect 1853 6563 1919 6566
rect 2037 6626 2103 6629
rect 5390 6626 5396 6628
rect 2037 6624 5396 6626
rect 2037 6568 2042 6624
rect 2098 6568 5396 6624
rect 2037 6566 5396 6568
rect 2037 6563 2103 6566
rect 5390 6564 5396 6566
rect 5460 6564 5466 6628
rect 6142 6560 6462 6561
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 6495 6462 6496
rect 11340 6560 11660 6561
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 6495 11660 6496
rect 16538 6560 16858 6561
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 6495 16858 6496
rect 2773 6492 2839 6493
rect 2773 6488 2820 6492
rect 2884 6490 2890 6492
rect 3785 6490 3851 6493
rect 3918 6490 3924 6492
rect 2773 6432 2778 6488
rect 2773 6428 2820 6432
rect 2884 6430 2930 6490
rect 3785 6488 3924 6490
rect 3785 6432 3790 6488
rect 3846 6432 3924 6488
rect 3785 6430 3924 6432
rect 2884 6428 2890 6430
rect 2773 6427 2839 6428
rect 3785 6427 3851 6430
rect 3918 6428 3924 6430
rect 3988 6428 3994 6492
rect 1577 6354 1643 6357
rect 15745 6354 15811 6357
rect 1577 6352 15811 6354
rect 1577 6296 1582 6352
rect 1638 6296 15750 6352
rect 15806 6296 15811 6352
rect 1577 6294 15811 6296
rect 1577 6291 1643 6294
rect 15745 6291 15811 6294
rect 0 6218 800 6248
rect 2773 6218 2839 6221
rect 0 6216 2839 6218
rect 0 6160 2778 6216
rect 2834 6160 2839 6216
rect 0 6158 2839 6160
rect 0 6128 800 6158
rect 2773 6155 2839 6158
rect 3417 6218 3483 6221
rect 20069 6218 20135 6221
rect 3417 6216 20135 6218
rect 3417 6160 3422 6216
rect 3478 6160 20074 6216
rect 20130 6160 20135 6216
rect 3417 6158 20135 6160
rect 3417 6155 3483 6158
rect 20069 6155 20135 6158
rect 3325 6084 3391 6085
rect 3325 6082 3372 6084
rect 3280 6080 3372 6082
rect 3280 6024 3330 6080
rect 3280 6022 3372 6024
rect 3325 6020 3372 6022
rect 3436 6020 3442 6084
rect 3325 6019 3391 6020
rect 3543 6016 3863 6017
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3543 5951 3863 5952
rect 8741 6016 9061 6017
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 5951 9061 5952
rect 13939 6016 14259 6017
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 5951 14259 5952
rect 19137 6016 19457 6017
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 5951 19457 5952
rect 974 5884 980 5948
rect 1044 5946 1050 5948
rect 1577 5946 1643 5949
rect 3233 5946 3299 5949
rect 1044 5944 1643 5946
rect 1044 5888 1582 5944
rect 1638 5888 1643 5944
rect 1044 5886 1643 5888
rect 1044 5884 1050 5886
rect 1577 5883 1643 5886
rect 2270 5944 3299 5946
rect 2270 5888 3238 5944
rect 3294 5888 3299 5944
rect 2270 5886 3299 5888
rect 0 5810 800 5840
rect 2270 5810 2330 5886
rect 3233 5883 3299 5886
rect 4286 5884 4292 5948
rect 4356 5946 4362 5948
rect 4613 5946 4679 5949
rect 4981 5948 5047 5949
rect 4981 5946 5028 5948
rect 4356 5944 4679 5946
rect 4356 5888 4618 5944
rect 4674 5888 4679 5944
rect 4356 5886 4679 5888
rect 4936 5944 5028 5946
rect 4936 5888 4986 5944
rect 4936 5886 5028 5888
rect 4356 5884 4362 5886
rect 4613 5883 4679 5886
rect 4981 5884 5028 5886
rect 5092 5884 5098 5948
rect 5349 5946 5415 5949
rect 8293 5946 8359 5949
rect 5349 5944 8359 5946
rect 5349 5888 5354 5944
rect 5410 5888 8298 5944
rect 8354 5888 8359 5944
rect 5349 5886 8359 5888
rect 4981 5883 5047 5884
rect 5349 5883 5415 5886
rect 8293 5883 8359 5886
rect 0 5750 2330 5810
rect 2497 5810 2563 5813
rect 18689 5810 18755 5813
rect 2497 5808 18755 5810
rect 2497 5752 2502 5808
rect 2558 5752 18694 5808
rect 18750 5752 18755 5808
rect 2497 5750 18755 5752
rect 0 5720 800 5750
rect 2497 5747 2563 5750
rect 18689 5747 18755 5750
rect 2037 5674 2103 5677
rect 7557 5674 7623 5677
rect 2037 5672 7623 5674
rect 2037 5616 2042 5672
rect 2098 5616 7562 5672
rect 7618 5616 7623 5672
rect 2037 5614 7623 5616
rect 2037 5611 2103 5614
rect 7557 5611 7623 5614
rect 1025 5538 1091 5541
rect 4613 5538 4679 5541
rect 1025 5536 4679 5538
rect 1025 5480 1030 5536
rect 1086 5480 4618 5536
rect 4674 5480 4679 5536
rect 1025 5478 4679 5480
rect 1025 5475 1091 5478
rect 4613 5475 4679 5478
rect 6142 5472 6462 5473
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 5407 6462 5408
rect 11340 5472 11660 5473
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 5407 11660 5408
rect 16538 5472 16858 5473
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 5407 16858 5408
rect 1301 5404 1367 5405
rect 1301 5402 1348 5404
rect 1256 5400 1348 5402
rect 1256 5344 1306 5400
rect 1256 5342 1348 5344
rect 1301 5340 1348 5342
rect 1412 5340 1418 5404
rect 2037 5402 2103 5405
rect 2037 5400 6010 5402
rect 2037 5344 2042 5400
rect 2098 5344 6010 5400
rect 2037 5342 6010 5344
rect 1301 5339 1367 5340
rect 2037 5339 2103 5342
rect 0 5266 800 5296
rect 1393 5266 1459 5269
rect 0 5264 1459 5266
rect 0 5208 1398 5264
rect 1454 5208 1459 5264
rect 0 5206 1459 5208
rect 0 5176 800 5206
rect 1393 5203 1459 5206
rect 2497 5266 2563 5269
rect 3877 5266 3943 5269
rect 4102 5266 4108 5268
rect 2497 5264 2790 5266
rect 2497 5208 2502 5264
rect 2558 5208 2790 5264
rect 2497 5206 2790 5208
rect 2497 5203 2563 5206
rect 2730 5130 2790 5206
rect 3877 5264 4108 5266
rect 3877 5208 3882 5264
rect 3938 5208 4108 5264
rect 3877 5206 4108 5208
rect 3877 5203 3943 5206
rect 4102 5204 4108 5206
rect 4172 5204 4178 5268
rect 5950 5266 6010 5342
rect 17953 5266 18019 5269
rect 5950 5264 18019 5266
rect 5950 5208 17958 5264
rect 18014 5208 18019 5264
rect 5950 5206 18019 5208
rect 17953 5203 18019 5206
rect 20805 5130 20871 5133
rect 2730 5128 20871 5130
rect 2730 5072 20810 5128
rect 20866 5072 20871 5128
rect 2730 5070 20871 5072
rect 20805 5067 20871 5070
rect 3543 4928 3863 4929
rect 0 4858 800 4888
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 4863 3863 4864
rect 8741 4928 9061 4929
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 4863 9061 4864
rect 13939 4928 14259 4929
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 4863 14259 4864
rect 19137 4928 19457 4929
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 4863 19457 4864
rect 2773 4858 2839 4861
rect 0 4856 2839 4858
rect 0 4800 2778 4856
rect 2834 4800 2839 4856
rect 0 4798 2839 4800
rect 0 4768 800 4798
rect 2773 4795 2839 4798
rect 1577 4722 1643 4725
rect 11053 4722 11119 4725
rect 1577 4720 11119 4722
rect 1577 4664 1582 4720
rect 1638 4664 11058 4720
rect 11114 4664 11119 4720
rect 1577 4662 11119 4664
rect 1577 4659 1643 4662
rect 11053 4659 11119 4662
rect 1577 4586 1643 4589
rect 8293 4586 8359 4589
rect 1577 4584 8359 4586
rect 1577 4528 1582 4584
rect 1638 4528 8298 4584
rect 8354 4528 8359 4584
rect 1577 4526 8359 4528
rect 1577 4523 1643 4526
rect 8293 4523 8359 4526
rect 0 4450 800 4480
rect 1853 4450 1919 4453
rect 0 4448 1919 4450
rect 0 4392 1858 4448
rect 1914 4392 1919 4448
rect 0 4390 1919 4392
rect 0 4360 800 4390
rect 1853 4387 1919 4390
rect 6142 4384 6462 4385
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 4319 6462 4320
rect 11340 4384 11660 4385
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 4319 11660 4320
rect 16538 4384 16858 4385
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 4319 16858 4320
rect 933 4042 999 4045
rect 3233 4042 3299 4045
rect 933 4040 3299 4042
rect 933 3984 938 4040
rect 994 3984 3238 4040
rect 3294 3984 3299 4040
rect 933 3982 3299 3984
rect 933 3979 999 3982
rect 3233 3979 3299 3982
rect 0 3906 800 3936
rect 2221 3906 2287 3909
rect 0 3904 2287 3906
rect 0 3848 2226 3904
rect 2282 3848 2287 3904
rect 0 3846 2287 3848
rect 0 3816 800 3846
rect 2221 3843 2287 3846
rect 3543 3840 3863 3841
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 3775 3863 3776
rect 8741 3840 9061 3841
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 3775 9061 3776
rect 13939 3840 14259 3841
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 3775 14259 3776
rect 19137 3840 19457 3841
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 3775 19457 3776
rect 1945 3634 2011 3637
rect 4521 3634 4587 3637
rect 1945 3632 4587 3634
rect 1945 3576 1950 3632
rect 2006 3576 4526 3632
rect 4582 3576 4587 3632
rect 1945 3574 4587 3576
rect 1945 3571 2011 3574
rect 4521 3571 4587 3574
rect 0 3498 800 3528
rect 2221 3498 2287 3501
rect 0 3496 2287 3498
rect 0 3440 2226 3496
rect 2282 3440 2287 3496
rect 0 3438 2287 3440
rect 0 3408 800 3438
rect 2221 3435 2287 3438
rect 6142 3296 6462 3297
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 3231 6462 3232
rect 11340 3296 11660 3297
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 3231 11660 3232
rect 16538 3296 16858 3297
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 3231 16858 3232
rect 0 2954 800 2984
rect 2773 2954 2839 2957
rect 0 2952 2839 2954
rect 0 2896 2778 2952
rect 2834 2896 2839 2952
rect 0 2894 2839 2896
rect 0 2864 800 2894
rect 2773 2891 2839 2894
rect 3543 2752 3863 2753
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2687 3863 2688
rect 8741 2752 9061 2753
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2687 9061 2688
rect 13939 2752 14259 2753
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2687 14259 2688
rect 19137 2752 19457 2753
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2687 19457 2688
rect 0 2546 800 2576
rect 2773 2546 2839 2549
rect 0 2544 2839 2546
rect 0 2488 2778 2544
rect 2834 2488 2839 2544
rect 0 2486 2839 2488
rect 0 2456 800 2486
rect 2773 2483 2839 2486
rect 6142 2208 6462 2209
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2143 6462 2144
rect 11340 2208 11660 2209
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2143 11660 2144
rect 16538 2208 16858 2209
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2143 16858 2144
rect 0 2002 800 2032
rect 3049 2002 3115 2005
rect 0 2000 3115 2002
rect 0 1944 3054 2000
rect 3110 1944 3115 2000
rect 0 1942 3115 1944
rect 0 1912 800 1942
rect 3049 1939 3115 1942
rect 0 1594 800 1624
rect 3969 1594 4035 1597
rect 0 1592 4035 1594
rect 0 1536 3974 1592
rect 4030 1536 4035 1592
rect 0 1534 4035 1536
rect 0 1504 800 1534
rect 3969 1531 4035 1534
rect 0 1050 800 1080
rect 3233 1050 3299 1053
rect 0 1048 3299 1050
rect 0 992 3238 1048
rect 3294 992 3299 1048
rect 0 990 3299 992
rect 0 960 800 990
rect 3233 987 3299 990
rect 0 642 800 672
rect 2865 642 2931 645
rect 0 640 2931 642
rect 0 584 2870 640
rect 2926 584 2931 640
rect 0 582 2931 584
rect 0 552 800 582
rect 2865 579 2931 582
rect 0 234 800 264
rect 2773 234 2839 237
rect 0 232 2839 234
rect 0 176 2778 232
rect 2834 176 2839 232
rect 0 174 2839 176
rect 0 144 800 174
rect 2773 171 2839 174
<< via3 >>
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 8524 20300 8588 20364
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 5028 19348 5092 19412
rect 6684 19348 6748 19412
rect 15148 19348 15212 19412
rect 16068 19408 16132 19412
rect 16068 19352 16082 19408
rect 16082 19352 16132 19408
rect 16068 19348 16132 19352
rect 16988 19408 17052 19412
rect 16988 19352 17002 19408
rect 17002 19352 17052 19408
rect 16988 19348 17052 19352
rect 19932 19348 19996 19412
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 4476 18804 4540 18868
rect 5948 18804 6012 18868
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 4292 18124 4356 18188
rect 4844 17988 4908 18052
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 17172 18124 17236 18188
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 5948 17504 6012 17508
rect 5948 17448 5962 17504
rect 5962 17448 6012 17504
rect 5948 17444 6012 17448
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 5948 16492 6012 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 1716 15328 1780 15332
rect 1716 15272 1766 15328
rect 1766 15272 1780 15328
rect 1716 15268 1780 15272
rect 2084 15328 2148 15332
rect 2084 15272 2134 15328
rect 2134 15272 2148 15328
rect 2084 15268 2148 15272
rect 19748 15268 19812 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 1164 14996 1228 15060
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 980 14316 1044 14380
rect 3924 14180 3988 14244
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 2636 13636 2700 13700
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 4476 13500 4540 13564
rect 4108 13364 4172 13428
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 15148 12684 15212 12748
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 1348 12004 1412 12068
rect 3188 12276 3252 12340
rect 6684 12276 6748 12340
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 3372 11596 3436 11660
rect 17172 11732 17236 11796
rect 5948 11460 6012 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 4292 10644 4356 10708
rect 16068 10508 16132 10572
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 1716 9480 1780 9484
rect 1716 9424 1730 9480
rect 1730 9424 1780 9480
rect 1716 9420 1780 9424
rect 4292 9420 4356 9484
rect 8524 9420 8588 9484
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 2084 8664 2148 8668
rect 2084 8608 2098 8664
rect 2098 8608 2148 8664
rect 2084 8604 2148 8608
rect 16988 8332 17052 8396
rect 2636 8196 2700 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 1348 7788 1412 7852
rect 5396 7788 5460 7852
rect 1348 7652 1412 7716
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 4844 7516 4908 7580
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 3188 6836 3252 6900
rect 1164 6700 1228 6764
rect 19932 6700 19996 6764
rect 5396 6564 5460 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 2820 6488 2884 6492
rect 2820 6432 2834 6488
rect 2834 6432 2884 6488
rect 2820 6428 2884 6432
rect 3924 6428 3988 6492
rect 3372 6080 3436 6084
rect 3372 6024 3386 6080
rect 3386 6024 3436 6080
rect 3372 6020 3436 6024
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 980 5884 1044 5948
rect 4292 5884 4356 5948
rect 5028 5944 5092 5948
rect 5028 5888 5042 5944
rect 5042 5888 5092 5944
rect 5028 5884 5092 5888
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 1348 5400 1412 5404
rect 1348 5344 1362 5400
rect 1362 5344 1412 5400
rect 1348 5340 1412 5344
rect 4108 5204 4172 5268
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
<< metal4 >>
rect 3543 20160 3863 20720
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3543 19072 3863 20096
rect 6142 20704 6462 20720
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 8523 20364 8589 20365
rect 8523 20300 8524 20364
rect 8588 20300 8589 20364
rect 8523 20299 8589 20300
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 5027 19412 5093 19413
rect 5027 19348 5028 19412
rect 5092 19348 5093 19412
rect 5027 19347 5093 19348
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3543 17984 3863 19008
rect 4475 18868 4541 18869
rect 4475 18804 4476 18868
rect 4540 18804 4541 18868
rect 4475 18803 4541 18804
rect 4291 18188 4357 18189
rect 4291 18124 4292 18188
rect 4356 18124 4357 18188
rect 4291 18123 4357 18124
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3543 16896 3863 17920
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 1715 15332 1781 15333
rect 1715 15268 1716 15332
rect 1780 15268 1781 15332
rect 1715 15267 1781 15268
rect 2083 15332 2149 15333
rect 2083 15268 2084 15332
rect 2148 15268 2149 15332
rect 2083 15267 2149 15268
rect 1163 15060 1229 15061
rect 1163 14996 1164 15060
rect 1228 14996 1229 15060
rect 1163 14995 1229 14996
rect 979 14380 1045 14381
rect 979 14316 980 14380
rect 1044 14316 1045 14380
rect 979 14315 1045 14316
rect 982 5949 1042 14315
rect 1166 6765 1226 14995
rect 1347 12068 1413 12069
rect 1347 12004 1348 12068
rect 1412 12004 1413 12068
rect 1347 12003 1413 12004
rect 1350 7853 1410 12003
rect 1718 9485 1778 15267
rect 1715 9484 1781 9485
rect 1715 9420 1716 9484
rect 1780 9420 1781 9484
rect 1715 9419 1781 9420
rect 2086 8669 2146 15267
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 2635 13700 2701 13701
rect 2635 13636 2636 13700
rect 2700 13636 2701 13700
rect 2635 13635 2701 13636
rect 2083 8668 2149 8669
rect 2083 8604 2084 8668
rect 2148 8604 2149 8668
rect 2083 8603 2149 8604
rect 2638 8261 2698 13635
rect 3543 13632 3863 14656
rect 3923 14244 3989 14245
rect 3923 14180 3924 14244
rect 3988 14180 3989 14244
rect 3923 14179 3989 14180
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3187 12340 3253 12341
rect 3187 12276 3188 12340
rect 3252 12276 3253 12340
rect 3187 12275 3253 12276
rect 2635 8260 2701 8261
rect 2635 8196 2636 8260
rect 2700 8196 2701 8260
rect 2635 8195 2701 8196
rect 1347 7852 1413 7853
rect 1347 7788 1348 7852
rect 1412 7788 1413 7852
rect 1347 7787 1413 7788
rect 1347 7716 1413 7717
rect 1347 7652 1348 7716
rect 1412 7652 1413 7716
rect 1347 7651 1413 7652
rect 1163 6764 1229 6765
rect 1163 6700 1164 6764
rect 1228 6700 1229 6764
rect 1163 6699 1229 6700
rect 979 5948 1045 5949
rect 979 5884 980 5948
rect 1044 5884 1045 5948
rect 979 5883 1045 5884
rect 1350 5405 1410 7651
rect 3190 6901 3250 12275
rect 3371 11660 3437 11661
rect 3371 11596 3372 11660
rect 3436 11596 3437 11660
rect 3371 11595 3437 11596
rect 3187 6900 3253 6901
rect 3187 6836 3188 6900
rect 3252 6836 3253 6900
rect 3187 6835 3253 6836
rect 3374 6085 3434 11595
rect 3543 11456 3863 12480
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3543 8192 3863 9216
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3371 6084 3437 6085
rect 3371 6020 3372 6084
rect 3436 6020 3437 6084
rect 3371 6019 3437 6020
rect 3543 6016 3863 7040
rect 3926 6493 3986 14179
rect 4107 13428 4173 13429
rect 4107 13364 4108 13428
rect 4172 13364 4173 13428
rect 4107 13363 4173 13364
rect 3923 6492 3989 6493
rect 3923 6428 3924 6492
rect 3988 6428 3989 6492
rect 3923 6427 3989 6428
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 1347 5404 1413 5405
rect 1347 5340 1348 5404
rect 1412 5340 1413 5404
rect 1347 5339 1413 5340
rect 3543 4928 3863 5952
rect 4110 5269 4170 13363
rect 4294 10709 4354 18123
rect 4478 13565 4538 18803
rect 4843 18052 4909 18053
rect 4843 17988 4844 18052
rect 4908 17988 4909 18052
rect 4843 17987 4909 17988
rect 4475 13564 4541 13565
rect 4475 13500 4476 13564
rect 4540 13500 4541 13564
rect 4475 13499 4541 13500
rect 4291 10708 4357 10709
rect 4291 10644 4292 10708
rect 4356 10644 4357 10708
rect 4291 10643 4357 10644
rect 4291 9484 4357 9485
rect 4291 9420 4292 9484
rect 4356 9420 4357 9484
rect 4291 9419 4357 9420
rect 4294 5949 4354 9419
rect 4846 7581 4906 17987
rect 4843 7580 4909 7581
rect 4843 7516 4844 7580
rect 4908 7516 4909 7580
rect 4843 7515 4909 7516
rect 5030 5949 5090 19347
rect 5947 18868 6013 18869
rect 5947 18804 5948 18868
rect 6012 18804 6013 18868
rect 5947 18803 6013 18804
rect 5950 17509 6010 18803
rect 6142 18528 6462 19552
rect 6683 19412 6749 19413
rect 6683 19348 6684 19412
rect 6748 19348 6749 19412
rect 6683 19347 6749 19348
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 5947 17508 6013 17509
rect 5947 17444 5948 17508
rect 6012 17444 6013 17508
rect 5947 17443 6013 17444
rect 5950 16557 6010 17443
rect 6142 17440 6462 18464
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 5947 16556 6013 16557
rect 5947 16492 5948 16556
rect 6012 16492 6013 16556
rect 5947 16491 6013 16492
rect 5950 11525 6010 16491
rect 6142 16352 6462 17376
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6686 12341 6746 19347
rect 6683 12340 6749 12341
rect 6683 12276 6684 12340
rect 6748 12276 6749 12340
rect 6683 12275 6749 12276
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 5947 11524 6013 11525
rect 5947 11460 5948 11524
rect 6012 11460 6013 11524
rect 5947 11459 6013 11460
rect 6142 10912 6462 11936
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 8526 9485 8586 20299
rect 8741 20160 9061 20720
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8523 9484 8589 9485
rect 8523 9420 8524 9484
rect 8588 9420 8589 9484
rect 8523 9419 8589 9420
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 5395 7852 5461 7853
rect 5395 7788 5396 7852
rect 5460 7788 5461 7852
rect 5395 7787 5461 7788
rect 5398 6629 5458 7787
rect 6142 7648 6462 8672
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 5395 6628 5461 6629
rect 5395 6564 5396 6628
rect 5460 6564 5461 6628
rect 5395 6563 5461 6564
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 4291 5948 4357 5949
rect 4291 5884 4292 5948
rect 4356 5884 4357 5948
rect 4291 5883 4357 5884
rect 5027 5948 5093 5949
rect 5027 5884 5028 5948
rect 5092 5884 5093 5948
rect 5027 5883 5093 5884
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 4107 5268 4173 5269
rect 4107 5204 4108 5268
rect 4172 5204 4173 5268
rect 4107 5203 4173 5204
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 3543 2128 3863 2688
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 6142 2208 6462 3232
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 6142 2128 6462 2144
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8741 2752 9061 3776
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 2128 9061 2688
rect 11340 20704 11660 20720
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11340 12000 11660 13024
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 11340 2208 11660 3232
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 11340 2128 11660 2144
rect 13939 20160 14259 20720
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 16538 20704 16858 20720
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 16067 19412 16133 19413
rect 16067 19348 16068 19412
rect 16132 19348 16133 19412
rect 16067 19347 16133 19348
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13939 16896 14259 17920
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 15150 12749 15210 19347
rect 15147 12748 15213 12749
rect 15147 12684 15148 12748
rect 15212 12684 15213 12748
rect 15147 12683 15213 12684
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 16070 10573 16130 19347
rect 16538 18528 16858 19552
rect 19137 20160 19457 20720
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 16987 19412 17053 19413
rect 16987 19348 16988 19412
rect 17052 19348 17053 19412
rect 16987 19347 17053 19348
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16538 17440 16858 18464
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16538 10912 16858 11936
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16067 10572 16133 10573
rect 16067 10508 16068 10572
rect 16132 10508 16133 10572
rect 16067 10507 16133 10508
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 13939 6016 14259 7040
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 13939 3840 14259 4864
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 13939 2752 14259 3776
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 2128 14259 2688
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16538 8736 16858 9760
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16990 8397 17050 19347
rect 19137 19072 19457 20096
rect 19931 19412 19997 19413
rect 19931 19348 19932 19412
rect 19996 19348 19997 19412
rect 19931 19347 19997 19348
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 17171 18188 17237 18189
rect 17171 18124 17172 18188
rect 17236 18124 17237 18188
rect 17171 18123 17237 18124
rect 17174 11797 17234 18123
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19747 15332 19813 15333
rect 19747 15268 19748 15332
rect 19812 15268 19813 15332
rect 19747 15267 19813 15268
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 17171 11796 17237 11797
rect 17171 11732 17172 11796
rect 17236 11732 17237 11796
rect 17171 11731 17237 11732
rect 19137 11456 19457 12480
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19137 9280 19457 10304
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 16987 8396 17053 8397
rect 16987 8332 16988 8396
rect 17052 8332 17053 8396
rect 16987 8331 17053 8332
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 2128 16858 2144
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19750 6578 19810 15267
rect 19934 6765 19994 19347
rect 19931 6764 19997 6765
rect 19931 6700 19932 6764
rect 19996 6700 19997 6764
rect 19931 6699 19997 6700
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 2128 19457 2688
<< via4 >>
rect 2734 6492 2970 6578
rect 2734 6428 2820 6492
rect 2820 6428 2884 6492
rect 2884 6428 2970 6492
rect 2734 6342 2970 6428
rect 19662 6342 19898 6578
<< metal5 >>
rect 2692 6578 19940 6620
rect 2692 6342 2734 6578
rect 2970 6342 19662 6578
rect 19898 6342 19940 6578
rect 2692 6300 19940 6342
use sky130_fd_sc_hd__diode_2  ANTENNA__077__A .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 3404 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1649977179
transform -1 0 19412 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A
timestamp 1649977179
transform -1 0 19872 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1649977179
transform -1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A
timestamp 1649977179
transform -1 0 20976 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 5060 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 6532 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 5888 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 4140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 4876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 5796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5980 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 20332 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 20792 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 21068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 20424 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 2484 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 5060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 3312 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 4140 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_1.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 2760 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 5888 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5060 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_3.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 10304 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 8280 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 7912 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_5.mux_l1_in_2__A1
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11408 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10856 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_7.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_11.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_13.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9016 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_15.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_17.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_19.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 11132 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_21.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_27.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_29.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_31.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_33.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 5244 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_35.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 3496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_37.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 4048 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_left_track_39.mux_l2_in_0__S
timestamp 1649977179
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16744 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 14260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_0.mux_l1_in_2__A0
timestamp 1649977179
transform -1 0 14260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 20792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 20240 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 21160 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_2.mux_l2_in_1__A1
timestamp 1649977179
transform -1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 9936 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 17572 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_4.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 10580 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 8464 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A0
timestamp 1649977179
transform 1 0 5888 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_6.mux_l1_in_1__A1
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_8.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_10.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 10120 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_12.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 15088 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 16836 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_14.mux_l1_in_0__A1
timestamp 1649977179
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 16928 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_16.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 16836 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_18.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 17848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_20.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 21160 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A0
timestamp 1649977179
transform -1 0 21160 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_22.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 18676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_24.mux_l1_in_1__A1
timestamp 1649977179
transform -1 0 19228 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A0
timestamp 1649977179
transform 1 0 15548 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_mux_top_track_26.mux_l1_in_0__A1
timestamp 1649977179
transform -1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output60_A
timestamp 1649977179
transform -1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_prog_clk_0_FTB00_A
timestamp 1649977179
transform -1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 1649977179
transform 1 0 4324 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39
timestamp 1649977179
transform 1 0 4692 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_118
timestamp 1649977179
transform 1 0 11960 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_122
timestamp 1649977179
transform 1 0 12328 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 1649977179
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_13
timestamp 1649977179
transform 1 0 2300 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_19
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_23
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_27
timestamp 1649977179
transform 1 0 3588 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_31
timestamp 1649977179
transform 1 0 3956 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_35
timestamp 1649977179
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1649977179
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_19
timestamp 1649977179
transform 1 0 2852 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_23
timestamp 1649977179
transform 1 0 3220 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_31
timestamp 1649977179
transform 1 0 3956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_35
timestamp 1649977179
transform 1 0 4324 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_39
timestamp 1649977179
transform 1 0 4692 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_63
timestamp 1649977179
transform 1 0 6900 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_75 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8004 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_17
timestamp 1649977179
transform 1 0 2668 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_21
timestamp 1649977179
transform 1 0 3036 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_25
timestamp 1649977179
transform 1 0 3404 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 1649977179
transform 1 0 4140 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37
timestamp 1649977179
transform 1 0 4508 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_4_6
timestamp 1649977179
transform 1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_11
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_20
timestamp 1649977179
transform 1 0 2944 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1649977179
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_35
timestamp 1649977179
transform 1 0 4324 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_39
timestamp 1649977179
transform 1 0 4692 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_43
timestamp 1649977179
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_55
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_6
timestamp 1649977179
transform 1 0 1656 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_11
timestamp 1649977179
transform 1 0 2116 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_16
timestamp 1649977179
transform 1 0 2576 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_20
timestamp 1649977179
transform 1 0 2944 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_24
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_28
timestamp 1649977179
transform 1 0 3680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_32
timestamp 1649977179
transform 1 0 4048 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_40
timestamp 1649977179
transform 1 0 4784 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_44
timestamp 1649977179
transform 1 0 5152 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_213
timestamp 1649977179
transform 1 0 20700 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_216
timestamp 1649977179
transform 1 0 20976 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_222
timestamp 1649977179
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 1649977179
transform 1 0 1656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_11
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_16
timestamp 1649977179
transform 1 0 2576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_21
timestamp 1649977179
transform 1 0 3036 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_25
timestamp 1649977179
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_31
timestamp 1649977179
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_35
timestamp 1649977179
transform 1 0 4324 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_39
timestamp 1649977179
transform 1 0 4692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_43
timestamp 1649977179
transform 1 0 5060 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_47
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_51
timestamp 1649977179
transform 1 0 5796 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_55
timestamp 1649977179
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_59
timestamp 1649977179
transform 1 0 6532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_71
timestamp 1649977179
transform 1 0 7636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_205
timestamp 1649977179
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_214
timestamp 1649977179
transform 1 0 20792 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1649977179
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_6
timestamp 1649977179
transform 1 0 1656 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_11
timestamp 1649977179
transform 1 0 2116 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_16
timestamp 1649977179
transform 1 0 2576 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_21
timestamp 1649977179
transform 1 0 3036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_26
timestamp 1649977179
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_30
timestamp 1649977179
transform 1 0 3864 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_34
timestamp 1649977179
transform 1 0 4232 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_38
timestamp 1649977179
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_41
timestamp 1649977179
transform 1 0 4876 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_7_45
timestamp 1649977179
transform 1 0 5244 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_52
timestamp 1649977179
transform 1 0 5888 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1649977179
transform 1 0 6532 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_63
timestamp 1649977179
transform 1 0 6900 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_71
timestamp 1649977179
transform 1 0 7636 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_76
timestamp 1649977179
transform 1 0 8096 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_92
timestamp 1649977179
transform 1 0 9568 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_104
timestamp 1649977179
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_209
timestamp 1649977179
transform 1 0 20332 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_221
timestamp 1649977179
transform 1 0 21436 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_6
timestamp 1649977179
transform 1 0 1656 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_11
timestamp 1649977179
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_16
timestamp 1649977179
transform 1 0 2576 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_21
timestamp 1649977179
transform 1 0 3036 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 1649977179
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_31
timestamp 1649977179
transform 1 0 3956 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_42
timestamp 1649977179
transform 1 0 4968 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_46
timestamp 1649977179
transform 1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_56
timestamp 1649977179
transform 1 0 6256 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_60
timestamp 1649977179
transform 1 0 6624 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_63
timestamp 1649977179
transform 1 0 6900 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_87
timestamp 1649977179
transform 1 0 9108 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_99
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_111
timestamp 1649977179
transform 1 0 11316 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_123
timestamp 1649977179
transform 1 0 12420 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1649977179
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_204
timestamp 1649977179
transform 1 0 19872 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_216
timestamp 1649977179
transform 1 0 20976 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_222
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_13
timestamp 1649977179
transform 1 0 2300 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_18
timestamp 1649977179
transform 1 0 2760 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_22
timestamp 1649977179
transform 1 0 3128 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_26
timestamp 1649977179
transform 1 0 3496 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_31
timestamp 1649977179
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_49
timestamp 1649977179
transform 1 0 5612 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_53
timestamp 1649977179
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_73
timestamp 1649977179
transform 1 0 7820 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_85
timestamp 1649977179
transform 1 0 8924 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_96
timestamp 1649977179
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_100
timestamp 1649977179
transform 1 0 10304 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_200
timestamp 1649977179
transform 1 0 19504 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_9_204
timestamp 1649977179
transform 1 0 19872 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_216
timestamp 1649977179
transform 1 0 20976 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_222
timestamp 1649977179
transform 1 0 21528 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_5
timestamp 1649977179
transform 1 0 1564 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_10
timestamp 1649977179
transform 1 0 2024 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_26
timestamp 1649977179
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_32
timestamp 1649977179
transform 1 0 4048 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_43
timestamp 1649977179
transform 1 0 5060 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_61
timestamp 1649977179
transform 1 0 6716 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_82
timestamp 1649977179
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_94
timestamp 1649977179
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_104
timestamp 1649977179
transform 1 0 10672 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_116
timestamp 1649977179
transform 1 0 11776 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_128
timestamp 1649977179
transform 1 0 12880 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_194
timestamp 1649977179
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_199
timestamp 1649977179
transform 1 0 19412 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_211
timestamp 1649977179
transform 1 0 20516 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_6
timestamp 1649977179
transform 1 0 1656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1649977179
transform 1 0 2116 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_16
timestamp 1649977179
transform 1 0 2576 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_21
timestamp 1649977179
transform 1 0 3036 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 1649977179
transform 1 0 6072 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_60
timestamp 1649977179
transform 1 0 6624 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_11_73
timestamp 1649977179
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_91
timestamp 1649977179
transform 1 0 9476 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_101
timestamp 1649977179
transform 1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_109
timestamp 1649977179
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_6
timestamp 1649977179
transform 1 0 1656 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_12_26
timestamp 1649977179
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_32
timestamp 1649977179
transform 1 0 4048 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_43
timestamp 1649977179
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_54
timestamp 1649977179
transform 1 0 6072 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_76
timestamp 1649977179
transform 1 0 8096 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_81
timestamp 1649977179
transform 1 0 8556 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_94
timestamp 1649977179
transform 1 0 9752 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_104
timestamp 1649977179
transform 1 0 10672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_108
timestamp 1649977179
transform 1 0 11040 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_112
timestamp 1649977179
transform 1 0 11408 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_124
timestamp 1649977179
transform 1 0 12512 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_136
timestamp 1649977179
transform 1 0 13616 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1649977179
transform 1 0 1748 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_17
timestamp 1649977179
transform 1 0 2668 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_29
timestamp 1649977179
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_34
timestamp 1649977179
transform 1 0 4232 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_50
timestamp 1649977179
transform 1 0 5704 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_54
timestamp 1649977179
transform 1 0 6072 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_63
timestamp 1649977179
transform 1 0 6900 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_101
timestamp 1649977179
transform 1 0 10396 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_109
timestamp 1649977179
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_129
timestamp 1649977179
transform 1 0 12972 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_139
timestamp 1649977179
transform 1 0 13892 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 1649977179
transform 1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_155
timestamp 1649977179
transform 1 0 15364 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_159
timestamp 1649977179
transform 1 0 15732 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_14_6
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_38
timestamp 1649977179
transform 1 0 4600 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 1649977179
transform 1 0 5060 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 1649977179
transform 1 0 8648 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_94
timestamp 1649977179
transform 1 0 9752 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_98
timestamp 1649977179
transform 1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_132
timestamp 1649977179
transform 1 0 13248 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_147
timestamp 1649977179
transform 1 0 14628 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_156
timestamp 1649977179
transform 1 0 15456 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_178
timestamp 1649977179
transform 1 0 17480 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_188
timestamp 1649977179
transform 1 0 18400 0 1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_33
timestamp 1649977179
transform 1 0 4140 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_44
timestamp 1649977179
transform 1 0 5152 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_54
timestamp 1649977179
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_60
timestamp 1649977179
transform 1 0 6624 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_71
timestamp 1649977179
transform 1 0 7636 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_97
timestamp 1649977179
transform 1 0 10028 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_100
timestamp 1649977179
transform 1 0 10304 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_110
timestamp 1649977179
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_126
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_144
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1649977179
transform 1 0 15364 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 1649977179
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_185
timestamp 1649977179
transform 1 0 18124 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_197
timestamp 1649977179
transform 1 0 19228 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_209
timestamp 1649977179
transform 1 0 20332 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_221
timestamp 1649977179
transform 1 0 21436 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 1649977179
transform 1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_33
timestamp 1649977179
transform 1 0 4140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_44
timestamp 1649977179
transform 1 0 5152 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_55
timestamp 1649977179
transform 1 0 6164 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_73
timestamp 1649977179
transform 1 0 7820 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_78
timestamp 1649977179
transform 1 0 8280 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_82
timestamp 1649977179
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_94
timestamp 1649977179
transform 1 0 9752 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_16_114
timestamp 1649977179
transform 1 0 11592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_138
timestamp 1649977179
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_150
timestamp 1649977179
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_154
timestamp 1649977179
transform 1 0 15272 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_16_174
timestamp 1649977179
transform 1 0 17112 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_185
timestamp 1649977179
transform 1 0 18124 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_16_190
timestamp 1649977179
transform 1 0 18584 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_6
timestamp 1649977179
transform 1 0 1656 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_11
timestamp 1649977179
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_16
timestamp 1649977179
transform 1 0 2576 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_21
timestamp 1649977179
transform 1 0 3036 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_26
timestamp 1649977179
transform 1 0 3496 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_44
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1649977179
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_66
timestamp 1649977179
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_84
timestamp 1649977179
transform 1 0 8832 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_88
timestamp 1649977179
transform 1 0 9200 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_99
timestamp 1649977179
transform 1 0 10212 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 1649977179
transform 1 0 11224 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_135
timestamp 1649977179
transform 1 0 13524 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_164
timestamp 1649977179
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_171
timestamp 1649977179
transform 1 0 16836 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 1649977179
transform 1 0 17204 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_192
timestamp 1649977179
transform 1 0 18768 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_17_202
timestamp 1649977179
transform 1 0 19688 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_216
timestamp 1649977179
transform 1 0 20976 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_221
timestamp 1649977179
transform 1 0 21436 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 1649977179
transform 1 0 1656 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_11
timestamp 1649977179
transform 1 0 2116 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_16
timestamp 1649977179
transform 1 0 2576 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_21
timestamp 1649977179
transform 1 0 3036 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_26
timestamp 1649977179
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1649977179
transform 1 0 4048 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_52
timestamp 1649977179
transform 1 0 5888 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_70
timestamp 1649977179
transform 1 0 7544 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_81
timestamp 1649977179
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_89
timestamp 1649977179
transform 1 0 9292 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1649977179
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_110
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1649977179
transform 1 0 12972 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_138
timestamp 1649977179
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_160
timestamp 1649977179
transform 1 0 15824 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_170
timestamp 1649977179
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_187
timestamp 1649977179
transform 1 0 18308 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_191
timestamp 1649977179
transform 1 0 18676 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_206
timestamp 1649977179
transform 1 0 20056 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_218
timestamp 1649977179
transform 1 0 21160 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_222
timestamp 1649977179
transform 1 0 21528 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_12
timestamp 1649977179
transform 1 0 2208 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_17
timestamp 1649977179
transform 1 0 2668 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_22
timestamp 1649977179
transform 1 0 3128 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_32
timestamp 1649977179
transform 1 0 4048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1649977179
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_65
timestamp 1649977179
transform 1 0 7084 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_83
timestamp 1649977179
transform 1 0 8740 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1649977179
transform 1 0 10396 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_110
timestamp 1649977179
transform 1 0 11224 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_139
timestamp 1649977179
transform 1 0 13892 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_143
timestamp 1649977179
transform 1 0 14260 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 1649977179
transform 1 0 15640 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_163
timestamp 1649977179
transform 1 0 16100 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_171
timestamp 1649977179
transform 1 0 16836 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_175
timestamp 1649977179
transform 1 0 17204 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_192
timestamp 1649977179
transform 1 0 18768 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_197
timestamp 1649977179
transform 1 0 19228 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_221
timestamp 1649977179
transform 1 0 21436 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_6
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_11
timestamp 1649977179
transform 1 0 2116 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_16
timestamp 1649977179
transform 1 0 2576 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_33
timestamp 1649977179
transform 1 0 4140 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_51
timestamp 1649977179
transform 1 0 5796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_62
timestamp 1649977179
transform 1 0 6808 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_72
timestamp 1649977179
transform 1 0 7728 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_82
timestamp 1649977179
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_89
timestamp 1649977179
transform 1 0 9292 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_99
timestamp 1649977179
transform 1 0 10212 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_126
timestamp 1649977179
transform 1 0 12696 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 1649977179
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_143
timestamp 1649977179
transform 1 0 14260 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 1649977179
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_164
timestamp 1649977179
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_174
timestamp 1649977179
transform 1 0 17112 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_186
timestamp 1649977179
transform 1 0 18216 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_191
timestamp 1649977179
transform 1 0 18676 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_205
timestamp 1649977179
transform 1 0 19964 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_217
timestamp 1649977179
transform 1 0 21068 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_7
timestamp 1649977179
transform 1 0 1748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_21_14
timestamp 1649977179
transform 1 0 2392 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_19
timestamp 1649977179
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_24
timestamp 1649977179
transform 1 0 3312 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_35
timestamp 1649977179
transform 1 0 4324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_60
timestamp 1649977179
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_72
timestamp 1649977179
transform 1 0 7728 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_83
timestamp 1649977179
transform 1 0 8740 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_101
timestamp 1649977179
transform 1 0 10396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_106
timestamp 1649977179
transform 1 0 10856 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1649977179
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_122
timestamp 1649977179
transform 1 0 12328 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_127
timestamp 1649977179
transform 1 0 12788 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_145
timestamp 1649977179
transform 1 0 14444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_178
timestamp 1649977179
transform 1 0 17480 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_196
timestamp 1649977179
transform 1 0 19136 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_206
timestamp 1649977179
transform 1 0 20056 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_210
timestamp 1649977179
transform 1 0 20424 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_214
timestamp 1649977179
transform 1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_218
timestamp 1649977179
transform 1 0 21160 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_221
timestamp 1649977179
transform 1 0 21436 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_26
timestamp 1649977179
transform 1 0 3496 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_45
timestamp 1649977179
transform 1 0 5244 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_55
timestamp 1649977179
transform 1 0 6164 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_73
timestamp 1649977179
transform 1 0 7820 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_78
timestamp 1649977179
transform 1 0 8280 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 1649977179
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_96
timestamp 1649977179
transform 1 0 9936 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_114
timestamp 1649977179
transform 1 0 11592 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_136
timestamp 1649977179
transform 1 0 13616 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_150
timestamp 1649977179
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_155
timestamp 1649977179
transform 1 0 15364 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_22_175
timestamp 1649977179
transform 1 0 17204 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_186
timestamp 1649977179
transform 1 0 18216 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1649977179
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_205
timestamp 1649977179
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_213
timestamp 1649977179
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_217
timestamp 1649977179
transform 1 0 21068 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_7
timestamp 1649977179
transform 1 0 1748 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_13
timestamp 1649977179
transform 1 0 2300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_17
timestamp 1649977179
transform 1 0 2668 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_34
timestamp 1649977179
transform 1 0 4232 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_23_54
timestamp 1649977179
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_60
timestamp 1649977179
transform 1 0 6624 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_64
timestamp 1649977179
transform 1 0 6992 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_98
timestamp 1649977179
transform 1 0 10120 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_110
timestamp 1649977179
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_122
timestamp 1649977179
transform 1 0 12328 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_127
timestamp 1649977179
transform 1 0 12788 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_139
timestamp 1649977179
transform 1 0 13892 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1649977179
transform 1 0 15548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_165
timestamp 1649977179
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_178
timestamp 1649977179
transform 1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_182
timestamp 1649977179
transform 1 0 17848 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 1649977179
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_210
timestamp 1649977179
transform 1 0 20424 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_214
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_218
timestamp 1649977179
transform 1 0 21160 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_7
timestamp 1649977179
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_13
timestamp 1649977179
transform 1 0 2300 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_19
timestamp 1649977179
transform 1 0 2852 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_33
timestamp 1649977179
transform 1 0 4140 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_43
timestamp 1649977179
transform 1 0 5060 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_76
timestamp 1649977179
transform 1 0 8096 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 1649977179
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_101
timestamp 1649977179
transform 1 0 10396 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_108
timestamp 1649977179
transform 1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_120
timestamp 1649977179
transform 1 0 12144 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_125
timestamp 1649977179
transform 1 0 12604 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 1649977179
transform 1 0 13800 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_152
timestamp 1649977179
transform 1 0 15088 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_156
timestamp 1649977179
transform 1 0 15456 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1649977179
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_206
timestamp 1649977179
transform 1 0 20056 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_210
timestamp 1649977179
transform 1 0 20424 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_214
timestamp 1649977179
transform 1 0 20792 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_218
timestamp 1649977179
transform 1 0 21160 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_222
timestamp 1649977179
transform 1 0 21528 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_7
timestamp 1649977179
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_13
timestamp 1649977179
transform 1 0 2300 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_19
timestamp 1649977179
transform 1 0 2852 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_25
timestamp 1649977179
transform 1 0 3404 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_29
timestamp 1649977179
transform 1 0 3772 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_50
timestamp 1649977179
transform 1 0 5704 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 1649977179
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_66
timestamp 1649977179
transform 1 0 7176 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_71
timestamp 1649977179
transform 1 0 7636 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_104
timestamp 1649977179
transform 1 0 10672 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_109
timestamp 1649977179
transform 1 0 11132 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_129
timestamp 1649977179
transform 1 0 12972 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_140
timestamp 1649977179
transform 1 0 13984 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1649977179
transform 1 0 14996 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_155
timestamp 1649977179
transform 1 0 15364 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_166
timestamp 1649977179
transform 1 0 16376 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_185
timestamp 1649977179
transform 1 0 18124 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_210
timestamp 1649977179
transform 1 0 20424 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_214
timestamp 1649977179
transform 1 0 20792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_218
timestamp 1649977179
transform 1 0 21160 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1649977179
transform 1 0 1748 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_38
timestamp 1649977179
transform 1 0 4600 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_57
timestamp 1649977179
transform 1 0 6348 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_67
timestamp 1649977179
transform 1 0 7268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_78
timestamp 1649977179
transform 1 0 8280 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_82
timestamp 1649977179
transform 1 0 8648 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_101
timestamp 1649977179
transform 1 0 10396 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_106
timestamp 1649977179
transform 1 0 10856 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_110
timestamp 1649977179
transform 1 0 11224 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1649977179
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_131
timestamp 1649977179
transform 1 0 13156 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1649977179
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_26_157
timestamp 1649977179
transform 1 0 15548 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_168
timestamp 1649977179
transform 1 0 16560 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_172
timestamp 1649977179
transform 1 0 16928 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_190
timestamp 1649977179
transform 1 0 18584 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 1649977179
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_206
timestamp 1649977179
transform 1 0 20056 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_216
timestamp 1649977179
transform 1 0 20976 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_9
timestamp 1649977179
transform 1 0 1932 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_20
timestamp 1649977179
transform 1 0 2944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_38
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_44
timestamp 1649977179
transform 1 0 5152 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_54
timestamp 1649977179
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_61
timestamp 1649977179
transform 1 0 6716 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_79
timestamp 1649977179
transform 1 0 8372 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_83
timestamp 1649977179
transform 1 0 8740 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_87
timestamp 1649977179
transform 1 0 9108 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_98
timestamp 1649977179
transform 1 0 10120 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1649977179
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1649977179
transform 1 0 11776 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_127
timestamp 1649977179
transform 1 0 12788 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_138
timestamp 1649977179
transform 1 0 13800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_148
timestamp 1649977179
transform 1 0 14720 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_159
timestamp 1649977179
transform 1 0 15732 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_166
timestamp 1649977179
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_177
timestamp 1649977179
transform 1 0 17388 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_199
timestamp 1649977179
transform 1 0 19412 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_203
timestamp 1649977179
transform 1 0 19780 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_221
timestamp 1649977179
transform 1 0 21436 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_6
timestamp 1649977179
transform 1 0 1656 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_16
timestamp 1649977179
transform 1 0 2576 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_26
timestamp 1649977179
transform 1 0 3496 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_45
timestamp 1649977179
transform 1 0 5244 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_58
timestamp 1649977179
transform 1 0 6440 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_28_71
timestamp 1649977179
transform 1 0 7636 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_82
timestamp 1649977179
transform 1 0 8648 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_104
timestamp 1649977179
transform 1 0 10672 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_122
timestamp 1649977179
transform 1 0 12328 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_138
timestamp 1649977179
transform 1 0 13800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_150
timestamp 1649977179
transform 1 0 14904 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_178
timestamp 1649977179
transform 1 0 17480 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_183
timestamp 1649977179
transform 1 0 17940 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_194
timestamp 1649977179
transform 1 0 18952 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_200
timestamp 1649977179
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_205
timestamp 1649977179
transform 1 0 19964 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_210
timestamp 1649977179
transform 1 0 20424 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_215
timestamp 1649977179
transform 1 0 20884 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_220
timestamp 1649977179
transform 1 0 21344 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_5
timestamp 1649977179
transform 1 0 1564 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_25
timestamp 1649977179
transform 1 0 3404 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1649977179
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_61
timestamp 1649977179
transform 1 0 6716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_65
timestamp 1649977179
transform 1 0 7084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1649977179
transform 1 0 8648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_94
timestamp 1649977179
transform 1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_98
timestamp 1649977179
transform 1 0 10120 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1649977179
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_131
timestamp 1649977179
transform 1 0 13156 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1649977179
transform 1 0 14168 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_147
timestamp 1649977179
transform 1 0 14628 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_159
timestamp 1649977179
transform 1 0 15732 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_164
timestamp 1649977179
transform 1 0 16192 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_29_185
timestamp 1649977179
transform 1 0 18124 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_195
timestamp 1649977179
transform 1 0 19044 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_200
timestamp 1649977179
transform 1 0 19504 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_210
timestamp 1649977179
transform 1 0 20424 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_215
timestamp 1649977179
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_221
timestamp 1649977179
transform 1 0 21436 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_5
timestamp 1649977179
transform 1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_26
timestamp 1649977179
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_33
timestamp 1649977179
transform 1 0 4140 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_44
timestamp 1649977179
transform 1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_62
timestamp 1649977179
transform 1 0 6808 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_72
timestamp 1649977179
transform 1 0 7728 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_82
timestamp 1649977179
transform 1 0 8648 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_87
timestamp 1649977179
transform 1 0 9108 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_98
timestamp 1649977179
transform 1 0 10120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_102
timestamp 1649977179
transform 1 0 10488 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1649977179
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_115
timestamp 1649977179
transform 1 0 11684 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_125
timestamp 1649977179
transform 1 0 12604 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_135
timestamp 1649977179
transform 1 0 13524 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_160
timestamp 1649977179
transform 1 0 15824 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_169
timestamp 1649977179
transform 1 0 16652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_178
timestamp 1649977179
transform 1 0 17480 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_183
timestamp 1649977179
transform 1 0 17940 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_188
timestamp 1649977179
transform 1 0 18400 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_193
timestamp 1649977179
transform 1 0 18860 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_200
timestamp 1649977179
transform 1 0 19504 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_205
timestamp 1649977179
transform 1 0 19964 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_214
timestamp 1649977179
transform 1 0 20792 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_220
timestamp 1649977179
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_13
timestamp 1649977179
transform 1 0 2300 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_32
timestamp 1649977179
transform 1 0 4048 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_38
timestamp 1649977179
transform 1 0 4600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_42
timestamp 1649977179
transform 1 0 4968 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_52
timestamp 1649977179
transform 1 0 5888 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_63
timestamp 1649977179
transform 1 0 6900 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1649977179
transform 1 0 7912 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1649977179
transform 1 0 8924 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_89
timestamp 1649977179
transform 1 0 9292 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 1649977179
transform 1 0 10856 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_110
timestamp 1649977179
transform 1 0 11224 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_124
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_130
timestamp 1649977179
transform 1 0 13064 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_135
timestamp 1649977179
transform 1 0 13524 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_140
timestamp 1649977179
transform 1 0 13984 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_144
timestamp 1649977179
transform 1 0 14352 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_154
timestamp 1649977179
transform 1 0 15272 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_159
timestamp 1649977179
transform 1 0 15732 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1649977179
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_172
timestamp 1649977179
transform 1 0 16928 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_177
timestamp 1649977179
transform 1 0 17388 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_182
timestamp 1649977179
transform 1 0 17848 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_187
timestamp 1649977179
transform 1 0 18308 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_192
timestamp 1649977179
transform 1 0 18768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_197
timestamp 1649977179
transform 1 0 19228 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_202
timestamp 1649977179
transform 1 0 19688 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_31_210
timestamp 1649977179
transform 1 0 20424 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 1649977179
transform 1 0 20976 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_221
timestamp 1649977179
transform 1 0 21436 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_14
timestamp 1649977179
transform 1 0 2392 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_26
timestamp 1649977179
transform 1 0 3496 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_45
timestamp 1649977179
transform 1 0 5244 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_32_64
timestamp 1649977179
transform 1 0 6992 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_82
timestamp 1649977179
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_95
timestamp 1649977179
transform 1 0 9844 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_113
timestamp 1649977179
transform 1 0 11500 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_123
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_138
timestamp 1649977179
transform 1 0 13800 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_144
timestamp 1649977179
transform 1 0 14352 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_149
timestamp 1649977179
transform 1 0 14812 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_154
timestamp 1649977179
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_160
timestamp 1649977179
transform 1 0 15824 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_169
timestamp 1649977179
transform 1 0 16652 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_175
timestamp 1649977179
transform 1 0 17204 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_180
timestamp 1649977179
transform 1 0 17664 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_184
timestamp 1649977179
transform 1 0 18032 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_190
timestamp 1649977179
transform 1 0 18584 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_194
timestamp 1649977179
transform 1 0 18952 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_199
timestamp 1649977179
transform 1 0 19412 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_14
timestamp 1649977179
transform 1 0 2392 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_26
timestamp 1649977179
transform 1 0 3496 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_43
timestamp 1649977179
transform 1 0 5060 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1649977179
transform 1 0 6532 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_73
timestamp 1649977179
transform 1 0 7820 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_82
timestamp 1649977179
transform 1 0 8648 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1649977179
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_33_109
timestamp 1649977179
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_33_121
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_127
timestamp 1649977179
transform 1 0 12788 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_135
timestamp 1649977179
transform 1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_139
timestamp 1649977179
transform 1 0 13892 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_145
timestamp 1649977179
transform 1 0 14444 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_151
timestamp 1649977179
transform 1 0 14996 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_157
timestamp 1649977179
transform 1 0 15548 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1649977179
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_173
timestamp 1649977179
transform 1 0 17020 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1649977179
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_185
timestamp 1649977179
transform 1 0 18124 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_191
timestamp 1649977179
transform 1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_195
timestamp 1649977179
transform 1 0 19044 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_201
timestamp 1649977179
transform 1 0 19596 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_207
timestamp 1649977179
transform 1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_221
timestamp 1649977179
transform 1 0 21436 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 8832 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 13984 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  _068_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 3864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1649977179
transform -1 0 2576 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1649977179
transform 1 0 6440 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1649977179
transform 1 0 4784 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1649977179
transform -1 0 2116 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1649977179
transform -1 0 1748 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1649977179
transform -1 0 2116 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1649977179
transform -1 0 3496 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1649977179
transform 1 0 13248 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1649977179
transform -1 0 3036 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1649977179
transform -1 0 4692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1649977179
transform 1 0 14996 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1649977179
transform 1 0 18492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1649977179
transform 1 0 16008 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1649977179
transform 1 0 17572 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1649977179
transform 1 0 19412 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1649977179
transform 1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1649977179
transform 1 0 20608 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform 1 0 19688 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1649977179
transform 1 0 18584 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform 1 0 20148 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1649977179
transform 1 0 20148 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform 1 0 21160 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1649977179
transform 1 0 21068 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 18952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1649977179
transform -1 0 19504 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1649977179
transform -1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 20792 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1649977179
transform 1 0 20976 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_mem_left_track_1.prog_clk .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13616 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform -1 0 7084 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform -1 0 9660 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform -1 0 12236 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_mem_left_track_1.prog_clk
timestamp 1649977179
transform 1 0 15640 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12604 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1649977179
transform -1 0 8188 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1649977179
transform 1 0 6992 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1649977179
transform -1 0 8648 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1649977179
transform 1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold7
timestamp 1649977179
transform -1 0 7084 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1649977179
transform 1 0 14720 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold9
timestamp 1649977179
transform 1 0 13156 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold10
timestamp 1649977179
transform -1 0 6164 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1649977179
transform 1 0 12788 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1649977179
transform -1 0 17112 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1649977179
transform 1 0 9476 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1649977179
transform -1 0 10396 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1649977179
transform -1 0 6072 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1649977179
transform -1 0 7728 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1649977179
transform 1 0 17664 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1649977179
transform 1 0 10304 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1649977179
transform 1 0 9936 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1649977179
transform 1 0 13984 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1649977179
transform -1 0 13524 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1649977179
transform 1 0 9016 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1649977179
transform 1 0 3956 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1649977179
transform -1 0 8648 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1649977179
transform -1 0 4048 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold27
timestamp 1649977179
transform -1 0 14996 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold28
timestamp 1649977179
transform 1 0 16744 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold29
timestamp 1649977179
transform 1 0 20240 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold30
timestamp 1649977179
transform -1 0 2484 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold31
timestamp 1649977179
transform -1 0 8648 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold32
timestamp 1649977179
transform 1 0 19320 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold33
timestamp 1649977179
transform 1 0 18952 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold34
timestamp 1649977179
transform 1 0 11684 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold35
timestamp 1649977179
transform -1 0 11316 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold36
timestamp 1649977179
transform -1 0 2484 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold37
timestamp 1649977179
transform -1 0 3496 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold38
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold39
timestamp 1649977179
transform -1 0 3404 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold40
timestamp 1649977179
transform -1 0 5060 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold41
timestamp 1649977179
transform 1 0 19872 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold42
timestamp 1649977179
transform -1 0 6072 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold43
timestamp 1649977179
transform 1 0 16744 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold44
timestamp 1649977179
transform -1 0 11224 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold45
timestamp 1649977179
transform -1 0 3496 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold46
timestamp 1649977179
transform 1 0 18308 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold47
timestamp 1649977179
transform -1 0 12512 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold48
timestamp 1649977179
transform -1 0 6072 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold49
timestamp 1649977179
transform 1 0 13156 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold50
timestamp 1649977179
transform 1 0 6716 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold51
timestamp 1649977179
transform 1 0 6532 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold52
timestamp 1649977179
transform -1 0 9936 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold53
timestamp 1649977179
transform 1 0 1932 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold54
timestamp 1649977179
transform -1 0 2576 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold55
timestamp 1649977179
transform 1 0 5520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold56
timestamp 1649977179
transform -1 0 8648 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold57
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold58
timestamp 1649977179
transform 1 0 2668 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold59
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold60
timestamp 1649977179
transform 1 0 9936 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold61
timestamp 1649977179
transform -1 0 15088 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform 1 0 21160 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 2116 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform -1 0 1656 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform -1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1656 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 2116 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 4232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 1656 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 2576 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 2576 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 1656 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 3496 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 3036 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 2116 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 2576 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1649977179
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 3036 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 4140 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 8004 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1649977179
transform -1 0 8648 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1649977179
transform -1 0 9108 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform 1 0 20148 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1649977179
transform 1 0 10764 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 19228 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1649977179
transform 1 0 17112 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 16008 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform -1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 14352 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 12512 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 1656 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform -1 0 4140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform -1 0 2852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 12328 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 12512 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform -1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1649977179
transform -1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input45
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input46
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input47
timestamp 1649977179
transform -1 0 2300 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input48
timestamp 1649977179
transform -1 0 3404 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input49
timestamp 1649977179
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input50
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1649977179
transform 1 0 4232 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1649977179
transform -1 0 2300 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input54
timestamp 1649977179
transform -1 0 2392 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input55
timestamp 1649977179
transform -1 0 2392 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input56
timestamp 1649977179
transform 1 0 2576 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1649977179
transform -1 0 3496 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform 1 0 3772 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1649977179
transform -1 0 21436 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18124 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4140 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_1.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 3312 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2024 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 3220 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_3.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 4140 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5244 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_5.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7176 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 9476 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_7.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 7084 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7820 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_9.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 7360 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7268 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_11.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_13.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10396 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_15.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9200 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 10856 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_17.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 11500 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_19.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8648 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7176 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_21.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 8372 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 7084 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_23.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 7820 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 7544 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_25.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5152 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4416 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_27.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5796 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_29.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6072 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_31.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6072 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 5336 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_33.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 6992 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5244 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_35.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4048 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 5244 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_37.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 4600 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 2760 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_left_track_39.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 5244 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 21436 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_0.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 14076 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15548 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15088 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_2.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform -1 0 18124 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 15824 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 13156 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_4.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 10856 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11592 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_6.sky130_fd_sc_hd__dfxtp_1_2_
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 12972 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_8.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 11224 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 10120 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_10.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_12.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 12880 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_14.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 15824 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 14720 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_16.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 14904 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 15732 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_18.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 18124 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 17112 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_20.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform -1 0 19412 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform 1 0 18492 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_22.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 18032 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 19136 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_24.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 17296 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_0_
timestamp 1649977179
transform -1 0 18768 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  mem_top_track_26.sky130_fd_sc_hd__dfxtp_1_1_
timestamp 1649977179
transform 1 0 15640 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_0_ .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4324 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_1_
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l1_in_2_
timestamp 1649977179
transform 1 0 2944 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l2_in_1_
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_1.mux_l2_in_1__124 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_1.mux_l3_in_0_
timestamp 1649977179
transform -1 0 2484 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_1.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_0_
timestamp 1649977179
transform 1 0 4876 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l1_in_1_
timestamp 1649977179
transform -1 0 5060 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_3.mux_l2_in_1__101
timestamp 1649977179
transform -1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l2_in_1_
timestamp 1649977179
transform 1 0 4140 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_3.mux_l3_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_3.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_1_
timestamp 1649977179
transform 1 0 8096 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l1_in_2_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7636 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_5.mux_l2_in_1__107
timestamp 1649977179
transform 1 0 8280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l2_in_1_
timestamp 1649977179
transform 1 0 6992 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_5.mux_l3_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_5.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3036 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9752 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l1_in_1_
timestamp 1649977179
transform -1 0 8096 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_7.mux_l2_in_1__108
timestamp 1649977179
transform 1 0 8372 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l2_in_1_
timestamp 1649977179
transform -1 0 6072 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_7.mux_l3_in_0_
timestamp 1649977179
transform 1 0 6256 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_7.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_9.mux_l1_in_1__109
timestamp 1649977179
transform 1 0 9016 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l1_in_1_
timestamp 1649977179
transform -1 0 7636 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_9.mux_l2_in_0_
timestamp 1649977179
transform 1 0 7728 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_9.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2760 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7912 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_11.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6900 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_11.mux_l2_in_0__125
timestamp 1649977179
transform 1 0 9016 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_11.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9660 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_13.mux_l2_in_0__126
timestamp 1649977179
transform 1 0 10856 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_13.mux_l2_in_0_
timestamp 1649977179
transform 1 0 9844 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_13.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l1_in_0_
timestamp 1649977179
transform -1 0 10120 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_15.mux_l2_in_0_
timestamp 1649977179
transform 1 0 10304 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_15.mux_l2_in_0__127
timestamp 1649977179
transform -1 0 10120 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_15.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2208 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l1_in_0_
timestamp 1649977179
transform -1 0 9844 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_17.mux_l2_in_0_
timestamp 1649977179
transform -1 0 10120 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_17.mux_l2_in_0__128
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_17.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12512 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l1_in_0_
timestamp 1649977179
transform 1 0 8096 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_19.mux_l2_in_0_
timestamp 1649977179
transform -1 0 7912 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_19.mux_l2_in_0__129
timestamp 1649977179
transform 1 0 17664 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_19.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7452 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_21.mux_l2_in_0_
timestamp 1649977179
transform 1 0 6808 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_21.mux_l2_in_0__130
timestamp 1649977179
transform 1 0 10580 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_21.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 3128 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l1_in_0_
timestamp 1649977179
transform 1 0 7268 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_23.mux_l2_in_0__131
timestamp 1649977179
transform 1 0 8004 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_23.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_23.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2024 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l1_in_1_
timestamp 1649977179
transform 1 0 5336 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_25.mux_l1_in_1__132
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_25.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4324 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_25.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2760 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_27.mux_l2_in_0__133
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_27.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4232 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_27.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l1_in_0_
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_29.mux_l2_in_0_
timestamp 1649977179
transform 1 0 4876 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_29.mux_l2_in_0__134
timestamp 1649977179
transform -1 0 2668 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_29.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5612 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_31.mux_l2_in_0_
timestamp 1649977179
transform 1 0 5060 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_31.mux_l2_in_0__102
timestamp 1649977179
transform -1 0 3496 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_31.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l1_in_0_
timestamp 1649977179
transform 1 0 5244 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_33.mux_l2_in_0_
timestamp 1649977179
transform -1 0 5152 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_33.mux_l2_in_0__103
timestamp 1649977179
transform -1 0 3496 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_33.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_35.mux_l2_in_0_
timestamp 1649977179
transform -1 0 3496 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_35.mux_l2_in_0__104
timestamp 1649977179
transform 1 0 10580 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_35.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 7636 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_37.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2116 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_37.mux_l2_in_0__105
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_37.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2116 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l1_in_0_
timestamp 1649977179
transform 1 0 3496 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_left_track_39.mux_l2_in_0_
timestamp 1649977179
transform 1 0 2668 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_left_track_39.mux_l2_in_0__106
timestamp 1649977179
transform -1 0 2392 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_left_track_39.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 2576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_0_
timestamp 1649977179
transform 1 0 13064 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_1_
timestamp 1649977179
transform 1 0 14168 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l1_in_2_
timestamp 1649977179
transform -1 0 13800 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13800 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_0.mux_l2_in_1__110
timestamp 1649977179
transform 1 0 15088 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l2_in_1_
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_0.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13984 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_0.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14812 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_0_
timestamp 1649977179
transform -1 0 15732 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l1_in_1_
timestamp 1649977179
transform 1 0 15732 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_0_
timestamp 1649977179
transform 1 0 14904 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_2.mux_l2_in_1__116
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l2_in_1_
timestamp 1649977179
transform -1 0 14904 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_2.mux_l3_in_0_
timestamp 1649977179
transform -1 0 15272 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_2.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18308 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_0_
timestamp 1649977179
transform 1 0 12972 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_1_
timestamp 1649977179
transform 1 0 13340 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l1_in_2_
timestamp 1649977179
transform 1 0 11960 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_0_
timestamp 1649977179
transform 1 0 12512 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l2_in_1_
timestamp 1649977179
transform -1 0 12604 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_4.mux_l2_in_1__121
timestamp 1649977179
transform 1 0 13524 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_4.mux_l3_in_0_
timestamp 1649977179
transform -1 0 13156 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_4.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13984 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11316 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l1_in_1_
timestamp 1649977179
transform 1 0 11316 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l2_in_1_
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_6.mux_l2_in_1__122
timestamp 1649977179
transform 1 0 12420 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_6.mux_l3_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_6.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_0_
timestamp 1649977179
transform 1 0 11776 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_8.mux_l1_in_1__123
timestamp 1649977179
transform 1 0 10948 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l1_in_1_
timestamp 1649977179
transform -1 0 10212 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_8.mux_l2_in_0_
timestamp 1649977179
transform -1 0 11224 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_8.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 15732 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l1_in_0_
timestamp 1649977179
transform -1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_10.mux_l2_in_0__111
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_10.mux_l2_in_0_
timestamp 1649977179
transform -1 0 13248 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_10.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 13800 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l1_in_0_
timestamp 1649977179
transform -1 0 14904 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_12.mux_l2_in_0__112
timestamp 1649977179
transform -1 0 13800 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_12.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15364 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_12.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 17940 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l1_in_0_
timestamp 1649977179
transform 1 0 15364 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_14.mux_l2_in_0__113
timestamp 1649977179
transform 1 0 15824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_14.mux_l2_in_0_
timestamp 1649977179
transform -1 0 15640 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_14.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19228 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l1_in_0_
timestamp 1649977179
transform -1 0 17480 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_16.mux_l2_in_0__114
timestamp 1649977179
transform -1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_16.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18216 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_16.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l1_in_0_
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_18.mux_l2_in_0__115
timestamp 1649977179
transform 1 0 16100 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_18.mux_l2_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_18.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform 1 0 21160 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_20.mux_l2_in_0__117
timestamp 1649977179
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_20.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18952 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_20.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19504 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l1_in_0_
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_22.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18492 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_22.mux_l2_in_0__118
timestamp 1649977179
transform 1 0 18400 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_22.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 19964 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_0_
timestamp 1649977179
transform 1 0 17480 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_24.mux_l1_in_1__119
timestamp 1649977179
transform -1 0 18676 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l1_in_1_
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_24.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18216 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_24.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 21068 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l1_in_0_
timestamp 1649977179
transform -1 0 16376 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__conb_1  mux_top_track_26.mux_l2_in_0__120
timestamp 1649977179
transform 1 0 18308 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  mux_top_track_26.mux_l2_in_0_
timestamp 1649977179
transform -1 0 18124 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  mux_top_track_26.sky130_fd_sc_hd__buf_4_0_
timestamp 1649977179
transform -1 0 18952 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output60 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11960 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output61
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output62
timestamp 1649977179
transform -1 0 2300 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output63
timestamp 1649977179
transform -1 0 2300 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output64
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1649977179
transform 1 0 1932 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1649977179
transform -1 0 1932 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1649977179
transform -1 0 5152 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1649977179
transform 1 0 6532 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1649977179
transform 1 0 8924 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1649977179
transform -1 0 1748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1649977179
transform -1 0 2300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1649977179
transform -1 0 2300 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1649977179
transform -1 0 3404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1649977179
transform 1 0 3036 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1649977179
transform -1 0 13524 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1649977179
transform -1 0 18676 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1649977179
transform -1 0 18584 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1649977179
transform -1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1649977179
transform -1 0 20148 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1649977179
transform 1 0 19596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1649977179
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1649977179
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1649977179
transform 1 0 20976 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1649977179
transform -1 0 20792 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1649977179
transform -1 0 14444 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1649977179
transform -1 0 14996 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1649977179
transform -1 0 15548 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1649977179
transform -1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1649977179
transform -1 0 15824 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output97
timestamp 1649977179
transform -1 0 17020 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1649977179
transform -1 0 17572 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform -1 0 17204 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform -1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  prog_clk_0_FTB00 .volare/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21436 0 1 19584
box -38 -48 1142 592
<< labels >>
rlabel metal4 s 6142 2128 6462 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 11340 2128 11660 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 16538 2128 16858 20720 6 VGND
port 0 nsew ground input
rlabel metal4 s 3543 2128 3863 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 8741 2128 9061 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 13939 2128 14259 20720 6 VPWR
port 1 nsew power input
rlabel metal4 s 19137 2128 19457 20720 6 VPWR
port 1 nsew power input
rlabel metal3 s 22200 11432 23000 11552 6 ccff_head
port 2 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 ccff_tail
port 3 nsew signal tristate
rlabel metal3 s 0 4360 800 4480 6 chanx_left_in[0]
port 4 nsew signal input
rlabel metal3 s 0 8984 800 9104 6 chanx_left_in[10]
port 5 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 chanx_left_in[11]
port 6 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 chanx_left_in[12]
port 7 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 chanx_left_in[13]
port 8 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 chanx_left_in[14]
port 9 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 chanx_left_in[15]
port 10 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 chanx_left_in[16]
port 11 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 chanx_left_in[17]
port 12 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 chanx_left_in[18]
port 13 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 chanx_left_in[19]
port 14 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 chanx_left_in[1]
port 15 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 chanx_left_in[2]
port 16 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 chanx_left_in[3]
port 17 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 chanx_left_in[4]
port 18 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 chanx_left_in[5]
port 19 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 chanx_left_in[6]
port 20 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 chanx_left_in[7]
port 21 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 chanx_left_in[8]
port 22 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 chanx_left_in[9]
port 23 nsew signal input
rlabel metal3 s 0 13744 800 13864 6 chanx_left_out[0]
port 24 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 chanx_left_out[10]
port 25 nsew signal tristate
rlabel metal3 s 0 18776 800 18896 6 chanx_left_out[11]
port 26 nsew signal tristate
rlabel metal3 s 0 19320 800 19440 6 chanx_left_out[12]
port 27 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 chanx_left_out[13]
port 28 nsew signal tristate
rlabel metal3 s 0 20272 800 20392 6 chanx_left_out[14]
port 29 nsew signal tristate
rlabel metal3 s 0 20680 800 20800 6 chanx_left_out[15]
port 30 nsew signal tristate
rlabel metal3 s 0 21224 800 21344 6 chanx_left_out[16]
port 31 nsew signal tristate
rlabel metal3 s 0 21632 800 21752 6 chanx_left_out[17]
port 32 nsew signal tristate
rlabel metal3 s 0 22176 800 22296 6 chanx_left_out[18]
port 33 nsew signal tristate
rlabel metal3 s 0 22584 800 22704 6 chanx_left_out[19]
port 34 nsew signal tristate
rlabel metal3 s 0 14152 800 14272 6 chanx_left_out[1]
port 35 nsew signal tristate
rlabel metal3 s 0 14560 800 14680 6 chanx_left_out[2]
port 36 nsew signal tristate
rlabel metal3 s 0 15104 800 15224 6 chanx_left_out[3]
port 37 nsew signal tristate
rlabel metal3 s 0 15512 800 15632 6 chanx_left_out[4]
port 38 nsew signal tristate
rlabel metal3 s 0 16056 800 16176 6 chanx_left_out[5]
port 39 nsew signal tristate
rlabel metal3 s 0 16464 800 16584 6 chanx_left_out[6]
port 40 nsew signal tristate
rlabel metal3 s 0 17008 800 17128 6 chanx_left_out[7]
port 41 nsew signal tristate
rlabel metal3 s 0 17416 800 17536 6 chanx_left_out[8]
port 42 nsew signal tristate
rlabel metal3 s 0 17960 800 18080 6 chanx_left_out[9]
port 43 nsew signal tristate
rlabel metal2 s 3882 22200 3938 23000 6 chany_top_in[0]
port 44 nsew signal input
rlabel metal2 s 8482 22200 8538 23000 6 chany_top_in[10]
port 45 nsew signal input
rlabel metal2 s 8942 22200 8998 23000 6 chany_top_in[11]
port 46 nsew signal input
rlabel metal2 s 9402 22200 9458 23000 6 chany_top_in[12]
port 47 nsew signal input
rlabel metal2 s 9862 22200 9918 23000 6 chany_top_in[13]
port 48 nsew signal input
rlabel metal2 s 10322 22200 10378 23000 6 chany_top_in[14]
port 49 nsew signal input
rlabel metal2 s 10782 22200 10838 23000 6 chany_top_in[15]
port 50 nsew signal input
rlabel metal2 s 11242 22200 11298 23000 6 chany_top_in[16]
port 51 nsew signal input
rlabel metal2 s 11702 22200 11758 23000 6 chany_top_in[17]
port 52 nsew signal input
rlabel metal2 s 12162 22200 12218 23000 6 chany_top_in[18]
port 53 nsew signal input
rlabel metal2 s 12622 22200 12678 23000 6 chany_top_in[19]
port 54 nsew signal input
rlabel metal2 s 4342 22200 4398 23000 6 chany_top_in[1]
port 55 nsew signal input
rlabel metal2 s 4802 22200 4858 23000 6 chany_top_in[2]
port 56 nsew signal input
rlabel metal2 s 5262 22200 5318 23000 6 chany_top_in[3]
port 57 nsew signal input
rlabel metal2 s 5722 22200 5778 23000 6 chany_top_in[4]
port 58 nsew signal input
rlabel metal2 s 6182 22200 6238 23000 6 chany_top_in[5]
port 59 nsew signal input
rlabel metal2 s 6642 22200 6698 23000 6 chany_top_in[6]
port 60 nsew signal input
rlabel metal2 s 7102 22200 7158 23000 6 chany_top_in[7]
port 61 nsew signal input
rlabel metal2 s 7562 22200 7618 23000 6 chany_top_in[8]
port 62 nsew signal input
rlabel metal2 s 8022 22200 8078 23000 6 chany_top_in[9]
port 63 nsew signal input
rlabel metal2 s 13082 22200 13138 23000 6 chany_top_out[0]
port 64 nsew signal tristate
rlabel metal2 s 17682 22200 17738 23000 6 chany_top_out[10]
port 65 nsew signal tristate
rlabel metal2 s 18142 22200 18198 23000 6 chany_top_out[11]
port 66 nsew signal tristate
rlabel metal2 s 18602 22200 18658 23000 6 chany_top_out[12]
port 67 nsew signal tristate
rlabel metal2 s 19062 22200 19118 23000 6 chany_top_out[13]
port 68 nsew signal tristate
rlabel metal2 s 19522 22200 19578 23000 6 chany_top_out[14]
port 69 nsew signal tristate
rlabel metal2 s 19982 22200 20038 23000 6 chany_top_out[15]
port 70 nsew signal tristate
rlabel metal2 s 20442 22200 20498 23000 6 chany_top_out[16]
port 71 nsew signal tristate
rlabel metal2 s 20902 22200 20958 23000 6 chany_top_out[17]
port 72 nsew signal tristate
rlabel metal2 s 21362 22200 21418 23000 6 chany_top_out[18]
port 73 nsew signal tristate
rlabel metal2 s 21822 22200 21878 23000 6 chany_top_out[19]
port 74 nsew signal tristate
rlabel metal2 s 13542 22200 13598 23000 6 chany_top_out[1]
port 75 nsew signal tristate
rlabel metal2 s 14002 22200 14058 23000 6 chany_top_out[2]
port 76 nsew signal tristate
rlabel metal2 s 14462 22200 14518 23000 6 chany_top_out[3]
port 77 nsew signal tristate
rlabel metal2 s 14922 22200 14978 23000 6 chany_top_out[4]
port 78 nsew signal tristate
rlabel metal2 s 15382 22200 15438 23000 6 chany_top_out[5]
port 79 nsew signal tristate
rlabel metal2 s 15842 22200 15898 23000 6 chany_top_out[6]
port 80 nsew signal tristate
rlabel metal2 s 16302 22200 16358 23000 6 chany_top_out[7]
port 81 nsew signal tristate
rlabel metal2 s 16762 22200 16818 23000 6 chany_top_out[8]
port 82 nsew signal tristate
rlabel metal2 s 17222 22200 17278 23000 6 chany_top_out[9]
port 83 nsew signal tristate
rlabel metal3 s 0 2456 800 2576 6 left_bottom_grid_pin_11_
port 84 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 left_bottom_grid_pin_13_
port 85 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 left_bottom_grid_pin_15_
port 86 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 left_bottom_grid_pin_17_
port 87 nsew signal input
rlabel metal3 s 0 144 800 264 6 left_bottom_grid_pin_1_
port 88 nsew signal input
rlabel metal3 s 0 552 800 672 6 left_bottom_grid_pin_3_
port 89 nsew signal input
rlabel metal3 s 0 960 800 1080 6 left_bottom_grid_pin_5_
port 90 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 left_bottom_grid_pin_7_
port 91 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 left_bottom_grid_pin_9_
port 92 nsew signal input
rlabel metal2 s 22282 22200 22338 23000 6 prog_clk_0_N_in
port 93 nsew signal input
rlabel metal2 s 202 22200 258 23000 6 top_left_grid_pin_42_
port 94 nsew signal input
rlabel metal2 s 662 22200 718 23000 6 top_left_grid_pin_43_
port 95 nsew signal input
rlabel metal2 s 1122 22200 1178 23000 6 top_left_grid_pin_44_
port 96 nsew signal input
rlabel metal2 s 1582 22200 1638 23000 6 top_left_grid_pin_45_
port 97 nsew signal input
rlabel metal2 s 2042 22200 2098 23000 6 top_left_grid_pin_46_
port 98 nsew signal input
rlabel metal2 s 2502 22200 2558 23000 6 top_left_grid_pin_47_
port 99 nsew signal input
rlabel metal2 s 2962 22200 3018 23000 6 top_left_grid_pin_48_
port 100 nsew signal input
rlabel metal2 s 3422 22200 3478 23000 6 top_left_grid_pin_49_
port 101 nsew signal input
rlabel metal2 s 22742 22200 22798 23000 6 top_right_grid_pin_1_
port 102 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 23000 23000
<< end >>
