magic
tech sky130A
magscale 1 2
timestamp 1650894385
<< obsli1 >>
rect 1104 2159 10856 11441
<< obsm1 >>
rect 750 2128 11210 11472
<< metal2 >>
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6734 0 6790 800
rect 8206 0 8262 800
rect 9678 0 9734 800
rect 11150 0 11206 800
<< obsm2 >>
rect 756 856 11204 11472
rect 866 800 2170 856
rect 2338 800 3642 856
rect 3810 800 5114 856
rect 5282 800 6678 856
rect 6846 800 8150 856
rect 8318 800 9622 856
rect 9790 800 11094 856
<< obsm3 >>
rect 2168 2143 9832 11457
<< metal4 >>
rect 2168 2128 2488 11472
rect 3392 2128 3712 11472
rect 4616 2128 4936 11472
rect 5840 2128 6160 11472
rect 7064 2128 7384 11472
rect 8288 2128 8608 11472
rect 9512 2128 9832 11472
<< labels >>
rlabel metal4 s 3392 2128 3712 11472 6 VGND
port 1 nsew ground input
rlabel metal4 s 5840 2128 6160 11472 6 VGND
port 1 nsew ground input
rlabel metal4 s 8288 2128 8608 11472 6 VGND
port 1 nsew ground input
rlabel metal4 s 2168 2128 2488 11472 6 VPWR
port 2 nsew power input
rlabel metal4 s 4616 2128 4936 11472 6 VPWR
port 2 nsew power input
rlabel metal4 s 7064 2128 7384 11472 6 VPWR
port 2 nsew power input
rlabel metal4 s 9512 2128 9832 11472 6 VPWR
port 2 nsew power input
rlabel metal2 s 754 0 810 800 6 x[0]
port 3 nsew signal output
rlabel metal2 s 2226 0 2282 800 6 x[1]
port 4 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 x[2]
port 5 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 x[3]
port 6 nsew signal output
rlabel metal2 s 6734 0 6790 800 6 x[4]
port 7 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 x[5]
port 8 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 x[6]
port 9 nsew signal output
rlabel metal2 s 11150 0 11206 800 6 x[7]
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 12000 14000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 113050
string GDS_FILE /home/karim/work/ef/clear-harden/openlane/tie_array/runs/22_04_25_15_46/results/signoff/tie_array.magic.gds
string GDS_START 23752
<< end >>

